// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_108 written by SynthGen on 2021/04/05 11:08:34
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_108 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n983, n995, n984, n974, n967, n1008, n962, n965,
 n1015, n993, n988, n981, n1003, n973, n989, n970,
 n1021, n1029, n1025, n1023, n1026, n1032, n1022, n1020,
 n1027, n1017, n1024, n1030, n1019, n1018, n1028, n1031);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n983, n995, n984, n974, n967, n1008, n962, n965,
 n1015, n993, n988, n981, n1003, n973, n989, n970,
 n1021, n1029, n1025, n1023, n1026, n1032, n1022, n1020,
 n1027, n1017, n1024, n1030, n1019, n1018, n1028, n1031;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n963, n964, n966, n968, n969, n971, n972,
 n975, n976, n977, n978, n979, n980, n982, n985,
 n986, n987, n990, n991, n992, n994, n996, n997,
 n998, n999, n1000, n1001, n1002, n1004, n1005, n1006,
 n1007, n1009, n1010, n1011, n1012, n1013, n1014, n1016;

not  g0 (n138, n7);
not  g1 (n109, n13);
buf  g2 (n79, n2);
buf  g3 (n64, n25);
buf  g4 (n99, n25);
not  g5 (n56, n4);
not  g6 (n67, n17);
buf  g7 (n40, n12);
buf  g8 (n103, n2);
buf  g9 (n121, n3);
buf  g10 (n115, n16);
buf  g11 (n135, n11);
not  g12 (n89, n27);
not  g13 (n52, n21);
not  g14 (n33, n17);
not  g15 (n133, n13);
buf  g16 (n34, n11);
not  g17 (n119, n5);
buf  g18 (n141, n9);
buf  g19 (n134, n20);
not  g20 (n118, n18);
buf  g21 (n108, n15);
not  g22 (n49, n19);
not  g23 (n57, n8);
not  g24 (n102, n7);
not  g25 (n116, n24);
buf  g26 (n75, n10);
buf  g27 (n36, n14);
not  g28 (n53, n1);
buf  g29 (n94, n6);
not  g30 (n85, n22);
buf  g31 (n107, n24);
not  g32 (n101, n15);
buf  g33 (n58, n10);
buf  g34 (n87, n15);
not  g35 (n143, n21);
not  g36 (n106, n14);
not  g37 (n100, n27);
buf  g38 (n93, n26);
not  g39 (n44, n6);
buf  g40 (n105, n18);
not  g41 (n110, n8);
buf  g42 (n111, n22);
buf  g43 (n77, n13);
buf  g44 (n68, n5);
not  g45 (n66, n2);
buf  g46 (n139, n28);
not  g47 (n114, n17);
not  g48 (n80, n1);
buf  g49 (n144, n25);
not  g50 (n126, n1);
buf  g51 (n54, n16);
buf  g52 (n86, n22);
not  g53 (n129, n23);
not  g54 (n39, n5);
buf  g55 (n62, n10);
not  g56 (n45, n15);
buf  g57 (n117, n24);
not  g58 (n69, n25);
not  g59 (n124, n21);
buf  g60 (n51, n2);
buf  g61 (n78, n26);
not  g62 (n43, n6);
not  g63 (n55, n8);
buf  g64 (n84, n6);
buf  g65 (n35, n18);
buf  g66 (n73, n27);
buf  g67 (n96, n16);
not  g68 (n104, n24);
buf  g69 (n70, n28);
not  g70 (n81, n10);
buf  g71 (n98, n14);
buf  g72 (n130, n22);
buf  g73 (n38, n26);
not  g74 (n48, n3);
not  g75 (n74, n9);
buf  g76 (n59, n3);
buf  g77 (n92, n8);
buf  g78 (n131, n4);
buf  g79 (n97, n17);
not  g80 (n60, n28);
not  g81 (n65, n12);
buf  g82 (n136, n12);
not  g83 (n132, n4);
not  g84 (n112, n12);
not  g85 (n137, n20);
not  g86 (n91, n11);
buf  g87 (n122, n4);
not  g88 (n127, n18);
not  g89 (n71, n13);
buf  g90 (n95, n20);
not  g91 (n123, n19);
not  g92 (n113, n9);
not  g93 (n42, n5);
not  g94 (n125, n14);
not  g95 (n47, n19);
buf  g96 (n140, n21);
not  g97 (n76, n1);
buf  g98 (n37, n23);
buf  g99 (n128, n11);
not  g100 (n41, n23);
buf  g101 (n142, n9);
buf  g102 (n72, n19);
buf  g103 (n61, n23);
not  g104 (n63, n26);
not  g105 (n46, n20);
buf  g106 (n120, n28);
buf  g107 (n88, n7);
buf  g108 (n90, n16);
not  g109 (n83, n7);
buf  g110 (n82, n27);
not  g111 (n50, n3);
buf  g112 (n236, n56);
buf  g113 (n201, n74);
not  g114 (n248, n58);
not  g115 (n149, n70);
not  g116 (n309, n75);
not  g117 (n184, n36);
buf  g118 (n209, n57);
buf  g119 (n171, n31);
buf  g120 (n163, n71);
buf  g121 (n237, n50);
buf  g122 (n241, n34);
not  g123 (n294, n52);
buf  g124 (n207, n64);
not  g125 (n316, n42);
buf  g126 (n159, n70);
not  g127 (n203, n45);
buf  g128 (n175, n49);
buf  g129 (n273, n39);
not  g130 (n205, n65);
buf  g131 (n307, n60);
not  g132 (n177, n29);
buf  g133 (n188, n66);
not  g134 (n311, n45);
not  g135 (n225, n41);
buf  g136 (n257, n60);
buf  g137 (n280, n62);
not  g138 (n252, n73);
buf  g139 (n187, n56);
buf  g140 (n238, n46);
not  g141 (n293, n61);
not  g142 (n224, n57);
buf  g143 (n227, n37);
not  g144 (n310, n44);
not  g145 (n290, n67);
buf  g146 (n214, n44);
not  g147 (n189, n34);
not  g148 (n244, n51);
not  g149 (n253, n65);
not  g150 (n314, n59);
not  g151 (n308, n50);
buf  g152 (n176, n76);
buf  g153 (n160, n36);
buf  g154 (n234, n44);
buf  g155 (n165, n72);
not  g156 (n230, n33);
not  g157 (n301, n35);
not  g158 (n212, n47);
buf  g159 (n157, n52);
buf  g160 (n202, n30);
buf  g161 (n170, n72);
not  g162 (n256, n59);
not  g163 (n263, n39);
not  g164 (n276, n48);
not  g165 (n279, n61);
not  g166 (n194, n69);
not  g167 (n216, n67);
buf  g168 (n195, n47);
not  g169 (n180, n70);
not  g170 (n231, n53);
not  g171 (n318, n66);
not  g172 (n199, n49);
buf  g173 (n173, n66);
not  g174 (n261, n40);
buf  g175 (n191, n69);
buf  g176 (n283, n68);
buf  g177 (n197, n68);
not  g178 (n255, n38);
not  g179 (n267, n49);
buf  g180 (n303, n37);
not  g181 (n297, n67);
not  g182 (n218, n31);
buf  g183 (n233, n55);
not  g184 (n295, n49);
not  g185 (n221, n30);
not  g186 (n240, n75);
not  g187 (n287, n68);
buf  g188 (n245, n43);
buf  g189 (n161, n34);
not  g190 (n289, n44);
not  g191 (n152, n37);
not  g192 (n148, n63);
buf  g193 (n223, n43);
buf  g194 (n264, n29);
not  g195 (n243, n33);
not  g196 (n168, n55);
buf  g197 (n247, n40);
not  g198 (n217, n74);
buf  g199 (n196, n46);
not  g200 (n183, n39);
buf  g201 (n271, n63);
not  g202 (n312, n47);
not  g203 (n299, n29);
not  g204 (n185, n41);
not  g205 (n158, n42);
not  g206 (n246, n62);
buf  g207 (n210, n62);
buf  g208 (n304, n73);
not  g209 (n296, n40);
not  g210 (n153, n38);
not  g211 (n292, n41);
not  g212 (n319, n60);
not  g213 (n146, n56);
buf  g214 (n232, n33);
not  g215 (n239, n69);
buf  g216 (n288, n64);
not  g217 (n269, n48);
not  g218 (n154, n38);
buf  g219 (n174, n41);
buf  g220 (n222, n71);
not  g221 (n182, n57);
buf  g222 (n250, n35);
buf  g223 (n274, n63);
not  g224 (n151, n51);
buf  g225 (n155, n58);
not  g226 (n179, n64);
not  g227 (n249, n74);
not  g228 (n313, n58);
not  g229 (n198, n34);
not  g230 (n254, n75);
not  g231 (n164, n76);
not  g232 (n204, n60);
buf  g233 (n228, n52);
not  g234 (n172, n58);
buf  g235 (n260, n55);
not  g236 (n282, n71);
not  g237 (n285, n54);
not  g238 (n259, n33);
not  g239 (n192, n55);
buf  g240 (n162, n59);
not  g241 (n178, n36);
buf  g242 (n278, n69);
buf  g243 (n169, n56);
buf  g244 (n281, n63);
buf  g245 (n229, n54);
not  g246 (n242, n45);
buf  g247 (n147, n50);
not  g248 (n150, n57);
buf  g249 (n206, n66);
not  g250 (n181, n75);
not  g251 (n235, n72);
not  g252 (n300, n48);
not  g253 (n302, n30);
not  g254 (n272, n53);
not  g255 (n305, n73);
buf  g256 (n298, n42);
not  g257 (n213, n53);
buf  g258 (n166, n61);
buf  g259 (n275, n71);
buf  g260 (n190, n76);
buf  g261 (n211, n48);
buf  g262 (n186, n46);
buf  g263 (n317, n61);
buf  g264 (n219, n35);
not  g265 (n167, n54);
buf  g266 (n268, n51);
not  g267 (n265, n67);
buf  g268 (n262, n62);
not  g269 (n277, n68);
not  g270 (n215, n35);
not  g271 (n270, n29);
not  g272 (n156, n70);
not  g273 (n258, n51);
buf  g274 (n145, n54);
buf  g275 (n284, n46);
buf  g276 (n266, n30);
not  g277 (n200, n53);
not  g278 (n291, n37);
not  g279 (n226, n74);
buf  g280 (n208, n39);
not  g281 (n251, n65);
not  g282 (n286, n31);
xor  g283 (n306, n65, n50, n47, n43);
or   g284 (n220, n38, n40, n45, n64);
and  g285 (n193, n52, n42, n31, n36);
and  g286 (n315, n73, n72, n43, n59);
buf  g287 (n326, n76);
not  g288 (n340, n89);
buf  g289 (n341, n32);
buf  g290 (n372, n82);
buf  g291 (n373, n153);
not  g292 (n338, n79);
not  g293 (n351, n83);
not  g294 (n357, n147);
not  g295 (n347, n148);
buf  g296 (n324, n85);
buf  g297 (n344, n80);
buf  g298 (n364, n147);
buf  g299 (n366, n150);
buf  g300 (n361, n146);
buf  g301 (n321, n80);
buf  g302 (n348, n90);
buf  g303 (n331, n152);
buf  g304 (n355, n148);
not  g305 (n346, n157);
not  g306 (n328, n150);
buf  g307 (n354, n158);
not  g308 (n369, n155);
buf  g309 (n362, n90);
not  g310 (n332, n84);
not  g311 (n322, n87);
not  g312 (n345, n149);
not  g313 (n367, n145);
not  g314 (n336, n152);
not  g315 (n333, n147);
buf  g316 (n356, n87);
buf  g317 (n334, n84);
not  g318 (n323, n88);
not  g319 (n327, n77);
buf  g320 (n353, n83);
xor  g321 (n339, n78, n85, n157, n82);
xor  g322 (n350, n86, n85, n90, n78);
or   g323 (n370, n153, n78, n149, n151);
or   g324 (n360, n152, n86, n158, n154);
nor  g325 (n337, n88, n79, n146, n150);
nor  g326 (n330, n77, n79, n89, n146);
and  g327 (n329, n150, n86, n148, n82);
nand g328 (n363, n149, n156, n32, n80);
xor  g329 (n371, n85, n87, n155, n156);
xnor g330 (n365, n151, n153, n82, n32);
xor  g331 (n352, n157, n87, n84, n86);
or   g332 (n359, n156, n80, n81, n153);
nor  g333 (n342, n83, n155, n88, n157);
xnor g334 (n358, n145, n151, n79, n89);
nand g335 (n349, n155, n146, n84, n154);
xnor g336 (n368, n77, n32, n152, n83);
and  g337 (n320, n154, n145);
and  g338 (n343, n149, n147, n81, n89);
nand g339 (n325, n148, n77, n88, n78);
or   g340 (n335, n151, n156, n81);
nor  g341 (n392, n231, n98, n286, n287);
nor  g342 (n466, n163, n367, n162, n263);
nor  g343 (n563, n252, n105, n279, n221);
xor  g344 (n494, n344, n320, n208, n197);
and  g345 (n385, n187, n301, n221, n322);
nand g346 (n401, n235, n160, n90, n335);
nor  g347 (n537, n214, n338, n168, n202);
and  g348 (n398, n356, n342, n159, n222);
and  g349 (n460, n188, n363, n258, n230);
xor  g350 (n473, n242, n300, n262, n299);
nand g351 (n582, n266, n284, n228, n257);
xnor g352 (n439, n359, n271, n246, n362);
xor  g353 (n569, n297, n358, n189, n343);
xor  g354 (n574, n256, n371, n205, n234);
nor  g355 (n374, n161, n244, n238, n357);
xor  g356 (n476, n225, n221, n170, n208);
xnor g357 (n549, n101, n333, n327, n366);
and  g358 (n532, n335, n345, n185);
xnor g359 (n454, n293, n211, n162, n183);
or   g360 (n554, n339, n234, n175, n344);
xnor g361 (n397, n220, n341, n257, n95);
xnor g362 (n464, n260, n293, n165, n249);
and  g363 (n526, n254, n282, n189, n372);
and  g364 (n493, n92, n104, n172, n325);
xnor g365 (n424, n265, n279, n270, n367);
or   g366 (n479, n283, n216, n351, n366);
nor  g367 (n525, n273, n203, n268, n289);
xor  g368 (n390, n263, n250, n99, n321);
and  g369 (n492, n286, n104, n255, n222);
nand g370 (n465, n295, n227, n324, n235);
nor  g371 (n380, n249, n373, n360, n351);
xor  g372 (n410, n277, n354, n326);
nor  g373 (n429, n176, n103, n178, n274);
nor  g374 (n388, n256, n217, n227, n94);
or   g375 (n575, n240, n286, n201, n190);
nor  g376 (n520, n252, n184, n201, n244);
nand g377 (n470, n249, n176, n167, n334);
xor  g378 (n430, n344, n92, n327, n196);
xnor g379 (n461, n187, n204, n279, n224);
nor  g380 (n522, n206, n241, n220, n356);
xnor g381 (n431, n358, n196, n233, n212);
xor  g382 (n440, n263, n264, n239, n329);
xnor g383 (n584, n260, n336, n178, n331);
nor  g384 (n434, n237, n202, n222, n219);
nor  g385 (n509, n238, n96, n171, n170);
and  g386 (n571, n100, n191, n371, n203);
nor  g387 (n472, n351, n192, n173, n199);
xnor g388 (n428, n105, n247, n365, n91);
and  g389 (n435, n371, n161, n207, n367);
or   g390 (n518, n162, n170, n248, n195);
xnor g391 (n417, n171, n355, n220, n227);
or   g392 (n394, n203, n100, n209, n350);
nor  g393 (n450, n96, n237, n101, n182);
xor  g394 (n572, n172, n360, n253, n273);
xnor g395 (n409, n186, n196, n370, n177);
xnor g396 (n570, n176, n210, n357, n213);
nand g397 (n540, n229, n93, n365, n176);
and  g398 (n497, n165, n99, n197, n181);
xnor g399 (n521, n188, n369, n248, n95);
xor  g400 (n421, n186, n321, n161, n267);
or   g401 (n527, n352, n253, n267, n167);
nor  g402 (n416, n288, n369, n229, n234);
or   g403 (n517, n270, n186, n329, n350);
nand g404 (n391, n213, n326, n246, n245);
nand g405 (n542, n241, n104, n197, n274);
and  g406 (n523, n357, n215, n206, n180);
xor  g407 (n568, n194, n179, n183, n331);
and  g408 (n487, n218, n284, n246, n223);
xor  g409 (n550, n216, n234, n262, n291);
nor  g410 (n387, n362, n361, n285, n298);
or   g411 (n507, n293, n346, n279, n189);
xnor g412 (n448, n183, n260, n103, n254);
nand g413 (n469, n338, n160, n295, n353);
nor  g414 (n573, n373, n275, n244, n247);
or   g415 (n412, n102, n102, n290, n297);
xnor g416 (n580, n226, n328, n200, n294);
nand g417 (n406, n106, n214, n293, n345);
or   g418 (n559, n240, n205, n213, n360);
nand g419 (n471, n182, n272, n276, n246);
xor  g420 (n558, n94, n327, n188, n259);
nor  g421 (n567, n186, n211, n350, n212);
nor  g422 (n411, n359, n265, n347, n276);
and  g423 (n415, n97, n353, n323);
nor  g424 (n543, n93, n320, n366, n262);
xnor g425 (n403, n332, n348, n273, n191);
or   g426 (n395, n346, n94, n248, n187);
xor  g427 (n578, n105, n261, n300);
xnor g428 (n566, n332, n237, n290, n236);
or   g429 (n586, n301, n224, n280, n294);
xor  g430 (n452, n93, n251, n165, n265);
or   g431 (n505, n269, n214, n288, n171);
nand g432 (n478, n177, n212, n240, n289);
xnor g433 (n519, n292, n256, n96, n209);
and  g434 (n539, n201, n251, n250, n180);
xnor g435 (n536, n289, n290, n258, n340);
xnor g436 (n457, n193, n181, n199, n368);
nor  g437 (n474, n239, n298, n178, n275);
and  g438 (n534, n346, n339, n277, n329);
nand g439 (n538, n292, n181, n320, n198);
xnor g440 (n496, n339, n103, n98, n324);
xnor g441 (n456, n224, n294, n288, n166);
xor  g442 (n477, n224, n231, n256, n207);
and  g443 (n407, n183, n171, n349, n282);
xor  g444 (n425, n272, n92, n239, n228);
xnor g445 (n515, n369, n164, n322, n163);
and  g446 (n581, n349, n335, n255, n269);
xnor g447 (n544, n91, n258, n361, n286);
and  g448 (n462, n221, n210, n295, n329);
nand g449 (n418, n179, n362, n225, n175);
nand g450 (n502, n218, n217, n258, n347);
xor  g451 (n548, n287, n164, n185, n91);
or   g452 (n447, n164, n352, n185, n95);
xnor g453 (n486, n346, n337, n267, n349);
or   g454 (n458, n344, n355, n188, n321);
or   g455 (n404, n297, n247, n202, n322);
nand g456 (n500, n252, n231, n208, n326);
xnor g457 (n400, n219, n98, n291, n184);
nand g458 (n378, n276, n97, n334, n338);
xnor g459 (n432, n101, n285, n358, n158);
or   g460 (n463, n217, n247, n180, n271);
nor  g461 (n459, n238, n206, n174, n324);
xnor g462 (n451, n349, n348, n193);
and  g463 (n414, n193, n323, n233, n200);
and  g464 (n511, n292, n264, n174, n260);
and  g465 (n506, n205, n225, n235, n105);
or   g466 (n490, n190, n272, n360, n270);
nand g467 (n579, n162, n160, n253, n191);
xnor g468 (n530, n177, n181, n274);
xor  g469 (n446, n192, n211, n275, n330);
and  g470 (n510, n368, n354, n259, n170);
nand g471 (n484, n180, n194, n354, n284);
nor  g472 (n485, n160, n270, n198, n169);
xor  g473 (n438, n241, n333, n331, n97);
xnor g474 (n442, n323, n253, n262, n372);
xnor g475 (n443, n348, n242, n281, n163);
or   g476 (n528, n192, n175, n216, n248);
and  g477 (n565, n207, n328, n332, n354);
xnor g478 (n386, n223, n353, n236, n102);
or   g479 (n557, n91, n226, n290, n163);
nand g480 (n503, n268, n272, n266, n365);
or   g481 (n427, n347, n284, n172, n254);
nand g482 (n408, n300, n194, n363, n100);
xor  g483 (n545, n366, n257, n294, n351);
or   g484 (n489, n343, n327, n371, n97);
nor  g485 (n501, n227, n191, n352, n177);
nor  g486 (n468, n232, n341, n277, n335);
xnor g487 (n504, n238, n173, n207, n276);
xnor g488 (n551, n337, n261, n356, n243);
nand g489 (n541, n363, n336, n198, n261);
xor  g490 (n512, n330, n340, n215, n295);
xnor g491 (n455, n242, n169, n283, n243);
or   g492 (n513, n209, n340, n266, n252);
and  g493 (n547, n325, n250, n179, n282);
xnor g494 (n377, n178, n300, n196, n245);
or   g495 (n482, n370, n368, n166, n299);
and  g496 (n382, n218, n232, n159, n211);
nand g497 (n585, n333, n231, n165, n195);
nor  g498 (n402, n357, n277, n330);
xnor g499 (n381, n283, n291, n200, n219);
nor  g500 (n546, n369, n159, n158, n278);
xor  g501 (n560, n265, n239, n102, n220);
nor  g502 (n552, n334, n200, n251, n223);
xnor g503 (n467, n281, n184, n208, n273);
xnor g504 (n524, n190, n296, n269, n99);
nor  g505 (n422, n280, n103, n267, n361);
xnor g506 (n498, n166, n331, n362, n278);
nor  g507 (n426, n226, n98, n337, n336);
or   g508 (n475, n218, n259, n281, n167);
nor  g509 (n413, n356, n347, n214, n199);
or   g510 (n583, n100, n343, n268, n249);
and  g511 (n531, n325, n182, n280, n301);
xor  g512 (n445, n173, n264, n228, n199);
and  g513 (n576, n106, n297, n202, n169);
and  g514 (n437, n350, n161, n174, n324);
nor  g515 (n379, n92, n187, n245, n296);
and  g516 (n556, n189, n298, n195, n179);
xor  g517 (n514, n332, n325, n172, n285);
xor  g518 (n553, n255, n225, n233, n264);
nor  g519 (n375, n278, n368, n203, n230);
nand g520 (n499, n341, n195, n372, n339);
nor  g521 (n533, n204, n345, n283, n173);
and  g522 (n577, n287, n242, n244, n229);
nor  g523 (n495, n93, n358, n359, n230);
and  g524 (n561, n323, n222, n226, n223);
xnor g525 (n433, n237, n299, n168);
nor  g526 (n420, n219, n321, n359, n236);
or   g527 (n516, n174, n182, n204, n250);
or   g528 (n376, n210, n287, n340, n99);
nand g529 (n396, n257, n328, n296, n301);
or   g530 (n384, n278, n236, n167, n291);
xnor g531 (n488, n364, n370, n210, n212);
and  g532 (n555, n364, n254, n104, n245);
and  g533 (n436, n363, n296, n343, n367);
and  g534 (n562, n280, n215, n201, n289);
or   g535 (n449, n364, n336, n164, n361);
and  g536 (n481, n342, n240, n185, n285);
xnor g537 (n441, n228, n204, n275, n190);
nor  g538 (n419, n230, n229, n106, n266);
xor  g539 (n405, n166, n251, n193, n235);
or   g540 (n480, n355, n334, n282, n106);
nand g541 (n508, n365, n168, n328, n213);
xnor g542 (n453, n184, n341, n271, n255);
or   g543 (n483, n232, n95, n281, n259);
nand g544 (n535, n370, n205, n337, n352);
xor  g545 (n564, n243, n192, n342, n241);
and  g546 (n389, n209, n197, n96, n269);
xor  g547 (n399, n159, n263, n292, n215);
and  g548 (n393, n271, n342, n338, n355);
xor  g549 (n444, n288, n243, n364, n168);
xnor g550 (n423, n217, n268, n94, n194);
nand g551 (n383, n175, n333, n322, n233);
and  g552 (n529, n169, n232, n216, n206);
xor  g553 (n491, n198, n298, n372, n101);
and  g554 (n588, n137, n123, n117, n107);
xnor g555 (n601, n140, n303, n138, n111);
xor  g556 (n634, n141, n142, n389, n388);
nor  g557 (n626, n118, n107, n378);
nor  g558 (n631, n374, n108, n139, n124);
nand g559 (n627, n308, n379, n113, n133);
xnor g560 (n608, n123, n136, n384);
xor  g561 (n617, n118, n130, n121, n132);
nand g562 (n600, n109, n117, n114, n144);
xor  g563 (n611, n119, n114, n115, n377);
and  g564 (n612, n383, n381, n129, n387);
xor  g565 (n591, n387, n389, n132, n382);
or   g566 (n622, n141, n122, n143, n134);
or   g567 (n638, n120, n113, n116);
or   g568 (n610, n373, n121, n141, n143);
xnor g569 (n596, n117, n381, n127, n302);
and  g570 (n616, n124, n390, n119, n111);
or   g571 (n615, n142, n378, n130, n144);
and  g572 (n613, n142, n120, n121, n375);
xnor g573 (n633, n380, n131, n109, n140);
nor  g574 (n614, n122, n127, n125, n120);
or   g575 (n603, n139, n382, n140, n129);
and  g576 (n624, n135, n304, n134);
xnor g577 (n595, n388, n305, n375, n306);
nor  g578 (n589, n379, n125, n138, n112);
xor  g579 (n618, n111, n376, n385, n108);
nor  g580 (n597, n140, n133, n387, n380);
nor  g581 (n598, n377, n116, n386, n118);
or   g582 (n635, n109, n304, n137, n302);
nor  g583 (n630, n131, n112, n136, n144);
and  g584 (n628, n128, n391, n118, n133);
xor  g585 (n606, n123, n133, n125, n115);
or   g586 (n623, n385, n114, n374, n143);
xor  g587 (n594, n392, n393, n109, n381);
or   g588 (n599, n135, n379, n386, n107);
or   g589 (n639, n302, n136, n305, n385);
nand g590 (n625, n113, n303, n115, n139);
nor  g591 (n643, n306, n134, n131, n121);
and  g592 (n632, n306, n127, n108, n117);
or   g593 (n605, n122, n384, n138, n391);
nor  g594 (n641, n393, n129, n144, n120);
nand g595 (n646, n123, n134, n124, n125);
and  g596 (n590, n374, n391, n305, n110);
nand g597 (n619, n132, n128, n384, n122);
or   g598 (n609, n138, n110);
xor  g599 (n587, n137, n130, n143, n111);
and  g600 (n604, n129, n141, n135, n132);
xnor g601 (n593, n377, n130, n142, n376);
nor  g602 (n620, n373, n128, n126, n107);
nor  g603 (n621, n112, n302, n392, n393);
and  g604 (n640, n306, n308, n376, n139);
nor  g605 (n602, n303, n116, n392);
and  g606 (n636, n307, n390, n112, n388);
nor  g607 (n637, n137, n108, n307, n126);
or   g608 (n642, n386, n380, n375, n115);
xor  g609 (n645, n127, n126, n128, n114);
xor  g610 (n607, n119, n307, n124);
or   g611 (n629, n304, n383, n135, n126);
xnor g612 (n644, n131, n119, n383, n303);
nand g613 (n592, n389, n305, n382, n390);
nor  g614 (n689, n506, n514, n641, n423);
and  g615 (n647, n471, n637, n483, n486);
and  g616 (n685, n414, n513, n638, n642);
nand g617 (n738, n473, n636, n618, n489);
and  g618 (n713, n631, n474, n587, n427);
nor  g619 (n711, n515, n415, n465, n495);
xnor g620 (n660, n466, n618, n460, n424);
and  g621 (n722, n615, n458, n400, n473);
nor  g622 (n726, n403, n441, n635, n447);
xnor g623 (n690, n628, n477, n482, n509);
nand g624 (n661, n512, n439, n508, n499);
xnor g625 (n762, n462, n402, n638, n454);
nand g626 (n686, n419, n504, n453, n628);
nor  g627 (n761, n644, n625, n433, n426);
or   g628 (n696, n401, n453, n633, n498);
and  g629 (n694, n626, n500, n408, n627);
nor  g630 (n702, n469, n631, n430, n496);
and  g631 (n718, n400, n398, n639, n600);
nand g632 (n715, n413, n616, n442, n395);
nor  g633 (n723, n466, n399, n487, n451);
xor  g634 (n719, n407, n437, n462, n409);
xor  g635 (n740, n633, n436, n416, n445);
and  g636 (n763, n414, n426, n646, n644);
or   g637 (n697, n464, n624, n427, n404);
or   g638 (n766, n462, n641, n629, n609);
xnor g639 (n760, n481, n464, n453, n411);
nand g640 (n683, n632, n514, n415, n399);
xor  g641 (n649, n505, n616, n633, n620);
nor  g642 (n650, n396, n405, n459, n408);
and  g643 (n730, n447, n505, n469, n606);
and  g644 (n734, n607, n611, n623, n429);
xnor g645 (n751, n412, n403, n442, n404);
nor  g646 (n669, n512, n394, n631, n448);
nor  g647 (n755, n455, n634, n470, n485);
xnor g648 (n680, n438, n417, n479, n461);
xnor g649 (n752, n646, n625, n424, n457);
nand g650 (n674, n490, n397, n604, n488);
or   g651 (n666, n446, n591, n449, n396);
xor  g652 (n733, n481, n640, n617, n509);
and  g653 (n692, n413, n494, n460, n467);
xor  g654 (n677, n418, n636, n610, n406);
or   g655 (n678, n439, n623, n498, n450);
nor  g656 (n721, n416, n460, n424, n643);
or   g657 (n758, n602, n507, n425, n464);
nand g658 (n743, n494, n411, n500, n432);
and  g659 (n688, n401, n456, n511, n399);
xor  g660 (n746, n434, n645, n478, n632);
nand g661 (n662, n430, n494, n440, n638);
xnor g662 (n684, n501, n483, n410, n403);
and  g663 (n695, n485, n476, n468, n472);
and  g664 (n732, n496, n489, n446, n415);
xnor g665 (n672, n433, n433, n506, n612);
nand g666 (n745, n432, n476, n640, n405);
or   g667 (n741, n617, n510, n469, n468);
or   g668 (n720, n482, n411, n475, n445);
nor  g669 (n705, n628, n637, n435, n630);
or   g670 (n747, n465, n436, n484, n430);
nand g671 (n764, n452, n402, n467, n438);
xor  g672 (n664, n620, n400, n452, n503);
and  g673 (n652, n497, n501, n639, n398);
xnor g674 (n671, n511, n467, n488, n624);
and  g675 (n725, n479, n444, n629, n515);
xnor g676 (n691, n429, n420, n491, n488);
or   g677 (n765, n414, n509, n504, n608);
or   g678 (n693, n613, n445, n443, n601);
and  g679 (n744, n419, n479, n629, n448);
and  g680 (n703, n404, n468, n642, n426);
nand g681 (n710, n487, n486, n471, n437);
nand g682 (n748, n508, n492, n420, n619);
nor  g683 (n735, n431, n417, n461, n475);
and  g684 (n653, n407, n487, n621, n425);
or   g685 (n727, n422, n516, n459, n496);
nand g686 (n739, n605, n478, n434, n410);
and  g687 (n708, n428, n484, n427, n497);
nand g688 (n731, n594, n474, n639, n499);
xnor g689 (n750, n516, n418, n480, n417);
nand g690 (n756, n626, n437, n413, n444);
xnor g691 (n757, n513, n431, n593, n483);
nor  g692 (n709, n428, n412, n635, n456);
and  g693 (n728, n492, n634, n420, n477);
xor  g694 (n753, n457, n472, n423, n493);
nor  g695 (n724, n441, n616, n619, n463);
xor  g696 (n673, n621, n595, n603, n480);
xor  g697 (n742, n407, n406, n397);
and  g698 (n654, n588, n421, n481, n627);
or   g699 (n670, n421, n449, n644, n475);
xnor g700 (n736, n642, n457, n500, n592);
and  g701 (n657, n508, n408, n435, n422);
xnor g702 (n767, n416, n598, n451, n432);
or   g703 (n679, n458, n491, n516, n625);
xor  g704 (n699, n503, n590, n472, n597);
xnor g705 (n648, n514, n515, n482, n440);
xnor g706 (n754, n495, n409, n618, n643);
and  g707 (n700, n505, n476, n627, n645);
xnor g708 (n704, n434, n645, n634, n635);
nand g709 (n769, n495, n619, n513, n493);
nand g710 (n681, n507, n589, n614, n395);
xor  g711 (n768, n470, n492, n622, n412);
and  g712 (n682, n405, n471, n502, n474);
nor  g713 (n701, n478, n466, n623, n396);
and  g714 (n712, n438, n461, n501, n439);
xor  g715 (n729, n443, n410, n621, n498);
and  g716 (n749, n441, n418, n463, n422);
nand g717 (n656, n506, n452, n394, n443);
xor  g718 (n698, n401, n473, n486, n429);
xor  g719 (n716, n599, n448, n491, n502);
xnor g720 (n668, n455, n409, n450, n398);
xnor g721 (n759, n512, n397, n626, n636);
xor  g722 (n737, n447, n622, n630);
or   g723 (n706, n449, n436, n395, n402);
or   g724 (n717, n641, n503, n423, n480);
nor  g725 (n651, n394, n510, n477, n490);
nor  g726 (n658, n643, n620, n617, n428);
xor  g727 (n675, n640, n507, n596, n450);
nor  g728 (n676, n630, n425, n490, n470);
nor  g729 (n655, n624, n419, n463, n431);
or   g730 (n667, n510, n502, n646, n485);
and  g731 (n665, n454, n465, n444, n440);
and  g732 (n714, n459, n435, n504, n637);
or   g733 (n663, n455, n451, n456, n632);
or   g734 (n707, n493, n489, n454, n446);
nand g735 (n659, n458, n497, n499, n646);
and  g736 (n687, n484, n442, n511, n421);
xnor g737 (n803, n662, n652, n550, n539);
and  g738 (n786, n656, n530, n544, n312);
xnor g739 (n770, n550, n525, n542, n310);
nand g740 (n814, n659, n309, n523, n539);
and  g741 (n798, n546, n657, n522, n553);
xor  g742 (n808, n532, n531, n310, n309);
xnor g743 (n774, n315, n546, n658, n653);
and  g744 (n818, n649, n311, n543, n538);
xnor g745 (n797, n318, n313, n517, n663);
nor  g746 (n791, n527, n656, n650, n318);
nand g747 (n776, n314, n521, n548, n522);
nor  g748 (n813, n548, n533, n524, n654);
or   g749 (n822, n551, n312, n533, n660);
xor  g750 (n821, n656, n520, n527, n537);
nand g751 (n800, n655, n316, n313, n518);
nand g752 (n819, n317, n316, n524, n526);
xnor g753 (n804, n552, n526, n535, n524);
xnor g754 (n795, n534, n521, n319, n529);
xnor g755 (n805, n540, n317, n517, n664);
nor  g756 (n809, n536, n310, n552, n663);
nor  g757 (n778, n309, n553, n542, n319);
nor  g758 (n772, n554, n552, n529, n541);
nand g759 (n801, n531, n523, n537, n659);
nand g760 (n812, n521, n314, n313, n317);
and  g761 (n815, n652, n527, n651, n543);
xor  g762 (n784, n538, n530, n650, n534);
nor  g763 (n782, n311, n551, n519, n663);
xor  g764 (n806, n548, n649, n523, n525);
xnor g765 (n777, n648, n313, n658, n517);
xor  g766 (n771, n520, n549, n661, n651);
xor  g767 (n810, n315, n551, n518, n664);
xnor g768 (n794, n547, n653, n309, n540);
or   g769 (n773, n647, n545, n314, n652);
or   g770 (n817, n531, n544, n519, n532);
or   g771 (n781, n650, n314, n648, n536);
nor  g772 (n799, n554, n311, n661, n310);
xor  g773 (n788, n541, n537, n520, n315);
nand g774 (n780, n528, n660, n544, n522);
xor  g775 (n787, n549, n662, n539, n533);
nand g776 (n796, n319, n316, n662, n317);
or   g777 (n775, n648, n664, n532, n545);
nand g778 (n807, n538, n655, n553, n312);
nor  g779 (n820, n655, n653, n316, n312);
xnor g780 (n802, n651, n542, n658, n545);
xor  g781 (n792, n308, n543, n525, n535);
or   g782 (n789, n536, n529, n318, n550);
xnor g783 (n793, n649, n540, n319, n530);
and  g784 (n816, n528, n547, n654, n519);
xnor g785 (n779, n534, n654, n549, n660);
xor  g786 (n785, n535, n308, n518, n657);
xnor g787 (n811, n659, n661, n318, n528);
xnor g788 (n783, n657, n547, n663, n541);
xor  g789 (n790, n546, n526, n315, n311);
or   g790 (n879, n756, n722, n686, n735);
or   g791 (n922, n666, n667, n745, n754);
or   g792 (n849, n708, n675, n792, n724);
and  g793 (n915, n787, n735, n786, n716);
nor  g794 (n888, n703, n708, n810, n681);
nand g795 (n917, n811, n687, n802, n715);
nor  g796 (n826, n698, n712, n711, n741);
xnor g797 (n855, n700, n698, n744, n799);
xnor g798 (n844, n797, n712, n739, n702);
xor  g799 (n851, n717, n733, n689, n696);
xor  g800 (n884, n741, n694, n690, n743);
and  g801 (n839, n780, n742, n665, n788);
nand g802 (n918, n674, n797, n677, n748);
xor  g803 (n951, n731, n822, n718, n805);
xnor g804 (n927, n796, n696, n693, n677);
or   g805 (n906, n821, n682, n758, n805);
xor  g806 (n866, n781, n756, n777, n740);
nand g807 (n882, n692, n794, n755, n723);
xnor g808 (n897, n697, n690, n692, n706);
xnor g809 (n824, n785, n750, n682, n678);
nor  g810 (n827, n750, n739, n734, n670);
nand g811 (n860, n707, n694, n708, n716);
xnor g812 (n935, n807, n797, n688, n668);
and  g813 (n941, n707, n729, n746, n820);
nand g814 (n905, n778, n816, n757, n722);
or   g815 (n853, n686, n758, n677, n554);
xnor g816 (n904, n808, n685, n720, n669);
xnor g817 (n894, n694, n714, n812, n735);
xor  g818 (n942, n725, n740, n822, n732);
nand g819 (n889, n686, n728, n802, n714);
xor  g820 (n933, n809, n679, n742);
nor  g821 (n911, n817, n807, n757, n753);
nor  g822 (n890, n748, n711, n710, n707);
xor  g823 (n937, n691, n677, n741, n814);
xnor g824 (n925, n761, n685, n759, n813);
xor  g825 (n896, n740, n770, n702, n795);
nand g826 (n945, n692, n819, n690, n801);
nor  g827 (n847, n743, n685, n681, n729);
xnor g828 (n886, n800, n712, n678);
xnor g829 (n932, n665, n753, n791, n754);
and  g830 (n944, n747, n700, n816, n775);
nor  g831 (n862, n808, n667, n799, n692);
xor  g832 (n828, n806, n708, n744, n805);
nor  g833 (n833, n798, n705, n714, n737);
and  g834 (n863, n752, n784, n710, n727);
or   g835 (n861, n671, n743, n820, n693);
or   g836 (n881, n815, n793, n666, n691);
nand g837 (n841, n796, n683, n666, n681);
nand g838 (n946, n738, n703, n801, n748);
nor  g839 (n876, n757, n710, n693, n745);
and  g840 (n920, n786, n670, n815, n725);
nand g841 (n830, n701, n746, n814, n713);
or   g842 (n891, n711, n789, n684, n822);
nor  g843 (n899, n814, n739, n785, n751);
and  g844 (n923, n734, n746, n803, n679);
xor  g845 (n865, n745, n779, n737, n756);
and  g846 (n854, n705, n720, n809, n678);
nor  g847 (n910, n718, n732, n706, n680);
xnor g848 (n936, n749, n690, n724, n803);
and  g849 (n838, n671, n761, n676, n701);
xor  g850 (n872, n669, n711, n792, n732);
or   g851 (n869, n821, n790, n689, n753);
and  g852 (n950, n800, n730, n746, n736);
xor  g853 (n870, n700, n725, n758, n670);
nand g854 (n850, n717, n669, n674, n703);
xor  g855 (n939, n697, n817, n705, n715);
nand g856 (n878, n666, n680, n817, n750);
or   g857 (n908, n713, n749, n790, n729);
xor  g858 (n912, n721, n723, n806, n755);
and  g859 (n947, n706, n678, n693, n731);
nor  g860 (n931, n796, n675, n757, n722);
nand g861 (n914, n755, n754, n813, n738);
xor  g862 (n929, n747, n799, n721, n774);
xor  g863 (n840, n679, n720, n758, n773);
xor  g864 (n864, n667, n696, n689, n819);
nand g865 (n856, n731, n810, n804, n709);
nand g866 (n832, n725, n728, n804, n760);
nand g867 (n877, n742, n710, n782, n680);
and  g868 (n919, n760, n787, n812, n815);
xor  g869 (n940, n555, n731, n719, n822);
nor  g870 (n857, n809, n751, n674, n795);
xor  g871 (n835, n668, n673, n709, n719);
and  g872 (n867, n801, n695, n776, n738);
xnor g873 (n949, n737, n730, n689, n771);
or   g874 (n837, n681, n787, n798, n716);
xor  g875 (n952, n740, n687, n807, n818);
nor  g876 (n842, n783, n688, n751, n744);
nand g877 (n825, n811, n716, n726, n680);
and  g878 (n934, n697, n672, n732, n727);
nand g879 (n913, n736, n700, n750, n794);
nand g880 (n858, n722, n713, n759, n715);
xnor g881 (n938, n811, n709, n726, n734);
nand g882 (n868, n791, n818, n738, n671);
xor  g883 (n901, n724, n672, n703, n682);
xnor g884 (n880, n793, n726, n665, n743);
xnor g885 (n895, n699, n694, n715, n792);
xnor g886 (n916, n676, n759, n679, n705);
nand g887 (n875, n665, n749, n686, n685);
and  g888 (n898, n744, n752, n719, n747);
nor  g889 (n836, n667, n727, n741, n795);
nor  g890 (n909, n816, n676, n752, n727);
or   g891 (n921, n687, n721, n723, n719);
xnor g892 (n883, n669, n818, n699, n674);
xnor g893 (n831, n704, n760, n672, n737);
xor  g894 (n924, n745, n684, n804, n736);
and  g895 (n885, n684, n717, n751, n696);
xor  g896 (n903, n709, n683, n707, n736);
xor  g897 (n874, n810, n726, n683, n701);
or   g898 (n902, n675, n733, n670, n739);
and  g899 (n859, n788, n793, n806, n704);
xor  g900 (n893, n794, n668, n821, n747);
or   g901 (n892, n702, n812, n756, n691);
xor  g902 (n846, n717, n672, n730, n706);
xor  g903 (n900, n668, n673, n555, n788);
xor  g904 (n907, n683, n753, n728, n760);
or   g905 (n871, n704, n755, n688, n759);
xor  g906 (n926, n664, n728, n704, n673);
xnor g907 (n948, n798, n718, n695, n721);
and  g908 (n829, n673, n702, n688, n808);
or   g909 (n823, n682, n733, n698, n752);
and  g910 (n873, n733, n803, n791, n800);
and  g911 (n928, n687, n713, n730, n749);
xor  g912 (n843, n684, n734, n714, n813);
xor  g913 (n930, n675, n695, n785, n697);
nand g914 (n943, n701, n790, n720, n786);
nor  g915 (n852, n729, n698, n699, n754);
or   g916 (n845, n789, n735, n819, n802);
xor  g917 (n848, n718, n691, n772, n724);
nand g918 (n887, n820, n723, n676, n695);
and  g919 (n834, n699, n789, n671, n748);
or   g920 (n986, n884, n846, n575, n870);
xnor g921 (n981, n570, n873, n574, n921);
nand g922 (n953, n557, n876, n887, n575);
and  g923 (n977, n583, n563, n561, n558);
or   g924 (n985, n569, n564, n582, n907);
and  g925 (n1016, n826, n577, n845, n561);
nor  g926 (n956, n575, n581, n933, n926);
or   g927 (n976, n763, n573, n909, n766);
and  g928 (n961, n901, n761, n769, n763);
and  g929 (n1015, n567, n580, n857, n934);
or   g930 (n975, n881, n922, n848, n912);
xnor g931 (n994, n880, n915, n584, n823);
xor  g932 (n968, n571, n866, n556, n768);
and  g933 (n1009, n847, n856, n767, n898);
nand g934 (n960, n904, n763, n581, n906);
xor  g935 (n969, n919, n852, n854, n829);
xor  g936 (n989, n916, n562, n878, n563);
nor  g937 (n963, n570, n578, n566, n894);
xnor g938 (n1012, n576, n902, n570, n765);
nand g939 (n980, n929, n564, n580, n882);
xor  g940 (n990, n763, n872, n889, n582);
nand g941 (n979, n581, n762, n936, n557);
or   g942 (n1003, n890, n908, n555, n586);
xor  g943 (n971, n913, n858, n865, n877);
and  g944 (n959, n874, n580, n843, n892);
and  g945 (n999, n766, n838, n582, n769);
xor  g946 (n972, n769, n886, n585, n861);
or   g947 (n974, n832, n840, n584, n879);
nand g948 (n1001, n565, n580, n576, n572);
or   g949 (n962, n769, n569, n911, n577);
nand g950 (n987, n577, n825, n574, n568);
nor  g951 (n992, n585, n875, n851, n841);
xnor g952 (n998, n586, n565, n867, n561);
nand g953 (n1014, n566, n583, n584, n850);
or   g954 (n1010, n920, n828, n765, n925);
xor  g955 (n983, n918, n842, n930, n579);
xor  g956 (n1000, n837, n849, n571, n556);
nand g957 (n993, n768, n905, n836, n834);
and  g958 (n973, n559, n869, n899, n768);
or   g959 (n1007, n917, n910, n578, n927);
or   g960 (n978, n827, n833, n764, n563);
xor  g961 (n958, n575, n767, n895, n853);
or   g962 (n982, n572, n762, n574, n585);
xnor g963 (n954, n583, n900, n767, n577);
or   g964 (n1008, n839, n871, n766, n562);
and  g965 (n964, n573, n558, n574, n893);
xor  g966 (n1013, n935, n585, n579, n573);
or   g967 (n1006, n560, n914, n924, n764);
xor  g968 (n984, n579, n586, n565, n923);
or   g969 (n996, n557, n768, n564, n576);
xor  g970 (n995, n888, n883, n859, n568);
nand g971 (n966, n566, n568, n558, n855);
nand g972 (n988, n560, n560, n762, n582);
and  g973 (n955, n586, n862, n864, n567);
xor  g974 (n1011, n824, n559, n860, n569);
and  g975 (n1005, n830, n584, n761, n767);
and  g976 (n1002, n764, n765, n932, n559);
and  g977 (n957, n903, n578, n572, n579);
or   g978 (n965, n571, n891, n765, n576);
xor  g979 (n1004, n844, n931, n764, n578);
and  g980 (n991, n567, n766, n573, n863);
nor  g981 (n997, n885, n581, n556, n868);
and  g982 (n970, n762, n928, n562, n896);
xor  g983 (n967, n897, n835, n831, n583);
xnor g984 (n1029, n1009, n943, n997, n972);
xnor g985 (n1028, n1005, n948, n940, n983);
nand g986 (n1021, n949, n992, n985, n971);
and  g987 (n1017, n952, n1002, n1012, n1010);
xor  g988 (n1022, n1000, n1013, n991, n1003);
and  g989 (n1025, n947, n976, n1016, n939);
xnor g990 (n1024, n979, n974, n1008, n998);
xnor g991 (n1020, n993, n975, n945, n987);
nor  g992 (n1027, n981, n951, n1015, n990);
xor  g993 (n1023, n1001, n946, n950, n984);
xor  g994 (n1018, n977, n1004, n986, n978);
or   g995 (n1032, n1014, n982, n995, n969);
or   g996 (n1031, n996, n989, n944, n988);
and  g997 (n1019, n999, n938, n942, n941);
and  g998 (n1026, n973, n994, n980, n1006);
nor  g999 (n1030, n1011, n937, n1007, n970);
endmodule
