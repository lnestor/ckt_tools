

module Stat_2188_30_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n1919,
  n1911,
  n1928,
  n1906,
  n1927,
  n1892,
  n1930,
  n1924,
  n1898,
  n1889,
  n1896,
  n1890,
  n1908,
  n1905,
  n1922,
  n1920,
  n1894,
  n1899,
  n1900,
  n1909,
  n1929,
  n1916,
  n1907,
  n1901,
  n1904,
  n1902,
  n1995,
  n1985,
  n1994,
  n1992,
  n1996,
  n2202,
  n2205,
  n2204,
  n2203
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1919;output n1911;output n1928;output n1906;output n1927;output n1892;output n1930;output n1924;output n1898;output n1889;output n1896;output n1890;output n1908;output n1905;output n1922;output n1920;output n1894;output n1899;output n1900;output n1909;output n1929;output n1916;output n1907;output n1901;output n1904;output n1902;output n1995;output n1985;output n1994;output n1992;output n1996;output n2202;output n2205;output n2204;output n2203;
  wire n18;wire n19;wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1891;wire n1893;wire n1895;wire n1897;wire n1903;wire n1910;wire n1912;wire n1913;wire n1914;wire n1915;wire n1917;wire n1918;wire n1921;wire n1923;wire n1925;wire n1926;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1993;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n76,
    n6
  );


  not
  g1
  (
    n49,
    n15
  );


  not
  g2
  (
    n25,
    n12
  );


  not
  g3
  (
    n55,
    n8
  );


  not
  g4
  (
    n65,
    n10
  );


  not
  g5
  (
    n63,
    n16
  );


  not
  g6
  (
    KeyWire_0_18,
    n13
  );


  buf
  g7
  (
    n19,
    n9
  );


  not
  g8
  (
    n47,
    n17
  );


  not
  g9
  (
    n35,
    n11
  );


  buf
  g10
  (
    n23,
    n2
  );


  buf
  g11
  (
    n57,
    n2
  );


  not
  g12
  (
    n38,
    n10
  );


  buf
  g13
  (
    n79,
    n3
  );


  not
  g14
  (
    n59,
    n9
  );


  not
  g15
  (
    n64,
    n3
  );


  not
  g16
  (
    n50,
    n13
  );


  not
  g17
  (
    n51,
    n4
  );


  not
  g18
  (
    n84,
    n10
  );


  not
  g19
  (
    n33,
    n8
  );


  not
  g20
  (
    n21,
    n6
  );


  not
  g21
  (
    n52,
    n3
  );


  buf
  g22
  (
    n44,
    n8
  );


  not
  g23
  (
    n27,
    n14
  );


  buf
  g24
  (
    n18,
    n10
  );


  buf
  g25
  (
    n69,
    n11
  );


  not
  g26
  (
    n77,
    n11
  );


  not
  g27
  (
    n30,
    n5
  );


  not
  g28
  (
    n32,
    n4
  );


  buf
  g29
  (
    n39,
    n3
  );


  not
  g30
  (
    n54,
    n5
  );


  not
  g31
  (
    n78,
    n2
  );


  not
  g32
  (
    n24,
    n6
  );


  not
  g33
  (
    n71,
    n1
  );


  buf
  g34
  (
    n37,
    n17
  );


  not
  g35
  (
    n70,
    n4
  );


  not
  g36
  (
    n83,
    n7
  );


  not
  g37
  (
    n29,
    n5
  );


  buf
  g38
  (
    n45,
    n12
  );


  not
  g39
  (
    n26,
    n7
  );


  buf
  g40
  (
    n53,
    n14
  );


  buf
  g41
  (
    n34,
    n9
  );


  buf
  g42
  (
    n82,
    n16
  );


  buf
  g43
  (
    n56,
    n11
  );


  buf
  g44
  (
    n61,
    n8
  );


  buf
  g45
  (
    n66,
    n5
  );


  not
  g46
  (
    n41,
    n6
  );


  buf
  g47
  (
    n42,
    n2
  );


  buf
  g48
  (
    n67,
    n13
  );


  buf
  g49
  (
    n36,
    n1
  );


  not
  g50
  (
    n40,
    n14
  );


  buf
  g51
  (
    n58,
    n14
  );


  not
  g52
  (
    n85,
    n17
  );


  not
  g53
  (
    n46,
    n16
  );


  not
  g54
  (
    n81,
    n4
  );


  not
  g55
  (
    KeyWire_0_13,
    n16
  );


  buf
  g56
  (
    n31,
    n7
  );


  buf
  g57
  (
    n80,
    n15
  );


  buf
  g58
  (
    n73,
    n9
  );


  buf
  g59
  (
    n75,
    n15
  );


  buf
  g60
  (
    n68,
    n17
  );


  buf
  g61
  (
    n60,
    n13
  );


  not
  g62
  (
    n28,
    n12
  );


  not
  g63
  (
    n43,
    n7
  );


  not
  g64
  (
    n74,
    n15
  );


  buf
  g65
  (
    n62,
    n1
  );


  buf
  g66
  (
    n20,
    n12
  );


  buf
  g67
  (
    n72,
    n1
  );


  not
  g68
  (
    n307,
    n66
  );


  not
  g69
  (
    n176,
    n83
  );


  buf
  g70
  (
    n119,
    n64
  );


  buf
  g71
  (
    n248,
    n19
  );


  buf
  g72
  (
    n88,
    n71
  );


  not
  g73
  (
    n212,
    n57
  );


  buf
  g74
  (
    n298,
    n69
  );


  buf
  g75
  (
    n208,
    n59
  );


  not
  g76
  (
    n209,
    n78
  );


  buf
  g77
  (
    n92,
    n38
  );


  buf
  g78
  (
    n200,
    n53
  );


  buf
  g79
  (
    n294,
    n44
  );


  buf
  g80
  (
    n252,
    n56
  );


  buf
  g81
  (
    n239,
    n78
  );


  buf
  g82
  (
    n346,
    n41
  );


  buf
  g83
  (
    n107,
    n68
  );


  buf
  g84
  (
    n115,
    n78
  );


  buf
  g85
  (
    n331,
    n25
  );


  not
  g86
  (
    n195,
    n52
  );


  buf
  g87
  (
    n242,
    n52
  );


  buf
  g88
  (
    n135,
    n53
  );


  buf
  g89
  (
    n321,
    n53
  );


  buf
  g90
  (
    KeyWire_0_7,
    n77
  );


  buf
  g91
  (
    n343,
    n76
  );


  buf
  g92
  (
    n123,
    n29
  );


  not
  g93
  (
    n339,
    n75
  );


  buf
  g94
  (
    n134,
    n51
  );


  not
  g95
  (
    n153,
    n57
  );


  buf
  g96
  (
    n259,
    n37
  );


  buf
  g97
  (
    n99,
    n43
  );


  buf
  g98
  (
    n150,
    n71
  );


  buf
  g99
  (
    n225,
    n18
  );


  not
  g100
  (
    n278,
    n72
  );


  buf
  g101
  (
    n311,
    n46
  );


  buf
  g102
  (
    n97,
    n84
  );


  not
  g103
  (
    n203,
    n81
  );


  buf
  g104
  (
    n261,
    n36
  );


  buf
  g105
  (
    n329,
    n63
  );


  not
  g106
  (
    n151,
    n74
  );


  not
  g107
  (
    n89,
    n57
  );


  not
  g108
  (
    n336,
    n38
  );


  buf
  g109
  (
    n93,
    n77
  );


  not
  g110
  (
    n280,
    n40
  );


  buf
  g111
  (
    n114,
    n43
  );


  buf
  g112
  (
    n273,
    n77
  );


  buf
  g113
  (
    n268,
    n37
  );


  buf
  g114
  (
    n341,
    n29
  );


  buf
  g115
  (
    n112,
    n56
  );


  buf
  g116
  (
    n183,
    n76
  );


  buf
  g117
  (
    n194,
    n38
  );


  buf
  g118
  (
    n265,
    n50
  );


  not
  g119
  (
    n223,
    n73
  );


  buf
  g120
  (
    n144,
    n35
  );


  not
  g121
  (
    n126,
    n41
  );


  buf
  g122
  (
    n215,
    n55
  );


  buf
  g123
  (
    n314,
    n71
  );


  not
  g124
  (
    n181,
    n37
  );


  not
  g125
  (
    n178,
    n36
  );


  not
  g126
  (
    n185,
    n26
  );


  not
  g127
  (
    n224,
    n63
  );


  not
  g128
  (
    n302,
    n32
  );


  buf
  g129
  (
    n309,
    n40
  );


  not
  g130
  (
    n148,
    n48
  );


  buf
  g131
  (
    n325,
    n43
  );


  not
  g132
  (
    n169,
    n66
  );


  not
  g133
  (
    n348,
    n22
  );


  not
  g134
  (
    n190,
    n54
  );


  not
  g135
  (
    n180,
    n42
  );


  not
  g136
  (
    n198,
    n60
  );


  buf
  g137
  (
    n269,
    n20
  );


  buf
  g138
  (
    n295,
    n68
  );


  buf
  g139
  (
    n320,
    n38
  );


  not
  g140
  (
    n274,
    n59
  );


  not
  g141
  (
    n304,
    n74
  );


  buf
  g142
  (
    n189,
    n51
  );


  buf
  g143
  (
    n262,
    n70
  );


  buf
  g144
  (
    n140,
    n33
  );


  buf
  g145
  (
    n202,
    n47
  );


  buf
  g146
  (
    n211,
    n41
  );


  buf
  g147
  (
    n221,
    n80
  );


  not
  g148
  (
    n167,
    n62
  );


  buf
  g149
  (
    n244,
    n74
  );


  not
  g150
  (
    n164,
    n25
  );


  not
  g151
  (
    n143,
    n61
  );


  not
  g152
  (
    n290,
    n18
  );


  buf
  g153
  (
    n324,
    n46
  );


  not
  g154
  (
    n338,
    n40
  );


  not
  g155
  (
    n187,
    n49
  );


  buf
  g156
  (
    n226,
    n27
  );


  not
  g157
  (
    n253,
    n24
  );


  not
  g158
  (
    n284,
    n63
  );


  buf
  g159
  (
    n227,
    n34
  );


  not
  g160
  (
    n258,
    n36
  );


  not
  g161
  (
    n102,
    n62
  );


  buf
  g162
  (
    n306,
    n84
  );


  not
  g163
  (
    n110,
    n81
  );


  buf
  g164
  (
    n130,
    n33
  );


  not
  g165
  (
    n206,
    n75
  );


  not
  g166
  (
    n175,
    n19
  );


  not
  g167
  (
    n249,
    n44
  );


  buf
  g168
  (
    n323,
    n81
  );


  not
  g169
  (
    n347,
    n70
  );


  not
  g170
  (
    n263,
    n79
  );


  not
  g171
  (
    n158,
    n34
  );


  buf
  g172
  (
    n147,
    n84
  );


  not
  g173
  (
    n305,
    n82
  );


  buf
  g174
  (
    n330,
    n67
  );


  not
  g175
  (
    n303,
    n45
  );


  not
  g176
  (
    n163,
    n60
  );


  not
  g177
  (
    n288,
    n58
  );


  buf
  g178
  (
    n218,
    n49
  );


  not
  g179
  (
    n219,
    n21
  );


  buf
  g180
  (
    n171,
    n61
  );


  buf
  g181
  (
    n308,
    n50
  );


  buf
  g182
  (
    n207,
    n52
  );


  buf
  g183
  (
    n335,
    n28
  );


  buf
  g184
  (
    n353,
    n85
  );


  buf
  g185
  (
    n316,
    n23
  );


  not
  g186
  (
    n356,
    n25
  );


  buf
  g187
  (
    n193,
    n45
  );


  buf
  g188
  (
    n201,
    n79
  );


  buf
  g189
  (
    n337,
    n48
  );


  buf
  g190
  (
    n94,
    n30
  );


  buf
  g191
  (
    KeyWire_0_19,
    n49
  );


  not
  g192
  (
    n111,
    n31
  );


  buf
  g193
  (
    n133,
    n85
  );


  not
  g194
  (
    n217,
    n21
  );


  not
  g195
  (
    n247,
    n24
  );


  buf
  g196
  (
    n138,
    n46
  );


  buf
  g197
  (
    n301,
    n47
  );


  buf
  g198
  (
    n255,
    n47
  );


  buf
  g199
  (
    n96,
    n19
  );


  buf
  g200
  (
    n214,
    n18
  );


  not
  g201
  (
    n136,
    n64
  );


  buf
  g202
  (
    n318,
    n85
  );


  not
  g203
  (
    n357,
    n27
  );


  not
  g204
  (
    n184,
    n33
  );


  buf
  g205
  (
    n222,
    n54
  );


  not
  g206
  (
    n254,
    n27
  );


  not
  g207
  (
    n299,
    n25
  );


  buf
  g208
  (
    n300,
    n85
  );


  buf
  g209
  (
    n128,
    n39
  );


  buf
  g210
  (
    n237,
    n22
  );


  buf
  g211
  (
    n245,
    n28
  );


  not
  g212
  (
    n101,
    n79
  );


  buf
  g213
  (
    n333,
    n51
  );


  not
  g214
  (
    n139,
    n44
  );


  buf
  g215
  (
    n205,
    n52
  );


  not
  g216
  (
    n313,
    n55
  );


  not
  g217
  (
    n327,
    n80
  );


  not
  g218
  (
    n129,
    n72
  );


  not
  g219
  (
    n162,
    n31
  );


  not
  g220
  (
    n270,
    n40
  );


  buf
  g221
  (
    n332,
    n55
  );


  buf
  g222
  (
    KeyWire_0_11,
    n80
  );


  buf
  g223
  (
    n326,
    n73
  );


  buf
  g224
  (
    n154,
    n82
  );


  buf
  g225
  (
    n354,
    n70
  );


  buf
  g226
  (
    n277,
    n39
  );


  not
  g227
  (
    n192,
    n36
  );


  not
  g228
  (
    n310,
    n68
  );


  buf
  g229
  (
    n334,
    n60
  );


  buf
  g230
  (
    n213,
    n60
  );


  buf
  g231
  (
    n186,
    n20
  );


  not
  g232
  (
    n235,
    n35
  );


  not
  g233
  (
    n345,
    n32
  );


  not
  g234
  (
    n116,
    n33
  );


  not
  g235
  (
    n272,
    n71
  );


  not
  g236
  (
    n236,
    n82
  );


  not
  g237
  (
    n246,
    n21
  );


  buf
  g238
  (
    n118,
    n22
  );


  buf
  g239
  (
    n267,
    n49
  );


  not
  g240
  (
    n243,
    n39
  );


  buf
  g241
  (
    n87,
    n54
  );


  not
  g242
  (
    n349,
    n29
  );


  buf
  g243
  (
    n233,
    n58
  );


  buf
  g244
  (
    n271,
    n69
  );


  not
  g245
  (
    n344,
    n74
  );


  not
  g246
  (
    n266,
    n83
  );


  not
  g247
  (
    n257,
    n75
  );


  buf
  g248
  (
    n106,
    n64
  );


  not
  g249
  (
    n287,
    n50
  );


  not
  g250
  (
    n121,
    n62
  );


  not
  g251
  (
    n315,
    n34
  );


  not
  g252
  (
    n355,
    n65
  );


  buf
  g253
  (
    n289,
    n20
  );


  not
  g254
  (
    n322,
    n83
  );


  not
  g255
  (
    n127,
    n83
  );


  not
  g256
  (
    n240,
    n78
  );


  buf
  g257
  (
    n103,
    n64
  );


  not
  g258
  (
    n250,
    n48
  );


  not
  g259
  (
    n312,
    n50
  );


  not
  g260
  (
    n160,
    n35
  );


  not
  g261
  (
    n231,
    n26
  );


  not
  g262
  (
    n131,
    n43
  );


  not
  g263
  (
    n152,
    n69
  );


  not
  g264
  (
    n196,
    n73
  );


  not
  g265
  (
    n238,
    n39
  );


  not
  g266
  (
    n292,
    n27
  );


  buf
  g267
  (
    n174,
    n54
  );


  buf
  g268
  (
    n228,
    n67
  );


  buf
  g269
  (
    n340,
    n29
  );


  buf
  g270
  (
    n229,
    n22
  );


  not
  g271
  (
    n165,
    n59
  );


  not
  g272
  (
    n275,
    n76
  );


  buf
  g273
  (
    n328,
    n77
  );


  not
  g274
  (
    n297,
    n67
  );


  not
  g275
  (
    n172,
    n65
  );


  buf
  g276
  (
    n122,
    n23
  );


  not
  g277
  (
    n161,
    n26
  );


  not
  g278
  (
    n342,
    n76
  );


  not
  g279
  (
    n155,
    n57
  );


  buf
  g280
  (
    n283,
    n28
  );


  not
  g281
  (
    n220,
    n73
  );


  buf
  g282
  (
    n145,
    n23
  );


  not
  g283
  (
    n241,
    n48
  );


  buf
  g284
  (
    n90,
    n67
  );


  buf
  g285
  (
    n98,
    n66
  );


  not
  g286
  (
    n170,
    n45
  );


  buf
  g287
  (
    n282,
    n31
  );


  buf
  g288
  (
    n109,
    n70
  );


  buf
  g289
  (
    n285,
    n30
  );


  not
  g290
  (
    n296,
    n65
  );


  buf
  g291
  (
    n108,
    n30
  );


  not
  g292
  (
    n156,
    n61
  );


  buf
  g293
  (
    n179,
    n47
  );


  buf
  g294
  (
    n197,
    n32
  );


  not
  g295
  (
    n113,
    n58
  );


  not
  g296
  (
    n142,
    n19
  );


  not
  g297
  (
    n166,
    n18
  );


  buf
  g298
  (
    n276,
    n63
  );


  not
  g299
  (
    n256,
    n80
  );


  not
  g300
  (
    n188,
    n32
  );


  buf
  g301
  (
    n146,
    n59
  );


  not
  g302
  (
    n286,
    n46
  );


  buf
  g303
  (
    n199,
    n28
  );


  not
  g304
  (
    n251,
    n56
  );


  buf
  g305
  (
    n157,
    n24
  );


  not
  g306
  (
    n168,
    n21
  );


  buf
  g307
  (
    n281,
    n55
  );


  buf
  g308
  (
    n100,
    n42
  );


  not
  g309
  (
    n137,
    n65
  );


  buf
  g310
  (
    n232,
    n58
  );


  not
  g311
  (
    n191,
    n34
  );


  buf
  g312
  (
    n104,
    n69
  );


  not
  g313
  (
    n124,
    n31
  );


  not
  g314
  (
    n351,
    n82
  );


  buf
  g315
  (
    n352,
    n61
  );


  not
  g316
  (
    n293,
    n37
  );


  not
  g317
  (
    n216,
    n23
  );


  not
  g318
  (
    n182,
    n56
  );


  not
  g319
  (
    n173,
    n53
  );


  not
  g320
  (
    n317,
    n24
  );


  buf
  g321
  (
    n204,
    n51
  );


  not
  g322
  (
    n230,
    n66
  );


  buf
  g323
  (
    n350,
    n62
  );


  not
  g324
  (
    n125,
    n81
  );


  not
  g325
  (
    n177,
    n84
  );


  not
  g326
  (
    n105,
    n42
  );


  buf
  g327
  (
    n141,
    n20
  );


  not
  g328
  (
    n210,
    n45
  );


  buf
  g329
  (
    n264,
    n41
  );


  not
  g330
  (
    n291,
    n79
  );


  buf
  g331
  (
    n132,
    n26
  );


  not
  g332
  (
    n260,
    n68
  );


  not
  g333
  (
    n117,
    n72
  );


  not
  g334
  (
    n319,
    n35
  );


  buf
  g335
  (
    n86,
    n72
  );


  not
  g336
  (
    n91,
    n75
  );


  not
  g337
  (
    n149,
    n42
  );


  buf
  g338
  (
    n95,
    n44
  );


  not
  g339
  (
    n159,
    n30
  );


  buf
  g340
  (
    n935,
    n177
  );


  not
  g341
  (
    n376,
    n272
  );


  not
  g342
  (
    n1166,
    n212
  );


  buf
  g343
  (
    n804,
    n142
  );


  not
  g344
  (
    n1189,
    n341
  );


  not
  g345
  (
    n921,
    n135
  );


  buf
  g346
  (
    n525,
    n217
  );


  not
  g347
  (
    n392,
    n196
  );


  buf
  g348
  (
    n941,
    n173
  );


  not
  g349
  (
    n1170,
    n292
  );


  buf
  g350
  (
    n1306,
    n221
  );


  buf
  g351
  (
    n491,
    n129
  );


  buf
  g352
  (
    n956,
    n325
  );


  buf
  g353
  (
    n817,
    n324
  );


  buf
  g354
  (
    n977,
    n226
  );


  buf
  g355
  (
    n918,
    n123
  );


  buf
  g356
  (
    n829,
    n162
  );


  not
  g357
  (
    n1262,
    n188
  );


  buf
  g358
  (
    n1136,
    n144
  );


  buf
  g359
  (
    n486,
    n312
  );


  buf
  g360
  (
    n1148,
    n332
  );


  not
  g361
  (
    n542,
    n119
  );


  not
  g362
  (
    n985,
    n144
  );


  not
  g363
  (
    n482,
    n165
  );


  buf
  g364
  (
    n961,
    n110
  );


  buf
  g365
  (
    n911,
    n329
  );


  not
  g366
  (
    n646,
    n339
  );


  not
  g367
  (
    n1362,
    n322
  );


  not
  g368
  (
    n791,
    n128
  );


  buf
  g369
  (
    n932,
    n149
  );


  not
  g370
  (
    n776,
    n161
  );


  not
  g371
  (
    n973,
    n98
  );


  not
  g372
  (
    n1358,
    n262
  );


  not
  g373
  (
    n898,
    n173
  );


  buf
  g374
  (
    n805,
    n214
  );


  not
  g375
  (
    n758,
    n142
  );


  not
  g376
  (
    n778,
    n241
  );


  buf
  g377
  (
    n936,
    n213
  );


  not
  g378
  (
    n1337,
    n290
  );


  not
  g379
  (
    n663,
    n190
  );


  not
  g380
  (
    n1131,
    n242
  );


  buf
  g381
  (
    n636,
    n113
  );


  not
  g382
  (
    n1308,
    n161
  );


  not
  g383
  (
    n1162,
    n145
  );


  not
  g384
  (
    n575,
    n227
  );


  not
  g385
  (
    n782,
    n214
  );


  buf
  g386
  (
    n1041,
    n213
  );


  not
  g387
  (
    n602,
    n228
  );


  buf
  g388
  (
    n1156,
    n113
  );


  buf
  g389
  (
    n1050,
    n155
  );


  not
  g390
  (
    n628,
    n115
  );


  buf
  g391
  (
    KeyWire_0_6,
    n185
  );


  not
  g392
  (
    n814,
    n204
  );


  not
  g393
  (
    KeyWire_0_31,
    n170
  );


  not
  g394
  (
    n780,
    n180
  );


  buf
  g395
  (
    n879,
    n298
  );


  buf
  g396
  (
    n1099,
    n167
  );


  not
  g397
  (
    n1333,
    n304
  );


  buf
  g398
  (
    n623,
    n154
  );


  not
  g399
  (
    n603,
    n273
  );


  buf
  g400
  (
    n1304,
    n277
  );


  not
  g401
  (
    n1270,
    n247
  );


  buf
  g402
  (
    n387,
    n243
  );


  not
  g403
  (
    n729,
    n246
  );


  not
  g404
  (
    n1251,
    n146
  );


  not
  g405
  (
    n893,
    n349
  );


  buf
  g406
  (
    n1079,
    n258
  );


  not
  g407
  (
    n1284,
    n155
  );


  buf
  g408
  (
    n1094,
    n202
  );


  not
  g409
  (
    n665,
    n152
  );


  not
  g410
  (
    n604,
    n153
  );


  buf
  g411
  (
    n1017,
    n345
  );


  not
  g412
  (
    n1240,
    n225
  );


  not
  g413
  (
    n933,
    n309
  );


  not
  g414
  (
    n1153,
    n195
  );


  not
  g415
  (
    n1159,
    n277
  );


  buf
  g416
  (
    n828,
    n167
  );


  buf
  g417
  (
    n582,
    n239
  );


  buf
  g418
  (
    n1207,
    n273
  );


  not
  g419
  (
    n620,
    n327
  );


  buf
  g420
  (
    n610,
    n265
  );


  buf
  g421
  (
    n966,
    n250
  );


  not
  g422
  (
    n1256,
    n261
  );


  buf
  g423
  (
    n1250,
    n166
  );


  not
  g424
  (
    n987,
    n295
  );


  not
  g425
  (
    n913,
    n308
  );


  not
  g426
  (
    n1070,
    n107
  );


  buf
  g427
  (
    n1291,
    n345
  );


  not
  g428
  (
    n1146,
    n163
  );


  buf
  g429
  (
    n710,
    n103
  );


  buf
  g430
  (
    n1283,
    n135
  );


  buf
  g431
  (
    n1003,
    n213
  );


  not
  g432
  (
    n470,
    n138
  );


  buf
  g433
  (
    n1255,
    n231
  );


  not
  g434
  (
    n1077,
    n89
  );


  buf
  g435
  (
    n1230,
    n347
  );


  buf
  g436
  (
    n1212,
    n337
  );


  buf
  g437
  (
    n407,
    n257
  );


  not
  g438
  (
    n381,
    n224
  );


  buf
  g439
  (
    n1025,
    n135
  );


  not
  g440
  (
    n450,
    n245
  );


  not
  g441
  (
    n1199,
    n86
  );


  not
  g442
  (
    n998,
    n294
  );


  not
  g443
  (
    n606,
    n237
  );


  buf
  g444
  (
    n592,
    n191
  );


  not
  g445
  (
    n1160,
    n298
  );


  not
  g446
  (
    n1062,
    n339
  );


  buf
  g447
  (
    n1059,
    n192
  );


  buf
  g448
  (
    n551,
    n303
  );


  buf
  g449
  (
    n594,
    n197
  );


  not
  g450
  (
    n437,
    n90
  );


  buf
  g451
  (
    n930,
    n234
  );


  not
  g452
  (
    n1368,
    n225
  );


  buf
  g453
  (
    n825,
    n280
  );


  buf
  g454
  (
    n666,
    n299
  );


  buf
  g455
  (
    n616,
    n288
  );


  not
  g456
  (
    n1098,
    n140
  );


  buf
  g457
  (
    n1219,
    n229
  );


  buf
  g458
  (
    n945,
    n324
  );


  not
  g459
  (
    n769,
    n120
  );


  buf
  g460
  (
    n990,
    n113
  );


  not
  g461
  (
    n1380,
    n272
  );


  buf
  g462
  (
    n1133,
    n86
  );


  buf
  g463
  (
    n1005,
    n216
  );


  not
  g464
  (
    n870,
    n167
  );


  not
  g465
  (
    n578,
    n176
  );


  buf
  g466
  (
    n746,
    n152
  );


  buf
  g467
  (
    n1247,
    n121
  );


  buf
  g468
  (
    n1272,
    n209
  );


  not
  g469
  (
    n652,
    n256
  );


  buf
  g470
  (
    n402,
    n339
  );


  not
  g471
  (
    n881,
    n350
  );


  buf
  g472
  (
    n757,
    n227
  );


  buf
  g473
  (
    n827,
    n91
  );


  buf
  g474
  (
    n1329,
    n245
  );


  buf
  g475
  (
    n1042,
    n253
  );


  buf
  g476
  (
    n970,
    n319
  );


  not
  g477
  (
    n873,
    n166
  );


  not
  g478
  (
    n1027,
    n189
  );


  buf
  g479
  (
    n896,
    n203
  );


  buf
  g480
  (
    n739,
    n154
  );


  not
  g481
  (
    n647,
    n274
  );


  buf
  g482
  (
    n656,
    n296
  );


  not
  g483
  (
    n1363,
    n263
  );


  not
  g484
  (
    n502,
    n232
  );


  not
  g485
  (
    n1327,
    n255
  );


  not
  g486
  (
    n607,
    n125
  );


  not
  g487
  (
    n454,
    n191
  );


  not
  g488
  (
    n438,
    n203
  );


  not
  g489
  (
    n971,
    n141
  );


  buf
  g490
  (
    n1158,
    n291
  );


  buf
  g491
  (
    n1246,
    n330
  );


  not
  g492
  (
    n489,
    n299
  );


  not
  g493
  (
    n609,
    n329
  );


  not
  g494
  (
    n1260,
    n289
  );


  buf
  g495
  (
    n810,
    n251
  );


  not
  g496
  (
    n587,
    n158
  );


  not
  g497
  (
    n877,
    n260
  );


  buf
  g498
  (
    n547,
    n288
  );


  buf
  g499
  (
    n528,
    n290
  );


  not
  g500
  (
    n1382,
    n160
  );


  not
  g501
  (
    n958,
    n158
  );


  buf
  g502
  (
    n1043,
    n333
  );


  buf
  g503
  (
    n1107,
    n89
  );


  not
  g504
  (
    n1374,
    n262
  );


  not
  g505
  (
    n513,
    n145
  );


  buf
  g506
  (
    n888,
    n280
  );


  not
  g507
  (
    n1319,
    n128
  );


  buf
  g508
  (
    n670,
    n264
  );


  not
  g509
  (
    n1195,
    n198
  );


  not
  g510
  (
    n382,
    n228
  );


  not
  g511
  (
    n1299,
    n348
  );


  not
  g512
  (
    n480,
    n299
  );


  not
  g513
  (
    n1209,
    n268
  );


  not
  g514
  (
    n978,
    n216
  );


  not
  g515
  (
    n458,
    n94
  );


  buf
  g516
  (
    n1048,
    n189
  );


  buf
  g517
  (
    n1378,
    n216
  );


  buf
  g518
  (
    n598,
    n132
  );


  buf
  g519
  (
    n1128,
    n139
  );


  not
  g520
  (
    n1175,
    n314
  );


  not
  g521
  (
    n484,
    n293
  );


  buf
  g522
  (
    n860,
    n115
  );


  buf
  g523
  (
    n940,
    n155
  );


  buf
  g524
  (
    n588,
    n122
  );


  buf
  g525
  (
    n546,
    n142
  );


  not
  g526
  (
    n1089,
    n95
  );


  not
  g527
  (
    n493,
    n263
  );


  not
  g528
  (
    n629,
    n221
  );


  buf
  g529
  (
    n537,
    n248
  );


  not
  g530
  (
    n1084,
    n278
  );


  buf
  g531
  (
    n612,
    n344
  );


  buf
  g532
  (
    n1091,
    n184
  );


  buf
  g533
  (
    n902,
    n97
  );


  not
  g534
  (
    n1036,
    n143
  );


  not
  g535
  (
    n1371,
    n192
  );


  not
  g536
  (
    n1085,
    n216
  );


  not
  g537
  (
    KeyWire_0_1,
    n183
  );


  buf
  g538
  (
    n1155,
    n250
  );


  not
  g539
  (
    n464,
    n283
  );


  not
  g540
  (
    n1102,
    n156
  );


  buf
  g541
  (
    n455,
    n224
  );


  buf
  g542
  (
    n643,
    n87
  );


  buf
  g543
  (
    n457,
    n267
  );


  buf
  g544
  (
    n723,
    n182
  );


  buf
  g545
  (
    n914,
    n214
  );


  not
  g546
  (
    n436,
    n110
  );


  not
  g547
  (
    n733,
    n303
  );


  buf
  g548
  (
    n1286,
    n308
  );


  buf
  g549
  (
    n763,
    n311
  );


  not
  g550
  (
    n874,
    n151
  );


  buf
  g551
  (
    n462,
    n306
  );


  not
  g552
  (
    n1228,
    n330
  );


  buf
  g553
  (
    n851,
    n350
  );


  buf
  g554
  (
    n713,
    n301
  );


  buf
  g555
  (
    n1068,
    n315
  );


  buf
  g556
  (
    n944,
    n266
  );


  buf
  g557
  (
    n989,
    n230
  );


  not
  g558
  (
    n1237,
    n279
  );


  buf
  g559
  (
    n712,
    n111
  );


  buf
  g560
  (
    n807,
    n91
  );


  buf
  g561
  (
    n1033,
    n94
  );


  not
  g562
  (
    n836,
    n240
  );


  not
  g563
  (
    n802,
    n174
  );


  not
  g564
  (
    n826,
    n289
  );


  not
  g565
  (
    n760,
    n264
  );


  buf
  g566
  (
    n658,
    n297
  );


  buf
  g567
  (
    n1058,
    n94
  );


  buf
  g568
  (
    n1346,
    n211
  );


  buf
  g569
  (
    n1002,
    n187
  );


  not
  g570
  (
    n1172,
    n181
  );


  not
  g571
  (
    n878,
    n277
  );


  buf
  g572
  (
    n1385,
    n272
  );


  buf
  g573
  (
    n899,
    n126
  );


  buf
  g574
  (
    n566,
    n214
  );


  buf
  g575
  (
    n808,
    n89
  );


  buf
  g576
  (
    n984,
    n168
  );


  not
  g577
  (
    n1309,
    n312
  );


  not
  g578
  (
    n649,
    n186
  );


  not
  g579
  (
    n1163,
    n157
  );


  buf
  g580
  (
    n813,
    n284
  );


  buf
  g581
  (
    n1197,
    n144
  );


  buf
  g582
  (
    n953,
    n88
  );


  not
  g583
  (
    n988,
    n318
  );


  buf
  g584
  (
    n524,
    n151
  );


  not
  g585
  (
    n1100,
    n134
  );


  not
  g586
  (
    n1145,
    n105
  );


  buf
  g587
  (
    n481,
    n265
  );


  not
  g588
  (
    n1258,
    n301
  );


  buf
  g589
  (
    n1072,
    n127
  );


  not
  g590
  (
    n1106,
    n245
  );


  buf
  g591
  (
    n752,
    n125
  );


  not
  g592
  (
    n1118,
    n118
  );


  not
  g593
  (
    n687,
    n233
  );


  buf
  g594
  (
    n522,
    n289
  );


  not
  g595
  (
    n1092,
    n269
  );


  buf
  g596
  (
    n1332,
    n110
  );


  not
  g597
  (
    n1294,
    n269
  );


  buf
  g598
  (
    n861,
    n157
  );


  buf
  g599
  (
    n815,
    n300
  );


  buf
  g600
  (
    n1387,
    n198
  );


  buf
  g601
  (
    n1113,
    n111
  );


  buf
  g602
  (
    n685,
    n305
  );


  not
  g603
  (
    n789,
    n321
  );


  not
  g604
  (
    n444,
    n250
  );


  buf
  g605
  (
    n679,
    n330
  );


  buf
  g606
  (
    n1220,
    n162
  );


  not
  g607
  (
    n573,
    n318
  );


  buf
  g608
  (
    n1035,
    n210
  );


  buf
  g609
  (
    KeyWire_0_24,
    n288
  );


  not
  g610
  (
    n391,
    n329
  );


  not
  g611
  (
    n377,
    n194
  );


  not
  g612
  (
    n749,
    n349
  );


  not
  g613
  (
    n714,
    n244
  );


  buf
  g614
  (
    n1295,
    n261
  );


  not
  g615
  (
    n580,
    n240
  );


  buf
  g616
  (
    n532,
    n246
  );


  not
  g617
  (
    n703,
    n259
  );


  buf
  g618
  (
    n765,
    n279
  );


  not
  g619
  (
    n1039,
    n95
  );


  buf
  g620
  (
    n1204,
    n251
  );


  not
  g621
  (
    n734,
    n348
  );


  not
  g622
  (
    n625,
    n274
  );


  buf
  g623
  (
    n473,
    n101
  );


  buf
  g624
  (
    n787,
    n278
  );


  buf
  g625
  (
    n1047,
    n139
  );


  not
  g626
  (
    n1190,
    n309
  );


  buf
  g627
  (
    n982,
    n218
  );


  not
  g628
  (
    n624,
    n236
  );


  buf
  g629
  (
    n1265,
    n323
  );


  buf
  g630
  (
    n1157,
    n310
  );


  buf
  g631
  (
    n891,
    n116
  );


  not
  g632
  (
    n1184,
    n116
  );


  not
  g633
  (
    n718,
    n327
  );


  not
  g634
  (
    n634,
    n255
  );


  not
  g635
  (
    n363,
    n133
  );


  buf
  g636
  (
    n835,
    n259
  );


  not
  g637
  (
    n567,
    n223
  );


  buf
  g638
  (
    n696,
    n314
  );


  not
  g639
  (
    n1046,
    n257
  );


  not
  g640
  (
    n853,
    n286
  );


  not
  g641
  (
    n1105,
    n235
  );


  buf
  g642
  (
    n880,
    n146
  );


  buf
  g643
  (
    n1292,
    n88
  );


  buf
  g644
  (
    n1021,
    n304
  );


  not
  g645
  (
    n1213,
    n97
  );


  buf
  g646
  (
    n919,
    n108
  );


  buf
  g647
  (
    n467,
    n161
  );


  not
  g648
  (
    n405,
    n148
  );


  buf
  g649
  (
    n980,
    n248
  );


  buf
  g650
  (
    n793,
    n145
  );


  not
  g651
  (
    n1132,
    n109
  );


  buf
  g652
  (
    n673,
    n212
  );


  not
  g653
  (
    n618,
    n177
  );


  not
  g654
  (
    n1009,
    n307
  );


  buf
  g655
  (
    n886,
    n96
  );


  buf
  g656
  (
    n1225,
    n262
  );


  not
  g657
  (
    n1242,
    n101
  );


  not
  g658
  (
    n1241,
    n204
  );


  buf
  g659
  (
    n1143,
    n231
  );


  buf
  g660
  (
    n715,
    n328
  );


  not
  g661
  (
    n463,
    n331
  );


  buf
  g662
  (
    n635,
    n274
  );


  buf
  g663
  (
    n740,
    n215
  );


  buf
  g664
  (
    n1305,
    n193
  );


  not
  g665
  (
    n736,
    n321
  );


  not
  g666
  (
    n380,
    n271
  );


  not
  g667
  (
    n964,
    n102
  );


  not
  g668
  (
    n654,
    n327
  );


  buf
  g669
  (
    n975,
    n87
  );


  not
  g670
  (
    n837,
    n287
  );


  not
  g671
  (
    n579,
    n261
  );


  buf
  g672
  (
    n1257,
    n221
  );


  buf
  g673
  (
    n1178,
    n219
  );


  not
  g674
  (
    n1124,
    n351
  );


  not
  g675
  (
    n617,
    n201
  );


  not
  g676
  (
    n1171,
    n114
  );


  not
  g677
  (
    n759,
    n229
  );


  not
  g678
  (
    n564,
    n313
  );


  not
  g679
  (
    n570,
    n148
  );


  not
  g680
  (
    n1310,
    n320
  );


  buf
  g681
  (
    n422,
    n335
  );


  buf
  g682
  (
    n526,
    n139
  );


  not
  g683
  (
    n840,
    n116
  );


  not
  g684
  (
    n699,
    n339
  );


  not
  g685
  (
    n386,
    n124
  );


  not
  g686
  (
    n1183,
    n169
  );


  buf
  g687
  (
    n1269,
    n141
  );


  not
  g688
  (
    n1114,
    n104
  );


  buf
  g689
  (
    n1187,
    n158
  );


  buf
  g690
  (
    n745,
    n295
  );


  buf
  g691
  (
    n426,
    n117
  );


  not
  g692
  (
    n1312,
    n184
  );


  not
  g693
  (
    n839,
    n277
  );


  buf
  g694
  (
    n1227,
    n224
  );


  buf
  g695
  (
    n499,
    n211
  );


  not
  g696
  (
    n931,
    n180
  );


  not
  g697
  (
    n1173,
    n104
  );


  not
  g698
  (
    n1116,
    n275
  );


  not
  g699
  (
    n995,
    n275
  );


  not
  g700
  (
    n927,
    n120
  );


  buf
  g701
  (
    n395,
    n294
  );


  buf
  g702
  (
    n1229,
    n342
  );


  not
  g703
  (
    n1315,
    n105
  );


  buf
  g704
  (
    KeyWire_0_21,
    n86
  );


  buf
  g705
  (
    n748,
    n301
  );


  not
  g706
  (
    n994,
    n319
  );


  not
  g707
  (
    n1108,
    n242
  );


  not
  g708
  (
    n1233,
    n340
  );


  buf
  g709
  (
    n1224,
    n112
  );


  not
  g710
  (
    n1115,
    n131
  );


  buf
  g711
  (
    n581,
    n302
  );


  buf
  g712
  (
    n417,
    n150
  );


  not
  g713
  (
    n1140,
    n168
  );


  not
  g714
  (
    n716,
    n202
  );


  not
  g715
  (
    n456,
    n293
  );


  buf
  g716
  (
    n706,
    n222
  );


  not
  g717
  (
    n479,
    n347
  );


  not
  g718
  (
    n1288,
    n285
  );


  not
  g719
  (
    n691,
    n306
  );


  buf
  g720
  (
    n969,
    n194
  );


  not
  g721
  (
    n447,
    n312
  );


  not
  g722
  (
    n1348,
    n291
  );


  not
  g723
  (
    n1210,
    n220
  );


  buf
  g724
  (
    n890,
    n338
  );


  buf
  g725
  (
    n514,
    n309
  );


  not
  g726
  (
    n585,
    n336
  );


  buf
  g727
  (
    n690,
    n333
  );


  not
  g728
  (
    n731,
    n282
  );


  buf
  g729
  (
    n468,
    n293
  );


  not
  g730
  (
    n800,
    n283
  );


  buf
  g731
  (
    n615,
    n230
  );


  buf
  g732
  (
    n571,
    n226
  );


  buf
  g733
  (
    n770,
    n230
  );


  not
  g734
  (
    n1277,
    n321
  );


  buf
  g735
  (
    n533,
    n171
  );


  buf
  g736
  (
    n1355,
    n124
  );


  buf
  g737
  (
    n697,
    n170
  );


  buf
  g738
  (
    n605,
    n182
  );


  buf
  g739
  (
    n419,
    n344
  );


  buf
  g740
  (
    n903,
    n345
  );


  buf
  g741
  (
    n680,
    n223
  );


  not
  g742
  (
    n675,
    n346
  );


  buf
  g743
  (
    n856,
    n129
  );


  not
  g744
  (
    n1066,
    n281
  );


  not
  g745
  (
    n859,
    n110
  );


  not
  g746
  (
    n809,
    n336
  );


  not
  g747
  (
    n997,
    n274
  );


  buf
  g748
  (
    n867,
    n87
  );


  not
  g749
  (
    n938,
    n159
  );


  buf
  g750
  (
    n1120,
    n220
  );


  not
  g751
  (
    n1038,
    n199
  );


  buf
  g752
  (
    n1142,
    n253
  );


  not
  g753
  (
    n857,
    n198
  );


  buf
  g754
  (
    n415,
    n152
  );


  not
  g755
  (
    n425,
    n207
  );


  buf
  g756
  (
    n767,
    n270
  );


  not
  g757
  (
    n981,
    n208
  );


  not
  g758
  (
    n1008,
    n178
  );


  not
  g759
  (
    n403,
    n156
  );


  not
  g760
  (
    n560,
    n252
  );


  buf
  g761
  (
    n671,
    n194
  );


  buf
  g762
  (
    n1064,
    n149
  );


  buf
  g763
  (
    n1336,
    n238
  );


  not
  g764
  (
    n901,
    n119
  );


  buf
  g765
  (
    n892,
    n350
  );


  not
  g766
  (
    n1375,
    n353
  );


  buf
  g767
  (
    n972,
    n282
  );


  buf
  g768
  (
    n872,
    n342
  );


  buf
  g769
  (
    n768,
    n280
  );


  buf
  g770
  (
    n926,
    n191
  );


  buf
  g771
  (
    n563,
    n230
  );


  buf
  g772
  (
    n1268,
    n302
  );


  buf
  g773
  (
    n474,
    n264
  );


  not
  g774
  (
    n1264,
    n164
  );


  buf
  g775
  (
    n1188,
    n182
  );


  buf
  g776
  (
    n1152,
    n246
  );


  buf
  g777
  (
    n889,
    n170
  );


  buf
  g778
  (
    n572,
    n178
  );


  buf
  g779
  (
    n488,
    n262
  );


  not
  g780
  (
    n370,
    n273
  );


  not
  g781
  (
    n820,
    n174
  );


  not
  g782
  (
    n421,
    n316
  );


  buf
  g783
  (
    n700,
    n132
  );


  buf
  g784
  (
    n601,
    n320
  );


  buf
  g785
  (
    n1314,
    n163
  );


  not
  g786
  (
    n883,
    n181
  );


  not
  g787
  (
    n1201,
    n300
  );


  buf
  g788
  (
    n1298,
    n280
  );


  not
  g789
  (
    n556,
    n106
  );


  buf
  g790
  (
    n843,
    n159
  );


  not
  g791
  (
    n1287,
    n350
  );


  buf
  g792
  (
    n507,
    n354
  );


  not
  g793
  (
    n631,
    n332
  );


  buf
  g794
  (
    n576,
    n241
  );


  not
  g795
  (
    n641,
    n136
  );


  not
  g796
  (
    n1364,
    n225
  );


  buf
  g797
  (
    n364,
    n239
  );


  not
  g798
  (
    n1279,
    n222
  );


  buf
  g799
  (
    n954,
    n137
  );


  buf
  g800
  (
    n414,
    n270
  );


  not
  g801
  (
    n637,
    n342
  );


  buf
  g802
  (
    n864,
    n185
  );


  buf
  g803
  (
    n367,
    n103
  );


  not
  g804
  (
    n627,
    n187
  );


  not
  g805
  (
    n411,
    n164
  );


  not
  g806
  (
    n952,
    n162
  );


  not
  g807
  (
    n897,
    n181
  );


  buf
  g808
  (
    n1231,
    n276
  );


  buf
  g809
  (
    n553,
    n311
  );


  not
  g810
  (
    n711,
    n223
  );


  buf
  g811
  (
    n957,
    n207
  );


  not
  g812
  (
    n1007,
    n234
  );


  not
  g813
  (
    n743,
    n172
  );


  buf
  g814
  (
    n781,
    n315
  );


  buf
  g815
  (
    n535,
    n175
  );


  not
  g816
  (
    n1326,
    n343
  );


  buf
  g817
  (
    n692,
    n90
  );


  buf
  g818
  (
    n949,
    n346
  );


  buf
  g819
  (
    n812,
    n336
  );


  buf
  g820
  (
    KeyWire_0_28,
    n344
  );


  not
  g821
  (
    n397,
    n292
  );


  not
  g822
  (
    n632,
    n93
  );


  not
  g823
  (
    n1370,
    n353
  );


  buf
  g824
  (
    n420,
    n167
  );


  buf
  g825
  (
    n429,
    n170
  );


  buf
  g826
  (
    n1141,
    n93
  );


  buf
  g827
  (
    n1330,
    n247
  );


  buf
  g828
  (
    KeyWire_0_26,
    n310
  );


  buf
  g829
  (
    n589,
    n176
  );


  not
  g830
  (
    n1061,
    n137
  );


  not
  g831
  (
    n1351,
    n268
  );


  not
  g832
  (
    n478,
    n106
  );


  buf
  g833
  (
    n369,
    n132
  );


  not
  g834
  (
    n920,
    n315
  );


  buf
  g835
  (
    n909,
    n221
  );


  not
  g836
  (
    n451,
    n96
  );


  buf
  g837
  (
    n569,
    n142
  );


  buf
  g838
  (
    n694,
    n139
  );


  not
  g839
  (
    n1129,
    n175
  );


  buf
  g840
  (
    n515,
    n96
  );


  not
  g841
  (
    n667,
    n173
  );


  buf
  g842
  (
    n494,
    n328
  );


  buf
  g843
  (
    n1119,
    n285
  );


  not
  g844
  (
    n471,
    n90
  );


  not
  g845
  (
    n393,
    n163
  );


  not
  g846
  (
    n1376,
    n193
  );


  not
  g847
  (
    n792,
    n152
  );


  not
  g848
  (
    KeyWire_0_22,
    n109
  );


  buf
  g849
  (
    n1232,
    n319
  );


  not
  g850
  (
    n432,
    n288
  );


  buf
  g851
  (
    n639,
    n125
  );


  not
  g852
  (
    n466,
    n195
  );


  buf
  g853
  (
    n1167,
    n261
  );


  not
  g854
  (
    n762,
    n344
  );


  buf
  g855
  (
    n678,
    n253
  );


  not
  g856
  (
    n1049,
    n147
  );


  not
  g857
  (
    n1016,
    n176
  );


  not
  g858
  (
    n593,
    n311
  );


  buf
  g859
  (
    n912,
    n106
  );


  not
  g860
  (
    n430,
    n187
  );


  not
  g861
  (
    n1096,
    n129
  );


  buf
  g862
  (
    n1367,
    n93
  );


  buf
  g863
  (
    n728,
    n317
  );


  not
  g864
  (
    n497,
    n240
  );


  not
  g865
  (
    n1365,
    n281
  );


  not
  g866
  (
    KeyWire_0_5,
    n276
  );


  not
  g867
  (
    n937,
    n209
  );


  buf
  g868
  (
    n841,
    n158
  );


  buf
  g869
  (
    n684,
    n197
  );


  not
  g870
  (
    n362,
    n100
  );


  buf
  g871
  (
    n830,
    n237
  );


  not
  g872
  (
    n1259,
    n324
  );


  not
  g873
  (
    n1243,
    n327
  );


  buf
  g874
  (
    n375,
    n222
  );


  not
  g875
  (
    n1023,
    n191
  );


  buf
  g876
  (
    n503,
    n99
  );


  buf
  g877
  (
    n1067,
    n303
  );


  not
  g878
  (
    n1275,
    n217
  );


  buf
  g879
  (
    n655,
    n219
  );


  buf
  g880
  (
    n950,
    n89
  );


  buf
  g881
  (
    n423,
    n204
  );


  buf
  g882
  (
    n764,
    n133
  );


  buf
  g883
  (
    n934,
    n298
  );


  buf
  g884
  (
    n709,
    n104
  );


  buf
  g885
  (
    n614,
    n267
  );


  not
  g886
  (
    n558,
    n117
  );


  buf
  g887
  (
    n1176,
    n112
  );


  buf
  g888
  (
    n983,
    n188
  );


  not
  g889
  (
    KeyWire_0_14,
    n107
  );


  buf
  g890
  (
    n500,
    n305
  );


  not
  g891
  (
    n705,
    n180
  );


  not
  g892
  (
    n396,
    n308
  );


  buf
  g893
  (
    n1032,
    n150
  );


  not
  g894
  (
    n1198,
    n94
  );


  buf
  g895
  (
    n534,
    n278
  );


  not
  g896
  (
    n1252,
    n123
  );


  buf
  g897
  (
    n409,
    n255
  );


  not
  g898
  (
    n552,
    n118
  );


  not
  g899
  (
    n947,
    n348
  );


  not
  g900
  (
    n738,
    n320
  );


  not
  g901
  (
    n986,
    n159
  );


  not
  g902
  (
    n445,
    n122
  );


  buf
  g903
  (
    n1248,
    n182
  );


  buf
  g904
  (
    n968,
    n213
  );


  buf
  g905
  (
    n1087,
    n92
  );


  buf
  g906
  (
    n1343,
    n257
  );


  not
  g907
  (
    n1109,
    n103
  );


  buf
  g908
  (
    n485,
    n200
  );


  not
  g909
  (
    n477,
    n156
  );


  buf
  g910
  (
    n1073,
    n105
  );


  buf
  g911
  (
    n1111,
    n168
  );


  buf
  g912
  (
    n442,
    n179
  );


  buf
  g913
  (
    n544,
    n270
  );


  not
  g914
  (
    n963,
    n114
  );


  buf
  g915
  (
    n1369,
    n260
  );


  not
  g916
  (
    n657,
    n341
  );


  buf
  g917
  (
    n822,
    n266
  );


  not
  g918
  (
    n400,
    n232
  );


  not
  g919
  (
    n1185,
    n177
  );


  not
  g920
  (
    n1313,
    n115
  );


  not
  g921
  (
    n541,
    n271
  );


  not
  g922
  (
    n755,
    n215
  );


  buf
  g923
  (
    n1101,
    n153
  );


  buf
  g924
  (
    n674,
    n334
  );


  buf
  g925
  (
    n465,
    n138
  );


  buf
  g926
  (
    n1253,
    n138
  );


  not
  g927
  (
    n907,
    n248
  );


  buf
  g928
  (
    n701,
    n102
  );


  buf
  g929
  (
    n461,
    n212
  );


  not
  g930
  (
    n1236,
    n279
  );


  buf
  g931
  (
    n378,
    n258
  );


  buf
  g932
  (
    n404,
    n266
  );


  not
  g933
  (
    n446,
    n236
  );


  not
  g934
  (
    n801,
    n314
  );


  not
  g935
  (
    n644,
    n90
  );


  buf
  g936
  (
    n508,
    n150
  );


  not
  g937
  (
    n516,
    n206
  );


  buf
  g938
  (
    n720,
    n116
  );


  buf
  g939
  (
    n518,
    n189
  );


  not
  g940
  (
    n773,
    n284
  );


  buf
  g941
  (
    n645,
    n302
  );


  not
  g942
  (
    n519,
    n151
  );


  buf
  g943
  (
    n595,
    n237
  );


  buf
  g944
  (
    n398,
    n238
  );


  not
  g945
  (
    n1097,
    n169
  );


  not
  g946
  (
    n529,
    n249
  );


  not
  g947
  (
    n1180,
    n249
  );


  buf
  g948
  (
    n1179,
    n99
  );


  buf
  g949
  (
    n788,
    n322
  );


  buf
  g950
  (
    n662,
    n296
  );


  not
  g951
  (
    n1044,
    n190
  );


  buf
  g952
  (
    n1080,
    n346
  );


  buf
  g953
  (
    n490,
    n303
  );


  not
  g954
  (
    n1297,
    n201
  );


  not
  g955
  (
    n1018,
    n172
  );


  buf
  g956
  (
    n521,
    n229
  );


  not
  g957
  (
    n695,
    n102
  );


  buf
  g958
  (
    n583,
    n325
  );


  not
  g959
  (
    n408,
    n151
  );


  not
  g960
  (
    n1263,
    n294
  );


  not
  g961
  (
    n869,
    n173
  );


  buf
  g962
  (
    n900,
    n330
  );


  not
  g963
  (
    n406,
    n117
  );


  buf
  g964
  (
    n959,
    n296
  );


  buf
  g965
  (
    n1071,
    n136
  );


  buf
  g966
  (
    n775,
    n335
  );


  buf
  g967
  (
    n1359,
    n186
  );


  not
  g968
  (
    n783,
    n275
  );


  buf
  g969
  (
    n1147,
    n301
  );


  not
  g970
  (
    n1063,
    n332
  );


  not
  g971
  (
    n1273,
    n337
  );


  buf
  g972
  (
    n1013,
    n269
  );


  not
  g973
  (
    n1081,
    n241
  );


  buf
  g974
  (
    n702,
    n291
  );


  buf
  g975
  (
    n1217,
    n197
  );


  buf
  g976
  (
    n1137,
    n343
  );


  buf
  g977
  (
    n424,
    n253
  );


  not
  g978
  (
    n708,
    n174
  );


  not
  g979
  (
    n688,
    n284
  );


  buf
  g980
  (
    n1356,
    n217
  );


  not
  g981
  (
    n794,
    n147
  );


  buf
  g982
  (
    n1121,
    n122
  );


  buf
  g983
  (
    n1103,
    n259
  );


  not
  g984
  (
    n871,
    n144
  );


  buf
  g985
  (
    n413,
    n189
  );


  not
  g986
  (
    n821,
    n209
  );


  not
  g987
  (
    n942,
    n352
  );


  not
  g988
  (
    n682,
    n120
  );


  buf
  g989
  (
    n999,
    n263
  );


  buf
  g990
  (
    n1037,
    n313
  );


  not
  g991
  (
    n1093,
    n199
  );


  buf
  g992
  (
    n545,
    n215
  );


  buf
  g993
  (
    n365,
    n346
  );


  buf
  g994
  (
    n668,
    n307
  );


  buf
  g995
  (
    n360,
    n322
  );


  buf
  g996
  (
    n885,
    n174
  );


  not
  g997
  (
    n1192,
    n217
  );


  buf
  g998
  (
    n721,
    n199
  );


  buf
  g999
  (
    n1117,
    n275
  );


  buf
  g1000
  (
    n619,
    n134
  );


  not
  g1001
  (
    n597,
    n210
  );


  not
  g1002
  (
    n664,
    n223
  );


  not
  g1003
  (
    n476,
    n338
  );


  buf
  g1004
  (
    n568,
    n194
  );


  not
  g1005
  (
    n1239,
    n307
  );


  buf
  g1006
  (
    n475,
    n291
  );


  not
  g1007
  (
    n418,
    n240
  );


  buf
  g1008
  (
    n1249,
    n306
  );


  not
  g1009
  (
    n979,
    n318
  );


  buf
  g1010
  (
    n726,
    n318
  );


  not
  g1011
  (
    n751,
    n266
  );


  not
  g1012
  (
    n577,
    n178
  );


  buf
  g1013
  (
    n741,
    n86
  );


  not
  g1014
  (
    n1206,
    n276
  );


  not
  g1015
  (
    n1169,
    n184
  );


  not
  g1016
  (
    n371,
    n271
  );


  buf
  g1017
  (
    n520,
    n172
  );


  buf
  g1018
  (
    n1082,
    n127
  );


  buf
  g1019
  (
    n523,
    n290
  );


  not
  g1020
  (
    n943,
    n202
  );


  buf
  g1021
  (
    n844,
    n98
  );


  buf
  g1022
  (
    n1357,
    n302
  );


  buf
  g1023
  (
    n472,
    n234
  );


  buf
  g1024
  (
    n928,
    n352
  );


  buf
  g1025
  (
    n555,
    n128
  );


  buf
  g1026
  (
    n967,
    n326
  );


  not
  g1027
  (
    n1208,
    n305
  );


  buf
  g1028
  (
    n753,
    n306
  );


  buf
  g1029
  (
    n1130,
    n155
  );


  buf
  g1030
  (
    n1164,
    n313
  );


  not
  g1031
  (
    n651,
    n203
  );


  not
  g1032
  (
    n1205,
    n149
  );


  buf
  g1033
  (
    n562,
    n164
  );


  buf
  g1034
  (
    KeyWire_0_3,
    n218
  );


  not
  g1035
  (
    n1366,
    n352
  );


  not
  g1036
  (
    n1377,
    n206
  );


  buf
  g1037
  (
    n895,
    n247
  );


  not
  g1038
  (
    n1028,
    n246
  );


  not
  g1039
  (
    n766,
    n146
  );


  buf
  g1040
  (
    n816,
    n212
  );


  buf
  g1041
  (
    n511,
    n263
  );


  buf
  g1042
  (
    n946,
    n177
  );


  not
  g1043
  (
    n510,
    n95
  );


  buf
  g1044
  (
    n848,
    n296
  );


  not
  g1045
  (
    n1218,
    n232
  );


  buf
  g1046
  (
    n1030,
    n140
  );


  not
  g1047
  (
    n1060,
    n292
  );


  not
  g1048
  (
    n1196,
    n297
  );


  not
  g1049
  (
    n730,
    n124
  );


  not
  g1050
  (
    n785,
    n238
  );


  buf
  g1051
  (
    n683,
    n328
  );


  not
  g1052
  (
    KeyWire_0_12,
    n160
  );


  buf
  g1053
  (
    n1222,
    n247
  );


  not
  g1054
  (
    n443,
    n243
  );


  not
  g1055
  (
    n1149,
    n100
  );


  buf
  g1056
  (
    n915,
    n314
  );


  buf
  g1057
  (
    n1266,
    n108
  );


  buf
  g1058
  (
    n653,
    n286
  );


  buf
  g1059
  (
    n1215,
    n186
  );


  buf
  g1060
  (
    n543,
    n140
  );


  buf
  g1061
  (
    n483,
    n111
  );


  not
  g1062
  (
    n747,
    n99
  );


  buf
  g1063
  (
    n428,
    n106
  );


  not
  g1064
  (
    n1090,
    n286
  );


  not
  g1065
  (
    n496,
    n184
  );


  not
  g1066
  (
    n366,
    n341
  );


  not
  g1067
  (
    n1354,
    n218
  );


  buf
  g1068
  (
    n469,
    n227
  );


  buf
  g1069
  (
    n1165,
    n92
  );


  not
  g1070
  (
    n845,
    n331
  );


  buf
  g1071
  (
    n1235,
    n196
  );


  not
  g1072
  (
    n440,
    n140
  );


  not
  g1073
  (
    n512,
    n333
  );


  buf
  g1074
  (
    n1321,
    n241
  );


  not
  g1075
  (
    n1316,
    n286
  );


  not
  g1076
  (
    n358,
    n343
  );


  buf
  g1077
  (
    n852,
    n265
  );


  not
  g1078
  (
    n1301,
    n103
  );


  buf
  g1079
  (
    n976,
    n245
  );


  buf
  g1080
  (
    n1276,
    n134
  );


  not
  g1081
  (
    n750,
    n233
  );


  not
  g1082
  (
    n1150,
    n326
  );


  not
  g1083
  (
    n790,
    n254
  );


  buf
  g1084
  (
    n550,
    n181
  );


  buf
  g1085
  (
    n724,
    n267
  );


  buf
  g1086
  (
    n622,
    n290
  );


  buf
  g1087
  (
    n1051,
    n300
  );


  buf
  g1088
  (
    n1174,
    n222
  );


  not
  g1089
  (
    n383,
    n281
  );


  buf
  g1090
  (
    n495,
    n153
  );


  not
  g1091
  (
    n744,
    n309
  );


  buf
  g1092
  (
    n1350,
    n294
  );


  buf
  g1093
  (
    n795,
    n257
  );


  not
  g1094
  (
    n756,
    n325
  );


  not
  g1095
  (
    n1193,
    n108
  );


  not
  g1096
  (
    n772,
    n111
  );


  not
  g1097
  (
    n1045,
    n141
  );


  not
  g1098
  (
    n803,
    n138
  );


  not
  g1099
  (
    n737,
    n252
  );


  buf
  g1100
  (
    n866,
    n313
  );


  not
  g1101
  (
    n584,
    n207
  );


  not
  g1102
  (
    n784,
    n131
  );


  buf
  g1103
  (
    n1056,
    n129
  );


  buf
  g1104
  (
    n1307,
    n125
  );


  buf
  g1105
  (
    n1139,
    n321
  );


  not
  g1106
  (
    n1234,
    n353
  );


  not
  g1107
  (
    n876,
    n204
  );


  buf
  g1108
  (
    n1203,
    n249
  );


  not
  g1109
  (
    n1076,
    n235
  );


  buf
  g1110
  (
    n906,
    n295
  );


  not
  g1111
  (
    n452,
    n244
  );


  not
  g1112
  (
    n385,
    n193
  );


  not
  g1113
  (
    n517,
    n287
  );


  not
  g1114
  (
    n799,
    n163
  );


  buf
  g1115
  (
    n924,
    n91
  );


  not
  g1116
  (
    n433,
    n145
  );


  not
  g1117
  (
    n1331,
    n201
  );


  not
  g1118
  (
    n1238,
    n352
  );


  buf
  g1119
  (
    n1361,
    n235
  );


  not
  g1120
  (
    n1135,
    n345
  );


  not
  g1121
  (
    n727,
    n218
  );


  not
  g1122
  (
    n818,
    n208
  );


  buf
  g1123
  (
    n548,
    n147
  );


  not
  g1124
  (
    n1078,
    n206
  );


  buf
  g1125
  (
    n608,
    n264
  );


  not
  g1126
  (
    n1001,
    n224
  );


  buf
  g1127
  (
    n965,
    n210
  );


  not
  g1128
  (
    n431,
    n124
  );


  buf
  g1129
  (
    n798,
    n136
  );


  not
  g1130
  (
    n591,
    n251
  );


  buf
  g1131
  (
    n894,
    n168
  );


  not
  g1132
  (
    n399,
    n126
  );


  not
  g1133
  (
    n611,
    n312
  );


  buf
  g1134
  (
    n991,
    n272
  );


  not
  g1135
  (
    n390,
    n154
  );


  not
  g1136
  (
    n882,
    n304
  );


  buf
  g1137
  (
    n1245,
    n338
  );


  not
  g1138
  (
    n1303,
    n118
  );


  buf
  g1139
  (
    n771,
    n200
  );


  buf
  g1140
  (
    n722,
    n267
  );


  not
  g1141
  (
    n372,
    n105
  );


  not
  g1142
  (
    n1057,
    n135
  );


  buf
  g1143
  (
    n368,
    n97
  );


  buf
  g1144
  (
    n460,
    n137
  );


  buf
  g1145
  (
    n1317,
    n119
  );


  not
  g1146
  (
    n1322,
    n342
  );


  not
  g1147
  (
    n434,
    n348
  );


  not
  g1148
  (
    n626,
    n175
  );


  buf
  g1149
  (
    n498,
    n353
  );


  buf
  g1150
  (
    n698,
    n310
  );


  not
  g1151
  (
    n1075,
    n164
  );


  not
  g1152
  (
    n1323,
    n98
  );


  not
  g1153
  (
    n993,
    n153
  );


  not
  g1154
  (
    n1014,
    n299
  );


  buf
  g1155
  (
    n427,
    n150
  );


  buf
  g1156
  (
    n1289,
    n278
  );


  buf
  g1157
  (
    n955,
    n317
  );


  buf
  g1158
  (
    n1341,
    n211
  );


  not
  g1159
  (
    n875,
    n316
  );


  not
  g1160
  (
    n509,
    n165
  );


  not
  g1161
  (
    n559,
    n258
  );


  buf
  g1162
  (
    n672,
    n130
  );


  buf
  g1163
  (
    n1381,
    n315
  );


  buf
  g1164
  (
    n1282,
    n297
  );


  buf
  g1165
  (
    n858,
    n141
  );


  buf
  g1166
  (
    n1015,
    n166
  );


  not
  g1167
  (
    KeyWire_0_20,
    n206
  );


  not
  g1168
  (
    n1010,
    n337
  );


  buf
  g1169
  (
    n659,
    n179
  );


  not
  g1170
  (
    n1372,
    n107
  );


  buf
  g1171
  (
    n539,
    n176
  );


  buf
  g1172
  (
    n540,
    n188
  );


  not
  g1173
  (
    n916,
    n233
  );


  buf
  g1174
  (
    n868,
    n109
  );


  buf
  g1175
  (
    n487,
    n143
  );


  not
  g1176
  (
    n586,
    n324
  );


  buf
  g1177
  (
    n811,
    n269
  );


  buf
  g1178
  (
    n1052,
    n128
  );


  not
  g1179
  (
    n832,
    n126
  );


  not
  g1180
  (
    n887,
    n161
  );


  buf
  g1181
  (
    n992,
    n220
  );


  not
  g1182
  (
    n633,
    n143
  );


  buf
  g1183
  (
    n854,
    n307
  );


  not
  g1184
  (
    n1360,
    n192
  );


  not
  g1185
  (
    n806,
    n284
  );


  not
  g1186
  (
    n960,
    n126
  );


  buf
  g1187
  (
    n1339,
    n179
  );


  not
  g1188
  (
    n922,
    n208
  );


  not
  g1189
  (
    n786,
    n121
  );


  not
  g1190
  (
    n1020,
    n130
  );


  buf
  g1191
  (
    n1340,
    n258
  );


  not
  g1192
  (
    n831,
    n308
  );


  not
  g1193
  (
    n908,
    n219
  );


  buf
  g1194
  (
    n492,
    n347
  );


  buf
  g1195
  (
    n1226,
    n323
  );


  buf
  g1196
  (
    n796,
    n205
  );


  not
  g1197
  (
    n1069,
    n169
  );


  not
  g1198
  (
    n779,
    n252
  );


  buf
  g1199
  (
    n774,
    n336
  );


  buf
  g1200
  (
    n669,
    n162
  );


  not
  g1201
  (
    n1384,
    n228
  );


  buf
  g1202
  (
    KeyWire_0_16,
    n154
  );


  buf
  g1203
  (
    n838,
    n220
  );


  not
  g1204
  (
    n439,
    n166
  );


  not
  g1205
  (
    n819,
    n268
  );


  buf
  g1206
  (
    n642,
    n317
  );


  buf
  g1207
  (
    n1386,
    n178
  );


  buf
  g1208
  (
    n536,
    n114
  );


  buf
  g1209
  (
    n905,
    n322
  );


  buf
  g1210
  (
    n640,
    n130
  );


  buf
  g1211
  (
    n1216,
    n349
  );


  not
  g1212
  (
    n1031,
    n100
  );


  not
  g1213
  (
    n884,
    n338
  );


  buf
  g1214
  (
    n681,
    n148
  );


  not
  g1215
  (
    n1244,
    n283
  );


  buf
  g1216
  (
    n1214,
    n132
  );


  not
  g1217
  (
    n416,
    n337
  );


  buf
  g1218
  (
    n1054,
    n254
  );


  buf
  g1219
  (
    n1211,
    n134
  );


  not
  g1220
  (
    n1300,
    n326
  );


  not
  g1221
  (
    n833,
    n268
  );


  not
  g1222
  (
    n565,
    n334
  );


  not
  g1223
  (
    n917,
    n236
  );


  not
  g1224
  (
    n686,
    n88
  );


  not
  g1225
  (
    n1154,
    n107
  );


  buf
  g1226
  (
    n650,
    n298
  );


  not
  g1227
  (
    n1024,
    n283
  );


  not
  g1228
  (
    n435,
    n183
  );


  buf
  g1229
  (
    n1280,
    n113
  );


  buf
  g1230
  (
    n735,
    n335
  );


  not
  g1231
  (
    n1151,
    n341
  );


  not
  g1232
  (
    n453,
    n333
  );


  buf
  g1233
  (
    n1095,
    n192
  );


  not
  g1234
  (
    n862,
    n239
  );


  buf
  g1235
  (
    n501,
    n148
  );


  buf
  g1236
  (
    n504,
    n172
  );


  not
  g1237
  (
    n1335,
    n250
  );


  buf
  g1238
  (
    n1000,
    n101
  );


  buf
  g1239
  (
    n689,
    n118
  );


  buf
  g1240
  (
    n1144,
    n149
  );


  not
  g1241
  (
    n574,
    n205
  );


  buf
  g1242
  (
    n1026,
    n93
  );


  buf
  g1243
  (
    n824,
    n98
  );


  buf
  g1244
  (
    n1202,
    n328
  );


  not
  g1245
  (
    n1293,
    n147
  );


  not
  g1246
  (
    n910,
    n92
  );


  buf
  g1247
  (
    n621,
    n202
  );


  not
  g1248
  (
    KeyWire_0_10,
    n254
  );


  buf
  g1249
  (
    n948,
    n203
  );


  not
  g1250
  (
    n996,
    n347
  );


  not
  g1251
  (
    n1125,
    n183
  );


  buf
  g1252
  (
    n1281,
    n131
  );


  not
  g1253
  (
    n929,
    n171
  );


  buf
  g1254
  (
    n359,
    n351
  );


  not
  g1255
  (
    n742,
    n285
  );


  buf
  g1256
  (
    n1352,
    n225
  );


  buf
  g1257
  (
    n725,
    n169
  );


  not
  g1258
  (
    n1338,
    n226
  );


  not
  g1259
  (
    n1383,
    n279
  );


  not
  g1260
  (
    n1182,
    n123
  );


  not
  g1261
  (
    n1221,
    n334
  );


  not
  g1262
  (
    n1285,
    n295
  );


  buf
  g1263
  (
    n1004,
    n205
  );


  not
  g1264
  (
    n1161,
    n160
  );


  not
  g1265
  (
    n707,
    n157
  );


  not
  g1266
  (
    n1342,
    n198
  );


  buf
  g1267
  (
    n717,
    n99
  );


  not
  g1268
  (
    n361,
    n320
  );


  buf
  g1269
  (
    n530,
    n185
  );


  buf
  g1270
  (
    n1290,
    n325
  );


  not
  g1271
  (
    n549,
    n260
  );


  buf
  g1272
  (
    n630,
    n289
  );


  buf
  g1273
  (
    n1006,
    n281
  );


  buf
  g1274
  (
    n1254,
    n108
  );


  not
  g1275
  (
    n1134,
    n200
  );


  not
  g1276
  (
    n842,
    n188
  );


  not
  g1277
  (
    n1271,
    n187
  );


  buf
  g1278
  (
    n1373,
    n340
  );


  not
  g1279
  (
    n834,
    n195
  );


  buf
  g1280
  (
    n648,
    n87
  );


  not
  g1281
  (
    n962,
    n235
  );


  not
  g1282
  (
    n373,
    n186
  );


  not
  g1283
  (
    n410,
    n316
  );


  buf
  g1284
  (
    n531,
    n136
  );


  buf
  g1285
  (
    n379,
    n114
  );


  not
  g1286
  (
    n1181,
    n285
  );


  buf
  g1287
  (
    n1186,
    n196
  );


  not
  g1288
  (
    KeyWire_0_0,
    n351
  );


  not
  g1289
  (
    n1019,
    n102
  );


  not
  g1290
  (
    n1110,
    n133
  );


  not
  g1291
  (
    n660,
    n239
  );


  buf
  g1292
  (
    n951,
    n133
  );


  buf
  g1293
  (
    n596,
    n317
  );


  not
  g1294
  (
    n704,
    n293
  );


  buf
  g1295
  (
    n1040,
    n156
  );


  buf
  g1296
  (
    KeyWire_0_25,
    n236
  );


  buf
  g1297
  (
    n1168,
    n287
  );


  buf
  g1298
  (
    n676,
    n137
  );


  not
  g1299
  (
    n1353,
    n255
  );


  not
  g1300
  (
    n412,
    n234
  );


  not
  g1301
  (
    n1123,
    n119
  );


  buf
  g1302
  (
    n863,
    n326
  );


  buf
  g1303
  (
    n1112,
    n300
  );


  not
  g1304
  (
    n1324,
    n226
  );


  buf
  g1305
  (
    n506,
    n282
  );


  not
  g1306
  (
    n1311,
    n109
  );


  buf
  g1307
  (
    n1379,
    n323
  );


  not
  g1308
  (
    n797,
    n332
  );


  buf
  g1309
  (
    n693,
    n210
  );


  not
  g1310
  (
    n600,
    n101
  );


  buf
  g1311
  (
    n849,
    n270
  );


  buf
  g1312
  (
    n538,
    n282
  );


  buf
  g1313
  (
    n1053,
    n157
  );


  buf
  g1314
  (
    n384,
    n242
  );


  buf
  g1315
  (
    n1302,
    n121
  );


  not
  g1316
  (
    n401,
    n92
  );


  not
  g1317
  (
    n1012,
    n160
  );


  buf
  g1318
  (
    n823,
    n244
  );


  buf
  g1319
  (
    n441,
    n143
  );


  not
  g1320
  (
    n1296,
    n231
  );


  buf
  g1321
  (
    n1055,
    n193
  );


  buf
  g1322
  (
    n1088,
    n244
  );


  not
  g1323
  (
    n923,
    n310
  );


  not
  g1324
  (
    n939,
    n211
  );


  not
  g1325
  (
    n855,
    n123
  );


  not
  g1326
  (
    n590,
    n340
  );


  not
  g1327
  (
    n613,
    n256
  );


  not
  g1328
  (
    n846,
    n121
  );


  not
  g1329
  (
    n1349,
    n190
  );


  buf
  g1330
  (
    n1074,
    n165
  );


  not
  g1331
  (
    n1177,
    n104
  );


  buf
  g1332
  (
    n1122,
    n243
  );


  buf
  g1333
  (
    n1267,
    n254
  );


  not
  g1334
  (
    n847,
    n159
  );


  buf
  g1335
  (
    n389,
    n229
  );


  buf
  g1336
  (
    n638,
    n238
  );


  buf
  g1337
  (
    n561,
    n265
  );


  not
  g1338
  (
    n1274,
    n112
  );


  buf
  g1339
  (
    n1223,
    n130
  );


  not
  g1340
  (
    n1083,
    n146
  );


  not
  g1341
  (
    n865,
    n197
  );


  buf
  g1342
  (
    n1138,
    n331
  );


  not
  g1343
  (
    n1011,
    n228
  );


  buf
  g1344
  (
    n1345,
    n242
  );


  not
  g1345
  (
    n1086,
    n329
  );


  buf
  g1346
  (
    n777,
    n127
  );


  not
  g1347
  (
    n1022,
    n311
  );


  not
  g1348
  (
    n1194,
    n304
  );


  buf
  g1349
  (
    n554,
    n201
  );


  not
  g1350
  (
    n527,
    n208
  );


  not
  g1351
  (
    n1347,
    n233
  );


  not
  g1352
  (
    n557,
    n97
  );


  buf
  g1353
  (
    n1104,
    n232
  );


  or
  g1354
  (
    n661,
    n199,
    n219
  );


  xnor
  g1355
  (
    n1200,
    n100,
    n96
  );


  or
  g1356
  (
    n974,
    n195,
    n183,
    n171
  );


  or
  g1357
  (
    n754,
    n185,
    n259,
    n251,
    n319
  );


  nor
  g1358
  (
    n1126,
    n340,
    n292,
    n243,
    n112
  );


  xor
  g1359
  (
    n1318,
    n354,
    n200,
    n91,
    n305
  );


  xnor
  g1360
  (
    n677,
    n115,
    n207,
    n179,
    n316
  );


  xor
  g1361
  (
    n374,
    n237,
    n351,
    n165,
    n252
  );


  nand
  g1362
  (
    n459,
    n343,
    n205,
    n331,
    n227
  );


  or
  g1363
  (
    n1261,
    n249,
    n256,
    n196
  );


  nand
  g1364
  (
    n1191,
    n120,
    n273,
    n287,
    n349
  );


  and
  g1365
  (
    n388,
    n297,
    n276,
    n95,
    n248
  );


  xor
  g1366
  (
    n394,
    n334,
    n209,
    n127,
    n215
  );


  or
  g1367
  (
    n449,
    n117,
    n260,
    n323,
    n271
  );


  nand
  g1368
  (
    n761,
    n335,
    n180,
    n175,
    n122
  );


  xor
  g1369
  (
    n1034,
    n88,
    n190,
    n131,
    n231
  );


  nor
  g1370
  (
    n1785,
    n830,
    n463,
    n454,
    n1042
  );


  nor
  g1371
  (
    n1704,
    n1306,
    n1333,
    n1161,
    n1271
  );


  xnor
  g1372
  (
    n1415,
    n1147,
    n1004,
    n1242,
    n1160
  );


  nand
  g1373
  (
    n1769,
    n1048,
    n598,
    n1231,
    n478
  );


  nor
  g1374
  (
    n1527,
    n1121,
    n1138,
    n1257
  );


  or
  g1375
  (
    n1768,
    n1111,
    n1127,
    n1233,
    n1309
  );


  or
  g1376
  (
    n1419,
    n604,
    n1196,
    n1101,
    n382
  );


  nor
  g1377
  (
    n1787,
    n1281,
    n1245,
    n1254,
    n971
  );


  nor
  g1378
  (
    n1761,
    n716,
    n1244,
    n1177,
    n1000
  );


  nand
  g1379
  (
    n1518,
    n1218,
    n1357,
    n1301,
    n1137
  );


  nor
  g1380
  (
    n1472,
    n641,
    n678,
    n1087,
    n1167
  );


  xor
  g1381
  (
    n1606,
    n1289,
    n1349,
    n1279,
    n1214
  );


  and
  g1382
  (
    n1800,
    n991,
    n1327,
    n1141,
    n812
  );


  xnor
  g1383
  (
    n1391,
    n596,
    n570,
    n1263,
    n379
  );


  xor
  g1384
  (
    n1741,
    n736,
    n1331,
    n1110,
    n1127
  );


  or
  g1385
  (
    n1426,
    n1126,
    n402,
    n939,
    n1249
  );


  nor
  g1386
  (
    n1566,
    n1314,
    n1284,
    n509,
    n1274
  );


  nand
  g1387
  (
    n1425,
    n913,
    n1292,
    n955,
    n1190
  );


  nand
  g1388
  (
    n1546,
    n1260,
    n1216,
    n1056,
    n1324
  );


  nor
  g1389
  (
    n1807,
    n1132,
    n1144,
    n1161,
    n1156
  );


  or
  g1390
  (
    n1418,
    n1162,
    n643,
    n1142,
    n1159
  );


  nor
  g1391
  (
    n1681,
    n1361,
    n1312,
    n1160,
    n1300
  );


  nor
  g1392
  (
    n1691,
    n629,
    n749,
    n865,
    n1305
  );


  nand
  g1393
  (
    n1408,
    n615,
    n1258,
    n1367,
    n1097
  );


  xor
  g1394
  (
    n1745,
    n1205,
    n1365,
    n1222,
    n593
  );


  or
  g1395
  (
    n1485,
    n1346,
    n961,
    n1143,
    n1099
  );


  nand
  g1396
  (
    n1455,
    n1354,
    n794,
    n1260,
    n1228
  );


  nor
  g1397
  (
    n1570,
    n920,
    n1188,
    n1285,
    n1168
  );


  or
  g1398
  (
    n1707,
    n1371,
    n1084,
    n1061,
    n1002
  );


  or
  g1399
  (
    n1664,
    n979,
    n1236,
    n1100,
    n1182
  );


  nand
  g1400
  (
    n1801,
    n690,
    n1314,
    n669,
    n782
  );


  and
  g1401
  (
    n1489,
    n633,
    n1106,
    n1316,
    n1332
  );


  or
  g1402
  (
    n1841,
    n1285,
    n1179,
    n765,
    n1154
  );


  xor
  g1403
  (
    n1411,
    n413,
    n1150,
    n1312,
    n1026
  );


  and
  g1404
  (
    n1648,
    n510,
    n572,
    n1243,
    n1255
  );


  xor
  g1405
  (
    n1647,
    n684,
    n1118,
    n504,
    n1337
  );


  or
  g1406
  (
    n1536,
    n1280,
    n1269,
    n619,
    n1317
  );


  or
  g1407
  (
    n1850,
    n653,
    n1222,
    n1169,
    n1213
  );


  xor
  g1408
  (
    n1557,
    n655,
    n996,
    n1188,
    n637
  );


  nand
  g1409
  (
    n1584,
    n1178,
    n1168,
    n1057,
    n1109
  );


  nor
  g1410
  (
    n1397,
    n1104,
    n431,
    n983,
    n1114
  );


  or
  g1411
  (
    n1817,
    n1160,
    n1199,
    n1241,
    n1251
  );


  xnor
  g1412
  (
    n1693,
    n1174,
    n1272,
    n826,
    n369
  );


  and
  g1413
  (
    n1456,
    n1068,
    n1368,
    n704,
    n1242
  );


  nor
  g1414
  (
    n1609,
    n1011,
    n1230,
    n1143,
    n1309
  );


  and
  g1415
  (
    n1798,
    n1136,
    n1216,
    n446,
    n1278
  );


  xnor
  g1416
  (
    n1400,
    n1172,
    n825,
    n417,
    n1347
  );


  or
  g1417
  (
    n1506,
    n998,
    n621,
    n1006,
    n1268
  );


  or
  g1418
  (
    n1396,
    n770,
    n1281,
    n1153,
    n1157
  );


  xor
  g1419
  (
    n1533,
    n1142,
    n470,
    n943,
    n1261
  );


  nand
  g1420
  (
    n1713,
    n1290,
    n456,
    n1102,
    n1137
  );


  nand
  g1421
  (
    n1569,
    n662,
    n657,
    n1210,
    n1261
  );


  nor
  g1422
  (
    n1795,
    n671,
    n1284,
    n1174,
    n1256
  );


  or
  g1423
  (
    n1619,
    n1095,
    n423,
    n1215,
    n1268
  );


  nor
  g1424
  (
    n1718,
    n459,
    n1093,
    n477,
    n1280
  );


  xor
  g1425
  (
    n1446,
    n1160,
    n1221,
    n1296,
    n1237
  );


  nand
  g1426
  (
    n1847,
    n952,
    n1105,
    n1175,
    n1349
  );


  and
  g1427
  (
    n1441,
    n1253,
    n776,
    n1290,
    n1353
  );


  xor
  g1428
  (
    n1572,
    n389,
    n828,
    n1198,
    n1152
  );


  and
  g1429
  (
    n1661,
    n1352,
    n519,
    n683,
    n914
  );


  nand
  g1430
  (
    KeyWire_0_17,
    n1158,
    n790,
    n1369,
    n910
  );


  or
  g1431
  (
    n1791,
    n1305,
    n808,
    n1263,
    n839
  );


  xnor
  g1432
  (
    n1702,
    n1177,
    n527,
    n857,
    n1352
  );


  xnor
  g1433
  (
    n1594,
    n1156,
    n1287,
    n1232,
    n987
  );


  nand
  g1434
  (
    n1593,
    n1200,
    n1134,
    n523,
    n969
  );


  and
  g1435
  (
    n1595,
    n701,
    n1369,
    n638,
    n626
  );


  or
  g1436
  (
    n1486,
    n1259,
    n855,
    n1336,
    n660
  );


  or
  g1437
  (
    n1488,
    n1246,
    n995,
    n766,
    n1279
  );


  and
  g1438
  (
    n1494,
    n1316,
    n823,
    n1335,
    n928
  );


  nor
  g1439
  (
    n1442,
    n1019,
    n1202,
    n1112,
    n1322
  );


  or
  g1440
  (
    n1708,
    n691,
    n1271,
    n618,
    n1291
  );


  nor
  g1441
  (
    n1508,
    n816,
    n805,
    n1197
  );


  and
  g1442
  (
    n1631,
    n760,
    n1153,
    n1330,
    n1193
  );


  and
  g1443
  (
    n1434,
    n911,
    n1164,
    n1176,
    n1202
  );


  nand
  g1444
  (
    n1514,
    n586,
    n1105,
    n1170,
    n727
  );


  or
  g1445
  (
    n1535,
    n868,
    n795,
    n726,
    n1230
  );


  nor
  g1446
  (
    n1436,
    n1370,
    n613,
    n1311,
    n1245
  );


  or
  g1447
  (
    n1476,
    n1104,
    n1351,
    n1349,
    n1237
  );


  xnor
  g1448
  (
    n1530,
    n1293,
    n1367,
    n600,
    n1355
  );


  nor
  g1449
  (
    n1592,
    n1322,
    n1267,
    n1093,
    n550
  );


  xnor
  g1450
  (
    n1459,
    n1041,
    n1211,
    n829,
    n1159
  );


  nand
  g1451
  (
    n1428,
    n849,
    n1345,
    n1059,
    n1154
  );


  nand
  g1452
  (
    n1410,
    n1205,
    n1207,
    n1256,
    n755
  );


  nand
  g1453
  (
    n1522,
    n611,
    n1353,
    n1173,
    n1228
  );


  nand
  g1454
  (
    n1440,
    n898,
    n1329,
    n1193,
    n1111
  );


  or
  g1455
  (
    n1790,
    n1370,
    n1334,
    n1188,
    n1283
  );


  nor
  g1456
  (
    n1427,
    n644,
    n564,
    n1266,
    n1073
  );


  xor
  g1457
  (
    n1484,
    n1186,
    n1348,
    n405,
    n1133
  );


  xnor
  g1458
  (
    n1607,
    n1051,
    n918,
    n894,
    n1171
  );


  xnor
  g1459
  (
    n1849,
    n1234,
    n1326,
    n1173,
    n1043
  );


  nand
  g1460
  (
    n1816,
    n1120,
    n867,
    n632,
    n1234
  );


  xor
  g1461
  (
    n1483,
    n566,
    n1323,
    n1218,
    n1304
  );


  xor
  g1462
  (
    n1412,
    n1131,
    n1138,
    n836,
    n674
  );


  nor
  g1463
  (
    n1452,
    n1235,
    n440,
    n709,
    n1150
  );


  nand
  g1464
  (
    n1602,
    n1128,
    n773,
    n958,
    n1172
  );


  xor
  g1465
  (
    n1828,
    n842,
    n1251,
    n436,
    n1180
  );


  nor
  g1466
  (
    n1635,
    n1247,
    n1243,
    n1211,
    n869
  );


  nand
  g1467
  (
    n1523,
    n1171,
    n1220,
    n1209,
    n1294
  );


  nand
  g1468
  (
    n1820,
    n1262,
    n468,
    n1104,
    n1148
  );


  xor
  g1469
  (
    n1669,
    n1369,
    n1202,
    n1204,
    n801
  );


  or
  g1470
  (
    n1689,
    n1157,
    n1358,
    n473,
    n1366
  );


  or
  g1471
  (
    n1844,
    n1158,
    n1174,
    n479,
    n515
  );


  xnor
  g1472
  (
    n1394,
    n1231,
    n1269,
    n1116,
    n1227
  );


  xnor
  g1473
  (
    n1480,
    n799,
    n410,
    n1132,
    n843
  );


  nor
  g1474
  (
    n1474,
    n1125,
    n1122,
    n1267,
    n851
  );


  or
  g1475
  (
    n1389,
    n1338,
    n1300,
    n1350,
    n1323
  );


  or
  g1476
  (
    n1388,
    n605,
    n1024,
    n597,
    n847
  );


  and
  g1477
  (
    n1525,
    n1050,
    n1283,
    n1149,
    n1366
  );


  nand
  g1478
  (
    n1782,
    n827,
    n1247,
    n1282,
    n1230
  );


  xnor
  g1479
  (
    n1615,
    n452,
    n1212,
    n1085,
    n1192
  );


  nand
  g1480
  (
    n1622,
    n383,
    n1308,
    n1244,
    n1258
  );


  xnor
  g1481
  (
    n1836,
    n1148,
    n798,
    n1241,
    n1347
  );


  xnor
  g1482
  (
    n1640,
    n1320,
    n437,
    n1103,
    n1219
  );


  nand
  g1483
  (
    n1773,
    n886,
    n927,
    n1232,
    n1327
  );


  nor
  g1484
  (
    n1601,
    n616,
    n1137,
    n984,
    n548
  );


  xnor
  g1485
  (
    n1751,
    n506,
    n524,
    n1337,
    n871
  );


  and
  g1486
  (
    n1392,
    n1266,
    n1296,
    n663,
    n1167
  );


  nand
  g1487
  (
    n1432,
    n1302,
    n480,
    n1158,
    n1094
  );


  nand
  g1488
  (
    n1654,
    n1246,
    n752,
    n994,
    n1032
  );


  xnor
  g1489
  (
    n1788,
    n1157,
    n743,
    n861,
    n1189
  );


  and
  g1490
  (
    n1403,
    n1328,
    n1189,
    n434,
    n1003
  );


  and
  g1491
  (
    n1822,
    n1343,
    n1287,
    n1362,
    n1270
  );


  nor
  g1492
  (
    n1470,
    n625,
    n485,
    n1259,
    n1258
  );


  xor
  g1493
  (
    n1805,
    n673,
    n821,
    n1233,
    n1321
  );


  nor
  g1494
  (
    n1517,
    n1197,
    n936,
    n1125,
    n730
  );


  and
  g1495
  (
    n1839,
    n1304,
    n1209,
    n1262,
    n528
  );


  xnor
  g1496
  (
    n1487,
    n1331,
    n1234,
    n1187,
    n1238
  );


  xor
  g1497
  (
    n1842,
    n1363,
    n1194,
    n1185,
    n1193
  );


  xor
  g1498
  (
    n1687,
    n1250,
    n1239,
    n1190,
    n1280
  );


  nand
  g1499
  (
    n1652,
    n1276,
    n1265,
    n972,
    n1175
  );


  xnor
  g1500
  (
    n1600,
    n870,
    n451,
    n785,
    n1318
  );


  nand
  g1501
  (
    n1598,
    n1120,
    n1105,
    n1200,
    n1214
  );


  or
  g1502
  (
    n1660,
    n1092,
    n1367,
    n1028,
    n1299
  );


  xor
  g1503
  (
    n1580,
    n1214,
    n556,
    n962,
    n555
  );


  or
  g1504
  (
    n1553,
    n1314,
    n1253,
    n1169,
    n1320
  );


  or
  g1505
  (
    n1815,
    n890,
    n1305,
    n1220,
    n1252
  );


  nor
  g1506
  (
    n1477,
    n1305,
    n450,
    n1236,
    n1156
  );


  and
  g1507
  (
    n1478,
    n1007,
    n1268,
    n1111,
    n1303
  );


  nor
  g1508
  (
    n1812,
    n1206,
    n1203,
    n1108,
    n1182
  );


  nor
  g1509
  (
    n1447,
    n1094,
    n1161,
    n1127,
    n1200
  );


  nor
  g1510
  (
    n1762,
    n989,
    n1370,
    n1103,
    n941
  );


  xor
  g1511
  (
    n1473,
    n393,
    n1198,
    n896,
    n1269
  );


  or
  g1512
  (
    n1588,
    n803,
    n1212,
    n1296,
    n1307
  );


  xor
  g1513
  (
    n1571,
    n1288,
    n1335,
    n1297,
    n975
  );


  xnor
  g1514
  (
    n1683,
    n1313,
    n416,
    n1117,
    n582
  );


  xnor
  g1515
  (
    n1405,
    n1113,
    n1241,
    n1311,
    n1152
  );


  xnor
  g1516
  (
    n1678,
    n1325,
    n837,
    n676,
    n668
  );


  and
  g1517
  (
    n1774,
    n374,
    n664,
    n1070,
    n491
  );


  nand
  g1518
  (
    n1611,
    n365,
    n1325,
    n1372,
    n1110
  );


  nor
  g1519
  (
    n1797,
    n1149,
    n1180,
    n1364,
    n1217
  );


  nand
  g1520
  (
    n1561,
    n1162,
    n1139,
    n1306,
    n1164
  );


  or
  g1521
  (
    n1448,
    n780,
    n1135,
    n1098,
    n1318
  );


  xor
  g1522
  (
    n1747,
    n1115,
    n1246,
    n1306,
    n1334
  );


  nand
  g1523
  (
    n1539,
    n1307,
    n1308,
    n841,
    n963
  );


  nand
  g1524
  (
    n1736,
    n1117,
    n1129,
    n1060,
    n1360
  );


  nand
  g1525
  (
    n1417,
    n1278,
    n1152,
    n1171,
    n1254
  );


  nand
  g1526
  (
    n1821,
    n507,
    n1112,
    n1210,
    n713
  );


  xnor
  g1527
  (
    n1433,
    n1152,
    n1195,
    n1090,
    n731
  );


  xor
  g1528
  (
    n1735,
    n769,
    n1126,
    n620,
    n697
  );


  and
  g1529
  (
    n1587,
    n1173,
    n522,
    n1274,
    n568
  );


  and
  g1530
  (
    n1776,
    n1332,
    n1205,
    n1243,
    n448
  );


  or
  g1531
  (
    n1639,
    n599,
    n442,
    n1075,
    n443
  );


  nand
  g1532
  (
    n1714,
    n1328,
    n756,
    n1221,
    n739
  );


  and
  g1533
  (
    n1690,
    n917,
    n1367,
    n1225,
    n1078
  );


  xnor
  g1534
  (
    n1748,
    n1183,
    n1360,
    n1315,
    n1119
  );


  or
  g1535
  (
    n1453,
    n916,
    n1355,
    n1132,
    n732
  );


  xor
  g1536
  (
    n1668,
    n679,
    n1142,
    n594,
    n601
  );


  and
  g1537
  (
    n1726,
    n1312,
    n1263,
    n1220,
    n1302
  );


  or
  g1538
  (
    n1458,
    n786,
    n409,
    n1344,
    n1203
  );


  and
  g1539
  (
    n1672,
    n647,
    n1179,
    n1275,
    n1103
  );


  xor
  g1540
  (
    n1491,
    n1156,
    n466,
    n1341,
    n724
  );


  nand
  g1541
  (
    n1722,
    n401,
    n761,
    n1102
  );


  nand
  g1542
  (
    n1764,
    n1297,
    n1338,
    n1301,
    n852
  );


  nor
  g1543
  (
    n1500,
    n1158,
    n1355,
    n1195,
    n419
  );


  nor
  g1544
  (
    n1610,
    n1221,
    n721,
    n1178,
    n1292
  );


  nor
  g1545
  (
    n1555,
    n542,
    n1236,
    n1337,
    n1302
  );


  or
  g1546
  (
    n1715,
    n976,
    n1319,
    n862,
    n1166
  );


  and
  g1547
  (
    n1549,
    n642,
    n1150,
    n584,
    n1183
  );


  nor
  g1548
  (
    n1402,
    n492,
    n1145,
    n859,
    n1244
  );


  nor
  g1549
  (
    n1576,
    n1229,
    n447,
    n1227,
    n521
  );


  xnor
  g1550
  (
    n1560,
    n547,
    n1322,
    n1315,
    n1141
  );


  nand
  g1551
  (
    n1445,
    n1308,
    n1249,
    n461,
    n1142
  );


  and
  g1552
  (
    n1780,
    n1199,
    n587,
    n878,
    n1125
  );


  xor
  g1553
  (
    n1772,
    n892,
    n1226,
    n789,
    n408
  );


  nor
  g1554
  (
    n1501,
    n1248,
    n552,
    n1301,
    n1184
  );


  nand
  g1555
  (
    n1651,
    n1351,
    n421,
    n1206,
    n418
  );


  nand
  g1556
  (
    n1573,
    n677,
    n1238,
    n490,
    n1088
  );


  or
  g1557
  (
    n1667,
    n986,
    n1109,
    n1134,
    n1096
  );


  xnor
  g1558
  (
    n1686,
    n973,
    n1124,
    n1128,
    n1222
  );


  xor
  g1559
  (
    n1632,
    n813,
    n1368,
    n1309,
    n1344
  );


  xnor
  g1560
  (
    n1665,
    n465,
    n503,
    n1226,
    n484
  );


  xor
  g1561
  (
    n1694,
    n1364,
    n1297,
    n1161,
    n1168
  );


  nor
  g1562
  (
    n1490,
    n453,
    n648,
    n525,
    n1067
  );


  and
  g1563
  (
    n1728,
    n1179,
    n1364,
    n494,
    n698
  );


  nor
  g1564
  (
    n1393,
    n1039,
    n1309,
    n1242,
    n1286
  );


  xor
  g1565
  (
    n1684,
    n809,
    n1239,
    n1114,
    n1098
  );


  or
  g1566
  (
    n1520,
    n1224,
    n905,
    n767,
    n646
  );


  and
  g1567
  (
    n1729,
    n1228,
    n1181,
    n1092,
    n1201
  );


  xor
  g1568
  (
    n1625,
    n1294,
    n1229,
    n1218,
    n1125
  );


  nor
  g1569
  (
    n1438,
    n1102,
    n493,
    n1344,
    n1271
  );


  and
  g1570
  (
    n1407,
    n1183,
    n802,
    n1186,
    n1106
  );


  or
  g1571
  (
    n1783,
    n1173,
    n1143,
    n1251,
    n1127
  );


  or
  g1572
  (
    n1467,
    n1008,
    n1233,
    n1219,
    n427
  );


  and
  g1573
  (
    n1528,
    n1005,
    n1213,
    n1112,
    n1217
  );


  xnor
  g1574
  (
    n1753,
    n921,
    n1304,
    n687,
    n1298
  );


  xnor
  g1575
  (
    n1830,
    n778,
    n1244,
    n705,
    n772
  );


  xnor
  g1576
  (
    n1789,
    n1069,
    n415,
    n1272,
    n1350
  );


  nand
  g1577
  (
    n1422,
    n1212,
    n476,
    n1225,
    n1119
  );


  nor
  g1578
  (
    n1597,
    n1135,
    n1353,
    n1076,
    n1295
  );


  nor
  g1579
  (
    n1495,
    n460,
    n1312,
    n627,
    n1340
  );


  nand
  g1580
  (
    n1786,
    n1054,
    n1198,
    n993,
    n583
  );


  nand
  g1581
  (
    n1818,
    n531,
    n1100,
    n1188,
    n1140
  );


  xnor
  g1582
  (
    n1511,
    n1313,
    n1047,
    n1273,
    n831
  );


  nand
  g1583
  (
    n1703,
    n1270,
    n1218,
    n1083,
    n1332
  );


  nor
  g1584
  (
    n1604,
    n1282,
    n1183,
    n551,
    n1185
  );


  xor
  g1585
  (
    n1605,
    n1126,
    n400,
    n422,
    n1129
  );


  xor
  g1586
  (
    n1471,
    n1133,
    n719,
    n1175,
    n696
  );


  nor
  g1587
  (
    n1519,
    n1252,
    n1233,
    n1146,
    n536
  );


  or
  g1588
  (
    n1548,
    n1217,
    n482,
    n1191,
    n901
  );


  xor
  g1589
  (
    n1540,
    n912,
    n1340,
    n608,
    n1122
  );


  xnor
  g1590
  (
    n1621,
    n609,
    n1287,
    n675,
    n738
  );


  nand
  g1591
  (
    n1613,
    n1162,
    n1261,
    n1205,
    n884
  );


  nor
  g1592
  (
    n1618,
    n1284,
    n1144,
    n1324,
    n1281
  );


  nor
  g1593
  (
    n1435,
    n1315,
    n1181,
    n1108,
    n1139
  );


  nor
  g1594
  (
    n1824,
    n703,
    n1163,
    n1192
  );


  and
  g1595
  (
    KeyWire_0_2,
    n889,
    n863,
    n540,
    n1308
  );


  xor
  g1596
  (
    n1556,
    n768,
    n1189,
    n720,
    n1187
  );


  nor
  g1597
  (
    n1450,
    n840,
    n589,
    n1146,
    n529
  );


  nor
  g1598
  (
    n1814,
    n1339,
    n650,
    n1187,
    n737
  );


  xor
  g1599
  (
    n1544,
    n1276,
    n777,
    n665,
    n1136
  );


  xor
  g1600
  (
    n1716,
    n1220,
    n1157,
    n1365,
    n1195
  );


  and
  g1601
  (
    n1696,
    n1317,
    n1170,
    n1017,
    n1302
  );


  nand
  g1602
  (
    n1579,
    n581,
    n1273,
    n1341,
    n1371
  );


  xnor
  g1603
  (
    n1803,
    n439,
    n1239,
    n1261,
    n1342
  );


  or
  g1604
  (
    n1843,
    n791,
    n513,
    n1264,
    n591
  );


  or
  g1605
  (
    n1832,
    n1315,
    n1333,
    n464,
    n628
  );


  xor
  g1606
  (
    n1463,
    n1318,
    n1286,
    n980,
    n1319
  );


  nor
  g1607
  (
    n1583,
    n824,
    n1365,
    n1336,
    n1366
  );


  nand
  g1608
  (
    n1591,
    n1323,
    n414,
    n924,
    n1185
  );


  nand
  g1609
  (
    n1732,
    n797,
    n1371,
    n1213,
    n1225
  );


  xor
  g1610
  (
    n1608,
    n1362,
    n923,
    n1252,
    n1178
  );


  or
  g1611
  (
    KeyWire_0_23,
    n1352,
    n1116,
    n1149,
    n999
  );


  xor
  g1612
  (
    n1804,
    n373,
    n533,
    n1206,
    n695
  );


  and
  g1613
  (
    n1835,
    n1091,
    n1022,
    n949,
    n712
  );


  xnor
  g1614
  (
    n1503,
    n1294,
    n1191,
    n1186,
    n1257
  );


  nand
  g1615
  (
    n1629,
    n763,
    n1115,
    n935,
    n1210
  );


  or
  g1616
  (
    n1794,
    n1291,
    n543,
    n1362,
    n854
  );


  or
  g1617
  (
    n1578,
    n946,
    n680,
    n428,
    n1106
  );


  nand
  g1618
  (
    KeyWire_0_15,
    n856,
    n1318,
    n1281,
    n449
  );


  xor
  g1619
  (
    n1742,
    n1177,
    n1222,
    n688,
    n1348
  );


  and
  g1620
  (
    n1406,
    n1275,
    n1101,
    n558,
    n406
  );


  xor
  g1621
  (
    n1829,
    n1333,
    n876,
    n1020,
    n1361
  );


  xnor
  g1622
  (
    n1521,
    n1206,
    n378,
    n559,
    n1168
  );


  nand
  g1623
  (
    n1796,
    n1093,
    n388,
    n1166,
    n1169
  );


  or
  g1624
  (
    n1757,
    n990,
    n634,
    n718,
    n957
  );


  xor
  g1625
  (
    n1481,
    n1262,
    n959,
    n1123,
    n1229
  );


  xnor
  g1626
  (
    n1655,
    n472,
    n750,
    n1278,
    n1129
  );


  xor
  g1627
  (
    n1740,
    n1231,
    n1094,
    n942,
    n534
  );


  xnor
  g1628
  (
    n1420,
    n1356,
    n1106,
    n1316,
    n945
  );


  xor
  g1629
  (
    n1603,
    n1351,
    n1130,
    n1226,
    n774
  );


  or
  g1630
  (
    n1825,
    n1314,
    n1191,
    n1320,
    n1234
  );


  xnor
  g1631
  (
    n1493,
    n1001,
    n934,
    n1155,
    n1124
  );


  or
  g1632
  (
    n1529,
    n1215,
    n1099,
    n895,
    n997
  );


  nor
  g1633
  (
    n1451,
    n981,
    n636,
    n1166,
    n1288
  );


  nand
  g1634
  (
    n1567,
    n746,
    n885,
    n1235,
    n1295
  );


  nand
  g1635
  (
    n1705,
    n1065,
    n764,
    n1029,
    n1303
  );


  nor
  g1636
  (
    n1793,
    n834,
    n891,
    n985,
    n640
  );


  nor
  g1637
  (
    n1706,
    n1113,
    n1289,
    n1283,
    n977
  );


  xnor
  g1638
  (
    n1444,
    n1209,
    n457,
    n1353,
    n489
  );


  or
  g1639
  (
    n1653,
    n445,
    n1194,
    n1260,
    n1117
  );


  xor
  g1640
  (
    n1515,
    n670,
    n1164,
    n1232,
    n1223
  );


  xnor
  g1641
  (
    n1831,
    n811,
    n820,
    n904,
    n1189
  );


  xnor
  g1642
  (
    n1675,
    n1204,
    n1131,
    n875,
    n645
  );


  or
  g1643
  (
    n1777,
    n1187,
    n929,
    n517,
    n1349
  );


  and
  g1644
  (
    n1721,
    n1255,
    n1298,
    n1342,
    n1359
  );


  nand
  g1645
  (
    n1827,
    n1249,
    n744,
    n1162,
    n1165
  );


  or
  g1646
  (
    n1416,
    n588,
    n1049,
    n967,
    n872
  );


  nand
  g1647
  (
    n1554,
    n1092,
    n1277,
    n1093,
    n887
  );


  xnor
  g1648
  (
    n1577,
    n745,
    n1130,
    n1303,
    n396
  );


  and
  g1649
  (
    n1826,
    n1174,
    n725,
    n1326,
    n411
  );


  nor
  g1650
  (
    n1811,
    n1240,
    n1124,
    n1119,
    n775
  );


  nor
  g1651
  (
    n1628,
    n565,
    n900,
    n500,
    n462
  );


  xor
  g1652
  (
    n1659,
    n1163,
    n498,
    n1251,
    n1235
  );


  nor
  g1653
  (
    n1547,
    n822,
    n1330,
    n1290,
    n1335
  );


  nand
  g1654
  (
    n1840,
    n800,
    n1147,
    n1316,
    n1242
  );


  nor
  g1655
  (
    n1504,
    n1329,
    n1207,
    n474,
    n1226
  );


  xor
  g1656
  (
    n1460,
    n1319,
    n728,
    n960,
    n1223
  );


  xnor
  g1657
  (
    n1763,
    n1283,
    n1199,
    n1110,
    n1196
  );


  and
  g1658
  (
    n1437,
    n1350,
    n1343,
    n1123,
    n925
  );


  nand
  g1659
  (
    n1677,
    n1155,
    n1052,
    n897,
    n1240
  );


  nand
  g1660
  (
    n1414,
    n1180,
    n1326,
    n1289,
    n381
  );


  xnor
  g1661
  (
    n1390,
    n1359,
    n1136,
    n1364,
    n1335
  );


  and
  g1662
  (
    n1692,
    n1329,
    n1201,
    n1207,
    n1223
  );


  xnor
  g1663
  (
    n1738,
    n1271,
    n1342,
    n1108,
    n1293
  );


  nor
  g1664
  (
    n1612,
    n873,
    n881,
    n1372,
    n1130
  );


  nor
  g1665
  (
    n1505,
    n360,
    n538,
    n1114,
    n1221
  );


  nor
  g1666
  (
    n1766,
    n1322,
    n853,
    n1149,
    n1223
  );


  xor
  g1667
  (
    n1663,
    n883,
    n617,
    n915,
    n362
  );


  xnor
  g1668
  (
    n1739,
    n759,
    n919,
    n1359,
    n932
  );


  nand
  g1669
  (
    n1617,
    n1053,
    n441,
    n1194,
    n1360
  );


  and
  g1670
  (
    n1475,
    n1292,
    n1328,
    n580,
    n1304
  );


  nand
  g1671
  (
    n1670,
    n433,
    n1195,
    n537,
    n420
  );


  nand
  g1672
  (
    n1509,
    n1245,
    n1339,
    n1098,
    n1211
  );


  or
  g1673
  (
    n1537,
    n1080,
    n1365,
    n1096,
    n1172
  );


  xor
  g1674
  (
    n1819,
    n363,
    n1278,
    n545,
    n1139
  );


  xor
  g1675
  (
    n1848,
    n520,
    n1331,
    n1167,
    n908
  );


  or
  g1676
  (
    n1720,
    n1184,
    n429,
    n903,
    n1082
  );


  nor
  g1677
  (
    n1676,
    n1096,
    n595,
    n1172,
    n1193
  );


  nor
  g1678
  (
    n1698,
    n1086,
    n1140,
    n733,
    n902
  );


  xnor
  g1679
  (
    n1754,
    n1131,
    n1135,
    n469,
    n931
  );


  xor
  g1680
  (
    n1709,
    n1362,
    n649,
    n699,
    n832
  );


  xnor
  g1681
  (
    n1585,
    n810,
    n781,
    n1307,
    n544
  );


  nand
  g1682
  (
    n1498,
    n1171,
    n1263,
    n514,
    n1337
  );


  nor
  g1683
  (
    n1642,
    n1151,
    n1370,
    n1181,
    n475
  );


  and
  g1684
  (
    n1737,
    n1358,
    n1204,
    n933
  );


  and
  g1685
  (
    n1623,
    n1345,
    n1134,
    n395,
    n530
  );


  xnor
  g1686
  (
    n1674,
    n1254,
    n1038,
    n432,
    n488
  );


  xor
  g1687
  (
    n1695,
    n1307,
    n610,
    n358,
    n1300
  );


  or
  g1688
  (
    n1449,
    n926,
    n1358,
    n1371,
    n864
  );


  xnor
  g1689
  (
    n1767,
    n1369,
    n1360,
    n1096,
    n1035
  );


  or
  g1690
  (
    n1563,
    n398,
    n1141,
    n386,
    n711
  );


  xnor
  g1691
  (
    n1778,
    n1296,
    n1138,
    n753,
    n1012
  );


  xor
  g1692
  (
    n1423,
    n968,
    n819,
    n992,
    n906
  );


  xnor
  g1693
  (
    n1759,
    n689,
    n1013,
    n685,
    n944
  );


  nand
  g1694
  (
    n1575,
    n1182,
    n1124,
    n1347,
    n481
  );


  nand
  g1695
  (
    n1744,
    n1266,
    n877,
    n1355,
    n686
  );


  nor
  g1696
  (
    n1545,
    n567,
    n771,
    n1293,
    n1289
  );


  nand
  g1697
  (
    n1626,
    n656,
    n835,
    n455,
    n954
  );


  nand
  g1698
  (
    n1688,
    n1363,
    n1077,
    n796,
    n505
  );


  xor
  g1699
  (
    n1499,
    n1260,
    n1175,
    n1203,
    n1167
  );


  xor
  g1700
  (
    n1837,
    n1286,
    n974,
    n784,
    n1122
  );


  xor
  g1701
  (
    n1599,
    n1297,
    n1252,
    n1231,
    n1256
  );


  or
  g1702
  (
    n1723,
    n1259,
    n1141,
    n1100,
    n1275
  );


  nor
  g1703
  (
    n1758,
    n1330,
    n590,
    n1139,
    n403
  );


  or
  g1704
  (
    n1550,
    n1121,
    n661,
    n1144,
    n1208
  );


  xor
  g1705
  (
    n1395,
    n1293,
    n1208,
    n1354,
    n359
  );


  nand
  g1706
  (
    n1649,
    n1295,
    n1118,
    n1238,
    n982
  );


  nor
  g1707
  (
    n1657,
    n1108,
    n399,
    n1361,
    n879
  );


  nand
  g1708
  (
    n1792,
    n1128,
    n1123,
    n1282,
    n1250
  );


  xor
  g1709
  (
    n1712,
    n1299,
    n1280,
    n1241,
    n1194
  );


  or
  g1710
  (
    n1620,
    n1217,
    n1203,
    n1184,
    n1151
  );


  nand
  g1711
  (
    n1466,
    n516,
    n1272,
    n1279,
    n1146
  );


  xor
  g1712
  (
    n1468,
    n1181,
    n438,
    n392,
    n1107
  );


  and
  g1713
  (
    n1513,
    n375,
    n1352,
    n1356,
    n1113
  );


  xor
  g1714
  (
    n1559,
    n1276,
    n546,
    n458,
    n532
  );


  nor
  g1715
  (
    n1710,
    n1300,
    n1133,
    n1250,
    n1324
  );


  xnor
  g1716
  (
    n1823,
    n787,
    n1290,
    n1248,
    n1055
  );


  xor
  g1717
  (
    n1671,
    n1185,
    n1107,
    n1109,
    n1286
  );


  nand
  g1718
  (
    n1541,
    n1303,
    n1136,
    n1273,
    n1255
  );


  xnor
  g1719
  (
    n1624,
    n511,
    n1338,
    n1282,
    n1116
  );


  xor
  g1720
  (
    n1656,
    n707,
    n1321,
    n734,
    n424
  );


  xnor
  g1721
  (
    n1534,
    n951,
    n1310,
    n788
  );


  xnor
  g1722
  (
    n1806,
    n1207,
    n1339,
    n1169,
    n635
  );


  and
  g1723
  (
    n1616,
    n1092,
    n1323,
    n1153,
    n573
  );


  or
  g1724
  (
    n1697,
    n860,
    n397,
    n1274,
    n1277
  );


  nor
  g1725
  (
    n1531,
    n747,
    n412,
    n639,
    n1295
  );


  xor
  g1726
  (
    n1646,
    n1240,
    n562,
    n1184,
    n1147
  );


  nand
  g1727
  (
    n1424,
    n708,
    n888,
    n1330,
    n557
  );


  nand
  g1728
  (
    n1409,
    n1327,
    n630,
    n1208,
    n623
  );


  xor
  g1729
  (
    n1666,
    n1118,
    n806,
    n1235,
    n1363
  );


  nor
  g1730
  (
    n1469,
    n1046,
    n576,
    n1201,
    n1147
  );


  xor
  g1731
  (
    n1496,
    n1145,
    n1199,
    n741,
    n1212
  );


  xnor
  g1732
  (
    n1641,
    n1228,
    n681,
    n579,
    n1232
  );


  nor
  g1733
  (
    n1552,
    n1224,
    n1333,
    n758,
    n1317
  );


  and
  g1734
  (
    n1700,
    n783,
    n1345,
    n377,
    n1198
  );


  or
  g1735
  (
    n1398,
    n1368,
    n754,
    n1179,
    n1287
  );


  and
  g1736
  (
    n1650,
    n735,
    n592,
    n1340,
    n1237
  );


  nor
  g1737
  (
    n1725,
    n1310,
    n366,
    n1357,
    n729
  );


  and
  g1738
  (
    n1512,
    n607,
    n1040,
    n1015,
    n1268
  );


  nand
  g1739
  (
    n1582,
    n1345,
    n1332,
    n858,
    n1166
  );


  nand
  g1740
  (
    n1638,
    n715,
    n1264,
    n1146,
    n1336
  );


  nor
  g1741
  (
    n1845,
    n1246,
    n1346,
    n1211,
    n1249
  );


  xor
  g1742
  (
    n1756,
    n1148,
    n1115,
    n838,
    n444
  );


  xor
  g1743
  (
    n1749,
    n1097,
    n1200,
    n1045,
    n1129
  );


  and
  g1744
  (
    n1562,
    n1227,
    n1247,
    n1010,
    n950
  );


  nand
  g1745
  (
    n1699,
    n407,
    n577,
    n723,
    n1101
  );


  and
  g1746
  (
    n1454,
    n1331,
    n1310,
    n714,
    n1306
  );


  xnor
  g1747
  (
    n1838,
    n1279,
    n1298,
    n1266,
    n1227
  );


  or
  g1748
  (
    n1808,
    n1237,
    n1342,
    n893,
    n1164
  );


  nor
  g1749
  (
    n1524,
    n1103,
    n1154,
    n1116,
    n1033
  );


  and
  g1750
  (
    n1543,
    n742,
    n1016,
    n940,
    n1097
  );


  or
  g1751
  (
    n1775,
    n1239,
    n1324,
    n1121,
    n1285
  );


  and
  g1752
  (
    n1662,
    n866,
    n964,
    n1170,
    n1265
  );


  or
  g1753
  (
    n1627,
    n1267,
    n1354,
    n1122,
    n1346
  );


  nand
  g1754
  (
    n1443,
    n1094,
    n1313,
    n1120,
    n624
  );


  nand
  g1755
  (
    n1630,
    n1341,
    n1128,
    n1118,
    n526
  );


  and
  g1756
  (
    n1701,
    n1269,
    n694,
    n394,
    n1357
  );


  and
  g1757
  (
    n1717,
    n1264,
    n497,
    n651,
    n1107
  );


  nor
  g1758
  (
    n1752,
    n487,
    n1121,
    n1270,
    n384
  );


  nand
  g1759
  (
    n1685,
    n1313,
    n779,
    n1213,
    n499
  );


  or
  g1760
  (
    n1637,
    n1356,
    n508,
    n1210,
    n1100
  );


  and
  g1761
  (
    n1526,
    n1191,
    n1177,
    n1334,
    n751
  );


  or
  g1762
  (
    n1429,
    n1285,
    n1265,
    n793,
    n814
  );


  nand
  g1763
  (
    n1644,
    n966,
    n850,
    n1104,
    n361
  );


  nand
  g1764
  (
    n1765,
    n1081,
    n682,
    n1190,
    n1143
  );


  and
  g1765
  (
    n1771,
    n502,
    n1074,
    n1197,
    n1110
  );


  xor
  g1766
  (
    n1614,
    n722,
    n380,
    n1137,
    n554
  );


  and
  g1767
  (
    n1634,
    n501,
    n1165,
    n1243,
    n1253
  );


  and
  g1768
  (
    KeyWire_0_4,
    n1119,
    n1123,
    n1201,
    n1348
  );


  or
  g1769
  (
    n1581,
    n1253,
    n804,
    n1257,
    n1354
  );


  or
  g1770
  (
    n1551,
    n425,
    n1329,
    n1256,
    n846
  );


  nand
  g1771
  (
    n1574,
    n1336,
    n1265,
    n1258,
    n953
  );


  or
  g1772
  (
    n1724,
    n1255,
    n654,
    n1111,
    n922
  );


  or
  g1773
  (
    n1809,
    n1044,
    n815,
    n1151,
    n938
  );


  or
  g1774
  (
    n1589,
    n541,
    n1062,
    n1267,
    n1063
  );


  xor
  g1775
  (
    n1482,
    n956,
    n700,
    n1334,
    n1097
  );


  nand
  g1776
  (
    n1431,
    n1131,
    n1163,
    n1112,
    n1030
  );


  nor
  g1777
  (
    n1658,
    n575,
    n391,
    n1262,
    n364
  );


  and
  g1778
  (
    n1439,
    n844,
    n1089,
    n1109,
    n1134
  );


  nand
  g1779
  (
    n1404,
    n435,
    n1326,
    n1180,
    n1071
  );


  or
  g1780
  (
    n1538,
    n1257,
    n1264,
    n1299,
    n1248
  );


  or
  g1781
  (
    n1401,
    n667,
    n483,
    n1215,
    n1275
  );


  nand
  g1782
  (
    n1734,
    n1159,
    n1216,
    n1064,
    n880
  );


  nor
  g1783
  (
    n1770,
    n1238,
    n486,
    n1259,
    n1176
  );


  nand
  g1784
  (
    n1399,
    n1344,
    n930,
    n1311,
    n518
  );


  and
  g1785
  (
    n1746,
    n1009,
    n606,
    n1132,
    n1145
  );


  xnor
  g1786
  (
    n1851,
    n372,
    n1163,
    n672,
    n1126
  );


  xor
  g1787
  (
    n1462,
    n1291,
    n1363,
    n1319,
    n1341
  );


  nand
  g1788
  (
    n1636,
    n1140,
    n571,
    n1095,
    n1037
  );


  xnor
  g1789
  (
    n1542,
    n1031,
    n807,
    n1170,
    n1190
  );


  or
  g1790
  (
    n1465,
    n1144,
    n1298,
    n1155,
    n471
  );


  nand
  g1791
  (
    n1502,
    n367,
    n1250,
    n578,
    n1159
  );


  or
  g1792
  (
    n1755,
    n1317,
    n1291,
    n988,
    n1292
  );


  nor
  g1793
  (
    n1633,
    n1130,
    n899,
    n1099,
    n1135
  );


  xnor
  g1794
  (
    n1532,
    n1165,
    n1095,
    n1327,
    n1196
  );


  xnor
  g1795
  (
    n1750,
    n833,
    n1245,
    n1288,
    n1357
  );


  xnor
  g1796
  (
    n1730,
    n512,
    n1192,
    n1270,
    n574
  );


  and
  g1797
  (
    n1461,
    n631,
    n1014,
    n1321,
    n1018
  );


  nor
  g1798
  (
    n1802,
    n706,
    n549,
    n1339,
    n1240
  );


  xnor
  g1799
  (
    n1731,
    n603,
    n1186,
    n702,
    n740
  );


  or
  g1800
  (
    n1430,
    n1209,
    n1214,
    n563,
    n1117
  );


  nor
  g1801
  (
    n1457,
    n1343,
    n1216,
    n1023,
    n1178
  );


  and
  g1802
  (
    KeyWire_0_29,
    n757,
    n1343,
    n569,
    n1301
  );


  xor
  g1803
  (
    n1596,
    n1236,
    n1277,
    n1272,
    n553
  );


  and
  g1804
  (
    n1781,
    n948,
    n561,
    n1099,
    n467
  );


  xnor
  g1805
  (
    n1711,
    n1150,
    n1219,
    n1072,
    n496
  );


  xnor
  g1806
  (
    n1799,
    n495,
    n748,
    n430,
    n387
  );


  and
  g1807
  (
    n1733,
    n1346,
    n1358,
    n1027,
    n1079
  );


  xor
  g1808
  (
    n1846,
    n1133,
    n1151,
    n1325,
    n792
  );


  xnor
  g1809
  (
    n1497,
    n909,
    n370,
    n390,
    n1176
  );


  nor
  g1810
  (
    n1810,
    n585,
    n1229,
    n1066,
    n1196
  );


  nor
  g1811
  (
    n1727,
    n1219,
    n1350,
    n1274,
    n404
  );


  and
  g1812
  (
    n1586,
    n1254,
    n1224,
    n693,
    n1148
  );


  xor
  g1813
  (
    n1464,
    n1340,
    n371,
    n602,
    n1284
  );


  nand
  g1814
  (
    n1760,
    n1348,
    n1247,
    n666,
    n848
  );


  xnor
  g1815
  (
    n1516,
    n1036,
    n817,
    n1356,
    n659
  );


  xor
  g1816
  (
    n1779,
    n1101,
    n426,
    n965,
    n1202
  );


  nand
  g1817
  (
    n1565,
    n1224,
    n1276,
    n560,
    n612
  );


  nor
  g1818
  (
    n1421,
    n622,
    n1359,
    n1107,
    n717
  );


  nand
  g1819
  (
    n1413,
    n937,
    n1105,
    n1321,
    n1368
  );


  or
  g1820
  (
    n1643,
    n1294,
    n1328,
    n845,
    n376
  );


  nand
  g1821
  (
    n1680,
    n882,
    n947,
    n1155,
    n1288
  );


  nor
  g1822
  (
    n1743,
    n1347,
    n1338,
    n1114,
    n692
  );


  xor
  g1823
  (
    n1510,
    n874,
    n1113,
    n1095,
    n385
  );


  and
  g1824
  (
    n1568,
    n1277,
    n818,
    n1225,
    n1120
  );


  or
  g1825
  (
    n1507,
    n1145,
    n1273,
    n658,
    n1154
  );


  nor
  g1826
  (
    n1682,
    n1021,
    n1230,
    n1325,
    n1311
  );


  or
  g1827
  (
    n1833,
    n1058,
    n1034,
    n762,
    n1215
  );


  nand
  g1828
  (
    n1564,
    n652,
    n1025,
    n978,
    n1320
  );


  nor
  g1829
  (
    n1834,
    n970,
    n1098,
    n1182,
    n1208
  );


  nand
  g1830
  (
    n1679,
    n1351,
    n1153,
    n1165,
    n1366
  );


  xnor
  g1831
  (
    n1813,
    n1361,
    n368,
    n1140,
    n710
  );


  xor
  g1832
  (
    n1719,
    n1115,
    n1176,
    n1299,
    n1248
  );


  and
  g1833
  (
    n1673,
    n539,
    n907,
    n614,
    n535
  );


  not
  g1834
  (
    n1865,
    n1404
  );


  buf
  g1835
  (
    n1862,
    n1405
  );


  buf
  g1836
  (
    n1852,
    n1407
  );


  not
  g1837
  (
    n1858,
    n1400
  );


  buf
  g1838
  (
    n1864,
    n1412
  );


  buf
  g1839
  (
    n1855,
    n1393
  );


  buf
  g1840
  (
    n1859,
    n1415
  );


  buf
  g1841
  (
    n1856,
    n1391
  );


  not
  g1842
  (
    n1863,
    n1395
  );


  not
  g1843
  (
    n1866,
    n1411
  );


  nor
  g1844
  (
    n1854,
    n1410,
    n1389,
    n1397,
    n1408
  );


  xor
  g1845
  (
    n1857,
    n1392,
    n1390,
    n1399,
    n1409
  );


  and
  g1846
  (
    n1853,
    n1417,
    n1398,
    n1413,
    n1388
  );


  and
  g1847
  (
    n1860,
    n1406,
    n1416,
    n1402,
    n1396
  );


  and
  g1848
  (
    n1861,
    n1414,
    n1403,
    n1401,
    n1394
  );


  buf
  g1849
  (
    n1881,
    n1862
  );


  not
  g1850
  (
    n1868,
    n1864
  );


  buf
  g1851
  (
    n1870,
    n1863
  );


  buf
  g1852
  (
    n1869,
    n1861
  );


  buf
  g1853
  (
    n1874,
    n1862
  );


  not
  g1854
  (
    n1885,
    n1863
  );


  not
  g1855
  (
    n1888,
    n1858
  );


  buf
  g1856
  (
    n1880,
    n1855
  );


  buf
  g1857
  (
    n1887,
    n1862
  );


  not
  g1858
  (
    n1873,
    n1864
  );


  not
  g1859
  (
    n1867,
    n1859
  );


  not
  g1860
  (
    n1871,
    n1856
  );


  not
  g1861
  (
    n1878,
    n1862
  );


  buf
  g1862
  (
    n1886,
    n1853
  );


  buf
  g1863
  (
    n1872,
    n1857
  );


  buf
  g1864
  (
    n1876,
    n1852
  );


  buf
  g1865
  (
    n1882,
    n1864
  );


  not
  g1866
  (
    n1884,
    n1863
  );


  not
  g1867
  (
    n1877,
    n1854
  );


  not
  g1868
  (
    n1883,
    n1864
  );


  not
  g1869
  (
    n1879,
    n1860
  );


  not
  g1870
  (
    n1875,
    n1863
  );


  nor
  g1871
  (
    n1896,
    n1466,
    n1871,
    n1465,
    n1515
  );


  or
  g1872
  (
    n1916,
    n1497,
    n1868,
    n1501,
    n1490
  );


  nor
  g1873
  (
    n1921,
    n1868,
    n1877,
    n1869,
    n1876
  );


  and
  g1874
  (
    n1912,
    n1873,
    n1874,
    n1536,
    n1486
  );


  xor
  g1875
  (
    n1923,
    n1427,
    n1453,
    n1418,
    n1428
  );


  xnor
  g1876
  (
    n1905,
    n1869,
    n1445,
    n1430,
    n1876
  );


  nand
  g1877
  (
    n1914,
    n1443,
    n1471,
    n1876,
    n1475
  );


  and
  g1878
  (
    n1920,
    n1477,
    n1871,
    n1875,
    n1434
  );


  and
  g1879
  (
    n1910,
    n1533,
    n1542,
    n1468,
    n1514
  );


  xor
  g1880
  (
    n1922,
    n1429,
    n1872,
    n1870,
    n1447
  );


  nand
  g1881
  (
    n1924,
    n1476,
    n1868,
    n1867,
    n1495
  );


  nor
  g1882
  (
    n1902,
    n1503,
    n1494,
    n1871,
    n1524
  );


  or
  g1883
  (
    n1913,
    n1457,
    n1874,
    n1472,
    n1869
  );


  xnor
  g1884
  (
    n1906,
    n1530,
    n1432,
    n1423,
    n1474
  );


  or
  g1885
  (
    n1901,
    n1499,
    n1870,
    n1451,
    n1534
  );


  xor
  g1886
  (
    n1911,
    n1543,
    n1518,
    n1446,
    n1437
  );


  xor
  g1887
  (
    n1889,
    n1875,
    n1482,
    n1450,
    n1425
  );


  or
  g1888
  (
    n1915,
    n1505,
    n1867,
    n1440
  );


  nand
  g1889
  (
    n1894,
    n1873,
    n1419,
    n1421,
    n1500
  );


  nor
  g1890
  (
    n1925,
    n1502,
    n1867,
    n1481,
    n1872
  );


  and
  g1891
  (
    n1898,
    n1877,
    n1422,
    n1492,
    n1522
  );


  xor
  g1892
  (
    n1917,
    n1467,
    n1876,
    n1875,
    n1458
  );


  xnor
  g1893
  (
    n1927,
    n1535,
    n1508,
    n1531,
    n1438
  );


  nand
  g1894
  (
    n1928,
    n1480,
    n1519,
    n1875,
    n1470
  );


  or
  g1895
  (
    n1897,
    n1869,
    n1491,
    n1461,
    n1511
  );


  and
  g1896
  (
    n1919,
    n1424,
    n1512,
    n1460,
    n1504
  );


  xnor
  g1897
  (
    n1892,
    n1479,
    n1527,
    n1442,
    n1473
  );


  xnor
  g1898
  (
    n1893,
    n1541,
    n1478,
    n1521,
    n1516
  );


  or
  g1899
  (
    n1929,
    n1431,
    n1469,
    n1513,
    n1452
  );


  xor
  g1900
  (
    n1895,
    n1462,
    n1456,
    n1444,
    n1420
  );


  and
  g1901
  (
    n1890,
    n1506,
    n1454,
    n1433,
    n1509
  );


  nor
  g1902
  (
    n1891,
    n1507,
    n1874,
    n1870,
    n1441
  );


  nand
  g1903
  (
    n1909,
    n1487,
    n1426,
    n1459,
    n1449
  );


  xnor
  g1904
  (
    n1908,
    n1874,
    n1523,
    n1498,
    n1529
  );


  xor
  g1905
  (
    n1918,
    n1870,
    n1872,
    n1510,
    n1488
  );


  nor
  g1906
  (
    n1907,
    n1539,
    n1528,
    n1871,
    n1496
  );


  and
  g1907
  (
    n1899,
    n1526,
    n1868,
    n1455,
    n1463
  );


  and
  g1908
  (
    n1904,
    n1520,
    n1485,
    n1872,
    n1532
  );


  nand
  g1909
  (
    n1903,
    n1517,
    n1464,
    n1493,
    n1540
  );


  xnor
  g1910
  (
    n1900,
    n1439,
    n1489,
    n1538,
    n1435
  );


  xor
  g1911
  (
    n1930,
    n1484,
    n1448,
    n1483,
    n1436
  );


  nor
  g1912
  (
    n1926,
    n1525,
    n1537,
    n1873
  );


  nand
  g1913
  (
    n1938,
    n1547,
    n1920,
    n1553,
    n1565
  );


  xnor
  g1914
  (
    n1937,
    n1566,
    n1563,
    n1552,
    n1562
  );


  nand
  g1915
  (
    n1931,
    n1918,
    n1551,
    n1554,
    n1546
  );


  xor
  g1916
  (
    n1932,
    n1559,
    n1557,
    n1919,
    n1560
  );


  nand
  g1917
  (
    n1936,
    n1550,
    n1545,
    n1549,
    n1922
  );


  nand
  g1918
  (
    n1933,
    n1555,
    n1561,
    n1921,
    n1564
  );


  and
  g1919
  (
    n1934,
    n1544,
    n1915,
    n1556,
    n1917
  );


  xor
  g1920
  (
    n1935,
    n1548,
    n1567,
    n1558,
    n1916
  );


  xnor
  g1921
  (
    n1944,
    n1883,
    n1883,
    n1879,
    n1881
  );


  and
  g1922
  (
    n1940,
    n1937,
    n1578,
    n1572,
    n1879
  );


  xnor
  g1923
  (
    n1951,
    n1583,
    n1882,
    n1587,
    n1879
  );


  nor
  g1924
  (
    n1945,
    n1586,
    n1937,
    n1931,
    n1579
  );


  and
  g1925
  (
    n1939,
    n1933,
    n1878,
    n1934,
    n1935
  );


  nand
  g1926
  (
    n1949,
    n1932,
    n1882,
    n1935,
    n1880
  );


  nor
  g1927
  (
    n1950,
    n1881,
    n1882,
    n1573,
    n1879
  );


  nand
  g1928
  (
    n1941,
    n1582,
    n1880,
    n1877
  );


  nand
  g1929
  (
    n1952,
    n1585,
    n1883,
    n1938,
    n1881
  );


  and
  g1930
  (
    n1953,
    n1580,
    n1937,
    n1936,
    n1880
  );


  or
  g1931
  (
    n1943,
    n1936,
    n1584,
    n1571,
    n1878
  );


  xor
  g1932
  (
    n1942,
    n1937,
    n1581,
    n1938
  );


  xor
  g1933
  (
    n1948,
    n1878,
    n1570,
    n1574,
    n1577
  );


  xnor
  g1934
  (
    n1946,
    n1882,
    n1877,
    n1576,
    n1878
  );


  nand
  g1935
  (
    n1947,
    n1881,
    n1569,
    n1568,
    n1575
  );


  nor
  g1936
  (
    n1955,
    n1595,
    n1591,
    n1948
  );


  xnor
  g1937
  (
    n1961,
    n1951,
    n1950,
    n1930
  );


  and
  g1938
  (
    n1964,
    n1376,
    n1939,
    n1372
  );


  xor
  g1939
  (
    n1957,
    n1600,
    n1378,
    n1373
  );


  nor
  g1940
  (
    n1963,
    n1601,
    n1375,
    n1923,
    n1592
  );


  and
  g1941
  (
    n1968,
    n1373,
    n1378,
    n1375,
    n1379
  );


  or
  g1942
  (
    n1974,
    n1594,
    n1945,
    n1377,
    n1589
  );


  nor
  g1943
  (
    n1969,
    n1590,
    n1593,
    n1952,
    n1376
  );


  nand
  g1944
  (
    n1967,
    n1602,
    n1377,
    n1952,
    n1374
  );


  nand
  g1945
  (
    n1962,
    n1949,
    n1375,
    n1951,
    n1378
  );


  and
  g1946
  (
    n1960,
    n1941,
    n1603,
    n1942,
    n1379
  );


  or
  g1947
  (
    n1959,
    n1377,
    n1588,
    n1376,
    n1926
  );


  xnor
  g1948
  (
    n1970,
    n1949,
    n1375,
    n1372,
    n1373
  );


  nand
  g1949
  (
    n1972,
    n1951,
    n1374,
    n1379,
    n1927
  );


  xor
  g1950
  (
    n1954,
    n1946,
    n1374,
    n1928,
    n1944
  );


  and
  g1951
  (
    n1958,
    n1950,
    n1377,
    n1943,
    n1924
  );


  xor
  g1952
  (
    n1966,
    n1950,
    n1599,
    n1597,
    n1373
  );


  xor
  g1953
  (
    n1956,
    n1929,
    n1950,
    n1947,
    n1952
  );


  nand
  g1954
  (
    n1971,
    n1952,
    n1376,
    n1380,
    n1596
  );


  or
  g1955
  (
    n1965,
    n1951,
    n1940,
    n1380,
    n1374
  );


  or
  g1956
  (
    n1973,
    n1598,
    n1379,
    n1378,
    n1925
  );


  nor
  g1957
  (
    n1976,
    n1954,
    n1608,
    n1604,
    n1606
  );


  xor
  g1958
  (
    n1975,
    n1955,
    n1607,
    n1609,
    n1605
  );


  xor
  g1959
  (
    n1982,
    n1622,
    n1623,
    n1381
  );


  or
  g1960
  (
    n1978,
    n1975,
    n1380,
    n1976,
    n1621
  );


  and
  g1961
  (
    n1980,
    n1620,
    n1381,
    n1618,
    n1625
  );


  and
  g1962
  (
    n1983,
    n1611,
    n1619,
    n1976,
    n1614
  );


  or
  g1963
  (
    n1979,
    n1975,
    n1975,
    n1381,
    n1613
  );


  nor
  g1964
  (
    KeyWire_0_9,
    n1615,
    n1381,
    n1610,
    n1617
  );


  nand
  g1965
  (
    n1981,
    n1616,
    n1976,
    n1975,
    n1624
  );


  nand
  g1966
  (
    KeyWire_0_30,
    n1382,
    n1380,
    n1612,
    n1976
  );


  buf
  g1967
  (
    n1986,
    n1628
  );


  buf
  g1968
  (
    n1996,
    n1978
  );


  buf
  g1969
  (
    n1993,
    n1977
  );


  not
  g1970
  (
    n1985,
    n1977
  );


  not
  g1971
  (
    n1992,
    n1980
  );


  not
  g1972
  (
    n1988,
    n1977
  );


  buf
  g1973
  (
    n1991,
    n1627
  );


  not
  g1974
  (
    n1995,
    n1630
  );


  or
  g1975
  (
    n1989,
    n1979,
    n1978
  );


  xor
  g1976
  (
    n1994,
    n1634,
    n1979,
    n1635,
    n1626
  );


  xor
  g1977
  (
    n1990,
    n1636,
    n1977,
    n1978,
    n1629
  );


  nand
  g1978
  (
    n1987,
    n1632,
    n1631,
    n1637,
    n1979
  );


  nand
  g1979
  (
    n1997,
    n1979,
    n1638,
    n1633,
    n1978
  );


  not
  g1980
  (
    n2000,
    n1992
  );


  buf
  g1981
  (
    n2002,
    n1991
  );


  not
  g1982
  (
    n1999,
    n1640
  );


  not
  g1983
  (
    n2001,
    n1639
  );


  or
  g1984
  (
    n1998,
    n1641,
    n1994,
    n1993,
    n1990
  );


  xnor
  g1985
  (
    n2004,
    n2001,
    n1980,
    n1981
  );


  nand
  g1986
  (
    n2003,
    n1982,
    n2000,
    n1980,
    n1999
  );


  and
  g1987
  (
    n2005,
    n1981,
    n1998,
    n1982
  );


  nand
  g1988
  (
    n2006,
    n1982,
    n1981,
    n354
  );


  xor
  g1989
  (
    n2007,
    n1643,
    n2004,
    n1645,
    n2003
  );


  nor
  g1990
  (
    n2008,
    n1644,
    n1642,
    n1646,
    n1382
  );


  xnor
  g1991
  (
    n2009,
    n1649,
    n1647,
    n1648,
    n2007
  );


  and
  g1992
  (
    n2011,
    n2009,
    n1655,
    n1653,
    n1650
  );


  or
  g1993
  (
    n2010,
    n1651,
    n1652,
    n2009,
    n1654
  );


  and
  g1994
  (
    n2018,
    n1662,
    n2011
  );


  nor
  g1995
  (
    n2012,
    n1658,
    n2010
  );


  nand
  g1996
  (
    n2016,
    n2011,
    n1660
  );


  xor
  g1997
  (
    n2017,
    n2010,
    n2011
  );


  nor
  g1998
  (
    n2019,
    n2011,
    n1663
  );


  xor
  g1999
  (
    n2013,
    n1657,
    n2010
  );


  nor
  g2000
  (
    n2014,
    n1656,
    n1661
  );


  xor
  g2001
  (
    n2015,
    n1659,
    n2010
  );


  not
  g2002
  (
    n2024,
    n1383
  );


  buf
  g2003
  (
    n2020,
    n2012
  );


  buf
  g2004
  (
    n2023,
    n1382
  );


  buf
  g2005
  (
    n2021,
    n2012
  );


  nand
  g2006
  (
    n2025,
    n1382,
    n2013,
    n2012
  );


  or
  g2007
  (
    n2022,
    n2012,
    n2013,
    n1383
  );


  xnor
  g2008
  (
    n2035,
    n1685,
    n1678,
    n1722,
    n1717
  );


  or
  g2009
  (
    n2038,
    n1723,
    n1668,
    n1711,
    n1699
  );


  xor
  g2010
  (
    n2044,
    n2024,
    n2021,
    n1714,
    n2020
  );


  nand
  g2011
  (
    n2042,
    n1708,
    n1680,
    n2022,
    n1709
  );


  or
  g2012
  (
    n2036,
    n1673,
    n1712,
    n1706,
    n1696
  );


  or
  g2013
  (
    n2037,
    n2023,
    n1718,
    n1689,
    n2022
  );


  nor
  g2014
  (
    n2028,
    n1674,
    n1666,
    n1690,
    n1693
  );


  or
  g2015
  (
    n2040,
    n1710,
    n2023,
    n1701,
    n1681
  );


  xor
  g2016
  (
    n2030,
    n1704,
    n2022,
    n1716,
    n2020
  );


  xor
  g2017
  (
    n2032,
    n1705,
    n1667,
    n1715,
    n1670
  );


  nand
  g2018
  (
    n2027,
    n1682,
    n1721,
    n1684,
    n1697
  );


  and
  g2019
  (
    n2029,
    n1695,
    n1692,
    n1686,
    n1687
  );


  or
  g2020
  (
    n2043,
    n2023,
    n1698,
    n1691,
    n1694
  );


  xor
  g2021
  (
    n2045,
    n2020,
    n2024,
    n2021,
    n1664
  );


  xnor
  g2022
  (
    n2033,
    n1665,
    n1700,
    n2021,
    n1676
  );


  or
  g2023
  (
    n2041,
    n1702,
    n1679,
    n1707,
    n2024
  );


  nand
  g2024
  (
    n2026,
    n1683,
    n1672,
    n1713,
    n1677
  );


  nand
  g2025
  (
    n2039,
    n1669,
    n1703,
    n2021,
    n2020
  );


  xnor
  g2026
  (
    n2034,
    n2023,
    n2024,
    n1671,
    n1675
  );


  xor
  g2027
  (
    n2031,
    n2022,
    n1719,
    n1720,
    n1688
  );


  and
  g2028
  (
    n2049,
    n2018,
    n1866
  );


  nor
  g2029
  (
    n2059,
    n2014,
    n2019,
    n2017,
    n1983
  );


  nor
  g2030
  (
    n2051,
    n2037,
    n1865,
    n1984,
    n2035
  );


  nand
  g2031
  (
    n2047,
    n1984,
    n2014,
    n2018,
    n2026
  );


  nand
  g2032
  (
    n2046,
    n2019,
    n2027,
    n2017,
    n2036
  );


  nand
  g2033
  (
    n2048,
    n1983,
    n2019,
    n1984
  );


  nor
  g2034
  (
    n2058,
    n2040,
    n1983,
    n2017,
    n1866
  );


  or
  g2035
  (
    n2054,
    n2014,
    n2015,
    n2016,
    n2013
  );


  and
  g2036
  (
    n2055,
    n2016,
    n2031,
    n2029,
    n2018
  );


  and
  g2037
  (
    n2060,
    n1983,
    n2034,
    n2013,
    n2017
  );


  xor
  g2038
  (
    n2050,
    n1865,
    n1866,
    n2032
  );


  nor
  g2039
  (
    n2056,
    n2030,
    n2039,
    n2028,
    n2014
  );


  xor
  g2040
  (
    n2057,
    n2038,
    n2015,
    n2041
  );


  nand
  g2041
  (
    n2052,
    n2018,
    n2033,
    n1865,
    n2016
  );


  xnor
  g2042
  (
    n2053,
    n1984,
    n2016,
    n2015,
    n1865
  );


  nor
  g2043
  (
    n2070,
    n1996,
    n2057,
    n1958
  );


  xor
  g2044
  (
    KeyWire_0_8,
    n1888,
    n2056,
    n2055
  );


  xor
  g2045
  (
    n2064,
    n2047,
    n1885,
    n2046,
    n1884
  );


  xor
  g2046
  (
    n2066,
    n1997,
    n2025,
    n2056,
    n1953
  );


  or
  g2047
  (
    n2071,
    n1959,
    n1887,
    n2025
  );


  nor
  g2048
  (
    n2077,
    n1888,
    n2057,
    n2054,
    n1953
  );


  and
  g2049
  (
    n2075,
    n2050,
    n1885,
    n1957,
    n1883
  );


  nor
  g2050
  (
    n2061,
    n1959,
    n1886,
    n1953,
    n2058
  );


  xnor
  g2051
  (
    n2063,
    n2052,
    n2059,
    n2054,
    n1886
  );


  nand
  g2052
  (
    n2068,
    n2054,
    n1888,
    n2056,
    n1959
  );


  xor
  g2053
  (
    n2069,
    n1958,
    n1958,
    n2055,
    n1885
  );


  nor
  g2054
  (
    n2067,
    n1886,
    n1959,
    n1938,
    n2025
  );


  and
  g2055
  (
    n2062,
    n1884,
    n1886,
    n1888,
    n1995
  );


  nand
  g2056
  (
    n2078,
    n2054,
    n2055,
    n1887,
    n1884
  );


  nor
  g2057
  (
    n2072,
    n2048,
    n2058,
    n1958
  );


  or
  g2058
  (
    KeyWire_0_27,
    n2049,
    n1885,
    n2025,
    n2058
  );


  xnor
  g2059
  (
    n2073,
    n2053,
    n1956,
    n1953,
    n2051
  );


  nor
  g2060
  (
    n2076,
    n2057,
    n1884,
    n2055,
    n1887
  );


  not
  g2061
  (
    n2097,
    n2064
  );


  not
  g2062
  (
    n2088,
    n2066
  );


  not
  g2063
  (
    n2096,
    n2063
  );


  or
  g2064
  (
    n2103,
    n2045,
    n1968,
    n1736,
    n1974
  );


  xnor
  g2065
  (
    n2091,
    n1969,
    n1962,
    n2062,
    n1970
  );


  nand
  g2066
  (
    n2107,
    n1727,
    n2065,
    n1730
  );


  or
  g2067
  (
    n2100,
    n1733,
    n1974,
    n1970
  );


  xor
  g2068
  (
    n2110,
    n1961,
    n1964,
    n1734,
    n2069
  );


  nor
  g2069
  (
    n2098,
    n1967,
    n1960,
    n2069,
    n2045
  );


  xor
  g2070
  (
    n2108,
    n2067,
    n1972,
    n1960,
    n2065
  );


  xnor
  g2071
  (
    n2101,
    n1961,
    n2069,
    n1970,
    n1968
  );


  nand
  g2072
  (
    n2094,
    n2042,
    n1729,
    n2061,
    n2043
  );


  xor
  g2073
  (
    n2109,
    n1971,
    n1964,
    n1963,
    n2070
  );


  xnor
  g2074
  (
    n2095,
    n2045,
    n2068,
    n2069,
    n2064
  );


  xor
  g2075
  (
    n2079,
    n2068,
    n1738,
    n1735,
    n1973
  );


  and
  g2076
  (
    n2102,
    n2066,
    n2067,
    n1966,
    n1968
  );


  nand
  g2077
  (
    n2083,
    n1725,
    n1966,
    n1963,
    n1967
  );


  nand
  g2078
  (
    n2082,
    n2061,
    n2067,
    n1973,
    n1960
  );


  xor
  g2079
  (
    n2085,
    n1732,
    n2068,
    n2061,
    n1961
  );


  xnor
  g2080
  (
    n2081,
    n1967,
    n1971,
    n1964,
    n1962
  );


  nand
  g2081
  (
    n2104,
    n1963,
    n1972,
    n1965,
    n1966
  );


  xnor
  g2082
  (
    n2105,
    n2062,
    n2062,
    n2045,
    n2066
  );


  xor
  g2083
  (
    n2086,
    n1971,
    n2044,
    n1731,
    n2063
  );


  nor
  g2084
  (
    n2089,
    n1969,
    n1961,
    n2063,
    n2061
  );


  nand
  g2085
  (
    n2087,
    n2065,
    n1726,
    n2063,
    n1965
  );


  or
  g2086
  (
    n2092,
    n1724,
    n1966,
    n1964,
    n2064
  );


  nor
  g2087
  (
    n2099,
    n2002,
    n1972,
    n1962,
    n2066
  );


  and
  g2088
  (
    n2084,
    n1962,
    n1968,
    n1965,
    n2064
  );


  or
  g2089
  (
    n2080,
    n1737,
    n1965,
    n2067,
    n2068
  );


  xnor
  g2090
  (
    n2090,
    n2062,
    n1971,
    n1969
  );


  and
  g2091
  (
    n2093,
    n1974,
    n1972,
    n1973,
    n1728
  );


  nand
  g2092
  (
    n2106,
    n1967,
    n1973,
    n1960,
    n1963
  );


  or
  g2093
  (
    n2116,
    n2060,
    n2090,
    n2059,
    n2107
  );


  or
  g2094
  (
    n2113,
    n2080,
    n2081,
    n1740,
    n2110
  );


  and
  g2095
  (
    n2114,
    n1974,
    n2102,
    n2079,
    n2094
  );


  and
  g2096
  (
    n2125,
    n2107,
    n2106,
    n355,
    n2060
  );


  nand
  g2097
  (
    n2111,
    n2106,
    n2110,
    n354,
    n2109
  );


  xor
  g2098
  (
    n2112,
    n2086,
    n2110,
    n2109,
    n2059
  );


  and
  g2099
  (
    n2118,
    n2083,
    n2099,
    n2089,
    n2107
  );


  xnor
  g2100
  (
    n2124,
    n2108,
    n2108,
    n2087,
    n2101
  );


  xor
  g2101
  (
    n2117,
    n2085,
    n2109,
    n1741,
    n2093
  );


  nor
  g2102
  (
    n2122,
    n1742,
    n2060,
    n2103,
    n2109
  );


  or
  g2103
  (
    n2119,
    n2092,
    n2006,
    n2097,
    n2084
  );


  or
  g2104
  (
    n2115,
    n2105,
    n2059,
    n2098,
    n2106
  );


  nor
  g2105
  (
    n2120,
    n2104,
    n2110,
    n2060,
    n2100
  );


  and
  g2106
  (
    n2121,
    n2006,
    n2107,
    n2088,
    n2108
  );


  nand
  g2107
  (
    n2126,
    n2082,
    n2091,
    n2108,
    n2106
  );


  nor
  g2108
  (
    n2123,
    n2096,
    n2095,
    n1739,
    n2005
  );


  nand
  g2109
  (
    n2140,
    n2075,
    n1386,
    n2078,
    n2122
  );


  nand
  g2110
  (
    n2145,
    n2077,
    n1385,
    n2073,
    n2118
  );


  xnor
  g2111
  (
    n2128,
    n2070,
    n2074,
    n2077,
    n2076
  );


  nand
  g2112
  (
    n2144,
    n2074,
    n2073,
    n2075,
    n2008
  );


  xnor
  g2113
  (
    n2132,
    n2120,
    n2076,
    n2122,
    n2072
  );


  xor
  g2114
  (
    n2127,
    n2072,
    n2078,
    n2121
  );


  and
  g2115
  (
    n2136,
    n1385,
    n2121,
    n2072,
    n2071
  );


  xor
  g2116
  (
    n2130,
    n2073,
    n1744,
    n2072,
    n1386
  );


  and
  g2117
  (
    n2146,
    n2070,
    n2070,
    n1745,
    n2075
  );


  nand
  g2118
  (
    n2141,
    n1743,
    n1387,
    n1385,
    n2073
  );


  xnor
  g2119
  (
    n2129,
    n1384,
    n2117,
    n2071
  );


  xnor
  g2120
  (
    n2139,
    n2114,
    n2121,
    n2115,
    n1384
  );


  xnor
  g2121
  (
    n2133,
    n2116,
    n2076,
    n1747,
    n1387
  );


  xor
  g2122
  (
    n2142,
    n1387,
    n2120,
    n2076,
    n2122
  );


  or
  g2123
  (
    n2135,
    n1384,
    n1384,
    n2078,
    n2074
  );


  and
  g2124
  (
    n2143,
    n1383,
    n2120,
    n2112,
    n2077
  );


  and
  g2125
  (
    n2138,
    n2071,
    n2122,
    n1383,
    n1387
  );


  xor
  g2126
  (
    n2134,
    n2113,
    n2111,
    n1386,
    n1746
  );


  xor
  g2127
  (
    n2137,
    n1385,
    n2074,
    n2119,
    n1386
  );


  nor
  g2128
  (
    n2131,
    n2120,
    n2078,
    n2077,
    n2075
  );


  nand
  g2129
  (
    n2168,
    n1809,
    n1768,
    n1760,
    n1804
  );


  xnor
  g2130
  (
    n2152,
    n1778,
    n1772,
    n1797,
    n1813
  );


  nor
  g2131
  (
    n2148,
    n1752,
    n1803,
    n2144,
    n2141
  );


  nor
  g2132
  (
    n2165,
    n1792,
    n1793,
    n1758,
    n1823
  );


  nand
  g2133
  (
    n2174,
    n2142,
    n1764,
    n1749,
    n1763
  );


  xor
  g2134
  (
    n2156,
    n1802,
    n1815,
    n1818,
    n1755
  );


  xor
  g2135
  (
    n2154,
    n1795,
    n1766,
    n2128,
    n1785
  );


  and
  g2136
  (
    n2150,
    n2143,
    n2138,
    n2142,
    n1820
  );


  or
  g2137
  (
    n2155,
    n1789,
    n1800,
    n1750,
    n2139
  );


  nor
  g2138
  (
    n2170,
    n2143,
    n1779,
    n1751,
    n1759
  );


  xnor
  g2139
  (
    n2160,
    n2136,
    n2144,
    n1774,
    n2142
  );


  or
  g2140
  (
    n2158,
    n2127,
    n1817,
    n1811,
    n2145
  );


  xor
  g2141
  (
    n2153,
    n1787,
    n1769,
    n2137,
    n1805
  );


  and
  g2142
  (
    n2163,
    n1828,
    n1821,
    n1794,
    n1829
  );


  or
  g2143
  (
    n2171,
    n1773,
    n1819,
    n2131,
    n1753
  );


  xnor
  g2144
  (
    n2173,
    n1765,
    n1806,
    n1814,
    n1824
  );


  xnor
  g2145
  (
    n2159,
    n2132,
    n2134,
    n1762,
    n1799
  );


  xor
  g2146
  (
    n2161,
    n1770,
    n2143,
    n2144,
    n1771
  );


  nand
  g2147
  (
    n2169,
    n2142,
    n1827,
    n2144,
    n1761
  );


  or
  g2148
  (
    n2157,
    n1756,
    n2129,
    n1801,
    n1775
  );


  and
  g2149
  (
    n2151,
    n1754,
    n1767,
    n1788,
    n1776
  );


  nor
  g2150
  (
    n2164,
    n1807,
    n1781,
    n1796,
    n1816
  );


  xnor
  g2151
  (
    n2149,
    n1798,
    n1783,
    n1830,
    n2130
  );


  or
  g2152
  (
    n2167,
    n1812,
    n1780,
    n1784,
    n1831
  );


  or
  g2153
  (
    n2147,
    n1748,
    n2133,
    n2143,
    n1786
  );


  xor
  g2154
  (
    n2166,
    n1810,
    n1808,
    n1782,
    n2135
  );


  or
  g2155
  (
    n2162,
    n1777,
    n1791,
    n1790,
    n1822
  );


  and
  g2156
  (
    n2172,
    n2140,
    n1757,
    n1826,
    n1825
  );


  nand
  g2157
  (
    n2188,
    n1837,
    n2123,
    n1844
  );


  and
  g2158
  (
    n2175,
    n2149,
    n1836,
    n1840,
    n2170
  );


  or
  g2159
  (
    n2178,
    n2161,
    n1838,
    n2165,
    n1847
  );


  or
  g2160
  (
    n2179,
    n2159,
    n2168,
    n2160,
    n1846
  );


  xnor
  g2161
  (
    n2183,
    n1839,
    n1845,
    n2154,
    n2171
  );


  and
  g2162
  (
    n2176,
    n2170,
    n2166,
    n1832,
    n2171
  );


  nand
  g2163
  (
    n2177,
    n2169,
    n2123,
    n2170,
    n2167
  );


  or
  g2164
  (
    n2185,
    n2148,
    n2125,
    n2170,
    n2163
  );


  xor
  g2165
  (
    n2182,
    n2147,
    n1843,
    n2124,
    n1833
  );


  xnor
  g2166
  (
    n2180,
    n1842,
    n1841,
    n2157,
    n2156
  );


  nor
  g2167
  (
    n2181,
    n2150,
    n1835,
    n2124,
    n2171
  );


  xor
  g2168
  (
    n2186,
    n2155,
    n2164,
    n2151,
    n2171
  );


  xnor
  g2169
  (
    n2187,
    n2123,
    n2124,
    n2153
  );


  nor
  g2170
  (
    n2184,
    n1834,
    n2152,
    n2162,
    n2158
  );


  xor
  g2171
  (
    n2198,
    n2125,
    n2174,
    n2173,
    n2177
  );


  or
  g2172
  (
    n2192,
    n2126,
    n1851,
    n2184,
    n2172
  );


  nand
  g2173
  (
    n2193,
    n355,
    n2174,
    n356,
    n2179
  );


  xnor
  g2174
  (
    n2201,
    n1850,
    n355,
    n1848,
    n2146
  );


  nand
  g2175
  (
    n2194,
    n2173,
    n2185,
    n356,
    n2175
  );


  and
  g2176
  (
    n2197,
    n2146,
    n355,
    n2174
  );


  or
  g2177
  (
    n2199,
    n2145,
    n1849,
    n2125,
    n2176
  );


  or
  g2178
  (
    n2196,
    n2172,
    n2146,
    n2178,
    n2188
  );


  xnor
  g2179
  (
    n2191,
    n2145,
    n2126
  );


  and
  g2180
  (
    n2200,
    n2125,
    n2173,
    n2172
  );


  and
  g2181
  (
    n2190,
    n2172,
    n2180,
    n2186,
    n356
  );


  nand
  g2182
  (
    n2189,
    n357,
    n2181,
    n356,
    n2146
  );


  nor
  g2183
  (
    n2195,
    n2145,
    n2182,
    n2187,
    n2183
  );


  xnor
  g2184
  (
    n2205,
    n2194,
    n357,
    n2195
  );


  or
  g2185
  (
    n2204,
    n2191,
    n2199,
    n2192,
    n2197
  );


  xor
  g2186
  (
    n2202,
    n357,
    n2200,
    n2193,
    n2196
  );


  nor
  g2187
  (
    n2203,
    n2198,
    n2201,
    n2190,
    n2189
  );


  xnor
  KeyGate_0_0
  (
    n1328,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1127,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1492,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1320,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1645,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n448,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1334,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n234,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n2074,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1977,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n732,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n279,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n505,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n48,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n925,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1479,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1029,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1590,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n22,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n120,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1278,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n904,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1344,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1558,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n850,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n719,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1065,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n2065,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n599,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n1784,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1984,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1325,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


