

module Stat_376_810
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n375,
  n377,
  n396,
  n386,
  n394,
  n380,
  n382,
  n374,
  n383,
  n384,
  n388,
  n392,
  n381,
  n390,
  n393,
  n395,
  n379,
  n389,
  n376,
  n378,
  n391,
  n385,
  n387,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n375;
  output n377;
  output n396;
  output n386;
  output n394;
  output n380;
  output n382;
  output n374;
  output n383;
  output n384;
  output n388;
  output n392;
  output n381;
  output n390;
  output n393;
  output n395;
  output n379;
  output n389;
  output n376;
  output n378;
  output n391;
  output n385;
  output n387;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n35,
    n1
  );


  not
  g1
  (
    n41,
    n5
  );


  not
  g2
  (
    n42,
    n5
  );


  buf
  g3
  (
    n34,
    n3
  );


  not
  g4
  (
    n26,
    n4
  );


  not
  g5
  (
    n23,
    n4
  );


  not
  g6
  (
    n27,
    n1
  );


  not
  g7
  (
    n40,
    n2
  );


  buf
  g8
  (
    n21,
    n5
  );


  not
  g9
  (
    n30,
    n1
  );


  not
  g10
  (
    n31,
    n3
  );


  not
  g11
  (
    n33,
    n3
  );


  buf
  g12
  (
    n29,
    n2
  );


  not
  g13
  (
    n38,
    n2
  );


  buf
  g14
  (
    n36,
    n4
  );


  not
  g15
  (
    n28,
    n6
  );


  buf
  g16
  (
    n24,
    n3
  );


  not
  g17
  (
    n39,
    n4
  );


  not
  g18
  (
    n32,
    n5
  );


  not
  g19
  (
    n22,
    n1
  );


  buf
  g20
  (
    n25,
    n6
  );


  buf
  g21
  (
    n37,
    n2
  );


  buf
  g22
  (
    n114,
    n16
  );


  not
  g23
  (
    n90,
    n38
  );


  buf
  g24
  (
    n69,
    n34
  );


  buf
  g25
  (
    n64,
    n10
  );


  buf
  g26
  (
    n53,
    n25
  );


  buf
  g27
  (
    KeyWire_0_11,
    n35
  );


  buf
  g28
  (
    n51,
    n32
  );


  not
  g29
  (
    n103,
    n22
  );


  buf
  g30
  (
    n126,
    n32
  );


  not
  g31
  (
    n87,
    n36
  );


  buf
  g32
  (
    n56,
    n40
  );


  buf
  g33
  (
    n98,
    n9
  );


  buf
  g34
  (
    n109,
    n40
  );


  not
  g35
  (
    n112,
    n8
  );


  not
  g36
  (
    n47,
    n11
  );


  buf
  g37
  (
    n127,
    n7
  );


  not
  g38
  (
    n116,
    n6
  );


  buf
  g39
  (
    KeyWire_0_1,
    n38
  );


  not
  g40
  (
    n75,
    n29
  );


  not
  g41
  (
    n128,
    n30
  );


  buf
  g42
  (
    n52,
    n27
  );


  buf
  g43
  (
    n46,
    n13
  );


  buf
  g44
  (
    n83,
    n23
  );


  not
  g45
  (
    n68,
    n29
  );


  buf
  g46
  (
    n118,
    n21
  );


  buf
  g47
  (
    KeyWire_0_10,
    n27
  );


  buf
  g48
  (
    n49,
    n7
  );


  buf
  g49
  (
    KeyWire_0_6,
    n31
  );


  not
  g50
  (
    n104,
    n41
  );


  buf
  g51
  (
    n106,
    n6
  );


  buf
  g52
  (
    n82,
    n26
  );


  buf
  g53
  (
    n85,
    n16
  );


  buf
  g54
  (
    n77,
    n23
  );


  buf
  g55
  (
    n92,
    n8
  );


  buf
  g56
  (
    n57,
    n34
  );


  not
  g57
  (
    n66,
    n33
  );


  not
  g58
  (
    n50,
    n25
  );


  not
  g59
  (
    n96,
    n9
  );


  not
  g60
  (
    n99,
    n31
  );


  not
  g61
  (
    n71,
    n17
  );


  buf
  g62
  (
    n59,
    n15
  );


  not
  g63
  (
    n120,
    n37
  );


  buf
  g64
  (
    n122,
    n10
  );


  not
  g65
  (
    n58,
    n29
  );


  buf
  g66
  (
    n55,
    n10
  );


  not
  g67
  (
    n70,
    n8
  );


  buf
  g68
  (
    n93,
    n36
  );


  not
  g69
  (
    n76,
    n33
  );


  buf
  g70
  (
    n100,
    n24
  );


  not
  g71
  (
    n124,
    n33
  );


  not
  g72
  (
    n62,
    n37
  );


  buf
  g73
  (
    n108,
    n15
  );


  buf
  g74
  (
    n45,
    n21
  );


  buf
  g75
  (
    n101,
    n41
  );


  buf
  g76
  (
    n67,
    n13
  );


  not
  g77
  (
    n48,
    n11
  );


  buf
  g78
  (
    n63,
    n28
  );


  not
  g79
  (
    n89,
    n34
  );


  buf
  g80
  (
    n73,
    n14
  );


  not
  g81
  (
    n65,
    n31
  );


  not
  g82
  (
    KeyWire_0_15,
    n28
  );


  buf
  g83
  (
    n61,
    n23
  );


  not
  g84
  (
    KeyWire_0_4,
    n12
  );


  buf
  g85
  (
    n88,
    n7
  );


  buf
  g86
  (
    n84,
    n17
  );


  buf
  g87
  (
    n72,
    n12
  );


  not
  g88
  (
    n95,
    n16
  );


  buf
  g89
  (
    n113,
    n41
  );


  not
  g90
  (
    n60,
    n12
  );


  buf
  g91
  (
    n94,
    n28
  );


  nand
  g92
  (
    n86,
    n30,
    n35
  );


  nand
  g93
  (
    n125,
    n25,
    n39,
    n23,
    n15
  );


  and
  g94
  (
    n110,
    n39,
    n12,
    n21,
    n27
  );


  xnor
  g95
  (
    n117,
    n24,
    n8,
    n35,
    n39
  );


  nand
  g96
  (
    n74,
    n33,
    n26,
    n35,
    n24
  );


  nor
  g97
  (
    n105,
    n11,
    n37,
    n7,
    n22
  );


  xor
  g98
  (
    n111,
    n11,
    n22,
    n14,
    n40
  );


  xnor
  g99
  (
    n81,
    n17,
    n31,
    n28,
    n38
  );


  or
  g100
  (
    n54,
    n21,
    n14,
    n39,
    n13
  );


  xnor
  g101
  (
    n91,
    n22,
    n38,
    n40,
    n14
  );


  xnor
  g102
  (
    n79,
    n32,
    n27,
    n41,
    n16
  );


  nand
  g103
  (
    n80,
    n42,
    n30,
    n29,
    n15
  );


  nand
  g104
  (
    n121,
    n30,
    n26,
    n36,
    n10
  );


  nand
  g105
  (
    n123,
    n42,
    n24,
    n17,
    n13
  );


  or
  g106
  (
    n115,
    n34,
    n37,
    n9,
    n32
  );


  nand
  g107
  (
    n78,
    n9,
    n26,
    n25,
    n36
  );


  not
  g108
  (
    n157,
    n50
  );


  buf
  g109
  (
    n154,
    n42
  );


  not
  g110
  (
    n135,
    n46
  );


  not
  g111
  (
    n147,
    n45
  );


  not
  g112
  (
    n143,
    n49
  );


  buf
  g113
  (
    n140,
    n48
  );


  buf
  g114
  (
    n139,
    n48
  );


  buf
  g115
  (
    n145,
    n43
  );


  not
  g116
  (
    n129,
    n49
  );


  buf
  g117
  (
    n144,
    n45
  );


  not
  g118
  (
    n141,
    n48
  );


  buf
  g119
  (
    n146,
    n47
  );


  buf
  g120
  (
    n148,
    n44
  );


  buf
  g121
  (
    n131,
    n45
  );


  not
  g122
  (
    n133,
    n50
  );


  not
  g123
  (
    n130,
    n47
  );


  not
  g124
  (
    n149,
    n47
  );


  buf
  g125
  (
    n137,
    n45
  );


  buf
  g126
  (
    n156,
    n43
  );


  not
  g127
  (
    n142,
    n49
  );


  buf
  g128
  (
    n138,
    n49
  );


  not
  g129
  (
    n153,
    n46
  );


  buf
  g130
  (
    KeyWire_0_9,
    n44
  );


  not
  g131
  (
    n132,
    n42
  );


  buf
  g132
  (
    n136,
    n48
  );


  buf
  g133
  (
    n150,
    n46
  );


  buf
  g134
  (
    n155,
    n47
  );


  or
  g135
  (
    n134,
    n43,
    n44
  );


  or
  g136
  (
    n151,
    n44,
    n43,
    n46
  );


  xnor
  g137
  (
    n182,
    n132,
    n58,
    n63,
    n60
  );


  and
  g138
  (
    n171,
    n66,
    n135,
    n52,
    n64
  );


  nor
  g139
  (
    n161,
    n54,
    n133,
    n64,
    n66
  );


  xnor
  g140
  (
    n173,
    n131,
    n53,
    n57,
    n52
  );


  xnor
  g141
  (
    n163,
    n61,
    n69,
    n51,
    n67
  );


  or
  g142
  (
    n169,
    n51,
    n67,
    n61,
    n62
  );


  nand
  g143
  (
    n183,
    n64,
    n68,
    n60,
    n70
  );


  xor
  g144
  (
    n177,
    n131,
    n54,
    n62,
    n70
  );


  nor
  g145
  (
    n164,
    n135,
    n134,
    n68,
    n132
  );


  or
  g146
  (
    n158,
    n71,
    n68,
    n70,
    n56
  );


  xor
  g147
  (
    n166,
    n71,
    n57,
    n51,
    n129
  );


  nand
  g148
  (
    n165,
    n50,
    n65,
    n62,
    n52
  );


  nor
  g149
  (
    n181,
    n55,
    n60,
    n135,
    n58
  );


  xnor
  g150
  (
    n178,
    n69,
    n53,
    n66,
    n61
  );


  xor
  g151
  (
    n175,
    n130,
    n70,
    n59,
    n65
  );


  and
  g152
  (
    n176,
    n68,
    n53,
    n60,
    n130
  );


  nor
  g153
  (
    n167,
    n65,
    n51,
    n59
  );


  and
  g154
  (
    n174,
    n129,
    n69,
    n133
  );


  nand
  g155
  (
    n185,
    n129,
    n56,
    n131,
    n63
  );


  and
  g156
  (
    n170,
    n131,
    n53,
    n134,
    n133
  );


  and
  g157
  (
    KeyWire_0_12,
    n57,
    n55,
    n135,
    n56
  );


  and
  g158
  (
    n162,
    n59,
    n132,
    n62
  );


  xnor
  g159
  (
    n160,
    n130,
    n67,
    n64,
    n54
  );


  xnor
  g160
  (
    n159,
    n57,
    n67,
    n66,
    n134
  );


  xnor
  g161
  (
    n180,
    n134,
    n133,
    n54,
    n61
  );


  nand
  g162
  (
    n179,
    n129,
    n63,
    n55,
    n58
  );


  xor
  g163
  (
    n168,
    n56,
    n130,
    n55,
    n63
  );


  nor
  g164
  (
    n184,
    n50,
    n58,
    n52,
    n65
  );


  nor
  g165
  (
    n254,
    n148,
    n163,
    n168,
    n81
  );


  xnor
  g166
  (
    n258,
    n173,
    n173,
    n178,
    n172
  );


  nor
  g167
  (
    n274,
    n79,
    n182,
    n111,
    n89
  );


  nor
  g168
  (
    n212,
    n87,
    n156,
    n89,
    n170
  );


  xnor
  g169
  (
    n219,
    n112,
    n153,
    n87,
    n121
  );


  xor
  g170
  (
    n238,
    n120,
    n152,
    n112,
    n139
  );


  nand
  g171
  (
    n232,
    n144,
    n99,
    n120,
    n149
  );


  nor
  g172
  (
    n277,
    n161,
    n115,
    n174,
    n88
  );


  nand
  g173
  (
    n222,
    n73,
    n80,
    n96,
    n103
  );


  xnor
  g174
  (
    n214,
    n101,
    n158,
    n179,
    n115
  );


  nor
  g175
  (
    n264,
    n103,
    n105,
    n145,
    n152
  );


  or
  g176
  (
    n231,
    n98,
    n136,
    n177,
    n117
  );


  xnor
  g177
  (
    n253,
    n154,
    n97,
    n86
  );


  and
  g178
  (
    KeyWire_0_0,
    n140,
    n180,
    n107,
    n143
  );


  nand
  g179
  (
    n196,
    n182,
    n103,
    n117,
    n84
  );


  nand
  g180
  (
    n281,
    n119,
    n139,
    n147
  );


  or
  g181
  (
    n227,
    n105,
    n176,
    n86,
    n112
  );


  xor
  g182
  (
    n249,
    n106,
    n165,
    n82
  );


  nand
  g183
  (
    n201,
    n146,
    n98,
    n176,
    n150
  );


  and
  g184
  (
    n272,
    n138,
    n102,
    n77,
    n164
  );


  nand
  g185
  (
    n263,
    n108,
    n162,
    n145,
    n85
  );


  nand
  g186
  (
    n209,
    n179,
    n153,
    n109,
    n94
  );


  nand
  g187
  (
    n270,
    n161,
    n150,
    n162,
    n72
  );


  nand
  g188
  (
    n218,
    n159,
    n160,
    n153,
    n180
  );


  xnor
  g189
  (
    n210,
    n92,
    n89,
    n74,
    n72
  );


  nor
  g190
  (
    n248,
    n145,
    n182,
    n146,
    n148
  );


  xnor
  g191
  (
    n188,
    n85,
    n101,
    n117,
    n81
  );


  xnor
  g192
  (
    n273,
    n166,
    n175,
    n75,
    n172
  );


  nor
  g193
  (
    n204,
    n82,
    n141,
    n94,
    n97
  );


  xor
  g194
  (
    n192,
    n138,
    n178,
    n91,
    n161
  );


  or
  g195
  (
    n225,
    n159,
    n166,
    n110,
    n73
  );


  nor
  g196
  (
    n194,
    n106,
    n175,
    n87,
    n92
  );


  xnor
  g197
  (
    n260,
    n137,
    n162,
    n150,
    n177
  );


  xor
  g198
  (
    n241,
    n83,
    n142,
    n100,
    n136
  );


  or
  g199
  (
    n268,
    n72,
    n156,
    n92,
    n181
  );


  xor
  g200
  (
    n276,
    n90,
    n180,
    n111,
    n96
  );


  nor
  g201
  (
    n186,
    n109,
    n156,
    n171,
    n94
  );


  xnor
  g202
  (
    n213,
    n114,
    n82,
    n76,
    n153
  );


  and
  g203
  (
    n187,
    n155,
    n148,
    n168,
    n88
  );


  xnor
  g204
  (
    n266,
    n119,
    n149,
    n151,
    n177
  );


  xnor
  g205
  (
    n262,
    n144,
    n143,
    n171,
    n95
  );


  nor
  g206
  (
    n257,
    n90,
    n169,
    n101,
    n149
  );


  xnor
  g207
  (
    n269,
    n172,
    n166,
    n176,
    n136
  );


  nor
  g208
  (
    KeyWire_0_7,
    n82,
    n163,
    n78,
    n152
  );


  nor
  g209
  (
    n252,
    n173,
    n107,
    n119,
    n168
  );


  nand
  g210
  (
    KeyWire_0_5,
    n77,
    n90,
    n174,
    n169
  );


  xor
  g211
  (
    n195,
    n73,
    n167,
    n144,
    n179
  );


  nand
  g212
  (
    n189,
    n106,
    n109,
    n77,
    n118
  );


  or
  g213
  (
    n226,
    n71,
    n109,
    n142,
    n80
  );


  nand
  g214
  (
    n245,
    n147,
    n98,
    n117,
    n79
  );


  and
  g215
  (
    n234,
    n154,
    n175,
    n116,
    n157
  );


  nor
  g216
  (
    n221,
    n141,
    n115,
    n140,
    n163
  );


  nand
  g217
  (
    n230,
    n78,
    n101,
    n179,
    n151
  );


  xor
  g218
  (
    n200,
    n172,
    n149,
    n157,
    n99
  );


  or
  g219
  (
    n228,
    n83,
    n102,
    n137,
    n118
  );


  xnor
  g220
  (
    n207,
    n83,
    n151,
    n140,
    n74
  );


  and
  g221
  (
    n240,
    n154,
    n142,
    n168,
    n84
  );


  or
  g222
  (
    n216,
    n108,
    n151,
    n100,
    n141
  );


  nor
  g223
  (
    n265,
    n155,
    n85,
    n99,
    n116
  );


  nor
  g224
  (
    n236,
    n100,
    n157,
    n139,
    n114
  );


  nand
  g225
  (
    n244,
    n112,
    n110,
    n143,
    n93
  );


  or
  g226
  (
    n250,
    n103,
    n102,
    n177,
    n96
  );


  nand
  g227
  (
    n246,
    n110,
    n155,
    n152,
    n76
  );


  xor
  g228
  (
    n235,
    n72,
    n75,
    n175,
    n99
  );


  xnor
  g229
  (
    n255,
    n97,
    n166,
    n178,
    n78
  );


  nand
  g230
  (
    n197,
    n174,
    n137,
    n181,
    n83
  );


  nand
  g231
  (
    n267,
    n88,
    n143,
    n97,
    n79
  );


  nor
  g232
  (
    n243,
    n78,
    n119,
    n77,
    n167
  );


  nand
  g233
  (
    n278,
    n167,
    n174,
    n95,
    n160
  );


  nor
  g234
  (
    n261,
    n104,
    n107,
    n162,
    n155
  );


  nand
  g235
  (
    n220,
    n161,
    n138,
    n95,
    n181
  );


  and
  g236
  (
    n237,
    n176,
    n160,
    n111,
    n102
  );


  nand
  g237
  (
    n202,
    n105,
    n170,
    n164,
    n169
  );


  xnor
  g238
  (
    n205,
    n156,
    n147,
    n120,
    n74
  );


  xor
  g239
  (
    n271,
    n159,
    n142,
    n84,
    n154
  );


  nor
  g240
  (
    n198,
    n105,
    n171,
    n120,
    n71
  );


  and
  g241
  (
    n206,
    n93,
    n173,
    n171,
    n164
  );


  xor
  g242
  (
    n279,
    n159,
    n91,
    n165,
    n104
  );


  nor
  g243
  (
    n211,
    n140,
    n74,
    n108,
    n178
  );


  nor
  g244
  (
    n256,
    n76,
    n157,
    n75,
    n96
  );


  or
  g245
  (
    n259,
    n80,
    n111,
    n150,
    n107
  );


  or
  g246
  (
    n223,
    n139,
    n88,
    n113,
    n75
  );


  nor
  g247
  (
    n217,
    n116,
    n114,
    n169,
    n136
  );


  nor
  g248
  (
    n193,
    n170,
    n163,
    n113,
    n137
  );


  or
  g249
  (
    n275,
    n181,
    n91,
    n87,
    n180
  );


  nor
  g250
  (
    n280,
    n160,
    n73,
    n92,
    n93
  );


  and
  g251
  (
    n203,
    n114,
    n80,
    n167,
    n121
  );


  xor
  g252
  (
    n224,
    n95,
    n108,
    n81,
    n89
  );


  xor
  g253
  (
    n251,
    n138,
    n110,
    n146,
    n104
  );


  or
  g254
  (
    n233,
    n145,
    n76,
    n118
  );


  xnor
  g255
  (
    n247,
    n84,
    n113,
    n115,
    n116
  );


  nor
  g256
  (
    n199,
    n94,
    n106,
    n93,
    n100
  );


  or
  g257
  (
    n190,
    n165,
    n148,
    n98,
    n91
  );


  nor
  g258
  (
    n208,
    n104,
    n146,
    n141,
    n170
  );


  xor
  g259
  (
    n239,
    n81,
    n85,
    n113,
    n86
  );


  and
  g260
  (
    KeyWire_0_14,
    n164,
    n144,
    n90,
    n79
  );


  xor
  g261
  (
    n288,
    n123,
    n183,
    n182
  );


  or
  g262
  (
    n284,
    n127,
    n193,
    n20
  );


  and
  g263
  (
    n297,
    n123,
    n185,
    n184
  );


  or
  g264
  (
    n293,
    n202,
    n185,
    n192
  );


  nor
  g265
  (
    n300,
    n124,
    n122,
    n205
  );


  nor
  g266
  (
    n305,
    n124,
    n206,
    n127
  );


  and
  g267
  (
    n302,
    n19,
    n122,
    n198
  );


  xnor
  g268
  (
    n290,
    n126,
    n191,
    n123
  );


  and
  g269
  (
    n296,
    n126,
    n184,
    n18
  );


  or
  g270
  (
    n291,
    n18,
    n183,
    n185
  );


  or
  g271
  (
    n283,
    n20,
    n199,
    n197
  );


  nand
  g272
  (
    n289,
    n125,
    n183,
    n123
  );


  nand
  g273
  (
    n285,
    n122,
    n125
  );


  xnor
  g274
  (
    n294,
    n124,
    n200,
    n187
  );


  xnor
  g275
  (
    n299,
    n185,
    n127,
    n121
  );


  and
  g276
  (
    n292,
    n18,
    n20,
    n201
  );


  nand
  g277
  (
    n298,
    n127,
    n184,
    n19
  );


  xor
  g278
  (
    n303,
    n121,
    n189,
    n19
  );


  nor
  g279
  (
    n301,
    n209,
    n128,
    n126
  );


  and
  g280
  (
    n286,
    n20,
    n194,
    n128,
    n196
  );


  xnor
  g281
  (
    n287,
    n184,
    n190,
    n204,
    n207
  );


  nand
  g282
  (
    n295,
    n186,
    n188,
    n125,
    n203
  );


  or
  g283
  (
    n304,
    n183,
    n122,
    n18,
    n208
  );


  and
  g284
  (
    n282,
    n124,
    n126,
    n19,
    n195
  );


  and
  g285
  (
    n356,
    n282,
    n267,
    n228,
    n225
  );


  nand
  g286
  (
    n361,
    n212,
    n295,
    n260,
    n244
  );


  xor
  g287
  (
    n316,
    n237,
    n236,
    n269,
    n233
  );


  nand
  g288
  (
    n344,
    n265,
    n266,
    n255,
    n237
  );


  and
  g289
  (
    n354,
    n277,
    n268,
    n291,
    n252
  );


  or
  g290
  (
    KeyWire_0_2,
    n287,
    n244,
    n238,
    n299
  );


  and
  g291
  (
    n318,
    n249,
    n272,
    n218,
    n232
  );


  and
  g292
  (
    n339,
    n263,
    n262,
    n261,
    n235
  );


  xnor
  g293
  (
    n352,
    n233,
    n292,
    n240,
    n210
  );


  and
  g294
  (
    n322,
    n246,
    n257,
    n298
  );


  nand
  g295
  (
    n321,
    n284,
    n288,
    n258,
    n245
  );


  nor
  g296
  (
    n331,
    n253,
    n234,
    n219,
    n265
  );


  nand
  g297
  (
    n338,
    n239,
    n294,
    n297,
    n264
  );


  xor
  g298
  (
    n306,
    n288,
    n246,
    n276,
    n279
  );


  nor
  g299
  (
    n360,
    n271,
    n275,
    n280,
    n293
  );


  nand
  g300
  (
    KeyWire_0_13,
    n299,
    n290,
    n278,
    n266
  );


  nand
  g301
  (
    n310,
    n251,
    n223,
    n261,
    n249
  );


  xnor
  g302
  (
    n317,
    n248,
    n250,
    n286,
    n236
  );


  xor
  g303
  (
    n340,
    n280,
    n226,
    n250,
    n295
  );


  xor
  g304
  (
    n342,
    n245,
    n277,
    n267,
    n299
  );


  xnor
  g305
  (
    n328,
    n248,
    n215,
    n250,
    n247
  );


  nand
  g306
  (
    n319,
    n260,
    n262,
    n279,
    n294
  );


  xnor
  g307
  (
    n308,
    n270,
    n261,
    n262,
    n296
  );


  or
  g308
  (
    n357,
    n273,
    n251,
    n233,
    n257
  );


  nand
  g309
  (
    n332,
    n276,
    n259,
    n247
  );


  or
  g310
  (
    n329,
    n281,
    n235,
    n222,
    n270
  );


  xnor
  g311
  (
    n337,
    n231,
    n238,
    n294,
    n276
  );


  xor
  g312
  (
    n370,
    n253,
    n296,
    n281,
    n234
  );


  nor
  g313
  (
    n362,
    n258,
    n272,
    n267,
    n276
  );


  or
  g314
  (
    n348,
    n247,
    n284,
    n274,
    n292
  );


  nor
  g315
  (
    n312,
    n271,
    n245,
    n231,
    n254
  );


  xor
  g316
  (
    n315,
    n293,
    n257,
    n263,
    n253
  );


  xnor
  g317
  (
    n311,
    n236,
    n292,
    n244,
    n278
  );


  nand
  g318
  (
    n327,
    n300,
    n252,
    n279,
    n258
  );


  nand
  g319
  (
    n335,
    n282,
    n285,
    n242,
    n243
  );


  nand
  g320
  (
    n324,
    n231,
    n291,
    n289,
    n288
  );


  xor
  g321
  (
    n349,
    n216,
    n269,
    n268,
    n283
  );


  xor
  g322
  (
    n347,
    n240,
    n259,
    n256,
    n264
  );


  xor
  g323
  (
    n334,
    n286,
    n286,
    n217,
    n249
  );


  and
  g324
  (
    n369,
    n275,
    n284,
    n285,
    n234
  );


  nand
  g325
  (
    n325,
    n295,
    n298,
    n291,
    n255
  );


  and
  g326
  (
    n345,
    n295,
    n269,
    n263,
    n232
  );


  xor
  g327
  (
    n351,
    n239,
    n214,
    n227,
    n241
  );


  and
  g328
  (
    n368,
    n298,
    n274,
    n275,
    n293
  );


  and
  g329
  (
    n314,
    n273,
    n256,
    n259,
    n220
  );


  xnor
  g330
  (
    n336,
    n261,
    n221,
    n290,
    n271
  );


  and
  g331
  (
    n373,
    n289,
    n285,
    n268,
    n284
  );


  nand
  g332
  (
    n323,
    n293,
    n294,
    n211,
    n277
  );


  nor
  g333
  (
    n367,
    n256,
    n238,
    n230,
    n289
  );


  and
  g334
  (
    n363,
    n242,
    n296,
    n292
  );


  nand
  g335
  (
    n350,
    n240,
    n263,
    n269,
    n264
  );


  xnor
  g336
  (
    n372,
    n241,
    n246,
    n289,
    n273
  );


  xor
  g337
  (
    n346,
    n291,
    n287,
    n282
  );


  nand
  g338
  (
    KeyWire_0_8,
    n273,
    n265,
    n213,
    n283
  );


  or
  g339
  (
    n320,
    n262,
    n275,
    n290,
    n255
  );


  and
  g340
  (
    n364,
    n251,
    n266,
    n268,
    n254
  );


  nand
  g341
  (
    n330,
    n297,
    n267,
    n288,
    n280
  );


  nor
  g342
  (
    n333,
    n271,
    n278,
    n266,
    n286
  );


  and
  g343
  (
    n309,
    n232,
    n260,
    n239,
    n243
  );


  nor
  g344
  (
    n307,
    n285,
    n229,
    n241,
    n299
  );


  xnor
  g345
  (
    n365,
    n257,
    n297,
    n237,
    n248
  );


  xnor
  g346
  (
    n371,
    n279,
    n242,
    n287,
    n283
  );


  xor
  g347
  (
    n326,
    n265,
    n264,
    n297,
    n252
  );


  nand
  g348
  (
    n358,
    n270,
    n281,
    n258,
    n224
  );


  or
  g349
  (
    n355,
    n270,
    n274,
    n243,
    n282
  );


  nand
  g350
  (
    n341,
    n280,
    n272,
    n260,
    n235
  );


  nor
  g351
  (
    n353,
    n283,
    n272,
    n254,
    n278
  );


  xnor
  g352
  (
    n313,
    n290,
    n274,
    n277,
    n281
  );


  nand
  g353
  (
    n387,
    n365,
    n332,
    n344,
    n329
  );


  xor
  g354
  (
    n374,
    n366,
    n363,
    n304,
    n319
  );


  or
  g355
  (
    n388,
    n304,
    n351,
    n373,
    n354
  );


  xor
  g356
  (
    n375,
    n346,
    n300,
    n350,
    n348
  );


  xnor
  g357
  (
    n396,
    n303,
    n317,
    n343,
    n304
  );


  or
  g358
  (
    KeyWire_0_3,
    n355,
    n301,
    n320,
    n328
  );


  xnor
  g359
  (
    n385,
    n342,
    n303,
    n324,
    n307
  );


  xor
  g360
  (
    n393,
    n358,
    n326,
    n335,
    n128
  );


  xor
  g361
  (
    n380,
    n341,
    n311,
    n340,
    n305
  );


  nor
  g362
  (
    n382,
    n314,
    n327,
    n301,
    n313
  );


  xnor
  g363
  (
    n384,
    n300,
    n306,
    n347,
    n337
  );


  nand
  g364
  (
    n376,
    n361,
    n356,
    n334,
    n302
  );


  xnor
  g365
  (
    n377,
    n300,
    n322,
    n318,
    n301
  );


  nor
  g366
  (
    n386,
    n304,
    n325,
    n352,
    n305
  );


  xor
  g367
  (
    n392,
    n370,
    n308,
    n364,
    n302
  );


  and
  g368
  (
    n394,
    n305,
    n331,
    n333,
    n362
  );


  xnor
  g369
  (
    n381,
    n353,
    n330,
    n316,
    n360
  );


  and
  g370
  (
    n390,
    n371,
    n310,
    n357,
    n338
  );


  and
  g371
  (
    n383,
    n368,
    n359,
    n303,
    n309
  );


  or
  g372
  (
    n379,
    n345,
    n303,
    n336,
    n321
  );


  nor
  g373
  (
    n395,
    n315,
    n301,
    n339,
    n302
  );


  nor
  g374
  (
    n389,
    n302,
    n312,
    n367,
    n372
  );


  and
  g375
  (
    n391,
    n305,
    n323,
    n369,
    n349
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n215,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n107,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n366,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n378,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n102,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n242,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n119,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n229,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n343,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n152,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n44,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n97,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n172,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n359,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n191,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n43,
    KeyNOTWire_0_15
  );


endmodule

