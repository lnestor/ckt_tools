

module Stat_1000_203
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n550,
  n622,
  n656,
  n640,
  n637,
  n620,
  n616,
  n638,
  n652,
  n641,
  n643,
  n621,
  n615,
  n624,
  n626,
  n639,
  n631,
  n979,
  n1008,
  n1000,
  n1006,
  n1013,
  n1025,
  n1016,
  n1022,
  n1024,
  n1011,
  n1021,
  n1012,
  n1032,
  n1031,
  n1030,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n550;output n622;output n656;output n640;output n637;output n620;output n616;output n638;output n652;output n641;output n643;output n621;output n615;output n624;output n626;output n639;output n631;output n979;output n1008;output n1000;output n1006;output n1013;output n1025;output n1016;output n1022;output n1024;output n1011;output n1021;output n1012;output n1032;output n1031;output n1030;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n617;wire n618;wire n619;wire n623;wire n625;wire n627;wire n628;wire n629;wire n630;wire n632;wire n633;wire n634;wire n635;wire n636;wire n642;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n653;wire n654;wire n655;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1007;wire n1009;wire n1010;wire n1014;wire n1015;wire n1017;wire n1018;wire n1019;wire n1020;wire n1023;wire n1026;wire n1027;wire n1028;wire n1029;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n41,
    n14
  );


  buf
  g1
  (
    n91,
    n9
  );


  buf
  g2
  (
    n40,
    n15
  );


  not
  g3
  (
    n83,
    n19
  );


  not
  g4
  (
    n68,
    n19
  );


  not
  g5
  (
    n62,
    n16
  );


  not
  g6
  (
    n48,
    n5
  );


  buf
  g7
  (
    n102,
    n11
  );


  buf
  g8
  (
    n38,
    n17
  );


  buf
  g9
  (
    n101,
    n20
  );


  buf
  g10
  (
    n100,
    n16
  );


  buf
  g11
  (
    n37,
    n6
  );


  not
  g12
  (
    n35,
    n12
  );


  buf
  g13
  (
    n36,
    n9
  );


  buf
  g14
  (
    n34,
    n19
  );


  not
  g15
  (
    n33,
    n21
  );


  not
  g16
  (
    n65,
    n20
  );


  not
  g17
  (
    n58,
    n17
  );


  not
  g18
  (
    n80,
    n8
  );


  buf
  g19
  (
    n39,
    n8
  );


  not
  g20
  (
    n97,
    n5
  );


  not
  g21
  (
    n77,
    n8
  );


  buf
  g22
  (
    n44,
    n11
  );


  buf
  g23
  (
    n94,
    n11
  );


  buf
  g24
  (
    n50,
    n21
  );


  buf
  g25
  (
    n89,
    n22
  );


  buf
  g26
  (
    n54,
    n17
  );


  not
  g27
  (
    n76,
    n4
  );


  not
  g28
  (
    n43,
    n7
  );


  buf
  g29
  (
    n99,
    n14
  );


  not
  g30
  (
    n66,
    n7
  );


  not
  g31
  (
    n86,
    n4
  );


  buf
  g32
  (
    n84,
    n10
  );


  buf
  g33
  (
    n90,
    n7
  );


  not
  g34
  (
    n63,
    n5
  );


  not
  g35
  (
    n64,
    n13
  );


  buf
  g36
  (
    n42,
    n17
  );


  buf
  g37
  (
    n46,
    n20
  );


  not
  g38
  (
    n98,
    n16
  );


  not
  g39
  (
    n78,
    n6
  );


  buf
  g40
  (
    n69,
    n2
  );


  buf
  g41
  (
    n71,
    n5
  );


  not
  g42
  (
    n74,
    n16
  );


  not
  g43
  (
    n67,
    n8
  );


  not
  g44
  (
    n45,
    n6
  );


  not
  g45
  (
    n49,
    n15
  );


  not
  g46
  (
    n47,
    n19
  );


  not
  g47
  (
    n85,
    n6
  );


  buf
  g48
  (
    n72,
    n12
  );


  not
  g49
  (
    n73,
    n22
  );


  buf
  g50
  (
    n51,
    n13
  );


  not
  g51
  (
    n53,
    n13
  );


  not
  g52
  (
    n95,
    n18
  );


  not
  g53
  (
    n82,
    n3
  );


  buf
  g54
  (
    n81,
    n20
  );


  not
  g55
  (
    n87,
    n14
  );


  not
  g56
  (
    n70,
    n4
  );


  buf
  g57
  (
    n59,
    n13
  );


  not
  g58
  (
    n104,
    n10
  );


  not
  g59
  (
    n56,
    n14
  );


  buf
  g60
  (
    n61,
    n12
  );


  buf
  g61
  (
    n103,
    n18
  );


  not
  g62
  (
    n96,
    n10
  );


  not
  g63
  (
    n57,
    n15
  );


  not
  g64
  (
    n93,
    n1
  );


  not
  g65
  (
    n55,
    n11
  );


  not
  g66
  (
    n79,
    n21
  );


  buf
  g67
  (
    n75,
    n9
  );


  not
  g68
  (
    n88,
    n15
  );


  buf
  g69
  (
    n52,
    n22
  );


  xnor
  g70
  (
    n60,
    n18,
    n18,
    n10,
    n9
  );


  xor
  g71
  (
    n92,
    n4,
    n12,
    n21,
    n7
  );


  buf
  g72
  (
    n196,
    n54
  );


  buf
  g73
  (
    n223,
    n63
  );


  not
  g74
  (
    n140,
    n49
  );


  buf
  g75
  (
    n216,
    n64
  );


  not
  g76
  (
    n284,
    n38
  );


  buf
  g77
  (
    n229,
    n34
  );


  buf
  g78
  (
    n277,
    n75
  );


  buf
  g79
  (
    n181,
    n38
  );


  buf
  g80
  (
    n156,
    n75
  );


  not
  g81
  (
    n226,
    n72
  );


  buf
  g82
  (
    n250,
    n46
  );


  buf
  g83
  (
    n221,
    n67
  );


  buf
  g84
  (
    n153,
    n63
  );


  not
  g85
  (
    n213,
    n63
  );


  buf
  g86
  (
    n279,
    n65
  );


  buf
  g87
  (
    n139,
    n59
  );


  not
  g88
  (
    n272,
    n73
  );


  not
  g89
  (
    n105,
    n70
  );


  not
  g90
  (
    n182,
    n56
  );


  not
  g91
  (
    n234,
    n71
  );


  buf
  g92
  (
    n138,
    n66
  );


  not
  g93
  (
    n188,
    n53
  );


  not
  g94
  (
    n168,
    n40
  );


  buf
  g95
  (
    n290,
    n37
  );


  not
  g96
  (
    n256,
    n48
  );


  buf
  g97
  (
    n253,
    n64
  );


  buf
  g98
  (
    n283,
    n35
  );


  not
  g99
  (
    n200,
    n65
  );


  buf
  g100
  (
    n254,
    n41
  );


  not
  g101
  (
    n113,
    n40
  );


  not
  g102
  (
    n195,
    n58
  );


  buf
  g103
  (
    n151,
    n39
  );


  not
  g104
  (
    n165,
    n47
  );


  not
  g105
  (
    n117,
    n73
  );


  buf
  g106
  (
    n269,
    n62
  );


  buf
  g107
  (
    n133,
    n50
  );


  not
  g108
  (
    n162,
    n68
  );


  buf
  g109
  (
    n131,
    n47
  );


  buf
  g110
  (
    n237,
    n78
  );


  not
  g111
  (
    n172,
    n62
  );


  not
  g112
  (
    n194,
    n59
  );


  buf
  g113
  (
    n235,
    n60
  );


  not
  g114
  (
    n210,
    n58
  );


  not
  g115
  (
    n218,
    n71
  );


  buf
  g116
  (
    n144,
    n68
  );


  buf
  g117
  (
    n110,
    n70
  );


  not
  g118
  (
    n289,
    n65
  );


  buf
  g119
  (
    n288,
    n71
  );


  buf
  g120
  (
    n246,
    n52
  );


  not
  g121
  (
    n108,
    n68
  );


  not
  g122
  (
    n219,
    n70
  );


  not
  g123
  (
    n189,
    n66
  );


  not
  g124
  (
    n285,
    n36
  );


  not
  g125
  (
    n228,
    n61
  );


  not
  g126
  (
    n201,
    n75
  );


  not
  g127
  (
    n206,
    n35
  );


  buf
  g128
  (
    n192,
    n51
  );


  not
  g129
  (
    n255,
    n37
  );


  buf
  g130
  (
    n114,
    n54
  );


  buf
  g131
  (
    n119,
    n76
  );


  not
  g132
  (
    n115,
    n50
  );


  not
  g133
  (
    n152,
    n41
  );


  buf
  g134
  (
    n247,
    n46
  );


  not
  g135
  (
    n170,
    n34
  );


  not
  g136
  (
    n106,
    n43
  );


  not
  g137
  (
    n273,
    n52
  );


  not
  g138
  (
    n262,
    n35
  );


  buf
  g139
  (
    n186,
    n66
  );


  not
  g140
  (
    n251,
    n62
  );


  not
  g141
  (
    n123,
    n62
  );


  buf
  g142
  (
    n267,
    n42
  );


  buf
  g143
  (
    n160,
    n33
  );


  buf
  g144
  (
    n190,
    n78
  );


  buf
  g145
  (
    n124,
    n40
  );


  not
  g146
  (
    n177,
    n67
  );


  not
  g147
  (
    n281,
    n79
  );


  buf
  g148
  (
    n149,
    n70
  );


  buf
  g149
  (
    n161,
    n64
  );


  not
  g150
  (
    n159,
    n77
  );


  buf
  g151
  (
    n282,
    n40
  );


  not
  g152
  (
    n164,
    n46
  );


  not
  g153
  (
    n230,
    n69
  );


  buf
  g154
  (
    n180,
    n37
  );


  not
  g155
  (
    n276,
    n36
  );


  buf
  g156
  (
    n122,
    n61
  );


  buf
  g157
  (
    n265,
    n59
  );


  buf
  g158
  (
    n109,
    n39
  );


  not
  g159
  (
    n154,
    n42
  );


  buf
  g160
  (
    n174,
    n55
  );


  buf
  g161
  (
    n214,
    n57
  );


  buf
  g162
  (
    n249,
    n44
  );


  not
  g163
  (
    n286,
    n56
  );


  not
  g164
  (
    n155,
    n57
  );


  buf
  g165
  (
    n121,
    n33
  );


  buf
  g166
  (
    n111,
    n69
  );


  buf
  g167
  (
    n143,
    n54
  );


  buf
  g168
  (
    n204,
    n48
  );


  not
  g169
  (
    n227,
    n74
  );


  not
  g170
  (
    n130,
    n56
  );


  not
  g171
  (
    n199,
    n58
  );


  not
  g172
  (
    n175,
    n41
  );


  not
  g173
  (
    n239,
    n58
  );


  buf
  g174
  (
    n211,
    n65
  );


  buf
  g175
  (
    n191,
    n78
  );


  buf
  g176
  (
    n187,
    n64
  );


  not
  g177
  (
    n112,
    n74
  );


  buf
  g178
  (
    n148,
    n45
  );


  buf
  g179
  (
    n236,
    n50
  );


  buf
  g180
  (
    n241,
    n56
  );


  buf
  g181
  (
    n163,
    n61
  );


  not
  g182
  (
    n193,
    n34
  );


  not
  g183
  (
    n127,
    n39
  );


  not
  g184
  (
    n268,
    n72
  );


  buf
  g185
  (
    n185,
    n59
  );


  buf
  g186
  (
    n260,
    n72
  );


  not
  g187
  (
    n135,
    n60
  );


  not
  g188
  (
    n176,
    n69
  );


  buf
  g189
  (
    n280,
    n77
  );


  buf
  g190
  (
    n274,
    n76
  );


  not
  g191
  (
    n134,
    n73
  );


  buf
  g192
  (
    n287,
    n75
  );


  buf
  g193
  (
    n157,
    n39
  );


  buf
  g194
  (
    n198,
    n55
  );


  buf
  g195
  (
    n118,
    n38
  );


  buf
  g196
  (
    n258,
    n73
  );


  not
  g197
  (
    n261,
    n36
  );


  not
  g198
  (
    n263,
    n42
  );


  not
  g199
  (
    n166,
    n55
  );


  buf
  g200
  (
    n145,
    n76
  );


  buf
  g201
  (
    n242,
    n35
  );


  not
  g202
  (
    n212,
    n63
  );


  buf
  g203
  (
    n183,
    n71
  );


  not
  g204
  (
    n184,
    n47
  );


  not
  g205
  (
    n128,
    n34
  );


  not
  g206
  (
    n203,
    n79
  );


  buf
  g207
  (
    n208,
    n78
  );


  buf
  g208
  (
    n142,
    n60
  );


  not
  g209
  (
    n270,
    n49
  );


  not
  g210
  (
    n120,
    n33
  );


  not
  g211
  (
    n179,
    n51
  );


  buf
  g212
  (
    n146,
    n61
  );


  not
  g213
  (
    n158,
    n53
  );


  buf
  g214
  (
    n173,
    n44
  );


  not
  g215
  (
    n126,
    n48
  );


  not
  g216
  (
    n107,
    n57
  );


  not
  g217
  (
    n264,
    n74
  );


  not
  g218
  (
    n178,
    n53
  );


  buf
  g219
  (
    n220,
    n77
  );


  buf
  g220
  (
    n125,
    n36
  );


  not
  g221
  (
    n243,
    n37
  );


  buf
  g222
  (
    n252,
    n66
  );


  buf
  g223
  (
    n238,
    n69
  );


  buf
  g224
  (
    n171,
    n76
  );


  buf
  g225
  (
    n244,
    n60
  );


  buf
  g226
  (
    n136,
    n38
  );


  not
  g227
  (
    n129,
    n41
  );


  not
  g228
  (
    n225,
    n74
  );


  not
  g229
  (
    n150,
    n43
  );


  not
  g230
  (
    n257,
    n47
  );


  not
  g231
  (
    n224,
    n72
  );


  not
  g232
  (
    n222,
    n48
  );


  buf
  g233
  (
    n275,
    n53
  );


  buf
  g234
  (
    n245,
    n45
  );


  not
  g235
  (
    n266,
    n33
  );


  not
  g236
  (
    n215,
    n43
  );


  not
  g237
  (
    n232,
    n67
  );


  buf
  g238
  (
    n132,
    n49
  );


  buf
  g239
  (
    n209,
    n49
  );


  buf
  g240
  (
    n248,
    n54
  );


  not
  g241
  (
    n207,
    n77
  );


  buf
  g242
  (
    n233,
    n46
  );


  buf
  g243
  (
    n231,
    n50
  );


  not
  g244
  (
    n205,
    n68
  );


  buf
  g245
  (
    n271,
    n67
  );


  not
  g246
  (
    n147,
    n51
  );


  not
  g247
  (
    n137,
    n57
  );


  not
  g248
  (
    n202,
    n52
  );


  not
  g249
  (
    n217,
    n51
  );


  not
  g250
  (
    n240,
    n44
  );


  buf
  g251
  (
    n259,
    n45
  );


  not
  g252
  (
    n197,
    n52
  );


  buf
  g253
  (
    n141,
    n45
  );


  buf
  g254
  (
    n278,
    n42
  );


  buf
  g255
  (
    n167,
    n44
  );


  buf
  g256
  (
    n116,
    n55
  );


  buf
  g257
  (
    n169,
    n43
  );


  buf
  g258
  (
    n338,
    n272
  );


  not
  g259
  (
    n349,
    n207
  );


  buf
  g260
  (
    n454,
    n98
  );


  not
  g261
  (
    n490,
    n80
  );


  not
  g262
  (
    n325,
    n105
  );


  not
  g263
  (
    n361,
    n189
  );


  buf
  g264
  (
    n434,
    n121
  );


  buf
  g265
  (
    n386,
    n164
  );


  buf
  g266
  (
    n462,
    n209
  );


  not
  g267
  (
    n380,
    n268
  );


  not
  g268
  (
    n491,
    n149
  );


  buf
  g269
  (
    n368,
    n194
  );


  buf
  g270
  (
    n427,
    n164
  );


  buf
  g271
  (
    n296,
    n144
  );


  not
  g272
  (
    n464,
    n272
  );


  not
  g273
  (
    n308,
    n171
  );


  not
  g274
  (
    n298,
    n239
  );


  buf
  g275
  (
    n399,
    n128
  );


  buf
  g276
  (
    n517,
    n229
  );


  buf
  g277
  (
    n457,
    n224
  );


  not
  g278
  (
    n404,
    n85
  );


  not
  g279
  (
    n449,
    n211
  );


  not
  g280
  (
    n385,
    n288
  );


  buf
  g281
  (
    n421,
    n175
  );


  buf
  g282
  (
    n416,
    n264
  );


  buf
  g283
  (
    n415,
    n170
  );


  buf
  g284
  (
    n396,
    n264
  );


  not
  g285
  (
    n480,
    n105
  );


  xor
  g286
  (
    n329,
    n117,
    n135,
    n150,
    n268
  );


  or
  g287
  (
    n374,
    n166,
    n118,
    n254,
    n240
  );


  or
  g288
  (
    n514,
    n185,
    n83,
    n285,
    n216
  );


  xnor
  g289
  (
    n486,
    n213,
    n263,
    n220,
    n212
  );


  xor
  g290
  (
    n458,
    n157,
    n168,
    n273,
    n281
  );


  xor
  g291
  (
    n388,
    n92,
    n275,
    n267,
    n274
  );


  nor
  g292
  (
    n472,
    n120,
    n286,
    n222,
    n202
  );


  xor
  g293
  (
    n412,
    n211,
    n261,
    n270,
    n93
  );


  nand
  g294
  (
    n419,
    n225,
    n165,
    n212,
    n248
  );


  nor
  g295
  (
    n305,
    n200,
    n282,
    n231,
    n111
  );


  and
  g296
  (
    n381,
    n171,
    n206,
    n179,
    n152
  );


  nor
  g297
  (
    n377,
    n232,
    n154,
    n220,
    n186
  );


  nor
  g298
  (
    n451,
    n132,
    n130,
    n180,
    n262
  );


  nand
  g299
  (
    n442,
    n191,
    n209,
    n178,
    n221
  );


  or
  g300
  (
    n471,
    n225,
    n192,
    n114,
    n91
  );


  xnor
  g301
  (
    n301,
    n113,
    n134,
    n287,
    n85
  );


  xor
  g302
  (
    n468,
    n285,
    n198,
    n194,
    n163
  );


  or
  g303
  (
    n474,
    n196,
    n152,
    n167,
    n226
  );


  xnor
  g304
  (
    n467,
    n116,
    n288,
    n139,
    n236
  );


  nand
  g305
  (
    n352,
    n216,
    n231,
    n154,
    n241
  );


  or
  g306
  (
    n379,
    n227,
    n186,
    n125,
    n163
  );


  nand
  g307
  (
    n513,
    n273,
    n180,
    n107,
    n199
  );


  nand
  g308
  (
    n369,
    n251,
    n218,
    n147,
    n124
  );


  nand
  g309
  (
    n346,
    n220,
    n217,
    n219,
    n157
  );


  xor
  g310
  (
    n433,
    n145,
    n134,
    n215,
    n148
  );


  xnor
  g311
  (
    n481,
    n258,
    n227,
    n214,
    n156
  );


  or
  g312
  (
    n351,
    n230,
    n184,
    n108,
    n208
  );


  and
  g313
  (
    n402,
    n121,
    n171,
    n149
  );


  xor
  g314
  (
    n477,
    n108,
    n218,
    n89,
    n169
  );


  nor
  g315
  (
    n487,
    n190,
    n162,
    n133,
    n112
  );


  and
  g316
  (
    n340,
    n247,
    n251,
    n266,
    n155
  );


  or
  g317
  (
    n339,
    n249,
    n90,
    n206,
    n137
  );


  or
  g318
  (
    n297,
    n178,
    n258,
    n105,
    n123
  );


  and
  g319
  (
    n398,
    n126,
    n110,
    n225
  );


  xnor
  g320
  (
    n510,
    n282,
    n258,
    n135,
    n259
  );


  and
  g321
  (
    n341,
    n247,
    n130,
    n174,
    n279
  );


  nand
  g322
  (
    n494,
    n140,
    n256,
    n187,
    n181
  );


  xor
  g323
  (
    n364,
    n245,
    n258,
    n242,
    n170
  );


  xor
  g324
  (
    n366,
    n269,
    n167,
    n82,
    n286
  );


  or
  g325
  (
    n470,
    n109,
    n252,
    n106,
    n84
  );


  nand
  g326
  (
    n327,
    n131,
    n275,
    n181,
    n215
  );


  nand
  g327
  (
    n429,
    n99,
    n82,
    n111,
    n184
  );


  xnor
  g328
  (
    n485,
    n200,
    n90,
    n158,
    n252
  );


  xor
  g329
  (
    n445,
    n127,
    n238,
    n138,
    n212
  );


  xor
  g330
  (
    n293,
    n254,
    n172,
    n263,
    n214
  );


  nand
  g331
  (
    n420,
    n264,
    n250,
    n184,
    n203
  );


  nor
  g332
  (
    n303,
    n148,
    n137,
    n142,
    n160
  );


  and
  g333
  (
    n432,
    n273,
    n153,
    n186,
    n84
  );


  xnor
  g334
  (
    n370,
    n198,
    n240,
    n280,
    n284
  );


  nand
  g335
  (
    n418,
    n143,
    n87,
    n129,
    n280
  );


  xnor
  g336
  (
    n410,
    n150,
    n83,
    n94,
    n114
  );


  nor
  g337
  (
    n446,
    n159,
    n199,
    n140,
    n182
  );


  or
  g338
  (
    n373,
    n119,
    n234,
    n225,
    n249
  );


  and
  g339
  (
    n306,
    n155,
    n245,
    n233,
    n195
  );


  or
  g340
  (
    n359,
    n133,
    n207,
    n289,
    n161
  );


  xnor
  g341
  (
    n372,
    n159,
    n120,
    n243,
    n228
  );


  and
  g342
  (
    n392,
    n281,
    n196,
    n213,
    n243
  );


  nand
  g343
  (
    n356,
    n276,
    n88,
    n132,
    n123
  );


  xnor
  g344
  (
    n319,
    n173,
    n250,
    n281,
    n120
  );


  and
  g345
  (
    n318,
    n213,
    n121,
    n232,
    n277
  );


  nand
  g346
  (
    n406,
    n118,
    n137,
    n90,
    n132
  );


  nand
  g347
  (
    n466,
    n205,
    n80,
    n237,
    n261
  );


  and
  g348
  (
    n507,
    n261,
    n217,
    n229,
    n277
  );


  nor
  g349
  (
    n300,
    n265,
    n274,
    n281,
    n257
  );


  xor
  g350
  (
    n417,
    n242,
    n264,
    n219,
    n216
  );


  xor
  g351
  (
    n328,
    n202,
    n189,
    n150,
    n149
  );


  or
  g352
  (
    n413,
    n214,
    n112,
    n176,
    n204
  );


  nand
  g353
  (
    n501,
    n223,
    n97,
    n252,
    n128
  );


  or
  g354
  (
    n342,
    n130,
    n157,
    n238,
    n197
  );


  or
  g355
  (
    n394,
    n126,
    n154,
    n249,
    n149
  );


  nand
  g356
  (
    n314,
    n106,
    n94,
    n211,
    n125
  );


  xor
  g357
  (
    n294,
    n110,
    n98,
    n164,
    n82
  );


  xor
  g358
  (
    n322,
    n245,
    n271,
    n199
  );


  and
  g359
  (
    n292,
    n266,
    n108,
    n253,
    n129
  );


  xnor
  g360
  (
    n358,
    n80,
    n93,
    n280,
    n250
  );


  nand
  g361
  (
    n335,
    n269,
    n96,
    n92,
    n197
  );


  xor
  g362
  (
    n321,
    n205,
    n165,
    n204,
    n162
  );


  or
  g363
  (
    n515,
    n162,
    n113,
    n129,
    n145
  );


  xor
  g364
  (
    n334,
    n263,
    n172,
    n202,
    n242
  );


  and
  g365
  (
    n407,
    n167,
    n141,
    n117,
    n289
  );


  or
  g366
  (
    n307,
    n254,
    n156,
    n183,
    n142
  );


  xor
  g367
  (
    n426,
    n95,
    n262,
    n176,
    n89
  );


  nor
  g368
  (
    n483,
    n236,
    n127,
    n224,
    n215
  );


  nand
  g369
  (
    n409,
    n231,
    n210,
    n271,
    n246
  );


  nor
  g370
  (
    n475,
    n205,
    n157,
    n244,
    n235
  );


  or
  g371
  (
    n465,
    n277,
    n211,
    n253,
    n250
  );


  xnor
  g372
  (
    n291,
    n134,
    n177,
    n228,
    n181
  );


  nor
  g373
  (
    n405,
    n213,
    n176,
    n147,
    n83
  );


  and
  g374
  (
    n367,
    n232,
    n216,
    n270
  );


  nand
  g375
  (
    n389,
    n161,
    n166,
    n153,
    n123
  );


  xnor
  g376
  (
    n363,
    n181,
    n151,
    n133,
    n201
  );


  nand
  g377
  (
    n503,
    n159,
    n139,
    n91,
    n146
  );


  or
  g378
  (
    n493,
    n219,
    n239,
    n185,
    n283
  );


  nand
  g379
  (
    n347,
    n136,
    n207,
    n197,
    n252
  );


  xor
  g380
  (
    n295,
    n284,
    n247,
    n248,
    n173
  );


  and
  g381
  (
    n443,
    n255,
    n151,
    n91,
    n210
  );


  nor
  g382
  (
    n505,
    n128,
    n248,
    n273,
    n203
  );


  xnor
  g383
  (
    n425,
    n162,
    n97,
    n239,
    n210
  );


  and
  g384
  (
    n344,
    n268,
    n166,
    n109,
    n283
  );


  xor
  g385
  (
    n400,
    n175,
    n197,
    n87,
    n231
  );


  xnor
  g386
  (
    n343,
    n266,
    n138,
    n272,
    n148
  );


  xnor
  g387
  (
    n489,
    n173,
    n90,
    n253,
    n230
  );


  xor
  g388
  (
    n492,
    n166,
    n165,
    n175,
    n170
  );


  nand
  g389
  (
    n350,
    n289,
    n190,
    n240,
    n127
  );


  nor
  g390
  (
    n383,
    n182,
    n283,
    n191,
    n256
  );


  xnor
  g391
  (
    n313,
    n188,
    n251,
    n164,
    n98
  );


  and
  g392
  (
    n357,
    n285,
    n265,
    n195,
    n95
  );


  xnor
  g393
  (
    n508,
    n269,
    n140,
    n236,
    n125
  );


  nand
  g394
  (
    n509,
    n112,
    n262,
    n278,
    n122
  );


  and
  g395
  (
    n378,
    n119,
    n218,
    n222,
    n247
  );


  xor
  g396
  (
    n430,
    n106,
    n260,
    n145,
    n238
  );


  xnor
  g397
  (
    n309,
    n208,
    n195,
    n259,
    n152
  );


  or
  g398
  (
    n436,
    n141,
    n208,
    n88,
    n260
  );


  or
  g399
  (
    n460,
    n141,
    n159,
    n185,
    n94
  );


  nand
  g400
  (
    n316,
    n99,
    n155,
    n108,
    n86
  );


  xnor
  g401
  (
    n362,
    n119,
    n86,
    n111,
    n263
  );


  and
  g402
  (
    n326,
    n278,
    n160,
    n212,
    n163
  );


  xnor
  g403
  (
    n497,
    n287,
    n168,
    n260,
    n232
  );


  nand
  g404
  (
    n384,
    n85,
    n81,
    n189,
    n287
  );


  xnor
  g405
  (
    n516,
    n142,
    n114,
    n185,
    n175
  );


  and
  g406
  (
    n302,
    n229,
    n98,
    n118,
    n122
  );


  or
  g407
  (
    n453,
    n131,
    n153,
    n201,
    n272
  );


  and
  g408
  (
    n304,
    n158,
    n173,
    n99,
    n182
  );


  xor
  g409
  (
    n376,
    n92,
    n126,
    n191,
    n113
  );


  xnor
  g410
  (
    n310,
    n81,
    n84,
    n223,
    n174
  );


  xnor
  g411
  (
    n439,
    n97,
    n100,
    n275,
    n143
  );


  xor
  g412
  (
    n324,
    n190,
    n84,
    n139,
    n244
  );


  and
  g413
  (
    n437,
    n158,
    n282,
    n136,
    n246
  );


  nor
  g414
  (
    n484,
    n246,
    n80,
    n187,
    n186
  );


  xnor
  g415
  (
    n375,
    n161,
    n177,
    n183,
    n286
  );


  xor
  g416
  (
    n441,
    n260,
    n183,
    n136,
    n178
  );


  and
  g417
  (
    n469,
    n191,
    n203,
    n178,
    n276
  );


  nor
  g418
  (
    n428,
    n163,
    n116,
    n93,
    n82
  );


  xnor
  g419
  (
    n431,
    n205,
    n248,
    n122,
    n237
  );


  xor
  g420
  (
    n337,
    n112,
    n274,
    n176,
    n168
  );


  or
  g421
  (
    n512,
    n198,
    n279,
    n244,
    n223
  );


  xor
  g422
  (
    n411,
    n141,
    n193,
    n243,
    n192
  );


  xnor
  g423
  (
    n479,
    n119,
    n276,
    n115,
    n184
  );


  nand
  g424
  (
    n482,
    n196,
    n135,
    n218,
    n131
  );


  xor
  g425
  (
    n456,
    n246,
    n96,
    n174,
    n160
  );


  nand
  g426
  (
    n511,
    n196,
    n288,
    n245,
    n267
  );


  nand
  g427
  (
    n382,
    n132,
    n138,
    n255,
    n267
  );


  and
  g428
  (
    n391,
    n279,
    n237,
    n137,
    n189
  );


  or
  g429
  (
    n390,
    n279,
    n148,
    n115,
    n128
  );


  or
  g430
  (
    n414,
    n187,
    n194,
    n215,
    n124
  );


  xnor
  g431
  (
    n403,
    n95,
    n204,
    n221,
    n188
  );


  and
  g432
  (
    n395,
    n249,
    n282,
    n115,
    n79
  );


  nand
  g433
  (
    n447,
    n156,
    n257,
    n129,
    n174
  );


  and
  g434
  (
    n498,
    n97,
    n105,
    n123,
    n136
  );


  or
  g435
  (
    n488,
    n193,
    n242,
    n114,
    n217
  );


  and
  g436
  (
    n435,
    n117,
    n224,
    n111,
    n251
  );


  nor
  g437
  (
    n355,
    n235,
    n190,
    n86,
    n152
  );


  or
  g438
  (
    n463,
    n241,
    n130,
    n228,
    n193
  );


  xnor
  g439
  (
    n299,
    n221,
    n262,
    n126,
    n256
  );


  nor
  g440
  (
    n478,
    n161,
    n131,
    n83,
    n203
  );


  xnor
  g441
  (
    n336,
    n88,
    n287,
    n169,
    n210
  );


  xor
  g442
  (
    n353,
    n233,
    n187,
    n86,
    n115
  );


  nand
  g443
  (
    n320,
    n100,
    n234,
    n142,
    n94
  );


  or
  g444
  (
    n504,
    n261,
    n234,
    n107,
    n116
  );


  nor
  g445
  (
    n459,
    n278,
    n202,
    n155,
    n228
  );


  nand
  g446
  (
    n444,
    n95,
    n199,
    n200,
    n234
  );


  and
  g447
  (
    n499,
    n284,
    n217,
    n167,
    n214
  );


  and
  g448
  (
    n496,
    n285,
    n280,
    n172,
    n222
  );


  xor
  g449
  (
    n330,
    n233,
    n198,
    n237,
    n206
  );


  nor
  g450
  (
    n397,
    n256,
    n150,
    n269,
    n177
  );


  or
  g451
  (
    n424,
    n89,
    n89,
    n156,
    n192
  );


  nand
  g452
  (
    n365,
    n99,
    n233,
    n107,
    n146
  );


  nand
  g453
  (
    n495,
    n183,
    n268,
    n227,
    n220
  );


  nor
  g454
  (
    n438,
    n201,
    n79,
    n92,
    n134
  );


  nand
  g455
  (
    n311,
    n81,
    n91,
    n139,
    n209
  );


  or
  g456
  (
    n371,
    n219,
    n271,
    n201,
    n179
  );


  xor
  g457
  (
    n450,
    n170,
    n172,
    n124,
    n188
  );


  nand
  g458
  (
    n333,
    n200,
    n106,
    n182,
    n226
  );


  nor
  g459
  (
    n440,
    n127,
    n276,
    n153,
    n259
  );


  xor
  g460
  (
    n401,
    n288,
    n122,
    n154,
    n87
  );


  nand
  g461
  (
    n452,
    n208,
    n144,
    n88,
    n147
  );


  nor
  g462
  (
    n354,
    n240,
    n143,
    n151
  );


  xnor
  g463
  (
    n506,
    n267,
    n124,
    n275,
    n144
  );


  or
  g464
  (
    n502,
    n116,
    n146,
    n235,
    n110
  );


  nor
  g465
  (
    n423,
    n206,
    n180,
    n169
  );


  or
  g466
  (
    n345,
    n192,
    n207,
    n179,
    n257
  );


  nor
  g467
  (
    n473,
    n257,
    n265,
    n284,
    n146
  );


  or
  g468
  (
    n387,
    n144,
    n277,
    n270,
    n117
  );


  or
  g469
  (
    n348,
    n243,
    n125,
    n235,
    n188
  );


  nor
  g470
  (
    n461,
    n209,
    n147,
    n239,
    n135
  );


  xnor
  g471
  (
    n323,
    n236,
    n118,
    n87,
    n81
  );


  nand
  g472
  (
    n331,
    n145,
    n244,
    n107,
    n113
  );


  and
  g473
  (
    n455,
    n238,
    n230,
    n177
  );


  and
  g474
  (
    n315,
    n93,
    n254,
    n195,
    n241
  );


  or
  g475
  (
    n500,
    n255,
    n283,
    n158,
    n168
  );


  nor
  g476
  (
    n448,
    n227,
    n194,
    n109,
    n133
  );


  or
  g477
  (
    n360,
    n179,
    n140,
    n169,
    n253
  );


  xor
  g478
  (
    n408,
    n241,
    n151,
    n286,
    n229
  );


  nand
  g479
  (
    n422,
    n266,
    n278,
    n121,
    n138
  );


  xnor
  g480
  (
    n317,
    n221,
    n96,
    n120,
    n274
  );


  xor
  g481
  (
    n476,
    n109,
    n193,
    n224,
    n222
  );


  xnor
  g482
  (
    n393,
    n259,
    n226,
    n160,
    n289
  );


  nor
  g483
  (
    n332,
    n265,
    n226,
    n255,
    n204
  );


  or
  g484
  (
    n312,
    n165,
    n85,
    n223,
    n96
  );


  buf
  g485
  (
    n547,
    n401
  );


  buf
  g486
  (
    n570,
    n295
  );


  not
  g487
  (
    n557,
    n292
  );


  not
  g488
  (
    n554,
    n485
  );


  nor
  g489
  (
    n533,
    n405,
    n406
  );


  xnor
  g490
  (
    n548,
    n344,
    n354,
    n316,
    n440
  );


  or
  g491
  (
    n528,
    n395,
    n412,
    n392,
    n384
  );


  nor
  g492
  (
    n560,
    n341,
    n375,
    n351,
    n389
  );


  nand
  g493
  (
    n546,
    n333,
    n298,
    n476,
    n414
  );


  xnor
  g494
  (
    n563,
    n457,
    n486,
    n449,
    n346
  );


  or
  g495
  (
    n550,
    n381,
    n368,
    n408,
    n294
  );


  xnor
  g496
  (
    n524,
    n312,
    n443,
    n420,
    n332
  );


  nand
  g497
  (
    n536,
    n437,
    n371,
    n398,
    n442
  );


  and
  g498
  (
    n559,
    n452,
    n355,
    n338,
    n369
  );


  and
  g499
  (
    n545,
    n478,
    n313,
    n309,
    n471
  );


  nand
  g500
  (
    n539,
    n446,
    n393,
    n422,
    n303
  );


  nand
  g501
  (
    n519,
    n315,
    n453,
    n349,
    n366
  );


  xnor
  g502
  (
    n543,
    n376,
    n320,
    n402,
    n424
  );


  nand
  g503
  (
    n525,
    n328,
    n467,
    n327,
    n466
  );


  nor
  g504
  (
    n555,
    n307,
    n318,
    n365,
    n324
  );


  nand
  g505
  (
    n542,
    n461,
    n435,
    n407,
    n374
  );


  nor
  g506
  (
    n556,
    n394,
    n329,
    n445,
    n396
  );


  xor
  g507
  (
    n562,
    n474,
    n441,
    n444,
    n310
  );


  nand
  g508
  (
    n537,
    n317,
    n464,
    n410,
    n431
  );


  xor
  g509
  (
    n531,
    n390,
    n308,
    n319,
    n339
  );


  nor
  g510
  (
    n569,
    n411,
    n475,
    n345,
    n304
  );


  xnor
  g511
  (
    n532,
    n300,
    n306,
    n387,
    n483
  );


  nand
  g512
  (
    n549,
    n469,
    n359,
    n334,
    n382
  );


  nand
  g513
  (
    n526,
    n472,
    n314,
    n348,
    n323
  );


  xor
  g514
  (
    n544,
    n372,
    n343,
    n330,
    n385
  );


  and
  g515
  (
    n566,
    n399,
    n347,
    n380,
    n409
  );


  nor
  g516
  (
    n538,
    n463,
    n311,
    n462,
    n356
  );


  xnor
  g517
  (
    n520,
    n415,
    n439,
    n326,
    n297
  );


  xnor
  g518
  (
    n567,
    n488,
    n425,
    n373,
    n379
  );


  xnor
  g519
  (
    n553,
    n403,
    n305,
    n477,
    n454
  );


  xnor
  g520
  (
    n568,
    n448,
    n352,
    n481,
    n299
  );


  xor
  g521
  (
    n530,
    n378,
    n342,
    n465,
    n426
  );


  or
  g522
  (
    n534,
    n337,
    n386,
    n302,
    n447
  );


  nand
  g523
  (
    n518,
    n450,
    n391,
    n357,
    n322
  );


  xor
  g524
  (
    n552,
    n388,
    n459,
    n423,
    n456
  );


  and
  g525
  (
    n541,
    n331,
    n336,
    n404,
    n479
  );


  xnor
  g526
  (
    n521,
    n416,
    n436,
    n480,
    n487
  );


  nand
  g527
  (
    n523,
    n360,
    n421,
    n484,
    n430
  );


  nor
  g528
  (
    n540,
    n301,
    n350,
    n361,
    n428
  );


  xor
  g529
  (
    n551,
    n468,
    n335,
    n353,
    n400
  );


  xnor
  g530
  (
    n564,
    n418,
    n362,
    n427,
    n417
  );


  and
  g531
  (
    n565,
    n434,
    n460,
    n429,
    n458
  );


  nor
  g532
  (
    n561,
    n364,
    n433,
    n291,
    n367
  );


  nand
  g533
  (
    n535,
    n482,
    n419,
    n293,
    n438
  );


  xor
  g534
  (
    n527,
    n377,
    n296,
    n432,
    n363
  );


  xor
  g535
  (
    n529,
    n451,
    n321,
    n325,
    n383
  );


  or
  g536
  (
    n558,
    n455,
    n397,
    n470,
    n358
  );


  xor
  g537
  (
    n522,
    n473,
    n370,
    n340,
    n413
  );


  buf
  g538
  (
    n579,
    n525
  );


  not
  g539
  (
    n594,
    n528
  );


  not
  g540
  (
    n595,
    n520
  );


  not
  g541
  (
    n576,
    n529
  );


  not
  g542
  (
    n572,
    n521
  );


  buf
  g543
  (
    n574,
    n530
  );


  not
  g544
  (
    n600,
    n523
  );


  not
  g545
  (
    n597,
    n522
  );


  not
  g546
  (
    n580,
    n522
  );


  not
  g547
  (
    n591,
    n527
  );


  buf
  g548
  (
    n577,
    n520
  );


  not
  g549
  (
    n585,
    n530
  );


  buf
  g550
  (
    n582,
    n527
  );


  not
  g551
  (
    n587,
    n530
  );


  not
  g552
  (
    n599,
    n518
  );


  buf
  g553
  (
    n584,
    n529
  );


  not
  g554
  (
    n601,
    n521
  );


  not
  g555
  (
    n596,
    n528
  );


  buf
  g556
  (
    n589,
    n529
  );


  not
  g557
  (
    n588,
    n524
  );


  buf
  g558
  (
    n598,
    n519
  );


  buf
  g559
  (
    n583,
    n525
  );


  buf
  g560
  (
    n581,
    n523
  );


  buf
  g561
  (
    n593,
    n526
  );


  buf
  g562
  (
    n590,
    n526
  );


  and
  g563
  (
    n592,
    n519,
    n529,
    n524
  );


  xnor
  g564
  (
    n578,
    n528,
    n521,
    n527,
    n530
  );


  nand
  g565
  (
    n573,
    n518,
    n520,
    n523,
    n526
  );


  and
  g566
  (
    n571,
    n525,
    n520,
    n524,
    n528
  );


  and
  g567
  (
    n586,
    n524,
    n527,
    n522,
    n525
  );


  nand
  g568
  (
    n575,
    n523,
    n526,
    n521,
    n522
  );


  not
  g569
  (
    n605,
    n535
  );


  not
  g570
  (
    n603,
    n533
  );


  buf
  g571
  (
    n608,
    n571
  );


  buf
  g572
  (
    n604,
    n532
  );


  buf
  g573
  (
    n607,
    n532
  );


  buf
  g574
  (
    n602,
    n535
  );


  nand
  g575
  (
    n610,
    n574,
    n533
  );


  xor
  g576
  (
    n613,
    n573,
    n535,
    n533,
    n574
  );


  xor
  g577
  (
    n612,
    n572,
    n571,
    n534,
    n531
  );


  xor
  g578
  (
    n606,
    n574,
    n532,
    n531
  );


  xnor
  g579
  (
    n609,
    n533,
    n572,
    n534
  );


  xnor
  g580
  (
    n614,
    n532,
    n573,
    n572
  );


  nor
  g581
  (
    n611,
    n534,
    n531,
    n572,
    n573
  );


  or
  g582
  (
    n623,
    n588,
    n602,
    n612,
    n540
  );


  nand
  g583
  (
    n648,
    n610,
    n538,
    n585,
    n595
  );


  xor
  g584
  (
    n634,
    n598,
    n603,
    n542,
    n594
  );


  xor
  g585
  (
    n619,
    n579,
    n610,
    n585,
    n611
  );


  and
  g586
  (
    n631,
    n594,
    n578,
    n577
  );


  nor
  g587
  (
    n620,
    n539,
    n578,
    n541,
    n612
  );


  xnor
  g588
  (
    n615,
    n595,
    n587,
    n609,
    n604
  );


  xor
  g589
  (
    n617,
    n606,
    n609,
    n593,
    n586
  );


  and
  g590
  (
    n650,
    n593,
    n606,
    n541,
    n598
  );


  and
  g591
  (
    AntiSAT_key_wire,
    n536,
    n582,
    n580,
    n606
  );


  or
  g592
  (
    n638,
    n598,
    n607,
    n583
  );


  or
  g593
  (
    n645,
    n598,
    n597,
    n605,
    n586
  );


  nand
  g594
  (
    n651,
    n593,
    n540,
    n577,
    n590
  );


  xor
  g595
  (
    n642,
    n575,
    n576,
    n581,
    n542
  );


  nand
  g596
  (
    n641,
    n539,
    n590,
    n608,
    n537
  );


  nor
  g597
  (
    n654,
    n587,
    n597,
    n581,
    n589
  );


  and
  g598
  (
    n630,
    n542,
    n612,
    n538,
    n611
  );


  xor
  g599
  (
    n621,
    n605,
    n588,
    n591,
    n595
  );


  xnor
  g600
  (
    n639,
    n593,
    n595,
    n604,
    n585
  );


  xnor
  g601
  (
    n632,
    n586,
    n536,
    n607,
    n603
  );


  nand
  g602
  (
    n633,
    n609,
    n592,
    n605,
    n604
  );


  xnor
  g603
  (
    n628,
    n608,
    n539,
    n579,
    n580
  );


  nor
  g604
  (
    n656,
    n596,
    n537,
    n592,
    n540
  );


  xor
  g605
  (
    n640,
    n589,
    n579,
    n584,
    n582
  );


  or
  g606
  (
    n625,
    n582,
    n603,
    n611,
    n538
  );


  or
  g607
  (
    n635,
    n604,
    n596,
    n581,
    n590
  );


  and
  g608
  (
    n637,
    n586,
    n591,
    n608,
    n540
  );


  nand
  g609
  (
    n644,
    n613,
    n575,
    n584,
    n576
  );


  nor
  g610
  (
    n616,
    n579,
    n603,
    n537,
    n612
  );


  xnor
  g611
  (
    n652,
    n587,
    n589,
    n577,
    n581
  );


  nand
  g612
  (
    n629,
    n541,
    n596,
    n542
  );


  nor
  g613
  (
    n653,
    n610,
    n541,
    n574,
    n577
  );


  xnor
  g614
  (
    n636,
    n607,
    n576,
    n592,
    n538
  );


  or
  g615
  (
    n646,
    n597,
    n588,
    n594,
    n606
  );


  nor
  g616
  (
    n618,
    n608,
    n537,
    n591,
    n578
  );


  nor
  g617
  (
    n647,
    n611,
    n535,
    n536,
    n594
  );


  xor
  g618
  (
    n627,
    n584,
    n575,
    n605,
    n607
  );


  and
  g619
  (
    n655,
    n589,
    n592,
    n597,
    n583
  );


  xor
  g620
  (
    n649,
    n582,
    n536,
    n591,
    n580
  );


  and
  g621
  (
    n626,
    n576,
    n583,
    n590,
    n580
  );


  nor
  g622
  (
    n643,
    n539,
    n587,
    n610,
    n575
  );


  or
  g623
  (
    n622,
    n585,
    n584,
    n588,
    n609
  );


  buf
  g624
  (
    n661,
    n643
  );


  buf
  g625
  (
    n664,
    n544
  );


  and
  g626
  (
    n659,
    n640,
    n544
  );


  nor
  g627
  (
    n663,
    n637,
    n645,
    n648
  );


  xor
  g628
  (
    n670,
    n543,
    n546,
    n544
  );


  and
  g629
  (
    n672,
    n614,
    n613,
    n543
  );


  and
  g630
  (
    n657,
    n651,
    n601,
    n599
  );


  xnor
  g631
  (
    n662,
    n546,
    n634,
    n545
  );


  nor
  g632
  (
    n674,
    n631,
    n546,
    n649
  );


  xnor
  g633
  (
    n660,
    n632,
    n543,
    n635
  );


  or
  g634
  (
    n673,
    n646,
    n642,
    n599
  );


  xnor
  g635
  (
    n669,
    n613,
    n600
  );


  nand
  g636
  (
    n668,
    n641,
    n601,
    n639
  );


  or
  g637
  (
    n667,
    n650,
    n638,
    n644
  );


  nand
  g638
  (
    n666,
    n636,
    n633,
    n599
  );


  nor
  g639
  (
    n665,
    n545,
    n543,
    n601
  );


  nor
  g640
  (
    n676,
    n600,
    n545
  );


  xor
  g641
  (
    n658,
    n546,
    n614,
    n600
  );


  nand
  g642
  (
    n671,
    n614,
    n647,
    n601
  );


  nand
  g643
  (
    n675,
    n613,
    n599,
    n614
  );


  or
  g644
  (
    n678,
    n663,
    n676
  );


  xor
  g645
  (
    n681,
    n659,
    n548,
    n100,
    n658
  );


  and
  g646
  (
    n680,
    n657,
    n490,
    n547,
    n658
  );


  xor
  g647
  (
    n690,
    n502,
    n663,
    n666,
    n662
  );


  nor
  g648
  (
    n684,
    n23,
    n661,
    n547,
    n492
  );


  nor
  g649
  (
    n704,
    n25,
    n669,
    n26,
    n654
  );


  and
  g650
  (
    n691,
    n670,
    n667,
    n661,
    n550
  );


  and
  g651
  (
    n708,
    n499,
    n672,
    n673,
    n494
  );


  and
  g652
  (
    n687,
    n25,
    n676,
    n496,
    n668
  );


  nand
  g653
  (
    n700,
    n663,
    n101,
    n500,
    n497
  );


  nor
  g654
  (
    n689,
    n662,
    n549,
    n674,
    n658
  );


  nor
  g655
  (
    n703,
    n103,
    n24,
    n673,
    n671
  );


  or
  g656
  (
    n713,
    n24,
    n670,
    n669,
    n22
  );


  xnor
  g657
  (
    n697,
    n666,
    n655,
    n550
  );


  and
  g658
  (
    n706,
    n23,
    n101,
    n668,
    n659
  );


  xnor
  g659
  (
    n696,
    n550,
    n661,
    n676,
    n675
  );


  xor
  g660
  (
    n695,
    n24,
    n661,
    n664
  );


  and
  g661
  (
    n711,
    n657,
    n665,
    n101,
    n674
  );


  or
  g662
  (
    n685,
    n674,
    n101,
    n548
  );


  xnor
  g663
  (
    n677,
    n26,
    n659,
    n504,
    n102
  );


  and
  g664
  (
    n688,
    n549,
    n652,
    n100,
    n23
  );


  or
  g665
  (
    n683,
    n666,
    n547,
    n676,
    n658
  );


  and
  g666
  (
    n702,
    n665,
    n489,
    n548,
    n503
  );


  and
  g667
  (
    n710,
    n671,
    n660,
    n495,
    n664
  );


  xnor
  g668
  (
    n679,
    n674,
    n549,
    n665,
    n671
  );


  and
  g669
  (
    n699,
    n26,
    n675,
    n670,
    n657
  );


  and
  g670
  (
    n701,
    n23,
    n491,
    n660,
    n673
  );


  nand
  g671
  (
    n692,
    n662,
    n672
  );


  xor
  g672
  (
    n705,
    n666,
    n663,
    n25,
    n669
  );


  or
  g673
  (
    n698,
    n24,
    n672,
    n656,
    n675
  );


  nor
  g674
  (
    n693,
    n102,
    n657,
    n653,
    n25
  );


  or
  g675
  (
    n694,
    n660,
    n670,
    n103,
    n668
  );


  or
  g676
  (
    n686,
    n660,
    n659,
    n501,
    n665
  );


  xor
  g677
  (
    n707,
    n549,
    n675,
    n102,
    n498
  );


  or
  g678
  (
    n682,
    n667,
    n547,
    n673,
    n103
  );


  and
  g679
  (
    n709,
    n102,
    n664,
    n667
  );


  nor
  g680
  (
    n712,
    n493,
    n668,
    n669,
    n671
  );


  buf
  g681
  (
    n718,
    n688
  );


  not
  g682
  (
    n747,
    n694
  );


  buf
  g683
  (
    n731,
    n686
  );


  buf
  g684
  (
    n735,
    n695
  );


  buf
  g685
  (
    n726,
    n682
  );


  buf
  g686
  (
    n716,
    n692
  );


  not
  g687
  (
    n715,
    n683
  );


  not
  g688
  (
    n737,
    n690
  );


  not
  g689
  (
    n740,
    n690
  );


  buf
  g690
  (
    n714,
    n684
  );


  buf
  g691
  (
    n725,
    n694
  );


  not
  g692
  (
    n732,
    n679
  );


  buf
  g693
  (
    n736,
    n679
  );


  not
  g694
  (
    n745,
    n680
  );


  not
  g695
  (
    n741,
    n691
  );


  buf
  g696
  (
    n748,
    n686
  );


  buf
  g697
  (
    n742,
    n677
  );


  not
  g698
  (
    n730,
    n678
  );


  buf
  g699
  (
    n743,
    n685
  );


  not
  g700
  (
    n746,
    n683
  );


  buf
  g701
  (
    n723,
    n681
  );


  buf
  g702
  (
    n717,
    n684
  );


  buf
  g703
  (
    n727,
    n689
  );


  buf
  g704
  (
    n721,
    n685
  );


  buf
  g705
  (
    n738,
    n693
  );


  buf
  g706
  (
    n733,
    n691
  );


  buf
  g707
  (
    n729,
    n687
  );


  not
  g708
  (
    n720,
    n680
  );


  not
  g709
  (
    n722,
    n687
  );


  not
  g710
  (
    n744,
    n682
  );


  buf
  g711
  (
    n728,
    n692
  );


  not
  g712
  (
    n749,
    n689
  );


  not
  g713
  (
    n734,
    n693
  );


  not
  g714
  (
    n739,
    n681
  );


  buf
  g715
  (
    n719,
    n688
  );


  not
  g716
  (
    n724,
    n678
  );


  nor
  g717
  (
    n753,
    n723,
    n708,
    n728
  );


  or
  g718
  (
    n784,
    n707,
    n746,
    n729,
    n559
  );


  or
  g719
  (
    n757,
    n710,
    n735,
    n704,
    n552
  );


  nand
  g720
  (
    n789,
    n712,
    n745,
    n735,
    n741
  );


  nand
  g721
  (
    n773,
    n734,
    n725,
    n556,
    n737
  );


  xor
  g722
  (
    n762,
    n554,
    n742,
    n719,
    n732
  );


  or
  g723
  (
    n794,
    n716,
    n698,
    n725,
    n746
  );


  or
  g724
  (
    n763,
    n731,
    n558,
    n709,
    n739
  );


  or
  g725
  (
    n801,
    n725,
    n740,
    n732,
    n743
  );


  xnor
  g726
  (
    n752,
    n560,
    n560,
    n742,
    n555
  );


  or
  g727
  (
    n797,
    n741,
    n718,
    n559,
    n748
  );


  xor
  g728
  (
    n769,
    n702,
    n730,
    n554,
    n700
  );


  nor
  g729
  (
    n798,
    n728,
    n711,
    n745,
    n727
  );


  xor
  g730
  (
    n778,
    n557,
    n551,
    n731,
    n727
  );


  and
  g731
  (
    n779,
    n747,
    n723,
    n749,
    n702
  );


  nor
  g732
  (
    n785,
    n714,
    n558,
    n715,
    n744
  );


  or
  g733
  (
    n782,
    n720,
    n749,
    n552,
    n719
  );


  nor
  g734
  (
    n800,
    n737,
    n700,
    n716,
    n710
  );


  xnor
  g735
  (
    n772,
    n728,
    n734,
    n557,
    n743
  );


  nand
  g736
  (
    n787,
    n727,
    n722,
    n555,
    n720
  );


  xor
  g737
  (
    n796,
    n738,
    n747,
    n708,
    n733
  );


  xnor
  g738
  (
    n765,
    n713,
    n747,
    n722,
    n736
  );


  xnor
  g739
  (
    n764,
    n723,
    n719,
    n714,
    n737
  );


  xnor
  g740
  (
    n771,
    n557,
    n727,
    n720,
    n705
  );


  and
  g741
  (
    n776,
    n722,
    n729,
    n740,
    n747
  );


  xnor
  g742
  (
    n802,
    n735,
    n714,
    n701,
    n712
  );


  xor
  g743
  (
    n760,
    n703,
    n715,
    n558,
    n722
  );


  xnor
  g744
  (
    n759,
    n733,
    n724,
    n706,
    n697
  );


  xor
  g745
  (
    n790,
    n699,
    n726,
    n555,
    n748
  );


  or
  g746
  (
    n770,
    n730,
    n743,
    n721,
    n749
  );


  xnor
  g747
  (
    n799,
    n717,
    n744,
    n552,
    n725
  );


  nand
  g748
  (
    n767,
    n717,
    n717,
    n704,
    n696
  );


  xor
  g749
  (
    n750,
    n729,
    n744,
    n558,
    n748
  );


  xor
  g750
  (
    n775,
    n744,
    n716,
    n717
  );


  or
  g751
  (
    n783,
    n554,
    n739,
    n553,
    n697
  );


  or
  g752
  (
    n792,
    n556,
    n742,
    n738,
    n731
  );


  xnor
  g753
  (
    n804,
    n559,
    n554,
    n557,
    n741
  );


  or
  g754
  (
    n803,
    n719,
    n748,
    n726,
    n745
  );


  nand
  g755
  (
    n755,
    n551,
    n721,
    n701,
    n740
  );


  xor
  g756
  (
    n788,
    n729,
    n706,
    n715,
    n734
  );


  and
  g757
  (
    n761,
    n738,
    n555,
    n724,
    n707
  );


  xnor
  g758
  (
    n756,
    n723,
    n734,
    n721,
    n735
  );


  nand
  g759
  (
    n795,
    n713,
    n741,
    n556,
    n718
  );


  nand
  g760
  (
    n786,
    n705,
    n721,
    n736,
    n738
  );


  xor
  g761
  (
    n780,
    n709,
    n740,
    n699,
    n718
  );


  xor
  g762
  (
    n766,
    n732,
    n746,
    n726,
    n724
  );


  nor
  g763
  (
    n768,
    n736,
    n746,
    n743,
    n726
  );


  and
  g764
  (
    n781,
    n715,
    n730,
    n737,
    n714
  );


  nand
  g765
  (
    n777,
    n736,
    n553,
    n731,
    n551
  );


  xnor
  g766
  (
    n791,
    n718,
    n698,
    n745,
    n739
  );


  nor
  g767
  (
    n793,
    n552,
    n553,
    n559,
    n711
  );


  nand
  g768
  (
    n758,
    n730,
    n695,
    n703,
    n733
  );


  and
  g769
  (
    n751,
    n553,
    n696,
    n733,
    n739
  );


  nor
  g770
  (
    n774,
    n720,
    n551,
    n728,
    n749
  );


  and
  g771
  (
    n754,
    n742,
    n556,
    n732,
    n724
  );


  not
  g772
  (
    n859,
    n797
  );


  not
  g773
  (
    n824,
    n790
  );


  not
  g774
  (
    n855,
    n795
  );


  not
  g775
  (
    n845,
    n791
  );


  buf
  g776
  (
    n808,
    n789
  );


  not
  g777
  (
    n850,
    n776
  );


  not
  g778
  (
    n838,
    n786
  );


  buf
  g779
  (
    n836,
    n793
  );


  buf
  g780
  (
    n854,
    n789
  );


  buf
  g781
  (
    n831,
    n804
  );


  not
  g782
  (
    n858,
    n802
  );


  not
  g783
  (
    n809,
    n797
  );


  not
  g784
  (
    n819,
    n765
  );


  not
  g785
  (
    n813,
    n789
  );


  buf
  g786
  (
    n844,
    n760
  );


  buf
  g787
  (
    n835,
    n770
  );


  buf
  g788
  (
    n846,
    n766
  );


  not
  g789
  (
    n842,
    n752
  );


  buf
  g790
  (
    n852,
    n795
  );


  not
  g791
  (
    n867,
    n787
  );


  not
  g792
  (
    n848,
    n782
  );


  not
  g793
  (
    n865,
    n799
  );


  not
  g794
  (
    n869,
    n751
  );


  buf
  g795
  (
    n832,
    n791
  );


  buf
  g796
  (
    n810,
    n788
  );


  buf
  g797
  (
    n833,
    n794
  );


  not
  g798
  (
    n805,
    n759
  );


  not
  g799
  (
    n834,
    n756
  );


  not
  g800
  (
    n823,
    n791
  );


  not
  g801
  (
    n806,
    n778
  );


  not
  g802
  (
    n829,
    n787
  );


  not
  g803
  (
    n821,
    n804
  );


  not
  g804
  (
    n856,
    n787
  );


  not
  g805
  (
    n870,
    n753
  );


  buf
  g806
  (
    n817,
    n802
  );


  not
  g807
  (
    n843,
    n803
  );


  buf
  g808
  (
    n847,
    n797
  );


  buf
  g809
  (
    n818,
    n773
  );


  not
  g810
  (
    n828,
    n803
  );


  buf
  g811
  (
    n820,
    n795
  );


  not
  g812
  (
    n851,
    n757
  );


  not
  g813
  (
    n866,
    n780
  );


  buf
  g814
  (
    n822,
    n771
  );


  buf
  g815
  (
    n830,
    n772
  );


  buf
  g816
  (
    n827,
    n799
  );


  buf
  g817
  (
    n807,
    n801
  );


  and
  g818
  (
    n853,
    n796,
    n804
  );


  xnor
  g819
  (
    n826,
    n800,
    n796,
    n783
  );


  nor
  g820
  (
    n814,
    n801,
    n798,
    n775
  );


  nor
  g821
  (
    n868,
    n785,
    n796,
    n800
  );


  or
  g822
  (
    n812,
    n763,
    n799,
    n769
  );


  nand
  g823
  (
    n825,
    n794,
    n801,
    n790
  );


  and
  g824
  (
    n839,
    n798,
    n794,
    n800
  );


  nor
  g825
  (
    n840,
    n802,
    n789,
    n755
  );


  nor
  g826
  (
    n863,
    n787,
    n801,
    n781
  );


  and
  g827
  (
    n849,
    n799,
    n790,
    n792
  );


  xnor
  g828
  (
    n864,
    n788,
    n777,
    n784
  );


  nor
  g829
  (
    n862,
    n758,
    n792,
    n795
  );


  xor
  g830
  (
    n815,
    n774,
    n792,
    n788
  );


  xor
  g831
  (
    n860,
    n767,
    n761,
    n792
  );


  and
  g832
  (
    n857,
    n794,
    n788,
    n798
  );


  xnor
  g833
  (
    n811,
    n754,
    n803,
    n796
  );


  nor
  g834
  (
    n837,
    n798,
    n793
  );


  xor
  g835
  (
    n861,
    n803,
    n802,
    n779
  );


  and
  g836
  (
    n871,
    n797,
    n800,
    n793
  );


  nand
  g837
  (
    n841,
    n791,
    n762,
    n764
  );


  or
  g838
  (
    n816,
    n790,
    n768,
    n804
  );


  buf
  g839
  (
    n887,
    n811
  );


  buf
  g840
  (
    n877,
    n813
  );


  buf
  g841
  (
    n875,
    n812
  );


  buf
  g842
  (
    n872,
    n811
  );


  not
  g843
  (
    n884,
    n807
  );


  not
  g844
  (
    n885,
    n805
  );


  not
  g845
  (
    n888,
    n808
  );


  buf
  g846
  (
    n890,
    n810
  );


  buf
  g847
  (
    n882,
    n808
  );


  buf
  g848
  (
    n876,
    n814
  );


  not
  g849
  (
    n891,
    n807
  );


  buf
  g850
  (
    n881,
    n809
  );


  not
  g851
  (
    n883,
    n808
  );


  not
  g852
  (
    n874,
    n806
  );


  or
  g853
  (
    n889,
    n807,
    n806,
    n805,
    n812
  );


  xor
  g854
  (
    n886,
    n810,
    n810,
    n811,
    n806
  );


  xor
  g855
  (
    n873,
    n807,
    n806,
    n812,
    n805
  );


  xnor
  g856
  (
    n879,
    n810,
    n813,
    n809
  );


  xor
  g857
  (
    n880,
    n813,
    n814,
    n811,
    n809
  );


  xor
  g858
  (
    n878,
    n812,
    n813,
    n805,
    n808
  );


  or
  g859
  (
    n971,
    n859,
    n818
  );


  xor
  g860
  (
    n918,
    n880,
    n888,
    n863,
    n846
  );


  and
  g861
  (
    n904,
    n847,
    n839,
    n816,
    n832
  );


  nor
  g862
  (
    n969,
    n838,
    n876,
    n883,
    n817
  );


  nand
  g863
  (
    n911,
    n814,
    n876,
    n840,
    n824
  );


  nor
  g864
  (
    n899,
    n883,
    n842,
    n853,
    n854
  );


  nor
  g865
  (
    n945,
    n837,
    n833,
    n850,
    n891
  );


  and
  g866
  (
    n928,
    n850,
    n890,
    n824,
    n836
  );


  nor
  g867
  (
    n946,
    n823,
    n882,
    n868,
    n855
  );


  and
  g868
  (
    n953,
    n819,
    n857,
    n861,
    n871
  );


  xnor
  g869
  (
    n898,
    n867,
    n857,
    n828,
    n849
  );


  or
  g870
  (
    n968,
    n858,
    n873,
    n881,
    n854
  );


  nor
  g871
  (
    n967,
    n863,
    n855,
    n833,
    n879
  );


  nor
  g872
  (
    n938,
    n848,
    n830,
    n815,
    n863
  );


  xor
  g873
  (
    n935,
    n835,
    n891,
    n877,
    n882
  );


  or
  g874
  (
    n936,
    n839,
    n821,
    n827,
    n814
  );


  or
  g875
  (
    n919,
    n875,
    n857,
    n852,
    n863
  );


  or
  g876
  (
    n939,
    n884,
    n845,
    n834,
    n829
  );


  xnor
  g877
  (
    n917,
    n820,
    n888,
    n827,
    n831
  );


  or
  g878
  (
    n940,
    n835,
    n846,
    n870,
    n887
  );


  xnor
  g879
  (
    n920,
    n837,
    n859,
    n832,
    n857
  );


  nor
  g880
  (
    n965,
    n862,
    n878,
    n821,
    n888
  );


  nor
  g881
  (
    n896,
    n841,
    n865,
    n844,
    n883
  );


  xnor
  g882
  (
    n970,
    n849,
    n844,
    n866,
    n840
  );


  xnor
  g883
  (
    n925,
    n824,
    n824,
    n855,
    n817
  );


  nor
  g884
  (
    n951,
    n861,
    n881,
    n828,
    n825
  );


  or
  g885
  (
    n895,
    n885,
    n831,
    n839,
    n891
  );


  nand
  g886
  (
    n916,
    n871,
    n836,
    n875,
    n822
  );


  or
  g887
  (
    n947,
    n871,
    n837,
    n846,
    n856
  );


  or
  g888
  (
    n892,
    n817,
    n831,
    n561,
    n877
  );


  xnor
  g889
  (
    n927,
    n822,
    n877,
    n886
  );


  nor
  g890
  (
    n963,
    n816,
    n860,
    n828,
    n858
  );


  nor
  g891
  (
    n921,
    n837,
    n832,
    n879
  );


  xnor
  g892
  (
    n934,
    n887,
    n889,
    n838,
    n848
  );


  xnor
  g893
  (
    n893,
    n838,
    n831,
    n834,
    n866
  );


  xnor
  g894
  (
    n931,
    n884,
    n889,
    n859,
    n870
  );


  xnor
  g895
  (
    n957,
    n873,
    n864,
    n880,
    n823
  );


  and
  g896
  (
    n933,
    n561,
    n890,
    n887,
    n816
  );


  nor
  g897
  (
    n960,
    n816,
    n886,
    n858,
    n855
  );


  and
  g898
  (
    n955,
    n841,
    n835,
    n843,
    n842
  );


  xnor
  g899
  (
    n948,
    n870,
    n820,
    n562,
    n832
  );


  nor
  g900
  (
    n929,
    n853,
    n826,
    n873,
    n877
  );


  xnor
  g901
  (
    n966,
    n885,
    n842,
    n852,
    n817
  );


  nor
  g902
  (
    n924,
    n838,
    n883,
    n833,
    n867
  );


  xnor
  g903
  (
    n894,
    n830,
    n875,
    n862,
    n815
  );


  or
  g904
  (
    n897,
    n849,
    n875,
    n818,
    n847
  );


  xor
  g905
  (
    n932,
    n872,
    n844,
    n876,
    n829
  );


  xnor
  g906
  (
    n942,
    n866,
    n836,
    n865,
    n864
  );


  xnor
  g907
  (
    n910,
    n868,
    n871,
    n872,
    n820
  );


  nor
  g908
  (
    n941,
    n818,
    n884,
    n890,
    n825
  );


  xnor
  g909
  (
    n937,
    n562,
    n851,
    n865,
    n849
  );


  and
  g910
  (
    n923,
    n826,
    n836,
    n835,
    n861
  );


  nand
  g911
  (
    n912,
    n868,
    n858,
    n840,
    n827
  );


  nand
  g912
  (
    n914,
    n820,
    n854,
    n822,
    n846
  );


  nand
  g913
  (
    n949,
    n815,
    n880,
    n827,
    n560
  );


  and
  g914
  (
    n913,
    n842,
    n885,
    n860,
    n847
  );


  xnor
  g915
  (
    n900,
    n865,
    n830,
    n822,
    n845
  );


  xnor
  g916
  (
    n902,
    n862,
    n825,
    n867
  );


  xnor
  g917
  (
    n952,
    n874,
    n874,
    n869,
    n882
  );


  xnor
  g918
  (
    n901,
    n885,
    n841,
    n850,
    n881
  );


  nand
  g919
  (
    n903,
    n869,
    n853,
    n889,
    n851
  );


  and
  g920
  (
    n950,
    n860,
    n828,
    n829,
    n834
  );


  xnor
  g921
  (
    n909,
    n826,
    n834,
    n853,
    n860
  );


  or
  g922
  (
    n905,
    n866,
    n845,
    n879,
    n561
  );


  nor
  g923
  (
    n962,
    n874,
    n862,
    n856,
    n864
  );


  xnor
  g924
  (
    n922,
    n874,
    n856,
    n888,
    n819
  );


  nand
  g925
  (
    n956,
    n852,
    n843,
    n818,
    n819
  );


  xnor
  g926
  (
    n944,
    n867,
    n560,
    n878,
    n861
  );


  nand
  g927
  (
    n958,
    n850,
    n876,
    n841,
    n823
  );


  or
  g928
  (
    n959,
    n848,
    n884,
    n881,
    n859
  );


  xnor
  g929
  (
    n915,
    n869,
    n856,
    n819,
    n891
  );


  and
  g930
  (
    n907,
    n873,
    n839,
    n840,
    n869
  );


  nor
  g931
  (
    n954,
    n844,
    n851,
    n829,
    n821
  );


  nand
  g932
  (
    n906,
    n826,
    n848,
    n886,
    n843
  );


  xor
  g933
  (
    n964,
    n889,
    n821,
    n854,
    n890
  );


  nor
  g934
  (
    n926,
    n878,
    n864,
    n872,
    n847
  );


  xnor
  g935
  (
    n930,
    n882,
    n830,
    n823,
    n845
  );


  nor
  g936
  (
    n961,
    n868,
    n878,
    n815,
    n870
  );


  xnor
  g937
  (
    n943,
    n851,
    n880,
    n872,
    n833
  );


  xor
  g938
  (
    n908,
    n561,
    n887,
    n843,
    n852
  );


  and
  g939
  (
    n984,
    n956,
    n562,
    n955
  );


  xnor
  g940
  (
    n973,
    n936,
    n919,
    n932,
    n940
  );


  xor
  g941
  (
    n991,
    n931,
    n908,
    n963,
    n926
  );


  xnor
  g942
  (
    n990,
    n944,
    n902,
    n918,
    n898
  );


  nand
  g943
  (
    n989,
    n943,
    n900,
    n892,
    n894
  );


  nor
  g944
  (
    n974,
    n962,
    n960,
    n964,
    n947
  );


  and
  g945
  (
    n985,
    n925,
    n895,
    n953,
    n945
  );


  nor
  g946
  (
    n977,
    n912,
    n927,
    n921,
    n924
  );


  and
  g947
  (
    n983,
    n933,
    n911,
    n958,
    n910
  );


  nand
  g948
  (
    n992,
    n906,
    n916,
    n913,
    n920
  );


  nor
  g949
  (
    n981,
    n960,
    n951,
    n939,
    n930
  );


  and
  g950
  (
    n975,
    n952,
    n923,
    n935,
    n962
  );


  xnor
  g951
  (
    n986,
    n948,
    n903,
    n961,
    n942
  );


  and
  g952
  (
    n982,
    n914,
    n962,
    n922,
    n949
  );


  nor
  g953
  (
    n976,
    n961,
    n907,
    n963,
    n959
  );


  xor
  g954
  (
    n972,
    n937,
    n899,
    n964,
    n901
  );


  xor
  g955
  (
    n988,
    n893,
    n904,
    n929,
    n946
  );


  or
  g956
  (
    n978,
    n928,
    n905,
    n962,
    n950
  );


  and
  g957
  (
    n979,
    n917,
    n896,
    n957,
    n963
  );


  and
  g958
  (
    n987,
    n909,
    n941,
    n938,
    n954
  );


  nand
  g959
  (
    n980,
    n897,
    n963,
    n934,
    n915
  );


  xor
  g960
  (
    n1010,
    n564,
    n968,
    n565,
    n103
  );


  xor
  g961
  (
    n1000,
    n983,
    n991,
    n565,
    n964
  );


  and
  g962
  (
    n1004,
    n990,
    n567,
    n976,
    n566
  );


  and
  g963
  (
    n1003,
    n967,
    n975,
    n992,
    n565
  );


  xnor
  g964
  (
    n996,
    n104,
    n971,
    n977,
    n979
  );


  and
  g965
  (
    n993,
    n563,
    n970,
    n985,
    n964
  );


  or
  g966
  (
    n1006,
    n104,
    n971,
    n965,
    n966
  );


  and
  g967
  (
    n1009,
    n970,
    n968,
    n563,
    n965
  );


  nand
  g968
  (
    n997,
    n987,
    n563,
    n970
  );


  or
  g969
  (
    n1008,
    n104,
    n967,
    n969,
    n968
  );


  nor
  g970
  (
    n999,
    n968,
    n988,
    n566,
    n981
  );


  xnor
  g971
  (
    n998,
    n966,
    n967,
    n566,
    n565
  );


  nor
  g972
  (
    n1001,
    n563,
    n965,
    n986,
    n564
  );


  xnor
  g973
  (
    n995,
    n967,
    n969,
    n971,
    n564
  );


  nor
  g974
  (
    n1007,
    n989,
    n980,
    n104,
    n973
  );


  and
  g975
  (
    n994,
    n971,
    n965,
    n982,
    n966
  );


  nand
  g976
  (
    n1005,
    n969,
    n966,
    n974,
    n978
  );


  nand
  g977
  (
    n1002,
    n564,
    n984,
    n969,
    n566
  );


  or
  g978
  (
    n1024,
    n511,
    n29,
    n31,
    n30
  );


  xnor
  g979
  (
    n1017,
    n569,
    n26,
    n31,
    n514
  );


  nand
  g980
  (
    n1012,
    n998,
    n32,
    n567,
    n1008
  );


  nand
  g981
  (
    n1023,
    n513,
    n30,
    n508
  );


  xnor
  g982
  (
    n1018,
    n27,
    n1006,
    n31,
    n28
  );


  nand
  g983
  (
    n1016,
    n515,
    n509,
    n997,
    n32
  );


  nor
  g984
  (
    n1015,
    n568,
    n27,
    n1004,
    n569
  );


  and
  g985
  (
    n1013,
    n568,
    n1001,
    n507,
    n1010
  );


  xor
  g986
  (
    n1022,
    n568,
    n1007,
    n28,
    n32
  );


  xnor
  g987
  (
    n1011,
    n512,
    n28,
    n999,
    n567
  );


  xnor
  g988
  (
    n1019,
    n31,
    n29,
    n32,
    n27
  );


  xnor
  g989
  (
    n1021,
    n1009,
    n1005,
    n996,
    n1003
  );


  nor
  g990
  (
    n1025,
    n506,
    n568,
    n1002,
    n29
  );


  nor
  g991
  (
    n1014,
    n28,
    n567,
    n505,
    n29
  );


  xor
  g992
  (
    n1020,
    n1000,
    n30,
    n510,
    n27
  );


  xnor
  g993
  (
    n1026,
    n569,
    n1024,
    n1022
  );


  and
  g994
  (
    n1027,
    n1020,
    n570,
    n1021
  );


  xnor
  g995
  (
    n1028,
    n569,
    n1019,
    n1023,
    n1025
  );


  nor
  g996
  (
    n1029,
    n1026,
    n570
  );


  or
  g997
  (
    n1031,
    n1027,
    n1029,
    n516,
    n1028
  );


  xnor
  g998
  (
    n1032,
    n517,
    n1029,
    n290
  );


  or
  g999
  (
    n1030,
    n1029,
    n290
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n624,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

