// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_489_535 written by SynthGen on 2021/05/24 19:47:35
module Stat_489_535( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25,
 n508, n492, n495, n490, n489, n496, n510, n507,
 n503, n491, n504, n514, n497, n505, n513, n494,
 n506, n500, n502, n512, n487, n509, n499, n498,
 n488, n501, n493, n511);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25;

output n508, n492, n495, n490, n489, n496, n510, n507,
 n503, n491, n504, n514, n497, n505, n513, n494,
 n506, n500, n502, n512, n487, n509, n499, n498,
 n488, n501, n493, n511;

wire n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486;

not  g0 (n97, n23);
buf  g1 (n101, n5);
not  g2 (n50, n18);
buf  g3 (n72, n5);
buf  g4 (n26, n6);
not  g5 (n34, n24);
not  g6 (n64, n25);
buf  g7 (n122, n14);
not  g8 (n56, n9);
not  g9 (n27, n23);
not  g10 (n109, n16);
buf  g11 (n114, n3);
not  g12 (n108, n5);
buf  g13 (n118, n16);
buf  g14 (n115, n1);
not  g15 (n43, n12);
buf  g16 (n52, n10);
not  g17 (n57, n22);
not  g18 (n41, n14);
not  g19 (n91, n14);
buf  g20 (n71, n7);
buf  g21 (n48, n9);
not  g22 (n106, n8);
not  g23 (n86, n25);
buf  g24 (n38, n21);
not  g25 (n53, n22);
buf  g26 (n47, n5);
not  g27 (n110, n1);
not  g28 (n42, n17);
buf  g29 (n55, n8);
not  g30 (n84, n16);
not  g31 (n94, n11);
not  g32 (n98, n16);
not  g33 (n61, n15);
not  g34 (n36, n14);
buf  g35 (n113, n18);
not  g36 (n74, n23);
buf  g37 (n104, n20);
buf  g38 (n121, n7);
not  g39 (n85, n23);
not  g40 (n105, n13);
buf  g41 (n81, n21);
not  g42 (n66, n10);
buf  g43 (n83, n4);
not  g44 (n70, n10);
buf  g45 (n30, n19);
buf  g46 (n111, n7);
buf  g47 (n68, n2);
buf  g48 (n73, n3);
not  g49 (n90, n11);
buf  g50 (n67, n24);
buf  g51 (n93, n6);
not  g52 (n82, n11);
buf  g53 (n87, n21);
not  g54 (n77, n1);
not  g55 (n120, n15);
buf  g56 (n116, n9);
not  g57 (n100, n4);
buf  g58 (n46, n7);
not  g59 (n95, n17);
not  g60 (n33, n18);
buf  g61 (n69, n19);
not  g62 (n60, n24);
buf  g63 (n79, n17);
buf  g64 (n99, n13);
buf  g65 (n102, n2);
buf  g66 (n89, n19);
not  g67 (n37, n13);
buf  g68 (n80, n25);
not  g69 (n39, n9);
not  g70 (n123, n17);
not  g71 (n112, n12);
buf  g72 (n92, n1);
buf  g73 (n32, n12);
not  g74 (n35, n22);
not  g75 (n45, n21);
buf  g76 (n62, n3);
buf  g77 (n125, n4);
not  g78 (n31, n10);
not  g79 (n78, n15);
buf  g80 (n51, n8);
buf  g81 (n65, n8);
buf  g82 (n75, n12);
not  g83 (n103, n25);
not  g84 (n44, n18);
buf  g85 (n96, n22);
buf  g86 (n58, n2);
buf  g87 (n54, n20);
buf  g88 (n76, n15);
not  g89 (n119, n4);
not  g90 (n29, n24);
buf  g91 (n59, n6);
buf  g92 (n107, n3);
not  g93 (n117, n6);
not  g94 (n40, n19);
buf  g95 (n88, n13);
not  g96 (n49, n20);
not  g97 (n28, n20);
not  g98 (n124, n11);
buf  g99 (n63, n2);
not  g100 (n216, n96);
buf  g101 (n179, n95);
buf  g102 (n270, n55);
buf  g103 (n231, n35);
not  g104 (n274, n33);
not  g105 (n271, n105);
not  g106 (n193, n101);
not  g107 (n161, n110);
not  g108 (n261, n52);
not  g109 (n176, n70);
not  g110 (n206, n84);
not  g111 (n165, n76);
buf  g112 (n152, n70);
not  g113 (n217, n83);
not  g114 (n214, n118);
buf  g115 (n177, n48);
not  g116 (n245, n108);
buf  g117 (n221, n89);
not  g118 (n131, n60);
not  g119 (n138, n38);
not  g120 (n196, n117);
not  g121 (n141, n123);
not  g122 (n126, n77);
buf  g123 (n247, n46);
buf  g124 (n254, n112);
not  g125 (n209, n88);
not  g126 (n192, n56);
not  g127 (n160, n117);
not  g128 (n218, n110);
not  g129 (n267, n35);
not  g130 (n148, n107);
buf  g131 (n255, n87);
not  g132 (n275, n113);
not  g133 (n129, n74);
not  g134 (n128, n85);
buf  g135 (n248, n44);
not  g136 (n240, n37);
buf  g137 (n151, n85);
not  g138 (n185, n61);
not  g139 (n205, n55);
not  g140 (n225, n52);
buf  g141 (n158, n80);
not  g142 (n145, n104);
buf  g143 (n210, n67);
buf  g144 (n224, n63);
buf  g145 (n219, n32);
buf  g146 (n264, n59);
not  g147 (n149, n122);
buf  g148 (n234, n116);
buf  g149 (n189, n32);
not  g150 (n220, n73);
not  g151 (n213, n56);
buf  g152 (n178, n42);
not  g153 (n139, n105);
not  g154 (n134, n51);
not  g155 (n146, n86);
not  g156 (n142, n41);
not  g157 (n182, n125);
buf  g158 (n239, n91);
buf  g159 (n170, n81);
not  g160 (n262, n110);
buf  g161 (n135, n93);
buf  g162 (n243, n110);
not  g163 (n187, n28);
not  g164 (n195, n26);
buf  g165 (n164, n108);
not  g166 (n207, n36);
buf  g167 (n252, n39);
buf  g168 (n166, n68);
buf  g169 (n222, n43);
not  g170 (n269, n89);
buf  g171 (n258, n46);
not  g172 (n265, n119);
buf  g173 (n150, n34);
or   g174 (n147, n40, n92);
xor  g175 (n136, n89, n66, n75, n79);
nand g176 (n184, n72, n39, n103, n107);
xnor g177 (n276, n120, n27, n111, n81);
nor  g178 (n186, n107, n34, n105, n59);
nand g179 (n257, n45, n115, n114);
or   g180 (n169, n119, n106, n72, n79);
nor  g181 (n223, n29, n64, n99, n82);
nand g182 (n143, n75, n80, n96, n91);
nor  g183 (n175, n81, n120, n79, n68);
and  g184 (n227, n54, n58, n86);
nand g185 (n171, n55, n53, n85, n107);
or   g186 (n235, n73, n97, n72, n76);
nor  g187 (n236, n102, n36, n120, n123);
and  g188 (n191, n50, n43, n62, n123);
or   g189 (n260, n44, n121, n94);
xor  g190 (n279, n121, n112, n60, n45);
or   g191 (n215, n37, n40, n82, n115);
xor  g192 (n268, n65, n50, n58, n69);
nor  g193 (n263, n90, n78, n29, n42);
and  g194 (n278, n102, n36, n90, n58);
xor  g195 (n156, n31, n115, n108, n104);
nor  g196 (n157, n47, n56, n101, n27);
xnor g197 (n155, n95, n93, n77, n79);
nor  g198 (n201, n76, n116, n92, n49);
and  g199 (n249, n42, n74, n90, n61);
or   g200 (n242, n43, n38, n90, n67);
xnor g201 (n266, n94, n73, n37, n33);
nor  g202 (n253, n91, n68, n71);
xor  g203 (n277, n84, n66, n34, n116);
xor  g204 (n163, n65, n109, n42, n27);
nor  g205 (n204, n74, n113, n88);
or   g206 (n140, n30, n69, n63, n53);
and  g207 (n256, n99, n59, n26, n30);
and  g208 (n172, n57, n31, n30, n41);
xnor g209 (n228, n32, n118, n49, n63);
xor  g210 (n246, n104, n43, n116, n118);
nor  g211 (n190, n106, n121, n113, n69);
or   g212 (n280, n38, n71, n95, n45);
and  g213 (n168, n64, n86, n87, n111);
nand g214 (n198, n66, n124, n54);
nand g215 (n244, n91, n75, n103, n84);
and  g216 (n183, n72, n33, n63, n39);
nand g217 (n154, n106, n92, n27, n67);
nor  g218 (n188, n64, n31, n36, n98);
and  g219 (n208, n125, n96, n109, n102);
or   g220 (n232, n122, n44, n124, n81);
or   g221 (n167, n46, n64, n55, n103);
and  g222 (n281, n97, n124, n111, n35);
xnor g223 (n137, n103, n97, n83, n123);
nor  g224 (n229, n28, n84, n113, n93);
xor  g225 (n199, n80, n61, n106, n82);
and  g226 (n194, n71, n65, n49, n96);
or   g227 (n238, n117, n109, n29, n87);
or   g228 (n251, n83, n50, n45, n112);
nor  g229 (n202, n62, n100, n52, n56);
and  g230 (n174, n39, n49, n51, n114);
xor  g231 (n162, n61, n98, n48, n99);
xnor g232 (n153, n46, n75, n37, n58);
and  g233 (n159, n26, n111, n100, n119);
nand g234 (n200, n53, n94, n80, n104);
nand g235 (n226, n101, n92, n89, n88);
or   g236 (n211, n119, n29, n66, n76);
nor  g237 (n132, n53, n48, n41, n95);
nand g238 (n130, n51, n109, n65, n54);
nor  g239 (n241, n69, n121, n100, n40);
xnor g240 (n197, n47, n78, n73, n122);
xor  g241 (n230, n41, n101, n32, n99);
xor  g242 (n237, n112, n74, n78, n54);
or   g243 (n203, n105, n59, n57, n50);
xor  g244 (n180, n62, n57, n51, n47);
and  g245 (n259, n125, n70, n48, n114);
or   g246 (n144, n82, n52, n60, n26);
xor  g247 (n133, n62, n30, n118, n77);
or   g248 (n250, n93, n108, n57, n71);
xnor g249 (n127, n100, n120, n78, n44);
nand g250 (n212, n38, n125, n85, n98);
xor  g251 (n233, n33, n47, n28, n60);
nor  g252 (n173, n28, n114, n83, n31);
or   g253 (n273, n70, n97, n98, n67);
xnor g254 (n181, n40, n35, n122, n102);
xnor g255 (n272, n87, n34, n77, n117);
xor  g256 (n302, n225, n218, n223, n193);
xor  g257 (n339, n225, n195, n263, n234);
nand g258 (n304, n134, n232, n171, n268);
nor  g259 (n287, n202, n242, n277, n214);
and  g260 (n394, n149, n191, n241, n180);
nand g261 (n321, n249, n201, n190, n257);
or   g262 (n355, n137, n273, n138, n200);
nor  g263 (n309, n141, n152, n210, n130);
nor  g264 (n317, n231, n247, n260, n137);
xor  g265 (n341, n216, n200, n146, n128);
and  g266 (n353, n159, n208, n199, n217);
xor  g267 (n319, n195, n163, n206, n147);
and  g268 (n306, n224, n180, n176, n202);
nand g269 (n376, n155, n145, n218, n167);
xnor g270 (n395, n182, n264, n192, n189);
or   g271 (n298, n221, n191, n151, n132);
and  g272 (n369, n185, n197, n141, n260);
xnor g273 (n359, n272, n272, n266, n274);
or   g274 (n337, n267, n211, n243, n227);
and  g275 (n311, n152, n272, n133, n233);
xnor g276 (n357, n247, n223, n204, n203);
nand g277 (n354, n247, n127, n212, n246);
or   g278 (n385, n214, n267, n183, n129);
nand g279 (n324, n270, n264, n278, n251);
nor  g280 (n331, n207, n213, n221, n181);
xnor g281 (n282, n193, n275, n248, n234);
or   g282 (n293, n147, n168, n252, n251);
xnor g283 (n351, n280, n160, n281, n153);
or   g284 (n368, n178, n194, n269, n163);
nand g285 (n398, n148, n252, n245, n166);
nor  g286 (n328, n270, n280, n164, n224);
and  g287 (n325, n217, n249, n171, n144);
and  g288 (n338, n207, n240, n187, n204);
nand g289 (n315, n181, n144, n174);
and  g290 (n292, n239, n235, n156, n212);
xor  g291 (n374, n196, n228, n256, n229);
xor  g292 (n362, n134, n254, n220, n135);
or   g293 (n314, n153, n258, n273, n178);
nand g294 (n387, n251, n195, n157, n196);
or   g295 (n379, n261, n145, n126, n191);
or   g296 (n386, n198, n273, n241, n259);
xnor g297 (n361, n225, n245, n184, n222);
nor  g298 (n390, n266, n205, n176, n206);
nor  g299 (n378, n183, n236, n259, n127);
or   g300 (n344, n211, n169, n255, n192);
or   g301 (n373, n208, n226, n209, n231);
nand g302 (n388, n140, n150, n215, n174);
xor  g303 (n358, n232, n190, n131, n235);
or   g304 (n397, n175, n230, n244, n243);
and  g305 (n366, n223, n153, n128, n269);
nand g306 (n389, n170, n276, n147, n186);
xnor g307 (n323, n219, n168, n265, n154);
and  g308 (n380, n215, n254, n207, n182);
xor  g309 (n286, n133, n239, n138, n271);
and  g310 (n305, n186, n242, n209, n263);
or   g311 (n329, n268, n237, n244, n136);
xor  g312 (n384, n260, n188, n184, n136);
xor  g313 (n318, n162, n219, n186, n210);
xnor g314 (n303, n198, n175, n154, n248);
or   g315 (n375, n131, n242, n279, n248);
or   g316 (n365, n255, n267, n228, n128);
xor  g317 (n347, n213, n150, n250, n240);
or   g318 (n313, n257, n148, n280, n182);
nand g319 (n392, n271, n196, n215, n243);
xnor g320 (n335, n236, n154, n270, n277);
and  g321 (n290, n268, n190, n137, n161);
or   g322 (n330, n226, n150, n224, n261);
xnor g323 (n346, n180, n158, n178, n262);
nor  g324 (n336, n149, n146, n173, n221);
nand g325 (n312, n141, n275, n143, n250);
xor  g326 (n334, n220, n140, n160);
nand g327 (n370, n143, n238, n135, n198);
and  g328 (n352, n155, n220, n240, n156);
xnor g329 (n364, n194, n271, n161, n266);
xnor g330 (n371, n170, n226, n232, n158);
xnor g331 (n297, n135, n250, n246, n278);
or   g332 (n342, n230, n143, n237, n199);
or   g333 (n345, n236, n152, n222, n206);
and  g334 (n301, n203, n192, n157, n262);
and  g335 (n288, n252, n139, n176, n126);
xor  g336 (n377, n214, n163, n173, n167);
or   g337 (n285, n205, n274, n139, n197);
xnor g338 (n340, n185, n205, n222, n166);
or   g339 (n350, n256, n245, n149, n162);
nor  g340 (n291, n218, n132, n217, n276);
nand g341 (n294, n263, n172, n193, n230);
nor  g342 (n327, n227, n256, n177, n139);
nand g343 (n299, n175, n281, n253, n187);
nand g344 (n381, n258, n168, n189, n201);
xor  g345 (n382, n167, n177, n127, n274);
or   g346 (n393, n254, n171, n203, n130);
nor  g347 (n296, n194, n211, n181, n136);
xnor g348 (n316, n142, n265, n155, n239);
xnor g349 (n308, n161, n156, n204, n238);
or   g350 (n372, n201, n159, n129, n188);
or   g351 (n343, n158, n189, n265, n133);
xnor g352 (n307, n162, n159, n157, n142);
and  g353 (n295, n183, n275, n202, n253);
or   g354 (n356, n172, n278, n165, n216);
and  g355 (n349, n165, n179, n258, n187);
xnor g356 (n360, n255, n238, n169, n166);
xnor g357 (n363, n235, n142, n148, n228);
xnor g358 (n348, n269, n213, n209, n165);
nand g359 (n310, n237, n179, n249, n129);
xor  g360 (n367, n216, n177, n231, n200);
nand g361 (n322, n145, n261, n281, n151);
nand g362 (n320, n208, n229, n227, n132);
nor  g363 (n383, n229, n257, n199, n233);
xor  g364 (n326, n219, n131, n184, n264);
nor  g365 (n333, n277, n144, n210, n276);
xor  g366 (n391, n130, n164, n279);
nor  g367 (n396, n138, n185, n188, n126);
or   g368 (n283, n212, n197, n262, n279);
nand g369 (n332, n172, n169, n134, n259);
xor  g370 (n300, n170, n246, n151, n173);
xor  g371 (n289, n241, n179, n233, n234);
or   g372 (n284, n253, n146, n244, n160);
nand g373 (n481, n321, n285, n334);
xnor g374 (n408, n284, n321, n319, n308);
xor  g375 (n474, n346, n331, n313, n339);
nand g376 (n456, n298, n325, n347, n394);
xnor g377 (n440, n380, n390, n326, n369);
nand g378 (n430, n342, n292, n318, n355);
nor  g379 (n421, n378, n283, n381, n302);
nor  g380 (n425, n320, n296, n338, n367);
xnor g381 (n470, n285, n337, n321, n318);
nand g382 (n410, n377, n391, n390, n358);
xnor g383 (n426, n380, n372, n362, n359);
nor  g384 (n455, n355, n301, n309, n371);
or   g385 (n483, n388, n290, n356);
xor  g386 (n448, n373, n350, n340, n284);
xor  g387 (n431, n341, n304, n300, n297);
xor  g388 (n459, n305, n390, n336, n386);
and  g389 (n458, n339, n305, n288, n333);
xor  g390 (n469, n320, n375, n326, n312);
and  g391 (n486, n357, n353, n324, n336);
or   g392 (n419, n389, n396, n316, n294);
xor  g393 (n452, n354, n353, n387, n314);
or   g394 (n471, n341, n318, n369, n328);
nor  g395 (n417, n303, n385, n351, n341);
nor  g396 (n438, n357, n391, n377, n375);
nor  g397 (n476, n290, n395, n315, n286);
xnor g398 (n433, n383, n364, n308, n327);
nand g399 (n467, n345, n307, n343, n309);
xor  g400 (n473, n346, n365, n301, n293);
or   g401 (n453, n362, n353, n380, n287);
nor  g402 (n401, n330, n322, n389, n357);
nand g403 (n485, n397, n387, n322, n367);
nand g404 (n449, n366, n368, n337, n398);
and  g405 (n444, n355, n310, n338, n361);
and  g406 (n437, n289, n311, n327, n329);
xor  g407 (n478, n289, n317, n284, n331);
xor  g408 (n484, n359, n291, n311, n345);
nor  g409 (n416, n366, n381, n297, n388);
and  g410 (n427, n373, n336, n326, n364);
xor  g411 (n441, n294, n371, n332, n282);
xor  g412 (n446, n356, n316, n317, n361);
or   g413 (n461, n297, n286, n396, n314);
xnor g414 (n429, n305, n323, n364, n375);
xor  g415 (n418, n367, n382, n343, n360);
nor  g416 (n402, n379, n330, n293, n352);
xor  g417 (n423, n313, n295, n389, n370);
xor  g418 (n405, n312, n383, n319, n330);
nand g419 (n466, n302, n323, n392, n344);
and  g420 (n413, n395, n288, n370, n302);
nor  g421 (n443, n317, n334, n290, n379);
and  g422 (n435, n361, n299, n301, n386);
xor  g423 (n428, n324, n393, n391, n329);
xnor g424 (n482, n300, n352, n371, n363);
or   g425 (n454, n315, n288, n351, n291);
nand g426 (n460, n366, n299, n370, n289);
or   g427 (n415, n328, n306, n325, n374);
and  g428 (n462, n300, n381, n382, n398);
xnor g429 (n479, n303, n287, n340, n360);
or   g430 (n465, n333, n349, n395, n348);
nor  g431 (n414, n382, n360, n379, n283);
xor  g432 (n457, n350, n335, n323, n307);
or   g433 (n472, n348, n308, n294, n368);
nand g434 (n403, n376, n311, n334, n392);
and  g435 (n439, n393, n307, n358, n304);
or   g436 (n409, n397, n335, n372, n342);
and  g437 (n468, n369, n329, n298, n363);
or   g438 (n436, n358, n292, n385, n392);
and  g439 (n407, n328, n310, n332, n384);
xnor g440 (n480, n298, n387, n348, n286);
nor  g441 (n399, n396, n349, n344, n338);
nand g442 (n442, n349, n374, n344, n324);
xor  g443 (n450, n282, n345, n394, n359);
xnor g444 (n424, n350, n388, n304, n282);
nor  g445 (n412, n339, n327, n312, n386);
nand g446 (n463, n303, n362, n296, n306);
nand g447 (n406, n397, n306, n347, n376);
and  g448 (n422, n295, n378, n374, n335);
and  g449 (n451, n291, n384, n365, n296);
and  g450 (n447, n313, n310, n346, n368);
nand g451 (n432, n337, n332, n285, n342);
nor  g452 (n464, n365, n299, n322, n340);
or   g453 (n420, n354, n287, n319, n295);
xor  g454 (n411, n343, n376, n385, n325);
or   g455 (n475, n363, n315, n331, n384);
nand g456 (n400, n373, n292, n394, n383);
nor  g457 (n434, n283, n293, n377, n351);
or   g458 (n477, n378, n393, n372, n354);
nor  g459 (n404, n398, n314, n333, n347);
or   g460 (n445, n316, n320, n309, n352);
nor  g461 (n491, n463, n486, n423, n411);
or   g462 (n501, n431, n449, n459, n479);
and  g463 (n496, n403, n414, n461, n484);
xnor g464 (n487, n478, n466, n400, n470);
and  g465 (n506, n438, n432, n480, n421);
xor  g466 (n489, n402, n478, n442, n457);
nor  g467 (n502, n462, n418, n467, n477);
xnor g468 (n505, n410, n477, n460, n441);
or   g469 (n493, n482, n426, n472, n476);
nor  g470 (n503, n446, n448, n399, n429);
xnor g471 (n510, n474, n475, n416, n479);
and  g472 (n492, n486, n484, n405, n427);
nor  g473 (n512, n435, n455, n422, n482);
xor  g474 (n509, n485, n482, n430, n480);
or   g475 (n511, n475, n484, n409, n445);
nor  g476 (n513, n420, n417, n454, n406);
and  g477 (n497, n465, n437, n483, n478);
or   g478 (n490, n443, n433, n444, n412);
xor  g479 (n498, n428, n456, n481, n485);
xnor g480 (n507, n479, n477, n476, n481);
or   g481 (n494, n483, n483, n485, n439);
nor  g482 (n500, n458, n404, n469, n481);
xnor g483 (n499, n425, n450, n436, n447);
xor  g484 (n488, n468, n419, n434, n415);
and  g485 (n495, n473, n424, n413, n464);
nor  g486 (n504, n486, n401, n476, n407);
and  g487 (n508, n471, n440, n451, n452);
nor  g488 (n514, n475, n408, n453, n480);
endmodule
