

module Stat_186_441
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n210,
  n217,
  n212,
  n213,
  n215,
  n207,
  n208,
  n209,
  n211,
  n204,
  n203,
  n214,
  n206,
  n202,
  n216,
  n205,
  n201,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;
  output n210;output n217;output n212;output n213;output n215;output n207;output n208;output n209;output n211;output n204;output n203;output n214;output n206;output n202;output n216;output n205;output n201;
  wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n72,
    n15
  );


  not
  g1
  (
    n54,
    n14
  );


  not
  g2
  (
    n79,
    n13
  );


  buf
  g3
  (
    n60,
    n14
  );


  not
  g4
  (
    n68,
    n1
  );


  not
  g5
  (
    n39,
    n7
  );


  not
  g6
  (
    n69,
    n19
  );


  buf
  g7
  (
    n52,
    n20
  );


  not
  g8
  (
    n81,
    n6
  );


  not
  g9
  (
    n64,
    n20
  );


  not
  g10
  (
    n87,
    n13
  );


  buf
  g11
  (
    n80,
    n10
  );


  not
  g12
  (
    n63,
    n2
  );


  buf
  g13
  (
    n62,
    n10
  );


  not
  g14
  (
    n85,
    n3
  );


  not
  g15
  (
    n33,
    n11
  );


  buf
  g16
  (
    n67,
    n21
  );


  not
  g17
  (
    n66,
    n6
  );


  not
  g18
  (
    n83,
    n5
  );


  buf
  g19
  (
    n53,
    n10
  );


  buf
  g20
  (
    n82,
    n5
  );


  buf
  g21
  (
    n55,
    n18
  );


  not
  g22
  (
    n58,
    n3
  );


  buf
  g23
  (
    n57,
    n8
  );


  buf
  g24
  (
    n43,
    n14
  );


  buf
  g25
  (
    n61,
    n20
  );


  not
  g26
  (
    n35,
    n4
  );


  not
  g27
  (
    n90,
    n9
  );


  buf
  g28
  (
    n47,
    n11
  );


  buf
  g29
  (
    n34,
    n19
  );


  not
  g30
  (
    n59,
    n13
  );


  buf
  g31
  (
    n42,
    n12
  );


  not
  g32
  (
    n94,
    n17
  );


  buf
  g33
  (
    n50,
    n8
  );


  buf
  g34
  (
    n40,
    n4
  );


  not
  g35
  (
    n92,
    n16
  );


  not
  g36
  (
    n71,
    n7
  );


  not
  g37
  (
    n91,
    n17
  );


  buf
  g38
  (
    n56,
    n11
  );


  buf
  g39
  (
    n32,
    n5
  );


  not
  g40
  (
    n49,
    n2
  );


  not
  g41
  (
    n44,
    n21
  );


  not
  g42
  (
    n48,
    n6
  );


  buf
  g43
  (
    n89,
    n7
  );


  buf
  g44
  (
    n74,
    n16
  );


  buf
  g45
  (
    n41,
    n4
  );


  buf
  g46
  (
    n70,
    n8
  );


  not
  g47
  (
    n51,
    n9
  );


  not
  g48
  (
    n86,
    n12
  );


  not
  g49
  (
    n36,
    n16
  );


  buf
  g50
  (
    n73,
    n9
  );


  buf
  g51
  (
    n38,
    n12
  );


  buf
  g52
  (
    n88,
    n3
  );


  buf
  g53
  (
    n78,
    n19
  );


  not
  g54
  (
    n46,
    n1
  );


  not
  g55
  (
    n65,
    n18
  );


  not
  g56
  (
    n76,
    n15
  );


  not
  g57
  (
    n75,
    n18
  );


  not
  g58
  (
    n45,
    n1
  );


  buf
  g59
  (
    n84,
    n21
  );


  not
  g60
  (
    n77,
    n2
  );


  buf
  g61
  (
    n93,
    n15
  );


  not
  g62
  (
    n37,
    n17
  );


  buf
  g63
  (
    n100,
    n43
  );


  not
  g64
  (
    n115,
    n37
  );


  not
  g65
  (
    n122,
    n36
  );


  buf
  g66
  (
    n130,
    n39
  );


  not
  g67
  (
    n116,
    n37
  );


  buf
  g68
  (
    n127,
    n34
  );


  buf
  g69
  (
    n97,
    n42
  );


  buf
  g70
  (
    n105,
    n43
  );


  buf
  g71
  (
    n107,
    n32
  );


  not
  g72
  (
    n118,
    n32
  );


  not
  g73
  (
    n106,
    n42
  );


  not
  g74
  (
    n99,
    n36
  );


  buf
  g75
  (
    n98,
    n37
  );


  not
  g76
  (
    n117,
    n39
  );


  not
  g77
  (
    n104,
    n38
  );


  not
  g78
  (
    n96,
    n33
  );


  not
  g79
  (
    n128,
    n40
  );


  buf
  g80
  (
    n113,
    n33
  );


  not
  g81
  (
    n129,
    n33
  );


  buf
  g82
  (
    n103,
    n41
  );


  not
  g83
  (
    n120,
    n44
  );


  not
  g84
  (
    n126,
    n32
  );


  not
  g85
  (
    n109,
    n41
  );


  not
  g86
  (
    n132,
    n34
  );


  not
  g87
  (
    n119,
    n36
  );


  not
  g88
  (
    n101,
    n35
  );


  not
  g89
  (
    n110,
    n40
  );


  buf
  g90
  (
    n121,
    n41
  );


  not
  g91
  (
    n95,
    n35
  );


  not
  g92
  (
    n111,
    n39
  );


  not
  g93
  (
    n131,
    n34
  );


  buf
  g94
  (
    n102,
    n40
  );


  not
  g95
  (
    n108,
    n42
  );


  buf
  g96
  (
    n124,
    n44
  );


  buf
  g97
  (
    n114,
    n35
  );


  not
  g98
  (
    n123,
    n38
  );


  not
  g99
  (
    n125,
    n43
  );


  not
  g100
  (
    n112,
    n38
  );


  and
  g101
  (
    n182,
    n125,
    n130,
    n106
  );


  nor
  g102
  (
    n141,
    n64,
    n65,
    n113
  );


  and
  g103
  (
    n144,
    n86,
    n124,
    n100
  );


  xnor
  g104
  (
    n147,
    n124,
    n92
  );


  and
  g105
  (
    n167,
    n66,
    n84
  );


  nand
  g106
  (
    n187,
    n27,
    n51,
    n26
  );


  nand
  g107
  (
    n161,
    n57,
    n83,
    n72
  );


  nand
  g108
  (
    n159,
    n66,
    n82,
    n93
  );


  or
  g109
  (
    n143,
    n28,
    n72,
    n69
  );


  and
  g110
  (
    n150,
    n116,
    n121,
    n85
  );


  xnor
  g111
  (
    n195,
    n85,
    n91,
    n67
  );


  xnor
  g112
  (
    n190,
    n25,
    n30,
    n24
  );


  nor
  g113
  (
    n181,
    n125,
    n31,
    n126
  );


  xnor
  g114
  (
    n135,
    n119,
    n50,
    n130
  );


  or
  g115
  (
    n173,
    n45,
    n48,
    n61
  );


  and
  g116
  (
    n200,
    n74,
    n47,
    n88
  );


  nor
  g117
  (
    n151,
    n124,
    n79,
    n76
  );


  nor
  g118
  (
    n192,
    n77,
    n125,
    n52
  );


  nand
  g119
  (
    n169,
    n128,
    n64,
    n89
  );


  and
  g120
  (
    n189,
    n80,
    n29,
    n107
  );


  nand
  g121
  (
    n138,
    n62,
    n26,
    n86
  );


  and
  g122
  (
    n148,
    n117,
    n55,
    n109
  );


  xnor
  g123
  (
    n186,
    n24,
    n131,
    n67
  );


  or
  g124
  (
    n133,
    n54,
    n118,
    n93,
    n22
  );


  or
  g125
  (
    n164,
    n59,
    n27,
    n91,
    n128
  );


  nand
  g126
  (
    n142,
    n79,
    n97,
    n61,
    n129
  );


  or
  g127
  (
    n156,
    n71,
    n26,
    n57,
    n48
  );


  and
  g128
  (
    n154,
    n47,
    n56,
    n126,
    n55
  );


  nor
  g129
  (
    n179,
    n63,
    n89,
    n120,
    n45
  );


  xnor
  g130
  (
    n145,
    n25,
    n51,
    n73,
    n102
  );


  and
  g131
  (
    n180,
    n132,
    n62,
    n50,
    n25
  );


  nand
  g132
  (
    n146,
    n55,
    n69,
    n128,
    n58
  );


  xor
  g133
  (
    n155,
    n90,
    n58,
    n28
  );


  and
  g134
  (
    n196,
    n110,
    n89,
    n94,
    n84
  );


  nor
  g135
  (
    n166,
    n60,
    n81,
    n119,
    n27
  );


  xor
  g136
  (
    n175,
    n105,
    n24,
    n29,
    n98
  );


  or
  g137
  (
    n198,
    n52,
    n75,
    n118,
    n90
  );


  nand
  g138
  (
    n171,
    n72,
    n85,
    n94,
    n46
  );


  xor
  g139
  (
    n165,
    n81,
    n53,
    n83,
    n63
  );


  and
  g140
  (
    n157,
    n101,
    n87,
    n28,
    n70
  );


  xor
  g141
  (
    n178,
    n87,
    n76,
    n78,
    n96
  );


  xnor
  g142
  (
    n152,
    n114,
    n60,
    n71,
    n126
  );


  or
  g143
  (
    n188,
    n80,
    n76,
    n49,
    n62
  );


  xnor
  g144
  (
    n149,
    n92,
    n70,
    n22,
    n60
  );


  nand
  g145
  (
    n136,
    n99,
    n95,
    n91,
    n77
  );


  or
  g146
  (
    n170,
    n83,
    n53,
    n49,
    n75
  );


  xor
  g147
  (
    n191,
    n81,
    n69,
    n23,
    n82
  );


  or
  g148
  (
    n177,
    n118,
    n31,
    n127,
    n54
  );


  or
  g149
  (
    n163,
    n74,
    n68,
    n50,
    n61
  );


  xor
  g150
  (
    n162,
    n121,
    n65,
    n123,
    n108
  );


  xor
  g151
  (
    n139,
    n74,
    n79,
    n87,
    n64
  );


  and
  g152
  (
    n172,
    n119,
    n123,
    n94,
    n77
  );


  and
  g153
  (
    n184,
    n73,
    n112,
    n51,
    n131
  );


  and
  g154
  (
    n193,
    n22,
    n127,
    n80,
    n88
  );


  nand
  g155
  (
    n197,
    n93,
    n129,
    n46,
    n66
  );


  or
  g156
  (
    n137,
    n103,
    n75,
    n23,
    n120
  );


  nand
  g157
  (
    n153,
    n56,
    n122,
    n59,
    n53
  );


  and
  g158
  (
    n134,
    n90,
    n78,
    n56,
    n132
  );


  nor
  g159
  (
    n176,
    n122,
    n29,
    n57,
    n54
  );


  nand
  g160
  (
    n183,
    n121,
    n46,
    n65,
    n82
  );


  xnor
  g161
  (
    n194,
    n78,
    n63,
    n30,
    n123
  );


  nor
  g162
  (
    n185,
    n68,
    n130,
    n122,
    n127
  );


  xor
  g163
  (
    n174,
    n132,
    n111,
    n70,
    n131
  );


  xnor
  g164
  (
    n168,
    n88,
    n47,
    n45,
    n104
  );


  nand
  g165
  (
    n199,
    n49,
    n129,
    n68,
    n48
  );


  nand
  g166
  (
    n158,
    n31,
    n52,
    n67,
    n23
  );


  nor
  g167
  (
    n140,
    n30,
    n44,
    n120,
    n73
  );


  nand
  g168
  (
    n160,
    n59,
    n86,
    n71,
    n115
  );


  xor
  g169
  (
    n210,
    n156,
    n190,
    n165,
    n171
  );


  or
  g170
  (
    n208,
    n177,
    n155,
    n135,
    n137
  );


  and
  g171
  (
    n206,
    n144,
    n138,
    n186,
    n136
  );


  or
  g172
  (
    n207,
    n147,
    n154,
    n134,
    n157
  );


  and
  g173
  (
    n211,
    n163,
    n170,
    n182,
    n193
  );


  nand
  g174
  (
    n201,
    n168,
    n162,
    n183,
    n166
  );


  nor
  g175
  (
    n209,
    n185,
    n188,
    n181,
    n194
  );


  xor
  g176
  (
    n215,
    n172,
    n152,
    n191,
    n141
  );


  xor
  g177
  (
    AntiSAT_key_wire,
    n169,
    n184,
    n133,
    n200
  );


  or
  g178
  (
    n214,
    n150,
    n195,
    n189,
    n196
  );


  nor
  g179
  (
    n212,
    n198,
    n173,
    n151,
    n160
  );


  and
  g180
  (
    n216,
    n179,
    n149,
    n153,
    n174
  );


  or
  g181
  (
    n203,
    n192,
    n175,
    n139,
    n159
  );


  or
  g182
  (
    n217,
    n164,
    n145,
    n161,
    n178
  );


  nand
  g183
  (
    n205,
    n143,
    n146,
    n167,
    n148
  );


  xor
  g184
  (
    n202,
    n176,
    n187,
    n142,
    n180
  );


  and
  g185
  (
    n204,
    n197,
    n199,
    n140,
    n158
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_0,
    keyIn_0_31,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_1,
    keyIn_0_32,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_2,
    keyIn_0_33,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_3,
    keyIn_0_34,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_4,
    keyIn_0_35,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_5,
    keyIn_0_36,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_6,
    keyIn_0_37,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_7,
    keyIn_0_38,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_8,
    keyIn_0_39,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_9,
    keyIn_0_40,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_10,
    keyIn_0_41,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_11,
    keyIn_0_42,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_12,
    keyIn_0_43,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_13,
    keyIn_0_44,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_14,
    keyIn_0_45,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_15,
    keyIn_0_46,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_16,
    keyIn_0_47,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_17,
    keyIn_0_48,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_18,
    keyIn_0_49,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_19,
    keyIn_0_50,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_20,
    keyIn_0_51,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_21,
    keyIn_0_52,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_22,
    keyIn_0_53,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_23,
    keyIn_0_54,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_24,
    keyIn_0_55,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_25,
    keyIn_0_56,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_26,
    keyIn_0_57,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_27,
    keyIn_0_58,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_28,
    keyIn_0_59,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_29,
    keyIn_0_60,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_30,
    keyIn_0_61,
    n31
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n213,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

