

module Stat_874_1512
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n697,
  n693,
  n706,
  n688,
  n719,
  n678,
  n671,
  n667,
  n708,
  n681,
  n672,
  n707,
  n710,
  n712,
  n684,
  n679,
  n774,
  n898,
  n895,
  n901,
  n902,
  n897,
  n899,
  n896,
  n903,
  n900,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;
  output n697;output n693;output n706;output n688;output n719;output n678;output n671;output n667;output n708;output n681;output n672;output n707;output n710;output n712;output n684;output n679;output n774;output n898;output n895;output n901;output n902;output n897;output n899;output n896;output n903;output n900;
  wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n668;wire n669;wire n670;wire n673;wire n674;wire n675;wire n676;wire n677;wire n680;wire n682;wire n683;wire n685;wire n686;wire n687;wire n689;wire n690;wire n691;wire n692;wire n694;wire n695;wire n696;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n709;wire n711;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n139,
    n25
  );


  not
  g1
  (
    n86,
    n7
  );


  buf
  g2
  (
    n53,
    n11
  );


  buf
  g3
  (
    n88,
    n5
  );


  not
  g4
  (
    n75,
    n24
  );


  not
  g5
  (
    n48,
    n26
  );


  buf
  g6
  (
    n34,
    n8
  );


  buf
  g7
  (
    n67,
    n2
  );


  buf
  g8
  (
    n122,
    n27
  );


  not
  g9
  (
    n84,
    n3
  );


  not
  g10
  (
    n61,
    n18
  );


  buf
  g11
  (
    n99,
    n25
  );


  buf
  g12
  (
    n140,
    n25
  );


  not
  g13
  (
    n108,
    n20
  );


  buf
  g14
  (
    n71,
    n10
  );


  not
  g15
  (
    n60,
    n14
  );


  buf
  g16
  (
    n134,
    n7
  );


  buf
  g17
  (
    n143,
    n20
  );


  buf
  g18
  (
    n79,
    n16
  );


  buf
  g19
  (
    n31,
    n20
  );


  buf
  g20
  (
    n104,
    n1
  );


  not
  g21
  (
    n126,
    n23
  );


  not
  g22
  (
    n144,
    n15
  );


  not
  g23
  (
    n54,
    n11
  );


  not
  g24
  (
    n73,
    n15
  );


  not
  g25
  (
    n128,
    n27
  );


  not
  g26
  (
    n70,
    n13
  );


  not
  g27
  (
    n107,
    n4
  );


  buf
  g28
  (
    n68,
    n7
  );


  buf
  g29
  (
    n120,
    n28
  );


  buf
  g30
  (
    n97,
    n8
  );


  not
  g31
  (
    n66,
    n28
  );


  buf
  g32
  (
    n38,
    n12
  );


  buf
  g33
  (
    n80,
    n8
  );


  buf
  g34
  (
    n83,
    n4
  );


  buf
  g35
  (
    n93,
    n16
  );


  not
  g36
  (
    n105,
    n16
  );


  not
  g37
  (
    n64,
    n15
  );


  buf
  g38
  (
    n117,
    n2
  );


  not
  g39
  (
    n131,
    n19
  );


  buf
  g40
  (
    n77,
    n13
  );


  not
  g41
  (
    n37,
    n2
  );


  not
  g42
  (
    n137,
    n6
  );


  not
  g43
  (
    n141,
    n9
  );


  not
  g44
  (
    n115,
    n18
  );


  not
  g45
  (
    n44,
    n12
  );


  not
  g46
  (
    n30,
    n22
  );


  not
  g47
  (
    n41,
    n29
  );


  buf
  g48
  (
    n135,
    n1
  );


  buf
  g49
  (
    n114,
    n26
  );


  buf
  g50
  (
    n133,
    n1
  );


  buf
  g51
  (
    n123,
    n6
  );


  buf
  g52
  (
    n45,
    n23
  );


  buf
  g53
  (
    n142,
    n11
  );


  buf
  g54
  (
    n96,
    n2
  );


  buf
  g55
  (
    n106,
    n17
  );


  not
  g56
  (
    n55,
    n19
  );


  not
  g57
  (
    n52,
    n19
  );


  not
  g58
  (
    n102,
    n26
  );


  buf
  g59
  (
    n58,
    n20
  );


  not
  g60
  (
    n69,
    n9
  );


  not
  g61
  (
    n65,
    n15
  );


  not
  g62
  (
    n116,
    n5
  );


  buf
  g63
  (
    n32,
    n7
  );


  not
  g64
  (
    n112,
    n22
  );


  not
  g65
  (
    n43,
    n28
  );


  buf
  g66
  (
    n74,
    n29
  );


  buf
  g67
  (
    n92,
    n14
  );


  not
  g68
  (
    n127,
    n17
  );


  buf
  g69
  (
    n101,
    n25
  );


  not
  g70
  (
    n138,
    n21
  );


  buf
  g71
  (
    n110,
    n24
  );


  not
  g72
  (
    n124,
    n9
  );


  not
  g73
  (
    n59,
    n29
  );


  not
  g74
  (
    n129,
    n4
  );


  not
  g75
  (
    n62,
    n4
  );


  buf
  g76
  (
    n85,
    n23
  );


  buf
  g77
  (
    n78,
    n17
  );


  not
  g78
  (
    n35,
    n9
  );


  buf
  g79
  (
    n130,
    n14
  );


  not
  g80
  (
    n121,
    n22
  );


  buf
  g81
  (
    n42,
    n12
  );


  not
  g82
  (
    n51,
    n14
  );


  buf
  g83
  (
    n50,
    n17
  );


  not
  g84
  (
    n98,
    n3
  );


  not
  g85
  (
    n103,
    n28
  );


  buf
  g86
  (
    n125,
    n27
  );


  buf
  g87
  (
    n113,
    n21
  );


  not
  g88
  (
    n109,
    n10
  );


  buf
  g89
  (
    n95,
    n24
  );


  not
  g90
  (
    n56,
    n22
  );


  not
  g91
  (
    n82,
    n3
  );


  not
  g92
  (
    n90,
    n5
  );


  buf
  g93
  (
    n57,
    n21
  );


  not
  g94
  (
    n33,
    n29
  );


  buf
  g95
  (
    n72,
    n12
  );


  not
  g96
  (
    n63,
    n11
  );


  buf
  g97
  (
    n46,
    n23
  );


  not
  g98
  (
    n94,
    n10
  );


  buf
  g99
  (
    n76,
    n19
  );


  not
  g100
  (
    n111,
    n13
  );


  buf
  g101
  (
    n89,
    n1
  );


  buf
  g102
  (
    n119,
    n6
  );


  buf
  g103
  (
    n145,
    n27
  );


  buf
  g104
  (
    n136,
    n18
  );


  not
  g105
  (
    n81,
    n5
  );


  buf
  g106
  (
    n91,
    n21
  );


  not
  g107
  (
    n39,
    n8
  );


  buf
  g108
  (
    n87,
    n10
  );


  not
  g109
  (
    n132,
    n13
  );


  not
  g110
  (
    n100,
    n3
  );


  not
  g111
  (
    n49,
    n26
  );


  not
  g112
  (
    n40,
    n24
  );


  not
  g113
  (
    n118,
    n18
  );


  buf
  g114
  (
    n47,
    n6
  );


  not
  g115
  (
    n36,
    n16
  );


  buf
  g116
  (
    n227,
    n97
  );


  not
  g117
  (
    n373,
    n92
  );


  buf
  g118
  (
    n369,
    n102
  );


  not
  g119
  (
    n270,
    n107
  );


  buf
  g120
  (
    n363,
    n65
  );


  not
  g121
  (
    n428,
    n75
  );


  not
  g122
  (
    n337,
    n83
  );


  not
  g123
  (
    n162,
    n32
  );


  not
  g124
  (
    n153,
    n32
  );


  buf
  g125
  (
    n241,
    n45
  );


  not
  g126
  (
    n311,
    n101
  );


  buf
  g127
  (
    n346,
    n58
  );


  not
  g128
  (
    n323,
    n84
  );


  buf
  g129
  (
    n249,
    n88
  );


  buf
  g130
  (
    n215,
    n104
  );


  buf
  g131
  (
    n397,
    n73
  );


  not
  g132
  (
    n156,
    n62
  );


  buf
  g133
  (
    n269,
    n69
  );


  buf
  g134
  (
    n423,
    n103
  );


  buf
  g135
  (
    n198,
    n78
  );


  buf
  g136
  (
    n429,
    n66
  );


  not
  g137
  (
    n348,
    n90
  );


  buf
  g138
  (
    n432,
    n94
  );


  buf
  g139
  (
    n309,
    n87
  );


  not
  g140
  (
    n217,
    n68
  );


  buf
  g141
  (
    n315,
    n74
  );


  not
  g142
  (
    n273,
    n63
  );


  buf
  g143
  (
    n155,
    n95
  );


  buf
  g144
  (
    n257,
    n61
  );


  not
  g145
  (
    n344,
    n96
  );


  not
  g146
  (
    n299,
    n91
  );


  buf
  g147
  (
    n419,
    n68
  );


  buf
  g148
  (
    n158,
    n43
  );


  buf
  g149
  (
    n292,
    n105
  );


  buf
  g150
  (
    n169,
    n65
  );


  buf
  g151
  (
    n178,
    n95
  );


  not
  g152
  (
    n338,
    n53
  );


  buf
  g153
  (
    n353,
    n86
  );


  not
  g154
  (
    n193,
    n77
  );


  not
  g155
  (
    n366,
    n52
  );


  buf
  g156
  (
    n226,
    n85
  );


  not
  g157
  (
    n418,
    n55
  );


  not
  g158
  (
    n167,
    n107
  );


  buf
  g159
  (
    n388,
    n100
  );


  not
  g160
  (
    n297,
    n79
  );


  not
  g161
  (
    n378,
    n87
  );


  buf
  g162
  (
    n426,
    n64
  );


  not
  g163
  (
    n285,
    n88
  );


  not
  g164
  (
    n176,
    n94
  );


  buf
  g165
  (
    n204,
    n96
  );


  not
  g166
  (
    n275,
    n105
  );


  buf
  g167
  (
    n367,
    n74
  );


  buf
  g168
  (
    n219,
    n64
  );


  buf
  g169
  (
    n197,
    n39
  );


  not
  g170
  (
    n345,
    n52
  );


  not
  g171
  (
    n194,
    n71
  );


  buf
  g172
  (
    n203,
    n109
  );


  not
  g173
  (
    n327,
    n98
  );


  not
  g174
  (
    n304,
    n65
  );


  buf
  g175
  (
    n164,
    n69
  );


  not
  g176
  (
    n268,
    n101
  );


  not
  g177
  (
    n320,
    n41
  );


  buf
  g178
  (
    n296,
    n70
  );


  not
  g179
  (
    n210,
    n54
  );


  not
  g180
  (
    n228,
    n51
  );


  not
  g181
  (
    n330,
    n52
  );


  not
  g182
  (
    n413,
    n83
  );


  buf
  g183
  (
    n416,
    n58
  );


  buf
  g184
  (
    n243,
    n88
  );


  buf
  g185
  (
    n370,
    n81
  );


  not
  g186
  (
    n212,
    n46
  );


  not
  g187
  (
    n175,
    n86
  );


  not
  g188
  (
    n308,
    n101
  );


  buf
  g189
  (
    n195,
    n43
  );


  buf
  g190
  (
    n393,
    n38
  );


  buf
  g191
  (
    n181,
    n102
  );


  not
  g192
  (
    n350,
    n51
  );


  buf
  g193
  (
    n191,
    n56
  );


  not
  g194
  (
    n160,
    n50
  );


  buf
  g195
  (
    n206,
    n79
  );


  not
  g196
  (
    n374,
    n106
  );


  not
  g197
  (
    n307,
    n51
  );


  buf
  g198
  (
    n154,
    n60
  );


  buf
  g199
  (
    n220,
    n47
  );


  buf
  g200
  (
    n364,
    n77
  );


  buf
  g201
  (
    n265,
    n82
  );


  buf
  g202
  (
    n360,
    n93
  );


  not
  g203
  (
    n216,
    n47
  );


  not
  g204
  (
    n261,
    n72
  );


  not
  g205
  (
    n358,
    n86
  );


  not
  g206
  (
    n400,
    n75
  );


  not
  g207
  (
    n317,
    n83
  );


  buf
  g208
  (
    n223,
    n99
  );


  buf
  g209
  (
    n151,
    n85
  );


  buf
  g210
  (
    n356,
    n70
  );


  buf
  g211
  (
    n161,
    n103
  );


  not
  g212
  (
    n385,
    n78
  );


  buf
  g213
  (
    n314,
    n67
  );


  not
  g214
  (
    n424,
    n45
  );


  not
  g215
  (
    n349,
    n73
  );


  not
  g216
  (
    n289,
    n63
  );


  buf
  g217
  (
    n406,
    n57
  );


  not
  g218
  (
    n229,
    n81
  );


  buf
  g219
  (
    n182,
    n83
  );


  not
  g220
  (
    n340,
    n76
  );


  buf
  g221
  (
    n371,
    n103
  );


  buf
  g222
  (
    n300,
    n35
  );


  buf
  g223
  (
    n278,
    n44
  );


  not
  g224
  (
    n322,
    n74
  );


  buf
  g225
  (
    n208,
    n30
  );


  buf
  g226
  (
    n224,
    n63
  );


  buf
  g227
  (
    n166,
    n97
  );


  buf
  g228
  (
    n386,
    n97
  );


  not
  g229
  (
    n382,
    n55
  );


  not
  g230
  (
    n282,
    n80
  );


  not
  g231
  (
    n173,
    n50
  );


  not
  g232
  (
    n359,
    n85
  );


  buf
  g233
  (
    n174,
    n80
  );


  not
  g234
  (
    n422,
    n64
  );


  not
  g235
  (
    n255,
    n62
  );


  not
  g236
  (
    n187,
    n76
  );


  not
  g237
  (
    n263,
    n71
  );


  buf
  g238
  (
    n379,
    n67
  );


  not
  g239
  (
    n427,
    n93
  );


  buf
  g240
  (
    n148,
    n56
  );


  buf
  g241
  (
    n389,
    n46
  );


  not
  g242
  (
    n368,
    n36
  );


  not
  g243
  (
    n329,
    n63
  );


  not
  g244
  (
    n365,
    n90
  );


  buf
  g245
  (
    n230,
    n77
  );


  buf
  g246
  (
    n202,
    n76
  );


  buf
  g247
  (
    n168,
    n98
  );


  buf
  g248
  (
    n399,
    n94
  );


  buf
  g249
  (
    n225,
    n96
  );


  buf
  g250
  (
    n339,
    n103
  );


  not
  g251
  (
    n242,
    n57
  );


  not
  g252
  (
    n211,
    n91
  );


  not
  g253
  (
    n313,
    n56
  );


  not
  g254
  (
    n172,
    n35
  );


  buf
  g255
  (
    n321,
    n81
  );


  buf
  g256
  (
    n411,
    n37
  );


  buf
  g257
  (
    n276,
    n89
  );


  buf
  g258
  (
    n417,
    n90
  );


  not
  g259
  (
    n325,
    n59
  );


  buf
  g260
  (
    n391,
    n58
  );


  not
  g261
  (
    n150,
    n55
  );


  not
  g262
  (
    n267,
    n69
  );


  not
  g263
  (
    n383,
    n52
  );


  not
  g264
  (
    n163,
    n80
  );


  not
  g265
  (
    n159,
    n99
  );


  buf
  g266
  (
    n306,
    n102
  );


  buf
  g267
  (
    n287,
    n66
  );


  buf
  g268
  (
    n234,
    n109
  );


  buf
  g269
  (
    n408,
    n78
  );


  not
  g270
  (
    n283,
    n59
  );


  not
  g271
  (
    n180,
    n31
  );


  not
  g272
  (
    n333,
    n51
  );


  buf
  g273
  (
    n362,
    n86
  );


  buf
  g274
  (
    n357,
    n89
  );


  not
  g275
  (
    n394,
    n59
  );


  buf
  g276
  (
    n252,
    n48
  );


  buf
  g277
  (
    n395,
    n49
  );


  buf
  g278
  (
    n171,
    n54
  );


  not
  g279
  (
    n213,
    n62
  );


  not
  g280
  (
    n240,
    n41
  );


  buf
  g281
  (
    n214,
    n71
  );


  buf
  g282
  (
    n403,
    n66
  );


  buf
  g283
  (
    n250,
    n96
  );


  buf
  g284
  (
    n341,
    n49
  );


  not
  g285
  (
    n256,
    n78
  );


  buf
  g286
  (
    n405,
    n75
  );


  not
  g287
  (
    n328,
    n68
  );


  buf
  g288
  (
    n401,
    n101
  );


  buf
  g289
  (
    n290,
    n38
  );


  not
  g290
  (
    n149,
    n61
  );


  not
  g291
  (
    n319,
    n108
  );


  buf
  g292
  (
    n375,
    n48
  );


  not
  g293
  (
    n258,
    n47
  );


  not
  g294
  (
    n284,
    n98
  );


  not
  g295
  (
    n396,
    n82
  );


  buf
  g296
  (
    n291,
    n48
  );


  not
  g297
  (
    n244,
    n82
  );


  not
  g298
  (
    n245,
    n44
  );


  not
  g299
  (
    n177,
    n39
  );


  buf
  g300
  (
    n146,
    n90
  );


  buf
  g301
  (
    n410,
    n49
  );


  buf
  g302
  (
    n336,
    n74
  );


  not
  g303
  (
    n351,
    n60
  );


  not
  g304
  (
    n310,
    n99
  );


  buf
  g305
  (
    n347,
    n40
  );


  not
  g306
  (
    n324,
    n95
  );


  buf
  g307
  (
    n205,
    n49
  );


  buf
  g308
  (
    n190,
    n92
  );


  buf
  g309
  (
    n390,
    n73
  );


  buf
  g310
  (
    n277,
    n79
  );


  buf
  g311
  (
    n185,
    n102
  );


  not
  g312
  (
    n233,
    n59
  );


  not
  g313
  (
    n326,
    n85
  );


  buf
  g314
  (
    n430,
    n62
  );


  buf
  g315
  (
    n231,
    n97
  );


  not
  g316
  (
    n152,
    n61
  );


  buf
  g317
  (
    n376,
    n100
  );


  not
  g318
  (
    n318,
    n46
  );


  not
  g319
  (
    n235,
    n95
  );


  not
  g320
  (
    n262,
    n48
  );


  buf
  g321
  (
    n165,
    n72
  );


  not
  g322
  (
    n239,
    n30
  );


  buf
  g323
  (
    n352,
    n105
  );


  buf
  g324
  (
    n218,
    n66
  );


  buf
  g325
  (
    n232,
    n84
  );


  not
  g326
  (
    n335,
    n108
  );


  not
  g327
  (
    n184,
    n73
  );


  buf
  g328
  (
    n279,
    n54
  );


  not
  g329
  (
    n259,
    n53
  );


  buf
  g330
  (
    n293,
    n68
  );


  not
  g331
  (
    n281,
    n104
  );


  not
  g332
  (
    n387,
    n100
  );


  not
  g333
  (
    n404,
    n98
  );


  not
  g334
  (
    n192,
    n34
  );


  not
  g335
  (
    n196,
    n76
  );


  not
  g336
  (
    n179,
    n88
  );


  not
  g337
  (
    n246,
    n93
  );


  not
  g338
  (
    n354,
    n60
  );


  buf
  g339
  (
    n207,
    n65
  );


  not
  g340
  (
    n274,
    n94
  );


  not
  g341
  (
    n407,
    n100
  );


  buf
  g342
  (
    n280,
    n46
  );


  not
  g343
  (
    n392,
    n104
  );


  not
  g344
  (
    n272,
    n108
  );


  not
  g345
  (
    n247,
    n99
  );


  buf
  g346
  (
    n409,
    n54
  );


  not
  g347
  (
    n209,
    n82
  );


  buf
  g348
  (
    n298,
    n58
  );


  not
  g349
  (
    n236,
    n91
  );


  buf
  g350
  (
    n361,
    n91
  );


  buf
  g351
  (
    n377,
    n84
  );


  not
  g352
  (
    n425,
    n70
  );


  buf
  g353
  (
    n305,
    n79
  );


  not
  g354
  (
    n286,
    n92
  );


  not
  g355
  (
    n238,
    n42
  );


  not
  g356
  (
    n221,
    n106
  );


  not
  g357
  (
    n316,
    n89
  );


  buf
  g358
  (
    n355,
    n106
  );


  buf
  g359
  (
    n186,
    n71
  );


  not
  g360
  (
    n271,
    n33
  );


  not
  g361
  (
    n157,
    n64
  );


  buf
  g362
  (
    n412,
    n92
  );


  not
  g363
  (
    n170,
    n57
  );


  not
  g364
  (
    n294,
    n50
  );


  buf
  g365
  (
    n342,
    n47
  );


  buf
  g366
  (
    n402,
    n31
  );


  buf
  g367
  (
    n312,
    n89
  );


  not
  g368
  (
    n201,
    n42
  );


  buf
  g369
  (
    n398,
    n80
  );


  buf
  g370
  (
    n301,
    n56
  );


  not
  g371
  (
    n248,
    n53
  );


  not
  g372
  (
    n237,
    n87
  );


  not
  g373
  (
    n334,
    n60
  );


  not
  g374
  (
    n266,
    n61
  );


  buf
  g375
  (
    n254,
    n53
  );


  not
  g376
  (
    n188,
    n40
  );


  buf
  g377
  (
    n260,
    n72
  );


  buf
  g378
  (
    n251,
    n67
  );


  buf
  g379
  (
    n183,
    n70
  );


  not
  g380
  (
    n332,
    n67
  );


  buf
  g381
  (
    n288,
    n55
  );


  buf
  g382
  (
    n380,
    n72
  );


  not
  g383
  (
    n421,
    n37
  );


  buf
  g384
  (
    n189,
    n105
  );


  not
  g385
  (
    n415,
    n104
  );


  not
  g386
  (
    n199,
    n87
  );


  buf
  g387
  (
    n200,
    n50
  );


  not
  g388
  (
    n384,
    n34
  );


  buf
  g389
  (
    n414,
    n81
  );


  not
  g390
  (
    n343,
    n106
  );


  buf
  g391
  (
    n431,
    n57
  );


  not
  g392
  (
    n420,
    n69
  );


  not
  g393
  (
    n303,
    n107
  );


  buf
  g394
  (
    n222,
    n75
  );


  buf
  g395
  (
    n147,
    n77
  );


  buf
  g396
  (
    n253,
    n108
  );


  buf
  g397
  (
    n302,
    n33
  );


  buf
  g398
  (
    n372,
    n93
  );


  buf
  g399
  (
    n331,
    n36
  );


  buf
  g400
  (
    n264,
    n107
  );


  buf
  g401
  (
    n381,
    n84
  );


  not
  g402
  (
    n295,
    n109
  );


  not
  g403
  (
    n508,
    n165
  );


  buf
  g404
  (
    n487,
    n297
  );


  buf
  g405
  (
    n500,
    n172
  );


  buf
  g406
  (
    n501,
    n200
  );


  not
  g407
  (
    n448,
    n305
  );


  not
  g408
  (
    n462,
    n337
  );


  buf
  g409
  (
    n496,
    n249
  );


  buf
  g410
  (
    n446,
    n404
  );


  buf
  g411
  (
    n482,
    n202
  );


  not
  g412
  (
    n435,
    n376
  );


  buf
  g413
  (
    n522,
    n394
  );


  not
  g414
  (
    n475,
    n227
  );


  not
  g415
  (
    n485,
    n329
  );


  not
  g416
  (
    n449,
    n392
  );


  buf
  g417
  (
    n472,
    n300
  );


  not
  g418
  (
    n516,
    n240
  );


  buf
  g419
  (
    n504,
    n235
  );


  not
  g420
  (
    n515,
    n197
  );


  not
  g421
  (
    n471,
    n324
  );


  buf
  g422
  (
    n458,
    n152
  );


  buf
  g423
  (
    n488,
    n217
  );


  buf
  g424
  (
    n512,
    n151
  );


  not
  g425
  (
    n503,
    n173
  );


  not
  g426
  (
    n489,
    n342
  );


  buf
  g427
  (
    n495,
    n354
  );


  buf
  g428
  (
    n447,
    n370
  );


  not
  g429
  (
    n442,
    n155
  );


  not
  g430
  (
    n465,
    n153
  );


  not
  g431
  (
    n524,
    n169
  );


  not
  g432
  (
    n511,
    n400
  );


  buf
  g433
  (
    n434,
    n257
  );


  not
  g434
  (
    n490,
    n391
  );


  not
  g435
  (
    n486,
    n352
  );


  buf
  g436
  (
    n478,
    n284
  );


  buf
  g437
  (
    n441,
    n243
  );


  or
  g438
  (
    n453,
    n228,
    n331,
    n383,
    n241
  );


  xnor
  g439
  (
    n521,
    n157,
    n167,
    n330,
    n348
  );


  xor
  g440
  (
    n466,
    n267,
    n275,
    n318,
    n160
  );


  and
  g441
  (
    n525,
    n283,
    n308,
    n378,
    n179
  );


  nand
  g442
  (
    n519,
    n381,
    n225,
    n256,
    n216
  );


  xnor
  g443
  (
    n520,
    n365,
    n213,
    n289,
    n203
  );


  or
  g444
  (
    n480,
    n338,
    n393,
    n280,
    n159
  );


  xnor
  g445
  (
    n497,
    n286,
    n347,
    n333,
    n168
  );


  nand
  g446
  (
    n473,
    n218,
    n315,
    n236,
    n294
  );


  nor
  g447
  (
    n491,
    n351,
    n343,
    n410,
    n328
  );


  and
  g448
  (
    n506,
    n199,
    n146,
    n210,
    n184
  );


  and
  g449
  (
    n499,
    n270,
    n185,
    n282,
    n192
  );


  nor
  g450
  (
    n477,
    n321,
    n224,
    n176,
    n373
  );


  or
  g451
  (
    n523,
    n317,
    n229,
    n411,
    n312
  );


  xnor
  g452
  (
    n439,
    n234,
    n369,
    n339,
    n209
  );


  or
  g453
  (
    n514,
    n340,
    n191,
    n412,
    n214
  );


  xnor
  g454
  (
    n509,
    n306,
    n367,
    n403,
    n353
  );


  and
  g455
  (
    n440,
    n389,
    n362,
    n287,
    n188
  );


  and
  g456
  (
    n481,
    n253,
    n296,
    n307,
    n345
  );


  xor
  g457
  (
    n502,
    n148,
    n162,
    n244,
    n149
  );


  xor
  g458
  (
    n470,
    n364,
    n279,
    n303,
    n374
  );


  nand
  g459
  (
    n474,
    n291,
    n368,
    n164,
    n208
  );


  nor
  g460
  (
    n498,
    n311,
    n226,
    n260,
    n258
  );


  or
  g461
  (
    n469,
    n246,
    n254,
    n237,
    n397
  );


  nor
  g462
  (
    n464,
    n302,
    n408,
    n174,
    n222
  );


  nand
  g463
  (
    n461,
    n183,
    n212,
    n268,
    n264
  );


  xor
  g464
  (
    n457,
    n207,
    n178,
    n401,
    n273
  );


  or
  g465
  (
    n510,
    n255,
    n299,
    n186,
    n147
  );


  and
  g466
  (
    n507,
    n310,
    n385,
    n193,
    n161
  );


  nand
  g467
  (
    n438,
    n301,
    n158,
    n319,
    n277
  );


  nor
  g468
  (
    n476,
    n251,
    n375,
    n320,
    n304
  );


  xor
  g469
  (
    n505,
    n390,
    n349,
    n344,
    n388
  );


  xnor
  g470
  (
    n452,
    n380,
    n327,
    n163,
    n262
  );


  or
  g471
  (
    n443,
    n361,
    n346,
    n395,
    n171
  );


  xnor
  g472
  (
    n437,
    n384,
    n154,
    n334,
    n233
  );


  nor
  g473
  (
    n451,
    n326,
    n215,
    n336,
    n285
  );


  or
  g474
  (
    n494,
    n177,
    n325,
    n156,
    n274
  );


  nor
  g475
  (
    n455,
    n316,
    n206,
    n314,
    n221
  );


  or
  g476
  (
    n484,
    n358,
    n298,
    n166,
    n363
  );


  or
  g477
  (
    n459,
    n407,
    n259,
    n189,
    n201
  );


  xor
  g478
  (
    n492,
    n292,
    n261,
    n360,
    n350
  );


  nor
  g479
  (
    n463,
    n371,
    n281,
    n295,
    n250
  );


  and
  g480
  (
    n513,
    n272,
    n205,
    n180,
    n396
  );


  xnor
  g481
  (
    n456,
    n196,
    n382,
    n323,
    n402
  );


  nor
  g482
  (
    n460,
    n290,
    n223,
    n187,
    n405
  );


  xor
  g483
  (
    n518,
    n252,
    n313,
    n355,
    n248
  );


  xor
  g484
  (
    n493,
    n211,
    n263,
    n341,
    n230
  );


  nand
  g485
  (
    n517,
    n288,
    n265,
    n231,
    n194
  );


  or
  g486
  (
    n467,
    n387,
    n238,
    n269,
    n175
  );


  and
  g487
  (
    n444,
    n195,
    n245,
    n398,
    n170
  );


  and
  g488
  (
    n479,
    n247,
    n204,
    n386,
    n219
  );


  nand
  g489
  (
    n468,
    n190,
    n181,
    n266,
    n379
  );


  xnor
  g490
  (
    n483,
    n278,
    n409,
    n372,
    n399
  );


  and
  g491
  (
    n454,
    n309,
    n322,
    n220,
    n242
  );


  nand
  g492
  (
    n433,
    n239,
    n335,
    n357,
    n182
  );


  and
  g493
  (
    n445,
    n356,
    n332,
    n359,
    n406
  );


  xor
  g494
  (
    n436,
    n366,
    n150,
    n293,
    n232
  );


  xor
  g495
  (
    n450,
    n276,
    n271,
    n377,
    n198
  );


  not
  g496
  (
    n530,
    n441
  );


  buf
  g497
  (
    n552,
    n458
  );


  not
  g498
  (
    n531,
    n434
  );


  not
  g499
  (
    n553,
    n437
  );


  not
  g500
  (
    n541,
    n445
  );


  not
  g501
  (
    n550,
    n433
  );


  buf
  g502
  (
    n546,
    n453
  );


  not
  g503
  (
    n533,
    n460
  );


  buf
  g504
  (
    n545,
    n451
  );


  buf
  g505
  (
    n544,
    n450
  );


  not
  g506
  (
    n534,
    n452
  );


  buf
  g507
  (
    n527,
    n439
  );


  not
  g508
  (
    n547,
    n449
  );


  buf
  g509
  (
    n529,
    n455
  );


  not
  g510
  (
    n535,
    n448
  );


  buf
  g511
  (
    n536,
    n442
  );


  buf
  g512
  (
    n526,
    n438
  );


  buf
  g513
  (
    n540,
    n457
  );


  not
  g514
  (
    n537,
    n443
  );


  not
  g515
  (
    n532,
    n446
  );


  buf
  g516
  (
    n528,
    n456
  );


  buf
  g517
  (
    n543,
    n436
  );


  buf
  g518
  (
    n549,
    n435
  );


  not
  g519
  (
    n542,
    n459
  );


  buf
  g520
  (
    n538,
    n454
  );


  not
  g521
  (
    n551,
    n444
  );


  buf
  g522
  (
    n539,
    n447
  );


  buf
  g523
  (
    n548,
    n440
  );


  buf
  g524
  (
    n604,
    n532
  );


  buf
  g525
  (
    n608,
    n526
  );


  not
  g526
  (
    n606,
    n465
  );


  buf
  g527
  (
    n624,
    n550
  );


  not
  g528
  (
    n584,
    n537
  );


  buf
  g529
  (
    n621,
    n550
  );


  buf
  g530
  (
    n600,
    n527
  );


  not
  g531
  (
    n562,
    n501
  );


  buf
  g532
  (
    n554,
    n540
  );


  not
  g533
  (
    n629,
    n530
  );


  not
  g534
  (
    n561,
    n544
  );


  buf
  g535
  (
    n610,
    n548
  );


  buf
  g536
  (
    n638,
    n553
  );


  not
  g537
  (
    n634,
    n505
  );


  not
  g538
  (
    n639,
    n548
  );


  not
  g539
  (
    n602,
    n539
  );


  buf
  g540
  (
    n581,
    n487
  );


  not
  g541
  (
    n628,
    n533
  );


  buf
  g542
  (
    n622,
    n545
  );


  buf
  g543
  (
    n616,
    n538
  );


  buf
  g544
  (
    n589,
    n529
  );


  buf
  g545
  (
    n583,
    n533
  );


  buf
  g546
  (
    n575,
    n532
  );


  not
  g547
  (
    n573,
    n547
  );


  buf
  g548
  (
    n594,
    n541
  );


  not
  g549
  (
    n559,
    n541
  );


  buf
  g550
  (
    n586,
    n468
  );


  buf
  g551
  (
    n570,
    n506
  );


  not
  g552
  (
    n617,
    n543
  );


  buf
  g553
  (
    n605,
    n464
  );


  not
  g554
  (
    n631,
    n528
  );


  not
  g555
  (
    n590,
    n508
  );


  not
  g556
  (
    n593,
    n542
  );


  buf
  g557
  (
    n627,
    n547
  );


  buf
  g558
  (
    n632,
    n546
  );


  not
  g559
  (
    n585,
    n486
  );


  not
  g560
  (
    n633,
    n529
  );


  buf
  g561
  (
    n613,
    n511
  );


  buf
  g562
  (
    n607,
    n537
  );


  not
  g563
  (
    n572,
    n531
  );


  buf
  g564
  (
    n595,
    n490
  );


  buf
  g565
  (
    n636,
    n540
  );


  not
  g566
  (
    n569,
    n502
  );


  not
  g567
  (
    n618,
    n507
  );


  not
  g568
  (
    n556,
    n551
  );


  not
  g569
  (
    n625,
    n489
  );


  not
  g570
  (
    n564,
    n550
  );


  not
  g571
  (
    n557,
    n545
  );


  not
  g572
  (
    n637,
    n539
  );


  not
  g573
  (
    n571,
    n552
  );


  not
  g574
  (
    n623,
    n533
  );


  not
  g575
  (
    n582,
    n504
  );


  not
  g576
  (
    n563,
    n479
  );


  not
  g577
  (
    n580,
    n532
  );


  buf
  g578
  (
    n574,
    n494
  );


  not
  g579
  (
    n560,
    n538
  );


  not
  g580
  (
    n598,
    n482
  );


  buf
  g581
  (
    n603,
    n531
  );


  not
  g582
  (
    n592,
    n549
  );


  not
  g583
  (
    n599,
    n538
  );


  or
  g584
  (
    n635,
    n536,
    n548
  );


  xor
  g585
  (
    n619,
    n534,
    n542
  );


  and
  g586
  (
    n566,
    n548,
    n534,
    n512,
    n474
  );


  and
  g587
  (
    n620,
    n526,
    n545,
    n499,
    n475
  );


  nor
  g588
  (
    n565,
    n551,
    n542,
    n498,
    n529
  );


  nor
  g589
  (
    n612,
    n540,
    n530,
    n527,
    n466
  );


  or
  g590
  (
    n588,
    n495,
    n528,
    n471,
    n552
  );


  xor
  g591
  (
    n640,
    n473,
    n492,
    n535,
    n484
  );


  and
  g592
  (
    n587,
    n467,
    n480,
    n528,
    n478
  );


  xnor
  g593
  (
    n596,
    n497,
    n549,
    n543,
    n493
  );


  or
  g594
  (
    n641,
    n500,
    n534,
    n543,
    n542
  );


  and
  g595
  (
    n611,
    n547,
    n526,
    n477,
    n536
  );


  xnor
  g596
  (
    n577,
    n462,
    n469,
    n531,
    n543
  );


  nor
  g597
  (
    n597,
    n539,
    n544,
    n528,
    n463
  );


  and
  g598
  (
    n630,
    n552,
    n540,
    n485,
    n546
  );


  or
  g599
  (
    n614,
    n546,
    n546,
    n551,
    n476
  );


  or
  g600
  (
    n576,
    n472,
    n541,
    n530,
    n536
  );


  xnor
  g601
  (
    n615,
    n545,
    n547,
    n481,
    n530
  );


  nand
  g602
  (
    n558,
    n527,
    n535,
    n483
  );


  xor
  g603
  (
    n591,
    n496,
    n553,
    n509
  );


  and
  g604
  (
    n626,
    n513,
    n503,
    n544,
    n537
  );


  or
  g605
  (
    n579,
    n533,
    n537,
    n539,
    n461
  );


  or
  g606
  (
    n555,
    n527,
    n553,
    n550,
    n538
  );


  or
  g607
  (
    n578,
    n549,
    n526,
    n510,
    n552
  );


  xor
  g608
  (
    n609,
    n535,
    n551,
    n532,
    n534
  );


  xor
  g609
  (
    n567,
    n488,
    n491,
    n531,
    n541
  );


  nor
  g610
  (
    n568,
    n510,
    n536,
    n529,
    n544
  );


  nor
  g611
  (
    n601,
    n470,
    n511,
    n512,
    n549
  );


  buf
  g612
  (
    n649,
    n564
  );


  buf
  g613
  (
    n653,
    n569
  );


  not
  g614
  (
    n651,
    n576
  );


  not
  g615
  (
    n647,
    n562
  );


  buf
  g616
  (
    n658,
    n561
  );


  buf
  g617
  (
    n646,
    n563
  );


  buf
  g618
  (
    n655,
    n568
  );


  buf
  g619
  (
    n650,
    n571
  );


  not
  g620
  (
    n644,
    n566
  );


  buf
  g621
  (
    n660,
    n578
  );


  buf
  g622
  (
    n642,
    n558
  );


  buf
  g623
  (
    n648,
    n567
  );


  buf
  g624
  (
    n663,
    n555
  );


  buf
  g625
  (
    n645,
    n556
  );


  not
  g626
  (
    n662,
    n570
  );


  buf
  g627
  (
    n664,
    n559
  );


  not
  g628
  (
    n656,
    n574
  );


  buf
  g629
  (
    n661,
    n572
  );


  not
  g630
  (
    n665,
    n560
  );


  not
  g631
  (
    n652,
    n573
  );


  buf
  g632
  (
    n659,
    n575
  );


  buf
  g633
  (
    n643,
    n557
  );


  not
  g634
  (
    n666,
    n565
  );


  buf
  g635
  (
    n654,
    n554
  );


  not
  g636
  (
    n657,
    n577
  );


  and
  g637
  (
    n685,
    n618,
    n617,
    n114,
    n654
  );


  nand
  g638
  (
    n684,
    n648,
    n122,
    n115,
    n126
  );


  nor
  g639
  (
    n669,
    n113,
    n131,
    n647,
    n115
  );


  xor
  g640
  (
    n692,
    n599,
    n118,
    n586,
    n115
  );


  xor
  g641
  (
    n708,
    n590,
    n127,
    n649,
    n664
  );


  nor
  g642
  (
    n691,
    n657,
    n645,
    n114,
    n580
  );


  or
  g643
  (
    n720,
    n616,
    n653,
    n110,
    n621
  );


  xnor
  g644
  (
    n697,
    n130,
    n124,
    n117,
    n661
  );


  and
  g645
  (
    n680,
    n661,
    n653,
    n125,
    n123
  );


  or
  g646
  (
    n671,
    n112,
    n116,
    n117,
    n649
  );


  xor
  g647
  (
    n667,
    n643,
    n656,
    n642,
    n608
  );


  xor
  g648
  (
    n695,
    n664,
    n121,
    n579,
    n657
  );


  nor
  g649
  (
    n674,
    n593,
    n111,
    n659,
    n613
  );


  xor
  g650
  (
    n681,
    n644,
    n659,
    n654,
    n120
  );


  and
  g651
  (
    n686,
    n119,
    n655,
    n649,
    n650
  );


  and
  g652
  (
    n703,
    n116,
    n119,
    n594,
    n661
  );


  xnor
  g653
  (
    n719,
    n598,
    n643,
    n656,
    n587
  );


  nand
  g654
  (
    n678,
    n606,
    n130,
    n658,
    n642
  );


  nor
  g655
  (
    n690,
    n655,
    n125,
    n127
  );


  xor
  g656
  (
    n713,
    n650,
    n129,
    n643,
    n648
  );


  xnor
  g657
  (
    n673,
    n646,
    n129,
    n120,
    n130
  );


  or
  g658
  (
    n698,
    n110,
    n600,
    n645,
    n610
  );


  nor
  g659
  (
    n693,
    n603,
    n646,
    n119,
    n662
  );


  and
  g660
  (
    n718,
    n650,
    n126,
    n648,
    n582
  );


  or
  g661
  (
    n710,
    n128,
    n126,
    n120,
    n123
  );


  and
  g662
  (
    n689,
    n124,
    n121,
    n644,
    n596
  );


  or
  g663
  (
    n668,
    n665,
    n661,
    n660,
    n664
  );


  xnor
  g664
  (
    n676,
    n653,
    n655,
    n658,
    n592
  );


  xor
  g665
  (
    n675,
    n123,
    n656,
    n647,
    n663
  );


  nand
  g666
  (
    n707,
    n654,
    n128,
    n116,
    n119
  );


  xnor
  g667
  (
    n709,
    n605,
    n646,
    n122,
    n652
  );


  xnor
  g668
  (
    n705,
    n646,
    n664,
    n657,
    n113
  );


  or
  g669
  (
    n694,
    n117,
    n124,
    n123,
    n112
  );


  or
  g670
  (
    n721,
    n116,
    n120,
    n117,
    n583
  );


  xnor
  g671
  (
    n679,
    n129,
    n647,
    n125,
    n591
  );


  or
  g672
  (
    n688,
    n653,
    n122,
    n658
  );


  nand
  g673
  (
    n722,
    n584,
    n619,
    n644,
    n642
  );


  nor
  g674
  (
    n704,
    n665,
    n662,
    n118,
    n648
  );


  and
  g675
  (
    n701,
    n601,
    n654,
    n651,
    n118
  );


  nand
  g676
  (
    n716,
    n659,
    n110,
    n589,
    n112
  );


  and
  g677
  (
    n677,
    n585,
    n659,
    n127,
    n651
  );


  nand
  g678
  (
    n711,
    n111,
    n125,
    n128,
    n122
  );


  xnor
  g679
  (
    n717,
    n130,
    n121,
    n112,
    n662
  );


  xor
  g680
  (
    n702,
    n114,
    n114,
    n113,
    n614
  );


  and
  g681
  (
    n672,
    n611,
    n660,
    n645,
    n655
  );


  nor
  g682
  (
    n696,
    n642,
    n115,
    n615,
    n650
  );


  nor
  g683
  (
    n682,
    n651,
    n663,
    n126,
    n607
  );


  and
  g684
  (
    AntiSAT_key_wire,
    n110,
    n121,
    n652,
    n609
  );


  or
  g685
  (
    n712,
    n662,
    n652,
    n111,
    n581
  );


  xnor
  g686
  (
    n714,
    n663,
    n128,
    n656,
    n643
  );


  xor
  g687
  (
    n699,
    n597,
    n129,
    n602,
    n612
  );


  or
  g688
  (
    n715,
    n109,
    n620,
    n657,
    n644
  );


  xnor
  g689
  (
    n687,
    n645,
    n647,
    n588,
    n660
  );


  xnor
  g690
  (
    n700,
    n665,
    n604,
    n595,
    n111
  );


  xor
  g691
  (
    n683,
    n118,
    n660,
    n651,
    n113
  );


  xnor
  g692
  (
    n670,
    n124,
    n649,
    n652,
    n663
  );


  buf
  g693
  (
    n729,
    n416
  );


  buf
  g694
  (
    n738,
    n719
  );


  not
  g695
  (
    n741,
    n693
  );


  buf
  g696
  (
    n757,
    n684
  );


  not
  g697
  (
    n746,
    n415
  );


  not
  g698
  (
    n726,
    n687
  );


  buf
  g699
  (
    n749,
    n429
  );


  not
  g700
  (
    n735,
    n709
  );


  buf
  g701
  (
    n756,
    n715
  );


  not
  g702
  (
    n739,
    n703
  );


  not
  g703
  (
    n758,
    n424
  );


  buf
  g704
  (
    n759,
    n713
  );


  buf
  g705
  (
    n762,
    n704
  );


  buf
  g706
  (
    n731,
    n422
  );


  buf
  g707
  (
    n744,
    n425
  );


  buf
  g708
  (
    n750,
    n718
  );


  not
  g709
  (
    n743,
    n711
  );


  buf
  g710
  (
    n728,
    n419
  );


  not
  g711
  (
    n727,
    n432
  );


  not
  g712
  (
    n725,
    n708
  );


  buf
  g713
  (
    n748,
    n417
  );


  not
  g714
  (
    n730,
    n685
  );


  not
  g715
  (
    n751,
    n418
  );


  buf
  g716
  (
    n752,
    n694
  );


  not
  g717
  (
    n732,
    n689
  );


  buf
  g718
  (
    n754,
    n430
  );


  buf
  g719
  (
    n740,
    n683
  );


  not
  g720
  (
    n733,
    n414
  );


  buf
  g721
  (
    n736,
    n720
  );


  buf
  g722
  (
    n742,
    n714
  );


  not
  g723
  (
    n753,
    n426
  );


  not
  g724
  (
    n737,
    n717
  );


  or
  g725
  (
    n747,
    n696,
    n427
  );


  nand
  g726
  (
    n761,
    n690,
    n721
  );


  or
  g727
  (
    n755,
    n712,
    n688,
    n707,
    n716
  );


  xnor
  g728
  (
    n724,
    n710,
    n428,
    n697,
    n692
  );


  xor
  g729
  (
    n734,
    n702,
    n413,
    n686,
    n700
  );


  nand
  g730
  (
    n745,
    n431,
    n420,
    n691,
    n699
  );


  nor
  g731
  (
    n723,
    n423,
    n421,
    n695,
    n722
  );


  xor
  g732
  (
    n760,
    n705,
    n701,
    n698,
    n706
  );


  buf
  g733
  (
    n764,
    n524
  );


  buf
  g734
  (
    n778,
    n734
  );


  not
  g735
  (
    n774,
    n517
  );


  not
  g736
  (
    n775,
    n732
  );


  or
  g737
  (
    n771,
    n735,
    n723
  );


  and
  g738
  (
    n773,
    n525,
    n731,
    n723,
    n518
  );


  or
  g739
  (
    n770,
    n734,
    n519,
    n523,
    n513
  );


  and
  g740
  (
    n763,
    n515,
    n724,
    n727,
    n521
  );


  and
  g741
  (
    n768,
    n525,
    n520,
    n523
  );


  nand
  g742
  (
    n777,
    n522,
    n516,
    n725
  );


  nor
  g743
  (
    n769,
    n730,
    n730,
    n522,
    n724
  );


  or
  g744
  (
    n766,
    n728,
    n731,
    n727,
    n729
  );


  nor
  g745
  (
    n772,
    n732,
    n518,
    n517,
    n729
  );


  or
  g746
  (
    n765,
    n728,
    n733,
    n514
  );


  xor
  g747
  (
    n767,
    n726,
    n524,
    n521,
    n515
  );


  xor
  g748
  (
    n776,
    n514,
    n519,
    n726,
    n516
  );


  buf
  g749
  (
    n788,
    n778
  );


  not
  g750
  (
    n791,
    n765
  );


  buf
  g751
  (
    n789,
    n665
  );


  not
  g752
  (
    n780,
    n666
  );


  buf
  g753
  (
    n779,
    n771
  );


  not
  g754
  (
    n781,
    n776
  );


  not
  g755
  (
    n782,
    n774
  );


  buf
  g756
  (
    n787,
    n764
  );


  buf
  g757
  (
    n783,
    n767
  );


  buf
  g758
  (
    n784,
    n766
  );


  nor
  g759
  (
    n792,
    n767,
    n768,
    n775
  );


  xor
  g760
  (
    n785,
    n772,
    n777,
    n774
  );


  xor
  g761
  (
    n790,
    n771,
    n769,
    n770,
    n773
  );


  nand
  g762
  (
    n786,
    n772,
    n778,
    n770,
    n766
  );


  nand
  g763
  (
    n793,
    n775,
    n769,
    n776,
    n773
  );


  buf
  g764
  (
    n803,
    n629
  );


  buf
  g765
  (
    n796,
    n782
  );


  buf
  g766
  (
    n797,
    n789
  );


  buf
  g767
  (
    n801,
    n780
  );


  buf
  g768
  (
    n799,
    n630
  );


  xnor
  g769
  (
    n794,
    n788,
    n785,
    n787
  );


  xor
  g770
  (
    n800,
    n626,
    n781,
    n627,
    n625
  );


  or
  g771
  (
    n798,
    n783,
    n623,
    n786,
    n779
  );


  and
  g772
  (
    n802,
    n622,
    n628,
    n634,
    n784
  );


  xnor
  g773
  (
    n795,
    n632,
    n631,
    n624,
    n633
  );


  buf
  g774
  (
    n814,
    n666
  );


  not
  g775
  (
    n811,
    n666
  );


  not
  g776
  (
    n804,
    n666
  );


  buf
  g777
  (
    n812,
    n798
  );


  buf
  g778
  (
    n805,
    n797
  );


  buf
  g779
  (
    n809,
    n803
  );


  not
  g780
  (
    n807,
    n796
  );


  buf
  g781
  (
    n808,
    n802
  );


  not
  g782
  (
    n810,
    n803
  );


  buf
  g783
  (
    n806,
    n794
  );


  xnor
  g784
  (
    n813,
    n800,
    n799,
    n801,
    n795
  );


  not
  g785
  (
    n820,
    n142
  );


  buf
  g786
  (
    n831,
    n140
  );


  buf
  g787
  (
    n830,
    n144
  );


  buf
  g788
  (
    n845,
    n135
  );


  not
  g789
  (
    n855,
    n138
  );


  not
  g790
  (
    n858,
    n136
  );


  buf
  g791
  (
    n849,
    n134
  );


  not
  g792
  (
    n827,
    n806
  );


  buf
  g793
  (
    n846,
    n139
  );


  not
  g794
  (
    n850,
    n137
  );


  buf
  g795
  (
    n816,
    n805
  );


  not
  g796
  (
    n822,
    n139
  );


  not
  g797
  (
    n842,
    n809
  );


  buf
  g798
  (
    n839,
    n142
  );


  not
  g799
  (
    n847,
    n805
  );


  buf
  g800
  (
    n825,
    n811
  );


  buf
  g801
  (
    n844,
    n811
  );


  buf
  g802
  (
    n837,
    n135
  );


  buf
  g803
  (
    n815,
    n810
  );


  not
  g804
  (
    n818,
    n805
  );


  not
  g805
  (
    n854,
    n131
  );


  buf
  g806
  (
    n843,
    n135
  );


  nor
  g807
  (
    n832,
    n134,
    n804,
    n639,
    n814
  );


  and
  g808
  (
    n828,
    n133,
    n807,
    n641,
    n637
  );


  and
  g809
  (
    n826,
    n806,
    n638,
    n808,
    n132
  );


  xnor
  g810
  (
    n841,
    n808,
    n143,
    n807,
    n813
  );


  and
  g811
  (
    n857,
    n137,
    n812,
    n131,
    n141
  );


  and
  g812
  (
    n824,
    n807,
    n636,
    n812,
    n141
  );


  or
  g813
  (
    n829,
    n145,
    n142,
    n136,
    n804
  );


  xor
  g814
  (
    n817,
    n144,
    n144,
    n808,
    n811
  );


  nand
  g815
  (
    n852,
    n806,
    n132,
    n811,
    n138
  );


  nand
  g816
  (
    n848,
    n145,
    n807,
    n138,
    n635
  );


  xnor
  g817
  (
    n819,
    n810,
    n141,
    n142,
    n143
  );


  nor
  g818
  (
    n856,
    n135,
    n814,
    n134
  );


  nand
  g819
  (
    n853,
    n809,
    n143,
    n132,
    n133
  );


  nand
  g820
  (
    n821,
    n805,
    n640,
    n140,
    n136
  );


  xor
  g821
  (
    n833,
    n813,
    n140,
    n136,
    n131
  );


  and
  g822
  (
    n838,
    n139,
    n804,
    n133,
    n143
  );


  xnor
  g823
  (
    n834,
    n132,
    n145,
    n140,
    n141
  );


  xnor
  g824
  (
    n836,
    n138,
    n139,
    n133,
    n134
  );


  xor
  g825
  (
    n851,
    n813,
    n145,
    n804,
    n809
  );


  nand
  g826
  (
    n840,
    n810,
    n812,
    n813
  );


  xnor
  g827
  (
    n823,
    n144,
    n810,
    n137,
    n814
  );


  nand
  g828
  (
    n835,
    n806,
    n809,
    n137,
    n808
  );


  nor
  g829
  (
    n886,
    n854,
    n856,
    n855,
    n739
  );


  nor
  g830
  (
    n891,
    n833,
    n853,
    n818,
    n836
  );


  nand
  g831
  (
    n870,
    n791,
    n790,
    n752,
    n745
  );


  xnor
  g832
  (
    n866,
    n738,
    n843,
    n739,
    n855
  );


  xor
  g833
  (
    n892,
    n753,
    n858,
    n845,
    n755
  );


  nor
  g834
  (
    n873,
    n828,
    n824,
    n842,
    n760
  );


  nand
  g835
  (
    n875,
    n842,
    n753,
    n793,
    n757
  );


  xor
  g836
  (
    n868,
    n837,
    n758,
    n848,
    n762
  );


  and
  g837
  (
    n879,
    n835,
    n749,
    n747,
    n851
  );


  xor
  g838
  (
    n859,
    n839,
    n762,
    n834,
    n847
  );


  nand
  g839
  (
    n889,
    n741,
    n841,
    n849,
    n847
  );


  xor
  g840
  (
    n894,
    n753,
    n737,
    n760,
    n762
  );


  xnor
  g841
  (
    n885,
    n754,
    n849,
    n748,
    n758
  );


  and
  g842
  (
    n874,
    n754,
    n845,
    n853,
    n762
  );


  nor
  g843
  (
    n887,
    n755,
    n851,
    n857,
    n756
  );


  or
  g844
  (
    n860,
    n756,
    n838,
    n852,
    n825
  );


  nand
  g845
  (
    n869,
    n822,
    n791,
    n761,
    n826
  );


  and
  g846
  (
    n871,
    n755,
    n817,
    n742,
    n738
  );


  nand
  g847
  (
    n881,
    n757,
    n848,
    n846,
    n735
  );


  nand
  g848
  (
    n888,
    n756,
    n736,
    n856,
    n754
  );


  nand
  g849
  (
    n862,
    n758,
    n743,
    n737,
    n854
  );


  nor
  g850
  (
    n882,
    n747,
    n753,
    n832,
    n793
  );


  xor
  g851
  (
    n872,
    n760,
    n746,
    n850,
    n841
  );


  and
  g852
  (
    n884,
    n740,
    n754,
    n759,
    n755
  );


  nor
  g853
  (
    n883,
    n815,
    n742,
    n740,
    n761
  );


  and
  g854
  (
    n867,
    n819,
    n745,
    n748,
    n756
  );


  and
  g855
  (
    n865,
    n844,
    n844,
    n750,
    n757
  );


  and
  g856
  (
    n864,
    n850,
    n758,
    n830,
    n816
  );


  or
  g857
  (
    n890,
    n820,
    n852,
    n761,
    n757
  );


  nand
  g858
  (
    n880,
    n761,
    n746,
    n858,
    n829
  );


  xor
  g859
  (
    n877,
    n750,
    n827,
    n846,
    n741
  );


  or
  g860
  (
    n878,
    n759,
    n792,
    n843
  );


  nand
  g861
  (
    n861,
    n751,
    n752,
    n823,
    n831
  );


  and
  g862
  (
    n863,
    n760,
    n736,
    n821,
    n751
  );


  and
  g863
  (
    n876,
    n744,
    n743,
    n840,
    n857
  );


  and
  g864
  (
    n893,
    n744,
    n749,
    n759
  );


  or
  g865
  (
    n896,
    n873,
    n859,
    n865,
    n892
  );


  nand
  g866
  (
    n901,
    n868,
    n862,
    n861,
    n880
  );


  nor
  g867
  (
    n895,
    n890,
    n881,
    n867,
    n879
  );


  xnor
  g868
  (
    n898,
    n876,
    n863,
    n885,
    n864
  );


  xnor
  g869
  (
    n897,
    n887,
    n872,
    n893,
    n869
  );


  xor
  g870
  (
    n899,
    n894,
    n884,
    n882,
    n886
  );


  xor
  g871
  (
    n900,
    n889,
    n866,
    n878,
    n883
  );


  nor
  g872
  (
    n902,
    n860,
    n877,
    n875,
    n891
  );


  xor
  g873
  (
    n903,
    n870,
    n871,
    n888,
    n874
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_29
  (
    gbar_input_0_0,
    keyIn_0_29,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_1,
    keyIn_0_30,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_2,
    keyIn_0_31,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_3,
    keyIn_0_32,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_4,
    keyIn_0_33,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_5,
    keyIn_0_34,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_6,
    keyIn_0_35,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_7,
    keyIn_0_36,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_8,
    keyIn_0_37,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_9,
    keyIn_0_38,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_10,
    keyIn_0_39,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_11,
    keyIn_0_40,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_12,
    keyIn_0_41,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_13,
    keyIn_0_42,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_14,
    keyIn_0_43,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_15,
    keyIn_0_44,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_16,
    keyIn_0_45,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_17,
    keyIn_0_46,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_18,
    keyIn_0_47,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_19,
    keyIn_0_48,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_20,
    keyIn_0_49,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_21,
    keyIn_0_50,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_22,
    keyIn_0_51,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_23,
    keyIn_0_52,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_24,
    keyIn_0_53,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_25,
    keyIn_0_54,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_26,
    keyIn_0_55,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_27,
    keyIn_0_56,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_28,
    keyIn_0_57,
    n29
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n706,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

