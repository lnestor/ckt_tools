// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_255_53 written by SynthGen on 2021/05/24 19:47:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_255_53 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28,
 n278, n282, n273, n275, n281, n274, n271, n270,
 n283, n267, n280, n276, n272, n277, n279, n269,
 n268);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28;

output n278, n282, n273, n275, n281, n274, n271, n270,
 n283, n267, n280, n276, n272, n277, n279, n269,
 n268;

wire n29, n30, n31, n32, n33, n34, n35, n36,
 n37, n38, n39, n40, n41, n42, n43, n44,
 n45, n46, n47, n48, n49, n50, n51, n52,
 n53, n54, n55, n56, n57, n58, n59, n60,
 n61, n62, n63, n64, n65, n66, n67, n68,
 n69, n70, n71, n72, n73, n74, n75, n76,
 n77, n78, n79, n80, n81, n82, n83, n84,
 n85, n86, n87, n88, n89, n90, n91, n92,
 n93, n94, n95, n96, n97, n98, n99, n100,
 n101, n102, n103, n104, n105, n106, n107, n108,
 n109, n110, n111, n112, n113, n114, n115, n116,
 n117, n118, n119, n120, n121, n122, n123, n124,
 n125, n126, n127, n128, n129, n130, n131, n132,
 n133, n134, n135, n136, n137, n138, n139, n140,
 n141, n142, n143, n144, n145, n146, n147, n148,
 n149, n150, n151, n152, n153, n154, n155, n156,
 n157, n158, n159, n160, n161, n162, n163, n164,
 n165, n166, n167, n168, n169, n170, n171, n172,
 n173, n174, n175, n176, n177, n178, n179, n180,
 n181, n182, n183, n184, n185, n186, n187, n188,
 n189, n190, n191, n192, n193, n194, n195, n196,
 n197, n198, n199, n200, n201, n202, n203, n204,
 n205, n206, n207, n208, n209, n210, n211, n212,
 n213, n214, n215, n216, n217, n218, n219, n220,
 n221, n222, n223, n224, n225, n226, n227, n228,
 n229, n230, n231, n232, n233, n234, n235, n236,
 n237, n238, n239, n240, n241, n242, n243, n244,
 n245, n246, n247, n248, n249, n250, n251, n252,
 n253, n254, n255, n256, n257, n258, n259, n260,
 n261, n262, n263, n264, n265, n266;

buf  g0 (n97, n16);
not  g1 (n56, n4);
buf  g2 (n71, n24);
not  g3 (n108, n11);
not  g4 (n95, n11);
not  g5 (n109, n1);
not  g6 (n39, n6);
buf  g7 (n76, n11);
buf  g8 (n82, n14);
not  g9 (n52, n7);
not  g10 (n69, n2);
buf  g11 (n54, n17);
not  g12 (n38, n18);
buf  g13 (n101, n16);
buf  g14 (n84, n19);
not  g15 (n66, n21);
not  g16 (n88, n12);
buf  g17 (n29, n19);
not  g18 (n55, n15);
buf  g19 (n100, n20);
buf  g20 (n121, n21);
not  g21 (n34, n4);
not  g22 (n94, n2);
buf  g23 (n91, n13);
buf  g24 (n92, n10);
not  g25 (n87, n8);
not  g26 (n120, n7);
not  g27 (n111, n23);
not  g28 (n107, n16);
buf  g29 (n67, n22);
buf  g30 (n90, n11);
buf  g31 (n46, n10);
buf  g32 (n78, n5);
buf  g33 (n114, n3);
buf  g34 (n93, n20);
buf  g35 (n89, n9);
not  g36 (n74, n23);
buf  g37 (n53, n13);
buf  g38 (n102, n10);
not  g39 (n86, n15);
buf  g40 (n48, n8);
buf  g41 (n116, n24);
not  g42 (n105, n9);
not  g43 (n117, n3);
buf  g44 (n79, n14);
buf  g45 (n42, n5);
not  g46 (n99, n15);
not  g47 (n85, n6);
buf  g48 (n70, n9);
not  g49 (n104, n21);
buf  g50 (n49, n23);
buf  g51 (n73, n2);
buf  g52 (n112, n13);
buf  g53 (n35, n16);
not  g54 (n44, n22);
buf  g55 (n63, n2);
buf  g56 (n59, n7);
buf  g57 (n68, n3);
buf  g58 (n119, n1);
not  g59 (n72, n4);
buf  g60 (n98, n20);
not  g61 (n106, n8);
buf  g62 (n58, n22);
not  g63 (n61, n12);
buf  g64 (n30, n21);
not  g65 (n40, n24);
not  g66 (n57, n18);
not  g67 (n43, n1);
not  g68 (n77, n13);
not  g69 (n33, n6);
buf  g70 (n60, n14);
buf  g71 (n45, n3);
buf  g72 (n75, n8);
not  g73 (n51, n23);
buf  g74 (n62, n5);
buf  g75 (n47, n1);
not  g76 (n32, n6);
not  g77 (n80, n12);
buf  g78 (n36, n14);
not  g79 (n118, n18);
buf  g80 (n65, n9);
buf  g81 (n123, n17);
not  g82 (n37, n20);
buf  g83 (n64, n17);
buf  g84 (n113, n17);
not  g85 (n96, n5);
buf  g86 (n50, n4);
not  g87 (n103, n15);
buf  g88 (n31, n7);
buf  g89 (n115, n18);
not  g90 (n81, n12);
not  g91 (n41, n19);
not  g92 (n110, n22);
buf  g93 (n122, n19);
buf  g94 (n83, n10);
buf  g95 (n127, n28);
buf  g96 (n142, n25);
not  g97 (n130, n27);
buf  g98 (n139, n28);
buf  g99 (n129, n36);
buf  g100 (n147, n30);
buf  g101 (n143, n36);
buf  g102 (n131, n37);
nor  g103 (n137, n32, n25, n26);
nand g104 (n146, n43, n30, n36, n39);
nor  g105 (n133, n34, n33, n28, n40);
nor  g106 (n126, n43, n42, n38, n32);
nand g107 (n141, n27, n36, n39, n33);
nor  g108 (n148, n41, n25, n29, n40);
xnor g109 (n124, n35, n38, n31, n25);
xor  g110 (n136, n26, n27, n42, n40);
and  g111 (n135, n31, n33, n35, n42);
xor  g112 (n134, n35, n33, n41, n37);
and  g113 (n125, n30, n27, n31, n28);
xor  g114 (n132, n26, n42, n34);
nor  g115 (n138, n26, n29, n37, n40);
xnor g116 (n140, n41, n29, n35, n32);
or   g117 (n144, n34, n39, n41);
or   g118 (n128, n37, n31, n32, n38);
or   g119 (n145, n24, n38, n30, n29);
or   g120 (n210, n99, n103, n139, n110);
xnor g121 (n185, n130, n72, n90, n65);
or   g122 (n163, n100, n89, n73);
xor  g123 (n230, n55, n64, n62, n110);
xor  g124 (n214, n96, n84, n54, n102);
xor  g125 (n176, n56, n145, n96, n132);
and  g126 (n245, n44, n74, n76, n97);
xnor g127 (n172, n51, n60, n113, n99);
or   g128 (n174, n140, n108, n58, n135);
xor  g129 (n239, n92, n49, n136, n73);
nand g130 (n223, n134, n81, n141, n147);
xor  g131 (n173, n80, n107, n126, n73);
xnor g132 (n234, n84, n61, n49, n75);
and  g133 (n192, n52, n138, n148, n77);
or   g134 (n206, n50, n55, n54, n131);
nand g135 (n161, n85, n57, n135, n77);
or   g136 (n227, n93, n107, n71, n85);
and  g137 (n217, n106, n75, n99, n83);
nor  g138 (n184, n81, n147, n105, n87);
xnor g139 (n237, n46, n64, n133, n68);
and  g140 (n205, n146, n93, n103, n77);
xor  g141 (n158, n43, n94, n148, n126);
or   g142 (n215, n58, n127, n131, n124);
xor  g143 (n156, n107, n61, n138, n76);
xnor g144 (n195, n143, n107, n88, n128);
xnor g145 (n167, n111, n91, n59, n70);
and  g146 (n218, n91, n101, n44, n85);
xnor g147 (n159, n105, n62, n118, n51);
nand g148 (n191, n68, n49, n73, n77);
and  g149 (n248, n134, n144, n63, n146);
xor  g150 (n232, n54, n95, n104, n91);
or   g151 (n168, n69, n82, n98, n115);
xor  g152 (n229, n112, n143, n89, n116);
nor  g153 (n196, n137, n67, n45, n47);
nand g154 (n231, n46, n106, n144, n48);
and  g155 (n243, n93, n109, n141, n81);
nor  g156 (n166, n114, n105, n93, n71);
xnor g157 (n233, n86, n86, n131, n84);
and  g158 (n194, n82, n56, n44);
xor  g159 (n154, n141, n55, n110, n135);
or   g160 (n212, n138, n60, n86, n134);
or   g161 (n189, n127, n53, n143, n141);
nand g162 (n221, n88, n48, n82, n142);
xnor g163 (n247, n79, n104, n66, n100);
xnor g164 (n193, n136, n124, n129, n70);
nor  g165 (n181, n102, n94, n126, n136);
xnor g166 (n164, n66, n125, n64, n144);
nor  g167 (n197, n86, n72, n88, n51);
nand g168 (n149, n74, n127, n52, n69);
xor  g169 (n236, n143, n78, n64, n115);
or   g170 (n208, n76, n59, n63, n67);
xnor g171 (n187, n65, n92, n117);
xnor g172 (n244, n106, n59, n111, n140);
xor  g173 (n207, n98, n81, n84, n75);
nand g174 (n213, n118, n87, n114, n103);
or   g175 (n235, n66, n43, n113, n108);
nor  g176 (n216, n139, n78, n72, n88);
or   g177 (n152, n116, n83, n58, n142);
xnor g178 (n182, n112, n60, n144, n50);
and  g179 (n201, n148, n114, n137, n145);
and  g180 (n175, n71, n58, n130, n101);
or   g181 (n183, n60, n55, n78, n98);
xor  g182 (n171, n50, n101, n96, n100);
xor  g183 (n186, n110, n130, n146, n95);
and  g184 (n169, n80, n138, n90, n116);
or   g185 (n170, n132, n148, n139, n67);
and  g186 (n180, n95, n63, n115, n65);
and  g187 (n240, n124, n46, n105, n133);
xor  g188 (n225, n100, n89, n83, n52);
xnor g189 (n203, n48, n132, n68, n79);
nand g190 (n199, n109, n114, n108, n146);
or   g191 (n211, n147, n62, n128, n54);
nand g192 (n228, n128, n112, n102, n56);
xor  g193 (n162, n59, n53, n101, n57);
nor  g194 (n160, n125, n70, n111, n131);
nor  g195 (n204, n117, n97, n52, n124);
or   g196 (n157, n98, n111, n104, n69);
xor  g197 (n224, n125, n91, n139, n102);
nand g198 (n202, n63, n94, n129, n45);
nor  g199 (n150, n126, n61, n116, n136);
and  g200 (n151, n99, n92, n133, n83);
nor  g201 (n209, n115, n95, n117);
xnor g202 (n246, n130, n128, n127, n67);
xor  g203 (n220, n108, n50, n90, n87);
xor  g204 (n155, n96, n145, n80, n113);
or   g205 (n177, n70, n97, n62, n104);
nor  g206 (n153, n90, n97, n133, n45);
nor  g207 (n179, n78, n140, n47, n75);
nand g208 (n200, n72, n142, n112, n45);
and  g209 (n219, n142, n71, n66, n82);
xnor g210 (n165, n132, n76, n51, n57);
nor  g211 (n222, n69, n44, n53, n61);
nor  g212 (n190, n79, n137, n145);
xor  g213 (n242, n47, n49, n103, n113);
xor  g214 (n241, n135, n65, n129, n87);
nor  g215 (n226, n47, n80, n106, n46);
or   g216 (n188, n48, n109, n85, n74);
xor  g217 (n238, n129, n147, n79, n57);
or   g218 (n198, n134, n140, n74, n94);
and  g219 (n178, n53, n125, n109, n68);
nor  g220 (n255, n204, n199, n171, n166);
xor  g221 (n250, n185, n120, n187, n167);
xor  g222 (n257, n183, n121, n150, n180);
nand g223 (n260, n121, n160, n118, n120);
or   g224 (n264, n168, n173, n205, n120);
nor  g225 (n251, n149, n184, n179, n174);
nand g226 (n266, n159, n152, n119, n155);
nor  g227 (n253, n172, n182, n203, n151);
nand g228 (n265, n177, n198, n197, n200);
nor  g229 (n259, n190, n119, n162, n206);
or   g230 (n263, n201, n119, n118, n164);
xor  g231 (n256, n161, n207, n153, n121);
nor  g232 (n254, n196, n194, n175, n202);
nor  g233 (n249, n163, n154, n188, n191);
xnor g234 (n262, n193, n119, n157, n158);
and  g235 (n261, n156, n165, n170, n120);
xnor g236 (n258, n192, n169, n178, n181);
nand g237 (n252, n189, n176, n186, n195);
nor  g238 (n276, n239, n211, n233, n250);
xor  g239 (n280, n231, n258, n236, n123);
nor  g240 (n281, n209, n253, n224, n234);
nand g241 (n282, n242, n266, n122);
nor  g242 (n277, n216, n251, n249, n208);
and  g243 (n269, n210, n227, n263, n246);
xnor g244 (n272, n232, n121, n123);
nor  g245 (n268, n237, n240, n256, n247);
and  g246 (n270, n254, n122, n264, n217);
nand g247 (n273, n228, n257, n212, n226);
and  g248 (n283, n265, n260, n219, n243);
nand g249 (n279, n241, n238, n220, n235);
xor  g250 (n274, n215, n259, n261, n218);
nor  g251 (n271, n222, n214, n122, n262);
xnor g252 (n278, n223, n255, n252, n230);
nand g253 (n267, n123, n225, n229, n221);
or   g254 (n275, n248, n213, n245, n244);
endmodule
