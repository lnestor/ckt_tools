

module Stat_1090_13_7
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n951,
  n954,
  n967,
  n936,
  n985,
  n995,
  n1087,
  n1086,
  n1085,
  n1079,
  n1073,
  n1092,
  n1093,
  n1094,
  n1100,
  n1098,
  n1110,
  n1113,
  n1114,
  n1111,
  n1112,
  n1109,
  n1115
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n951;output n954;output n967;output n936;output n985;output n995;output n1087;output n1086;output n1085;output n1079;output n1073;output n1092;output n1093;output n1094;output n1100;output n1098;output n1110;output n1113;output n1114;output n1111;output n1112;output n1109;output n1115;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n952;wire n953;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1088;wire n1089;wire n1090;wire n1091;wire n1095;wire n1096;wire n1097;wire n1099;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  not
  g0
  (
    n64,
    n14
  );


  buf
  g1
  (
    n55,
    n10
  );


  buf
  g2
  (
    n91,
    n12
  );


  not
  g3
  (
    n81,
    n2
  );


  not
  g4
  (
    n29,
    n8
  );


  not
  g5
  (
    n67,
    n15
  );


  not
  g6
  (
    n70,
    n17
  );


  not
  g7
  (
    n96,
    n19
  );


  buf
  g8
  (
    n60,
    n21
  );


  buf
  g9
  (
    n74,
    n15
  );


  buf
  g10
  (
    n109,
    n12
  );


  not
  g11
  (
    n101,
    n18
  );


  buf
  g12
  (
    n28,
    n4
  );


  not
  g13
  (
    n43,
    n18
  );


  not
  g14
  (
    n31,
    n4
  );


  buf
  g15
  (
    n41,
    n8
  );


  buf
  g16
  (
    KeyWire_0_63,
    n20
  );


  not
  g17
  (
    n52,
    n10
  );


  buf
  g18
  (
    n45,
    n16
  );


  buf
  g19
  (
    n59,
    n6
  );


  not
  g20
  (
    n88,
    n15
  );


  buf
  g21
  (
    n89,
    n3
  );


  buf
  g22
  (
    n75,
    n14
  );


  buf
  g23
  (
    KeyWire_0_40,
    n13
  );


  not
  g24
  (
    n39,
    n11
  );


  not
  g25
  (
    n26,
    n19
  );


  not
  g26
  (
    n76,
    n13
  );


  not
  g27
  (
    n40,
    n20
  );


  not
  g28
  (
    n83,
    n16
  );


  not
  g29
  (
    n87,
    n9
  );


  not
  g30
  (
    n35,
    n5
  );


  not
  g31
  (
    n48,
    n3
  );


  buf
  g32
  (
    n38,
    n22
  );


  buf
  g33
  (
    KeyWire_0_14,
    n18
  );


  buf
  g34
  (
    n42,
    n13
  );


  buf
  g35
  (
    n102,
    n1
  );


  not
  g36
  (
    n63,
    n6
  );


  not
  g37
  (
    n69,
    n17
  );


  buf
  g38
  (
    n84,
    n17
  );


  buf
  g39
  (
    n90,
    n7
  );


  not
  g40
  (
    n92,
    n8
  );


  buf
  g41
  (
    n95,
    n3
  );


  buf
  g42
  (
    n51,
    n4
  );


  not
  g43
  (
    n106,
    n14
  );


  not
  g44
  (
    n80,
    n18
  );


  not
  g45
  (
    n54,
    n19
  );


  not
  g46
  (
    n108,
    n2
  );


  buf
  g47
  (
    n94,
    n4
  );


  not
  g48
  (
    n103,
    n5
  );


  buf
  g49
  (
    n62,
    n9
  );


  not
  g50
  (
    n68,
    n21
  );


  buf
  g51
  (
    n72,
    n11
  );


  buf
  g52
  (
    n78,
    n9
  );


  buf
  g53
  (
    n93,
    n20
  );


  buf
  g54
  (
    n27,
    n10
  );


  not
  g55
  (
    KeyWire_0_22,
    n5
  );


  buf
  g56
  (
    n105,
    n19
  );


  buf
  g57
  (
    n37,
    n7
  );


  not
  g58
  (
    n46,
    n21
  );


  not
  g59
  (
    n71,
    n16
  );


  buf
  g60
  (
    n53,
    n3
  );


  buf
  g61
  (
    n82,
    n14
  );


  buf
  g62
  (
    n66,
    n21
  );


  buf
  g63
  (
    n50,
    n2
  );


  buf
  g64
  (
    n100,
    n16
  );


  buf
  g65
  (
    n65,
    n5
  );


  not
  g66
  (
    n49,
    n17
  );


  not
  g67
  (
    n44,
    n13
  );


  buf
  g68
  (
    n98,
    n15
  );


  not
  g69
  (
    n61,
    n7
  );


  buf
  g70
  (
    n79,
    n11
  );


  not
  g71
  (
    n73,
    n11
  );


  buf
  g72
  (
    n86,
    n8
  );


  buf
  g73
  (
    n32,
    n12
  );


  not
  g74
  (
    n57,
    n10
  );


  buf
  g75
  (
    n107,
    n7
  );


  not
  g76
  (
    n97,
    n9
  );


  not
  g77
  (
    n34,
    n2
  );


  not
  g78
  (
    n36,
    n20
  );


  not
  g79
  (
    n104,
    n12
  );


  buf
  g80
  (
    n30,
    n6
  );


  buf
  g81
  (
    n77,
    n1
  );


  buf
  g82
  (
    n33,
    n6
  );


  not
  g83
  (
    KeyWire_0_0,
    n1
  );


  buf
  g84
  (
    n172,
    n73
  );


  buf
  g85
  (
    n121,
    n24
  );


  buf
  g86
  (
    n187,
    n52
  );


  buf
  g87
  (
    n242,
    n35
  );


  not
  g88
  (
    n130,
    n56
  );


  not
  g89
  (
    n211,
    n33
  );


  buf
  g90
  (
    n258,
    n31
  );


  not
  g91
  (
    n301,
    n70
  );


  not
  g92
  (
    n192,
    n23
  );


  not
  g93
  (
    n141,
    n80
  );


  not
  g94
  (
    n292,
    n85
  );


  buf
  g95
  (
    KeyWire_0_24,
    n36
  );


  buf
  g96
  (
    n336,
    n88
  );


  not
  g97
  (
    n383,
    n95
  );


  not
  g98
  (
    n218,
    n59
  );


  not
  g99
  (
    n164,
    n73
  );


  buf
  g100
  (
    n232,
    n97
  );


  buf
  g101
  (
    KeyWire_0_53,
    n75
  );


  buf
  g102
  (
    n354,
    n81
  );


  buf
  g103
  (
    n436,
    n62
  );


  buf
  g104
  (
    n363,
    n87
  );


  buf
  g105
  (
    n259,
    n29
  );


  buf
  g106
  (
    n120,
    n53
  );


  buf
  g107
  (
    n197,
    n45
  );


  not
  g108
  (
    n288,
    n90
  );


  buf
  g109
  (
    n163,
    n33
  );


  not
  g110
  (
    n158,
    n73
  );


  not
  g111
  (
    n352,
    n62
  );


  not
  g112
  (
    n305,
    n48
  );


  buf
  g113
  (
    n329,
    n43
  );


  buf
  g114
  (
    n405,
    n87
  );


  buf
  g115
  (
    n194,
    n49
  );


  not
  g116
  (
    KeyWire_0_61,
    n89
  );


  buf
  g117
  (
    n170,
    n107
  );


  buf
  g118
  (
    KeyWire_0_3,
    n70
  );


  buf
  g119
  (
    n411,
    n29
  );


  not
  g120
  (
    n342,
    n50
  );


  not
  g121
  (
    n359,
    n86
  );


  buf
  g122
  (
    n313,
    n25
  );


  not
  g123
  (
    n371,
    n65
  );


  not
  g124
  (
    n268,
    n53
  );


  buf
  g125
  (
    n204,
    n62
  );


  not
  g126
  (
    KeyWire_0_49,
    n40
  );


  buf
  g127
  (
    n413,
    n53
  );


  buf
  g128
  (
    n118,
    n101
  );


  not
  g129
  (
    n429,
    n92
  );


  buf
  g130
  (
    n189,
    n79
  );


  buf
  g131
  (
    n276,
    n104
  );


  buf
  g132
  (
    n403,
    n93
  );


  not
  g133
  (
    n417,
    n86
  );


  not
  g134
  (
    n262,
    n59
  );


  not
  g135
  (
    n392,
    n36
  );


  not
  g136
  (
    KeyWire_0_43,
    n92
  );


  not
  g137
  (
    n142,
    n107
  );


  not
  g138
  (
    n186,
    n102
  );


  buf
  g139
  (
    n249,
    n81
  );


  buf
  g140
  (
    n365,
    n34
  );


  buf
  g141
  (
    n364,
    n31
  );


  buf
  g142
  (
    n202,
    n81
  );


  not
  g143
  (
    n348,
    n108
  );


  buf
  g144
  (
    KeyWire_0_41,
    n61
  );


  not
  g145
  (
    n428,
    n64
  );


  not
  g146
  (
    n122,
    n27
  );


  buf
  g147
  (
    n227,
    n42
  );


  buf
  g148
  (
    n291,
    n23
  );


  not
  g149
  (
    n302,
    n76
  );


  not
  g150
  (
    n128,
    n91
  );


  not
  g151
  (
    n331,
    n68
  );


  not
  g152
  (
    n117,
    n35
  );


  not
  g153
  (
    n287,
    n107
  );


  not
  g154
  (
    n212,
    n84
  );


  buf
  g155
  (
    n221,
    n94
  );


  buf
  g156
  (
    n119,
    n65
  );


  buf
  g157
  (
    n399,
    n60
  );


  not
  g158
  (
    n401,
    n34
  );


  buf
  g159
  (
    n112,
    n44
  );


  not
  g160
  (
    n304,
    n45
  );


  not
  g161
  (
    n433,
    n48
  );


  buf
  g162
  (
    n349,
    n86
  );


  buf
  g163
  (
    n230,
    n49
  );


  not
  g164
  (
    n239,
    n65
  );


  not
  g165
  (
    n283,
    n103
  );


  not
  g166
  (
    n214,
    n80
  );


  not
  g167
  (
    n271,
    n105
  );


  not
  g168
  (
    n357,
    n90
  );


  buf
  g169
  (
    n254,
    n39
  );


  not
  g170
  (
    n312,
    n49
  );


  buf
  g171
  (
    n133,
    n63
  );


  not
  g172
  (
    KeyWire_0_33,
    n95
  );


  buf
  g173
  (
    n224,
    n91
  );


  buf
  g174
  (
    n394,
    n28
  );


  buf
  g175
  (
    n309,
    n34
  );


  not
  g176
  (
    n389,
    n27
  );


  not
  g177
  (
    n184,
    n66
  );


  not
  g178
  (
    n215,
    n57
  );


  buf
  g179
  (
    n185,
    n54
  );


  not
  g180
  (
    n270,
    n34
  );


  buf
  g181
  (
    n297,
    n91
  );


  buf
  g182
  (
    n422,
    n102
  );


  not
  g183
  (
    n387,
    n46
  );


  buf
  g184
  (
    n161,
    n48
  );


  not
  g185
  (
    n370,
    n101
  );


  buf
  g186
  (
    KeyWire_0_30,
    n72
  );


  buf
  g187
  (
    n223,
    n78
  );


  not
  g188
  (
    n293,
    n105
  );


  buf
  g189
  (
    n376,
    n72
  );


  buf
  g190
  (
    n355,
    n67
  );


  buf
  g191
  (
    KeyWire_0_12,
    n61
  );


  not
  g192
  (
    n162,
    n77
  );


  not
  g193
  (
    n379,
    n39
  );


  not
  g194
  (
    n265,
    n32
  );


  buf
  g195
  (
    n237,
    n57
  );


  not
  g196
  (
    n166,
    n107
  );


  buf
  g197
  (
    n177,
    n94
  );


  not
  g198
  (
    n139,
    n26
  );


  buf
  g199
  (
    n395,
    n33
  );


  buf
  g200
  (
    n295,
    n82
  );


  not
  g201
  (
    n191,
    n95
  );


  buf
  g202
  (
    n248,
    n46
  );


  not
  g203
  (
    n427,
    n95
  );


  buf
  g204
  (
    n437,
    n41
  );


  not
  g205
  (
    n135,
    n100
  );


  not
  g206
  (
    n154,
    n71
  );


  buf
  g207
  (
    n247,
    n94
  );


  not
  g208
  (
    n178,
    n45
  );


  not
  g209
  (
    n384,
    n85
  );


  buf
  g210
  (
    n425,
    n83
  );


  buf
  g211
  (
    n386,
    n38
  );


  not
  g212
  (
    n207,
    n30
  );


  not
  g213
  (
    n334,
    n100
  );


  not
  g214
  (
    n374,
    n76
  );


  buf
  g215
  (
    n200,
    n104
  );


  not
  g216
  (
    n243,
    n73
  );


  buf
  g217
  (
    n167,
    n67
  );


  buf
  g218
  (
    n323,
    n63
  );


  buf
  g219
  (
    n285,
    n53
  );


  not
  g220
  (
    n426,
    n38
  );


  buf
  g221
  (
    n367,
    n106
  );


  not
  g222
  (
    n203,
    n68
  );


  buf
  g223
  (
    n174,
    n88
  );


  not
  g224
  (
    n353,
    n32
  );


  buf
  g225
  (
    n165,
    n69
  );


  not
  g226
  (
    n372,
    n46
  );


  buf
  g227
  (
    n205,
    n51
  );


  buf
  g228
  (
    n114,
    n98
  );


  not
  g229
  (
    n321,
    n36
  );


  buf
  g230
  (
    n303,
    n59
  );


  buf
  g231
  (
    n144,
    n28
  );


  buf
  g232
  (
    n256,
    n45
  );


  not
  g233
  (
    n198,
    n94
  );


  not
  g234
  (
    n216,
    n96
  );


  not
  g235
  (
    n327,
    n74
  );


  buf
  g236
  (
    n421,
    n108
  );


  buf
  g237
  (
    n317,
    n24
  );


  not
  g238
  (
    n281,
    n50
  );


  not
  g239
  (
    n308,
    n96
  );


  buf
  g240
  (
    n113,
    n83
  );


  buf
  g241
  (
    n140,
    n77
  );


  buf
  g242
  (
    n275,
    n71
  );


  not
  g243
  (
    n181,
    n83
  );


  buf
  g244
  (
    n241,
    n47
  );


  not
  g245
  (
    n326,
    n57
  );


  not
  g246
  (
    n390,
    n63
  );


  buf
  g247
  (
    KeyWire_0_57,
    n50
  );


  not
  g248
  (
    n388,
    n29
  );


  buf
  g249
  (
    KeyWire_0_13,
    n41
  );


  buf
  g250
  (
    n277,
    n93
  );


  not
  g251
  (
    n252,
    n43
  );


  buf
  g252
  (
    n307,
    n106
  );


  not
  g253
  (
    n233,
    n106
  );


  not
  g254
  (
    n138,
    n89
  );


  buf
  g255
  (
    n123,
    n69
  );


  not
  g256
  (
    n201,
    n26
  );


  not
  g257
  (
    n410,
    n75
  );


  buf
  g258
  (
    n406,
    n88
  );


  buf
  g259
  (
    n182,
    n56
  );


  buf
  g260
  (
    n314,
    n54
  );


  not
  g261
  (
    n324,
    n98
  );


  buf
  g262
  (
    n335,
    n64
  );


  not
  g263
  (
    n257,
    n39
  );


  not
  g264
  (
    n393,
    n74
  );


  buf
  g265
  (
    n131,
    n89
  );


  not
  g266
  (
    n213,
    n79
  );


  not
  g267
  (
    KeyWire_0_35,
    n48
  );


  buf
  g268
  (
    n377,
    n42
  );


  buf
  g269
  (
    n378,
    n99
  );


  buf
  g270
  (
    n206,
    n65
  );


  buf
  g271
  (
    n346,
    n58
  );


  buf
  g272
  (
    n310,
    n44
  );


  buf
  g273
  (
    KeyWire_0_58,
    n31
  );


  not
  g274
  (
    n136,
    n44
  );


  not
  g275
  (
    n290,
    n40
  );


  buf
  g276
  (
    n273,
    n49
  );


  not
  g277
  (
    n199,
    n82
  );


  not
  g278
  (
    n263,
    n51
  );


  buf
  g279
  (
    n345,
    n35
  );


  not
  g280
  (
    n325,
    n77
  );


  buf
  g281
  (
    n255,
    n52
  );


  not
  g282
  (
    n408,
    n76
  );


  buf
  g283
  (
    n173,
    n44
  );


  not
  g284
  (
    n179,
    n30
  );


  not
  g285
  (
    n315,
    n103
  );


  buf
  g286
  (
    n362,
    n93
  );


  buf
  g287
  (
    KeyWire_0_9,
    n64
  );


  not
  g288
  (
    n398,
    n23
  );


  not
  g289
  (
    n298,
    n79
  );


  buf
  g290
  (
    n402,
    n37
  );


  not
  g291
  (
    n296,
    n57
  );


  buf
  g292
  (
    n366,
    n96
  );


  not
  g293
  (
    n391,
    n28
  );


  buf
  g294
  (
    n344,
    n76
  );


  not
  g295
  (
    n412,
    n75
  );


  buf
  g296
  (
    n407,
    n37
  );


  not
  g297
  (
    n280,
    n42
  );


  buf
  g298
  (
    n409,
    n33
  );


  buf
  g299
  (
    n320,
    n87
  );


  not
  g300
  (
    n209,
    n24
  );


  not
  g301
  (
    n127,
    n56
  );


  buf
  g302
  (
    KeyWire_0_54,
    n41
  );


  not
  g303
  (
    n196,
    n61
  );


  buf
  g304
  (
    n319,
    n104
  );


  not
  g305
  (
    n152,
    n58
  );


  buf
  g306
  (
    n111,
    n37
  );


  buf
  g307
  (
    n159,
    n30
  );


  buf
  g308
  (
    n217,
    n27
  );


  buf
  g309
  (
    KeyWire_0_59,
    n71
  );


  buf
  g310
  (
    n322,
    n38
  );


  buf
  g311
  (
    n183,
    n41
  );


  not
  g312
  (
    n339,
    n83
  );


  buf
  g313
  (
    n431,
    n46
  );


  buf
  g314
  (
    n245,
    n97
  );


  not
  g315
  (
    n382,
    n42
  );


  not
  g316
  (
    n385,
    n24
  );


  not
  g317
  (
    n125,
    n99
  );


  buf
  g318
  (
    n361,
    n92
  );


  not
  g319
  (
    n358,
    n75
  );


  buf
  g320
  (
    n150,
    n103
  );


  buf
  g321
  (
    n396,
    n66
  );


  not
  g322
  (
    n360,
    n61
  );


  buf
  g323
  (
    n253,
    n100
  );


  not
  g324
  (
    n286,
    n69
  );


  buf
  g325
  (
    n330,
    n40
  );


  buf
  g326
  (
    n147,
    n78
  );


  buf
  g327
  (
    n180,
    n103
  );


  not
  g328
  (
    n251,
    n101
  );


  buf
  g329
  (
    n343,
    n99
  );


  not
  g330
  (
    n225,
    n50
  );


  not
  g331
  (
    KeyWire_0_17,
    n55
  );


  buf
  g332
  (
    n333,
    n100
  );


  not
  g333
  (
    n340,
    n106
  );


  buf
  g334
  (
    n278,
    n105
  );


  buf
  g335
  (
    n356,
    n52
  );


  buf
  g336
  (
    n146,
    n31
  );


  buf
  g337
  (
    n414,
    n97
  );


  not
  g338
  (
    n210,
    n80
  );


  not
  g339
  (
    n126,
    n56
  );


  buf
  g340
  (
    n220,
    n36
  );


  buf
  g341
  (
    n226,
    n60
  );


  not
  g342
  (
    n300,
    n30
  );


  buf
  g343
  (
    n155,
    n40
  );


  buf
  g344
  (
    n190,
    n38
  );


  not
  g345
  (
    n351,
    n85
  );


  not
  g346
  (
    n228,
    n82
  );


  not
  g347
  (
    n124,
    n68
  );


  buf
  g348
  (
    n350,
    n82
  );


  buf
  g349
  (
    n229,
    n63
  );


  buf
  g350
  (
    n269,
    n32
  );


  not
  g351
  (
    n416,
    n59
  );


  not
  g352
  (
    n264,
    n47
  );


  buf
  g353
  (
    n188,
    n26
  );


  buf
  g354
  (
    n424,
    n78
  );


  buf
  g355
  (
    n435,
    n58
  );


  not
  g356
  (
    n420,
    n98
  );


  not
  g357
  (
    KeyWire_0_31,
    n22
  );


  not
  g358
  (
    n267,
    n23
  );


  not
  g359
  (
    n438,
    n64
  );


  buf
  g360
  (
    n132,
    n104
  );


  buf
  g361
  (
    n260,
    n22
  );


  buf
  g362
  (
    n168,
    n81
  );


  not
  g363
  (
    n160,
    n80
  );


  not
  g364
  (
    n116,
    n52
  );


  buf
  g365
  (
    n115,
    n84
  );


  not
  g366
  (
    n231,
    n79
  );


  not
  g367
  (
    n151,
    n101
  );


  buf
  g368
  (
    n261,
    n86
  );


  not
  g369
  (
    n397,
    n96
  );


  buf
  g370
  (
    n208,
    n37
  );


  not
  g371
  (
    n432,
    n77
  );


  not
  g372
  (
    n419,
    n22
  );


  not
  g373
  (
    n418,
    n60
  );


  not
  g374
  (
    n272,
    n62
  );


  not
  g375
  (
    n415,
    n67
  );


  not
  g376
  (
    n153,
    n66
  );


  not
  g377
  (
    n246,
    n25
  );


  not
  g378
  (
    KeyWire_0_10,
    n28
  );


  buf
  g379
  (
    n318,
    n105
  );


  buf
  g380
  (
    n157,
    n39
  );


  buf
  g381
  (
    n240,
    n87
  );


  not
  g382
  (
    KeyWire_0_11,
    n93
  );


  not
  g383
  (
    n222,
    n88
  );


  not
  g384
  (
    n328,
    n29
  );


  not
  g385
  (
    n373,
    n66
  );


  not
  g386
  (
    n404,
    n51
  );


  not
  g387
  (
    n234,
    n74
  );


  not
  g388
  (
    n156,
    n90
  );


  buf
  g389
  (
    n193,
    n55
  );


  buf
  g390
  (
    KeyWire_0_44,
    n47
  );


  buf
  g391
  (
    n380,
    n67
  );


  buf
  g392
  (
    n434,
    n60
  );


  not
  g393
  (
    n284,
    n35
  );


  buf
  g394
  (
    n143,
    n72
  );


  buf
  g395
  (
    n238,
    n69
  );


  buf
  g396
  (
    n368,
    n58
  );


  buf
  g397
  (
    n176,
    n43
  );


  not
  g398
  (
    n381,
    n47
  );


  not
  g399
  (
    KeyWire_0_19,
    n89
  );


  xor
  g400
  (
    n299,
    n70,
    n84
  );


  nor
  g401
  (
    n134,
    n84,
    n68
  );


  xor
  g402
  (
    n306,
    n91,
    n26
  );


  and
  g403
  (
    n235,
    n90,
    n70
  );


  xnor
  g404
  (
    n338,
    n102,
    n97
  );


  xor
  g405
  (
    n369,
    n54,
    n55
  );


  or
  g406
  (
    n244,
    n32,
    n25
  );


  or
  g407
  (
    n169,
    n72,
    n27
  );


  xnor
  g408
  (
    n219,
    n78,
    n92
  );


  nor
  g409
  (
    n375,
    n85,
    n71
  );


  and
  g410
  (
    n423,
    n102,
    n54
  );


  xor
  g411
  (
    n110,
    n55,
    n98
  );


  and
  g412
  (
    n332,
    n51,
    n99
  );


  xnor
  g413
  (
    n171,
    n43,
    n74
  );


  buf
  g414
  (
    n482,
    n122
  );


  not
  g415
  (
    n499,
    n142
  );


  buf
  g416
  (
    n444,
    n119
  );


  buf
  g417
  (
    n502,
    n113
  );


  not
  g418
  (
    n442,
    n133
  );


  not
  g419
  (
    n460,
    n115
  );


  buf
  g420
  (
    n491,
    n114
  );


  not
  g421
  (
    n480,
    n115
  );


  buf
  g422
  (
    n454,
    n124
  );


  not
  g423
  (
    n500,
    n116
  );


  not
  g424
  (
    n488,
    n121
  );


  buf
  g425
  (
    n457,
    n138
  );


  buf
  g426
  (
    n472,
    n124
  );


  buf
  g427
  (
    n504,
    n128
  );


  buf
  g428
  (
    n485,
    n125
  );


  buf
  g429
  (
    n450,
    n109
  );


  buf
  g430
  (
    n486,
    n136
  );


  buf
  g431
  (
    n503,
    n118
  );


  not
  g432
  (
    n497,
    n133
  );


  not
  g433
  (
    n456,
    n129
  );


  not
  g434
  (
    n459,
    n131
  );


  buf
  g435
  (
    KeyWire_0_60,
    n136
  );


  buf
  g436
  (
    n467,
    n139
  );


  buf
  g437
  (
    n473,
    n117
  );


  buf
  g438
  (
    n496,
    n132
  );


  not
  g439
  (
    n477,
    n141
  );


  not
  g440
  (
    n483,
    n132
  );


  not
  g441
  (
    n458,
    n110
  );


  buf
  g442
  (
    n447,
    n118
  );


  buf
  g443
  (
    n495,
    n135
  );


  not
  g444
  (
    n484,
    n135
  );


  not
  g445
  (
    n498,
    n108
  );


  not
  g446
  (
    n466,
    n142
  );


  buf
  g447
  (
    n481,
    n117
  );


  not
  g448
  (
    n445,
    n123
  );


  buf
  g449
  (
    n505,
    n112
  );


  buf
  g450
  (
    n501,
    n120
  );


  buf
  g451
  (
    n479,
    n126
  );


  not
  g452
  (
    n474,
    n140
  );


  buf
  g453
  (
    n494,
    n141
  );


  buf
  g454
  (
    n471,
    n130
  );


  buf
  g455
  (
    n443,
    n139
  );


  buf
  g456
  (
    n493,
    n125
  );


  not
  g457
  (
    n455,
    n111
  );


  not
  g458
  (
    n478,
    n143
  );


  buf
  g459
  (
    KeyWire_0_16,
    n128
  );


  buf
  g460
  (
    n464,
    n134
  );


  not
  g461
  (
    n440,
    n112
  );


  buf
  g462
  (
    n453,
    n127
  );


  buf
  g463
  (
    n451,
    n122
  );


  not
  g464
  (
    n452,
    n137
  );


  not
  g465
  (
    KeyWire_0_39,
    n108
  );


  not
  g466
  (
    n461,
    n110
  );


  buf
  g467
  (
    n475,
    n123
  );


  not
  g468
  (
    n468,
    n109
  );


  not
  g469
  (
    n476,
    n114
  );


  buf
  g470
  (
    n490,
    n109
  );


  buf
  g471
  (
    n489,
    n121
  );


  buf
  g472
  (
    n492,
    n119
  );


  buf
  g473
  (
    n449,
    n111
  );


  buf
  g474
  (
    n470,
    n129
  );


  buf
  g475
  (
    n448,
    n109
  );


  not
  g476
  (
    n487,
    n116
  );


  buf
  g477
  (
    n507,
    n143
  );


  not
  g478
  (
    n446,
    n120
  );


  not
  g479
  (
    n441,
    n127
  );


  xor
  g480
  (
    n462,
    n131,
    n130,
    n138,
    n137
  );


  xnor
  g481
  (
    n506,
    n126,
    n140,
    n134,
    n113
  );


  and
  g482
  (
    n548,
    n227,
    n307,
    n258,
    n409
  );


  xnor
  g483
  (
    n626,
    n235,
    n322,
    n418,
    n165
  );


  xnor
  g484
  (
    n617,
    n417,
    n386,
    n346,
    n352
  );


  nand
  g485
  (
    n533,
    n155,
    n471,
    n246,
    n166
  );


  xor
  g486
  (
    n602,
    n190,
    n212,
    n159,
    n298
  );


  and
  g487
  (
    n607,
    n491,
    n222,
    n488,
    n228
  );


  nor
  g488
  (
    n714,
    n195,
    n366,
    n324,
    n394
  );


  and
  g489
  (
    n555,
    n471,
    n453,
    n473,
    n443
  );


  nor
  g490
  (
    KeyWire_0_1,
    n384,
    n280,
    n468,
    n452
  );


  xnor
  g491
  (
    n733,
    n180,
    n254,
    n372,
    n337
  );


  xnor
  g492
  (
    n690,
    n461,
    n314,
    n453,
    n457
  );


  nand
  g493
  (
    n509,
    n460,
    n171,
    n243,
    n175
  );


  nor
  g494
  (
    n670,
    n236,
    n155,
    n207,
    n405
  );


  nor
  g495
  (
    n575,
    n358,
    n300,
    n475,
    n466
  );


  and
  g496
  (
    n698,
    n460,
    n172,
    n189,
    n430
  );


  xor
  g497
  (
    n673,
    n451,
    n410,
    n496,
    n428
  );


  nor
  g498
  (
    n539,
    n371,
    n360,
    n467,
    n466
  );


  nand
  g499
  (
    n537,
    n448,
    n163,
    n276,
    n259
  );


  nor
  g500
  (
    n619,
    n398,
    n450,
    n286,
    n338
  );


  nand
  g501
  (
    n734,
    n198,
    n409,
    n260,
    n383
  );


  nand
  g502
  (
    n717,
    n177,
    n216,
    n387,
    n462
  );


  and
  g503
  (
    n701,
    n446,
    n476,
    n203,
    n422
  );


  nand
  g504
  (
    n597,
    n198,
    n272,
    n491,
    n154
  );


  and
  g505
  (
    n586,
    n441,
    n239,
    n334,
    n292
  );


  xnor
  g506
  (
    n572,
    n334,
    n443,
    n458,
    n424
  );


  xor
  g507
  (
    n704,
    n360,
    n421,
    n230,
    n486
  );


  xnor
  g508
  (
    n629,
    n371,
    n270,
    n174,
    n251
  );


  nor
  g509
  (
    n579,
    n409,
    n431,
    n379,
    n484
  );


  nor
  g510
  (
    n527,
    n178,
    n246,
    n395,
    n413
  );


  xnor
  g511
  (
    n729,
    n458,
    n255,
    n238,
    n332
  );


  xnor
  g512
  (
    n695,
    n197,
    n390,
    n209,
    n274
  );


  nor
  g513
  (
    n663,
    n472,
    n267,
    n367,
    n369
  );


  and
  g514
  (
    n675,
    n312,
    n442,
    n192,
    n456
  );


  xor
  g515
  (
    n551,
    n268,
    n263,
    n182,
    n399
  );


  xor
  g516
  (
    n642,
    n464,
    n189,
    n492,
    n465
  );


  xor
  g517
  (
    n705,
    n437,
    n318,
    n366,
    n497
  );


  or
  g518
  (
    n620,
    n384,
    n469,
    n414,
    n495
  );


  xnor
  g519
  (
    n563,
    n435,
    n384,
    n214,
    n221
  );


  nand
  g520
  (
    n712,
    n295,
    n417,
    n343,
    n487
  );


  xor
  g521
  (
    n651,
    n214,
    n380,
    n341
  );


  xnor
  g522
  (
    n656,
    n496,
    n422,
    n363,
    n485
  );


  nor
  g523
  (
    n638,
    n277,
    n206,
    n406,
    n209
  );


  nor
  g524
  (
    n585,
    n263,
    n450,
    n358,
    n422
  );


  nand
  g525
  (
    n599,
    n160,
    n475,
    n474,
    n248
  );


  xor
  g526
  (
    n685,
    n347,
    n336,
    n361,
    n230
  );


  xor
  g527
  (
    n576,
    n237,
    n388,
    n397,
    n419
  );


  xnor
  g528
  (
    n595,
    n204,
    n433,
    n311,
    n298
  );


  or
  g529
  (
    n552,
    n290,
    n389,
    n297,
    n277
  );


  and
  g530
  (
    n636,
    n495,
    n252,
    n481,
    n434
  );


  xor
  g531
  (
    n513,
    n250,
    n306,
    n441,
    n329
  );


  and
  g532
  (
    n658,
    n431,
    n483,
    n396,
    n356
  );


  xor
  g533
  (
    n627,
    n316,
    n382,
    n393,
    n491
  );


  or
  g534
  (
    n664,
    n375,
    n447,
    n220,
    n436
  );


  nand
  g535
  (
    KeyWire_0_18,
    n188,
    n259,
    n467,
    n368
  );


  or
  g536
  (
    n657,
    n219,
    n479,
    n380,
    n382
  );


  nand
  g537
  (
    n708,
    n478,
    n378,
    n161,
    n302
  );


  nor
  g538
  (
    n574,
    n335,
    n428,
    n351,
    n412
  );


  xnor
  g539
  (
    n608,
    n266,
    n185,
    n483,
    n370
  );


  xnor
  g540
  (
    n732,
    n315,
    n370,
    n455,
    n487
  );


  nand
  g541
  (
    n573,
    n358,
    n420,
    n157,
    n309
  );


  nand
  g542
  (
    n672,
    n423,
    n410,
    n448,
    n355
  );


  and
  g543
  (
    n542,
    n497,
    n221,
    n289,
    n449
  );


  xnor
  g544
  (
    KeyWire_0_47,
    n168,
    n229,
    n248,
    n428
  );


  xnor
  g545
  (
    n707,
    n301,
    n477,
    n284,
    n196
  );


  xor
  g546
  (
    n588,
    n485,
    n425,
    n351,
    n434
  );


  nand
  g547
  (
    n535,
    n270,
    n478,
    n442,
    n488
  );


  xnor
  g548
  (
    n655,
    n425,
    n476,
    n232,
    n379
  );


  nor
  g549
  (
    n521,
    n321,
    n394,
    n393,
    n454
  );


  nand
  g550
  (
    n606,
    n323,
    n415,
    n276,
    n336
  );


  nand
  g551
  (
    n616,
    n378,
    n383,
    n457,
    n473
  );


  xor
  g552
  (
    n697,
    n279,
    n333,
    n427,
    n493
  );


  xnor
  g553
  (
    n601,
    n147,
    n465,
    n493,
    n237
  );


  nand
  g554
  (
    n603,
    n285,
    n485,
    n477,
    n296
  );


  or
  g555
  (
    n643,
    n441,
    n399,
    n311,
    n426
  );


  or
  g556
  (
    n534,
    n164,
    n258,
    n326,
    n145
  );


  or
  g557
  (
    n683,
    n498,
    n245,
    n327,
    n308
  );


  nand
  g558
  (
    n634,
    n357,
    n151,
    n271,
    n402
  );


  nor
  g559
  (
    n684,
    n213,
    n443,
    n491,
    n279
  );


  nor
  g560
  (
    n645,
    n448,
    n453,
    n474,
    n480
  );


  xnor
  g561
  (
    n667,
    n488,
    n240,
    n312
  );


  nor
  g562
  (
    n665,
    n226,
    n482,
    n365,
    n372
  );


  nand
  g563
  (
    n621,
    n385,
    n406,
    n355,
    n348
  );


  nand
  g564
  (
    n728,
    n355,
    n472,
    n295,
    n167
  );


  and
  g565
  (
    n578,
    n208,
    n368,
    n484,
    n217
  );


  xnor
  g566
  (
    n727,
    n187,
    n173,
    n405,
    n249
  );


  and
  g567
  (
    n693,
    n328,
    n323,
    n489,
    n317
  );


  or
  g568
  (
    n677,
    n364,
    n460,
    n255,
    n400
  );


  and
  g569
  (
    n522,
    n353,
    n305,
    n360,
    n345
  );


  nor
  g570
  (
    n688,
    n390,
    n353,
    n444,
    n293
  );


  nand
  g571
  (
    n565,
    n219,
    n466,
    n208,
    n374
  );


  or
  g572
  (
    n512,
    n205,
    n460,
    n404,
    n158
  );


  nand
  g573
  (
    n628,
    n367,
    n418,
    n186,
    n271
  );


  xnor
  g574
  (
    n699,
    n436,
    n391,
    n363,
    n408
  );


  nand
  g575
  (
    n646,
    n383,
    n181,
    n424,
    n249
  );


  xor
  g576
  (
    KeyWire_0_20,
    n474,
    n199,
    n462,
    n241
  );


  and
  g577
  (
    KeyWire_0_46,
    n193,
    n188,
    n345,
    n365
  );


  xor
  g578
  (
    n523,
    n195,
    n490,
    n454,
    n257
  );


  xnor
  g579
  (
    n584,
    n477,
    n468,
    n315,
    n410
  );


  and
  g580
  (
    n709,
    n373,
    n456,
    n467,
    n375
  );


  or
  g581
  (
    n583,
    n496,
    n469,
    n166,
    n305
  );


  xor
  g582
  (
    n520,
    n185,
    n462,
    n489,
    n173
  );


  nor
  g583
  (
    n711,
    n446,
    n354,
    n339,
    n291
  );


  or
  g584
  (
    n678,
    n378,
    n256,
    n444,
    n294
  );


  nand
  g585
  (
    n696,
    n463,
    n475,
    n194,
    n450
  );


  or
  g586
  (
    n641,
    n403,
    n447,
    n152,
    n466
  );


  nand
  g587
  (
    n550,
    n223,
    n309,
    n488,
    n262
  );


  nand
  g588
  (
    n632,
    n398,
    n282,
    n180,
    n470
  );


  nand
  g589
  (
    n681,
    n341,
    n273,
    n275,
    n300
  );


  nand
  g590
  (
    n702,
    n470,
    n269,
    n416,
    n387
  );


  xnor
  g591
  (
    n553,
    n313,
    n327,
    n492,
    n342
  );


  nor
  g592
  (
    n689,
    n408,
    n447,
    n239,
    n455
  );


  nor
  g593
  (
    n682,
    n275,
    n474,
    n482,
    n478
  );


  xnor
  g594
  (
    n659,
    n423,
    n284,
    n338,
    n146
  );


  or
  g595
  (
    n605,
    n243,
    n395,
    n362,
    n350
  );


  or
  g596
  (
    n530,
    n184,
    n479,
    n339,
    n487
  );


  nand
  g597
  (
    n590,
    n489,
    n381,
    n184,
    n307
  );


  and
  g598
  (
    n631,
    n292,
    n191,
    n169,
    n144
  );


  nand
  g599
  (
    n594,
    n494,
    n303,
    n408,
    n216
  );


  xnor
  g600
  (
    n592,
    n415,
    n145,
    n200,
    n429
  );


  or
  g601
  (
    n660,
    n411,
    n423,
    n403,
    n459
  );


  or
  g602
  (
    n567,
    n201,
    n459,
    n165,
    n218
  );


  nor
  g603
  (
    n674,
    n283,
    n299,
    n459,
    n473
  );


  nand
  g604
  (
    n731,
    n494,
    n398,
    n417,
    n446
  );


  nand
  g605
  (
    n577,
    n479,
    n456,
    n233,
    n394
  );


  and
  g606
  (
    n524,
    n369,
    n446,
    n429,
    n196
  );


  nor
  g607
  (
    n547,
    n197,
    n349,
    n386,
    n396
  );


  and
  g608
  (
    n596,
    n310,
    n451,
    n485,
    n244
  );


  nor
  g609
  (
    n648,
    n340,
    n317,
    n183,
    n435
  );


  xnor
  g610
  (
    n554,
    n293,
    n489,
    n404,
    n169
  );


  xor
  g611
  (
    n723,
    n414,
    n345,
    n325,
    n273
  );


  and
  g612
  (
    n671,
    n452,
    n359,
    n306,
    n158
  );


  nor
  g613
  (
    n721,
    n178,
    n177,
    n455,
    n215
  );


  nor
  g614
  (
    n720,
    n181,
    n187,
    n340,
    n471
  );


  nand
  g615
  (
    KeyWire_0_7,
    n391,
    n391,
    n342,
    n413
  );


  nand
  g616
  (
    n730,
    n419,
    n430,
    n347,
    n242
  );


  and
  g617
  (
    n587,
    n154,
    n290,
    n401,
    n367
  );


  or
  g618
  (
    n703,
    n407,
    n234,
    n157,
    n469
  );


  xnor
  g619
  (
    n623,
    n302,
    n494,
    n463,
    n347
  );


  nand
  g620
  (
    n676,
    n244,
    n444,
    n234,
    n186
  );


  or
  g621
  (
    n679,
    n321,
    n365,
    n203,
    n457
  );


  xnor
  g622
  (
    n568,
    n151,
    n328,
    n288,
    n156
  );


  nand
  g623
  (
    n686,
    n388,
    n262,
    n356,
    n261
  );


  xnor
  g624
  (
    n538,
    n357,
    n326,
    n253,
    n418
  );


  nor
  g625
  (
    n560,
    n403,
    n433,
    n313,
    n261
  );


  xnor
  g626
  (
    n611,
    n220,
    n368,
    n250,
    n254
  );


  and
  g627
  (
    n719,
    n483,
    n150,
    n320,
    n470
  );


  xnor
  g628
  (
    n609,
    n170,
    n462,
    n236,
    n346
  );


  xor
  g629
  (
    n668,
    n395,
    n162,
    n445
  );


  xor
  g630
  (
    n716,
    n484,
    n458,
    n476,
    n294
  );


  xnor
  g631
  (
    n639,
    n411,
    n392,
    n468,
    n350
  );


  xnor
  g632
  (
    n625,
    n440,
    n372,
    n153,
    n480
  );


  nand
  g633
  (
    n581,
    n364,
    n172,
    n429,
    n451
  );


  and
  g634
  (
    n718,
    n451,
    n419,
    n264,
    n346
  );


  nor
  g635
  (
    n647,
    n461,
    n452,
    n457,
    n407
  );


  or
  g636
  (
    n680,
    n344,
    n303,
    n218,
    n393
  );


  nor
  g637
  (
    n525,
    n432,
    n217,
    n329,
    n453
  );


  nand
  g638
  (
    n564,
    n412,
    n260,
    n160,
    n389
  );


  nand
  g639
  (
    n556,
    n407,
    n150,
    n471,
    n440
  );


  xnor
  g640
  (
    n582,
    n411,
    n392,
    n448,
    n224
  );


  xnor
  g641
  (
    n528,
    n414,
    n426,
    n472,
    n454
  );


  nor
  g642
  (
    n561,
    n402,
    n445,
    n377,
    n331
  );


  nand
  g643
  (
    n591,
    n363,
    n385,
    n450,
    n228
  );


  and
  g644
  (
    n541,
    n364,
    n366,
    n447,
    n352
  );


  or
  g645
  (
    n562,
    n242,
    n374,
    n238,
    n149
  );


  and
  g646
  (
    n715,
    n392,
    n256,
    n461,
    n496
  );


  or
  g647
  (
    n543,
    n291,
    n204,
    n265,
    n373
  );


  nand
  g648
  (
    n669,
    n379,
    n473,
    n325,
    n434
  );


  nor
  g649
  (
    n508,
    n319,
    n406,
    n213,
    n486
  );


  and
  g650
  (
    n549,
    n475,
    n201,
    n421,
    n463
  );


  xnor
  g651
  (
    n624,
    n486,
    n484,
    n472,
    n490
  );


  nand
  g652
  (
    n559,
    n202,
    n426,
    n176,
    n210
  );


  nand
  g653
  (
    n516,
    n183,
    n399,
    n191,
    n229
  );


  xor
  g654
  (
    n517,
    n479,
    n331,
    n490,
    n389
  );


  and
  g655
  (
    n569,
    n330,
    n206,
    n171,
    n194
  );


  nand
  g656
  (
    n654,
    n288,
    n464,
    n495,
    n148
  );


  nor
  g657
  (
    n532,
    n163,
    n304,
    n436,
    n442
  );


  and
  g658
  (
    KeyWire_0_25,
    n387,
    n495,
    n281,
    n322
  );


  or
  g659
  (
    n630,
    n227,
    n382,
    n266,
    n476
  );


  xor
  g660
  (
    n615,
    n468,
    n352,
    n296,
    n465
  );


  nor
  g661
  (
    KeyWire_0_37,
    n224,
    n478,
    n449,
    n287
  );


  or
  g662
  (
    n598,
    n280,
    n212,
    n435,
    n497
  );


  and
  g663
  (
    n610,
    n497,
    n324,
    n350,
    n149
  );


  and
  g664
  (
    n511,
    n374,
    n304,
    n192,
    n445
  );


  and
  g665
  (
    n633,
    n480,
    n449,
    n318,
    n264
  );


  xnor
  g666
  (
    n531,
    n193,
    n467,
    n424,
    n267
  );


  or
  g667
  (
    n637,
    n354,
    n390,
    n376
  );


  or
  g668
  (
    n652,
    n148,
    n430,
    n179,
    n167
  );


  or
  g669
  (
    n518,
    n371,
    n458,
    n464,
    n356
  );


  nand
  g670
  (
    n725,
    n316,
    n175,
    n377,
    n482
  );


  nor
  g671
  (
    n713,
    n319,
    n415,
    n437,
    n349
  );


  nand
  g672
  (
    n613,
    n337,
    n153,
    n433,
    n477
  );


  xor
  g673
  (
    n600,
    n480,
    n376,
    n425,
    n152
  );


  and
  g674
  (
    n710,
    n493,
    n200,
    n357,
    n348
  );


  nand
  g675
  (
    KeyWire_0_62,
    n164,
    n274,
    n400,
    n226
  );


  xnor
  g676
  (
    n570,
    n440,
    n174,
    n452,
    n176
  );


  and
  g677
  (
    n649,
    n401,
    n247,
    n301,
    n369
  );


  xor
  g678
  (
    n724,
    n211,
    n272,
    n432,
    n421
  );


  xnor
  g679
  (
    n662,
    n146,
    n481,
    n205,
    n182
  );


  xnor
  g680
  (
    n515,
    n486,
    n483,
    n289,
    n416
  );


  xor
  g681
  (
    n589,
    n349,
    n241,
    n231,
    n225
  );


  nor
  g682
  (
    n692,
    n456,
    n487,
    n463,
    n359
  );


  xor
  g683
  (
    n546,
    n494,
    n332,
    n253,
    n490
  );


  or
  g684
  (
    n529,
    n459,
    n344,
    n493,
    n348
  );


  and
  g685
  (
    n614,
    n469,
    n375,
    n381,
    n416
  );


  xnor
  g686
  (
    n526,
    n449,
    n287,
    n335,
    n210
  );


  and
  g687
  (
    n635,
    n343,
    n354,
    n427,
    n361
  );


  nor
  g688
  (
    n514,
    n404,
    n147,
    n481,
    n297
  );


  or
  g689
  (
    n612,
    n190,
    n492,
    n359
  );


  nand
  g690
  (
    KeyWire_0_2,
    n308,
    n179,
    n373,
    n396
  );


  xnor
  g691
  (
    n726,
    n161,
    n235,
    n388,
    n233
  );


  xor
  g692
  (
    n540,
    n381,
    n257,
    n202,
    n268
  );


  xor
  g693
  (
    n661,
    n231,
    n432,
    n401,
    n370
  );


  and
  g694
  (
    n666,
    n251,
    n386,
    n420,
    n223
  );


  or
  g695
  (
    n571,
    n400,
    n431,
    n377,
    n281
  );


  or
  g696
  (
    n694,
    n144,
    n470,
    n353,
    n269
  );


  nor
  g697
  (
    n706,
    n285,
    n286,
    n252,
    n397
  );


  nand
  g698
  (
    n510,
    n314,
    n397,
    n245,
    n330
  );


  xor
  g699
  (
    n580,
    n247,
    n170,
    n278,
    n427
  );


  and
  g700
  (
    n545,
    n482,
    n412,
    n437,
    n225
  );


  or
  g701
  (
    n544,
    n405,
    n159,
    n455,
    n310
  );


  xnor
  g702
  (
    n691,
    n465,
    n351,
    n168,
    n362
  );


  and
  g703
  (
    n618,
    n207,
    n265,
    n283,
    n222
  );


  or
  g704
  (
    n687,
    n211,
    n461,
    n199,
    n464
  );


  xnor
  g705
  (
    n566,
    n413,
    n481,
    n362,
    n156
  );


  nand
  g706
  (
    n722,
    n420,
    n320,
    n282,
    n385
  );


  xor
  g707
  (
    n653,
    n215,
    n402,
    n454,
    n278
  );


  xor
  g708
  (
    n650,
    n299,
    n333,
    n361,
    n232
  );


  buf
  g709
  (
    n751,
    n552
  );


  not
  g710
  (
    n771,
    n531
  );


  buf
  g711
  (
    n806,
    n500
  );


  not
  g712
  (
    n826,
    n551
  );


  buf
  g713
  (
    n822,
    n499
  );


  not
  g714
  (
    n796,
    n594
  );


  buf
  g715
  (
    n818,
    n549
  );


  not
  g716
  (
    n799,
    n529
  );


  buf
  g717
  (
    n828,
    n540
  );


  buf
  g718
  (
    n768,
    n504
  );


  buf
  g719
  (
    KeyWire_0_34,
    n591
  );


  buf
  g720
  (
    n817,
    n572
  );


  not
  g721
  (
    n750,
    n571
  );


  buf
  g722
  (
    n765,
    n528
  );


  buf
  g723
  (
    n780,
    n559
  );


  buf
  g724
  (
    n807,
    n557
  );


  buf
  g725
  (
    n791,
    n501
  );


  buf
  g726
  (
    n821,
    n537
  );


  buf
  g727
  (
    n815,
    n592
  );


  not
  g728
  (
    n808,
    n588
  );


  buf
  g729
  (
    n805,
    n499
  );


  buf
  g730
  (
    n779,
    n595
  );


  not
  g731
  (
    n739,
    n516
  );


  not
  g732
  (
    n759,
    n565
  );


  buf
  g733
  (
    n823,
    n535
  );


  not
  g734
  (
    n777,
    n504
  );


  buf
  g735
  (
    n832,
    n498
  );


  not
  g736
  (
    n762,
    n592
  );


  not
  g737
  (
    n738,
    n526
  );


  not
  g738
  (
    n816,
    n590
  );


  buf
  g739
  (
    n735,
    n501
  );


  not
  g740
  (
    n764,
    n570
  );


  buf
  g741
  (
    n812,
    n518
  );


  not
  g742
  (
    n831,
    n505
  );


  buf
  g743
  (
    n819,
    n548
  );


  not
  g744
  (
    n802,
    n573
  );


  not
  g745
  (
    n769,
    n517
  );


  buf
  g746
  (
    n757,
    n577
  );


  buf
  g747
  (
    n781,
    n502
  );


  buf
  g748
  (
    n789,
    n595
  );


  not
  g749
  (
    KeyWire_0_32,
    n513
  );


  buf
  g750
  (
    KeyWire_0_23,
    n585
  );


  not
  g751
  (
    n784,
    n593
  );


  not
  g752
  (
    n801,
    n534
  );


  buf
  g753
  (
    n742,
    n515
  );


  not
  g754
  (
    n753,
    n576
  );


  buf
  g755
  (
    n811,
    n544
  );


  not
  g756
  (
    n813,
    n499
  );


  buf
  g757
  (
    n760,
    n568
  );


  buf
  g758
  (
    n736,
    n579
  );


  not
  g759
  (
    n798,
    n503
  );


  buf
  g760
  (
    n748,
    n527
  );


  not
  g761
  (
    n763,
    n566
  );


  not
  g762
  (
    n797,
    n580
  );


  buf
  g763
  (
    n790,
    n596
  );


  buf
  g764
  (
    n785,
    n499
  );


  buf
  g765
  (
    n756,
    n514
  );


  buf
  g766
  (
    n804,
    n547
  );


  not
  g767
  (
    n744,
    n587
  );


  buf
  g768
  (
    n824,
    n564
  );


  not
  g769
  (
    n761,
    n589
  );


  not
  g770
  (
    n800,
    n582
  );


  buf
  g771
  (
    n767,
    n530
  );


  not
  g772
  (
    n814,
    n539
  );


  buf
  g773
  (
    n745,
    n508
  );


  buf
  g774
  (
    n788,
    n522
  );


  buf
  g775
  (
    n783,
    n581
  );


  buf
  g776
  (
    n747,
    n546
  );


  buf
  g777
  (
    n752,
    n574
  );


  buf
  g778
  (
    n809,
    n503
  );


  not
  g779
  (
    n770,
    n498
  );


  buf
  g780
  (
    n829,
    n567
  );


  not
  g781
  (
    n740,
    n538
  );


  not
  g782
  (
    n772,
    n525
  );


  buf
  g783
  (
    n803,
    n584
  );


  not
  g784
  (
    n775,
    n560
  );


  not
  g785
  (
    n741,
    n502
  );


  not
  g786
  (
    n774,
    n561
  );


  buf
  g787
  (
    n794,
    n558
  );


  buf
  g788
  (
    n766,
    n586
  );


  buf
  g789
  (
    n792,
    n501
  );


  buf
  g790
  (
    KeyWire_0_48,
    n533
  );


  buf
  g791
  (
    n758,
    n532
  );


  not
  g792
  (
    n830,
    n554
  );


  not
  g793
  (
    n820,
    n502
  );


  not
  g794
  (
    n755,
    n500
  );


  buf
  g795
  (
    n810,
    n562
  );


  not
  g796
  (
    KeyWire_0_51,
    n498
  );


  or
  g797
  (
    n746,
    n500,
    n578,
    n521
  );


  or
  g798
  (
    KeyWire_0_45,
    n563,
    n583,
    n555,
    n500
  );


  xnor
  g799
  (
    n793,
    n519,
    n593,
    n509,
    n550
  );


  xor
  g800
  (
    n825,
    n594,
    n543,
    n512,
    n553
  );


  and
  g801
  (
    n776,
    n504,
    n541,
    n536,
    n511
  );


  and
  g802
  (
    n782,
    n503,
    n591,
    n569,
    n598
  );


  xnor
  g803
  (
    n786,
    n503,
    n523,
    n510,
    n556
  );


  nor
  g804
  (
    n773,
    n542,
    n545,
    n504,
    n502
  );


  or
  g805
  (
    n743,
    n501,
    n505,
    n597,
    n520
  );


  nor
  g806
  (
    n754,
    n597,
    n524,
    n596,
    n575
  );


  nand
  g807
  (
    n917,
    n670,
    n750,
    n645,
    n636
  );


  xor
  g808
  (
    n924,
    n738,
    n749,
    n748,
    n622
  );


  xnor
  g809
  (
    n896,
    n723,
    n688,
    n749,
    n745
  );


  or
  g810
  (
    n911,
    n643,
    n666,
    n615,
    n617
  );


  or
  g811
  (
    KeyWire_0_55,
    n763,
    n720,
    n633,
    n739
  );


  xnor
  g812
  (
    n843,
    n702,
    n759,
    n721,
    n602
  );


  nor
  g813
  (
    n916,
    n764,
    n679,
    n760,
    n615
  );


  nand
  g814
  (
    n910,
    n724,
    n635,
    n757,
    n640
  );


  xor
  g815
  (
    n913,
    n681,
    n600,
    n749,
    n689
  );


  or
  g816
  (
    n837,
    n606,
    n728,
    n629,
    n744
  );


  nand
  g817
  (
    n912,
    n664,
    n761,
    n738,
    n640
  );


  and
  g818
  (
    n897,
    n763,
    n719,
    n721,
    n685
  );


  nand
  g819
  (
    n833,
    n700,
    n743,
    n628,
    n680
  );


  xor
  g820
  (
    n909,
    n724,
    n656,
    n736,
    n698
  );


  xor
  g821
  (
    n844,
    n730,
    n634,
    n609,
    n742
  );


  xnor
  g822
  (
    n902,
    n650,
    n601,
    n738,
    n696
  );


  nand
  g823
  (
    n870,
    n762,
    n692,
    n718,
    n607
  );


  nor
  g824
  (
    n847,
    n703,
    n632,
    n655,
    n636
  );


  and
  g825
  (
    n845,
    n725,
    n618,
    n736,
    n737
  );


  nand
  g826
  (
    n838,
    n673,
    n742,
    n726,
    n626
  );


  and
  g827
  (
    n893,
    n708,
    n753,
    n674,
    n702
  );


  xnor
  g828
  (
    KeyWire_0_27,
    n758,
    n759,
    n627
  );


  nor
  g829
  (
    n901,
    n633,
    n750,
    n661,
    n706
  );


  nand
  g830
  (
    n883,
    n599,
    n688,
    n691,
    n755
  );


  or
  g831
  (
    n920,
    n647,
    n735,
    n687
  );


  xor
  g832
  (
    n905,
    n629,
    n614,
    n605,
    n665
  );


  or
  g833
  (
    n895,
    n759,
    n729,
    n723,
    n620
  );


  nand
  g834
  (
    n861,
    n747,
    n642,
    n611,
    n645
  );


  xor
  g835
  (
    KeyWire_0_26,
    n761,
    n706,
    n621,
    n616
  );


  and
  g836
  (
    n855,
    n726,
    n660,
    n739,
    n654
  );


  nand
  g837
  (
    n878,
    n651,
    n612,
    n755,
    n655
  );


  xor
  g838
  (
    n852,
    n701,
    n756,
    n639,
    n745
  );


  xnor
  g839
  (
    n835,
    n701,
    n753,
    n731,
    n754
  );


  xor
  g840
  (
    n879,
    n697,
    n714,
    n665,
    n760
  );


  xnor
  g841
  (
    n851,
    n749,
    n680,
    n664,
    n715
  );


  nand
  g842
  (
    n840,
    n674,
    n627,
    n695,
    n738
  );


  xnor
  g843
  (
    n860,
    n631,
    n671,
    n694,
    n697
  );


  xor
  g844
  (
    n839,
    n764,
    n741,
    n744,
    n761
  );


  nor
  g845
  (
    n846,
    n754,
    n656,
    n689,
    n637
  );


  xnor
  g846
  (
    n863,
    n746,
    n678,
    n657,
    n745
  );


  nand
  g847
  (
    n919,
    n630,
    n755,
    n682,
    n727
  );


  nor
  g848
  (
    n857,
    n614,
    n616,
    n761,
    n728
  );


  or
  g849
  (
    n859,
    n740,
    n662,
    n753,
    n644
  );


  and
  g850
  (
    n891,
    n722,
    n694,
    n716,
    n705
  );


  or
  g851
  (
    n894,
    n757,
    n696,
    n754,
    n676
  );


  and
  g852
  (
    KeyWire_0_42,
    n751,
    n606,
    n741,
    n619
  );


  xnor
  g853
  (
    n899,
    n603,
    n639,
    n744,
    n600
  );


  xor
  g854
  (
    n908,
    n602,
    n676,
    n763,
    n681
  );


  nand
  g855
  (
    n903,
    n653,
    n647,
    n707,
    n730
  );


  and
  g856
  (
    n906,
    n618,
    n675,
    n648,
    n630
  );


  nand
  g857
  (
    n925,
    n763,
    n686,
    n658,
    n736
  );


  nor
  g858
  (
    n834,
    n652,
    n659,
    n621,
    n745
  );


  and
  g859
  (
    n888,
    n719,
    n695,
    n740,
    n748
  );


  or
  g860
  (
    n876,
    n667,
    n747,
    n660,
    n693
  );


  xnor
  g861
  (
    KeyWire_0_8,
    n683,
    n757,
    n740,
    n670
  );


  xnor
  g862
  (
    n868,
    n741,
    n712,
    n609,
    n748
  );


  nor
  g863
  (
    n858,
    n746,
    n698,
    n760,
    n617
  );


  nor
  g864
  (
    n866,
    n741,
    n703,
    n682,
    n746
  );


  xnor
  g865
  (
    n842,
    n743,
    n705,
    n758,
    n649
  );


  xnor
  g866
  (
    n871,
    n710,
    n672,
    n671,
    n699
  );


  or
  g867
  (
    n927,
    n641,
    n743,
    n657,
    n685
  );


  xnor
  g868
  (
    n836,
    n711,
    n666,
    n679,
    n648
  );


  nand
  g869
  (
    n850,
    n663,
    n731,
    n644,
    n740
  );


  nor
  g870
  (
    n886,
    n661,
    n762,
    n687,
    n641
  );


  xor
  g871
  (
    n882,
    n699,
    n623,
    n752,
    n709
  );


  nor
  g872
  (
    n875,
    n603,
    n713,
    n725
  );


  and
  g873
  (
    n849,
    n622,
    n737,
    n746
  );


  nor
  g874
  (
    n862,
    n604,
    n608,
    n612,
    n631
  );


  xnor
  g875
  (
    n887,
    n620,
    n608,
    n653,
    n700
  );


  nand
  g876
  (
    n856,
    n711,
    n709,
    n737,
    n632
  );


  xnor
  g877
  (
    n884,
    n605,
    n751,
    n756,
    n684
  );


  and
  g878
  (
    n922,
    n684,
    n710,
    n754,
    n743
  );


  xnor
  g879
  (
    n907,
    n756,
    n613,
    n690,
    n729
  );


  or
  g880
  (
    n853,
    n717,
    n717,
    n718,
    n625
  );


  and
  g881
  (
    KeyWire_0_15,
    n750,
    n762,
    n611,
    n650
  );


  or
  g882
  (
    n872,
    n607,
    n654,
    n704,
    n643
  );


  nor
  g883
  (
    n864,
    n668,
    n646,
    n663,
    n625
  );


  and
  g884
  (
    n877,
    n764,
    n755,
    n712,
    n690
  );


  xor
  g885
  (
    n918,
    n601,
    n667,
    n757,
    n628
  );


  xnor
  g886
  (
    n900,
    n659,
    n683,
    n744,
    n715
  );


  xnor
  g887
  (
    n885,
    n649,
    n613,
    n691,
    n707
  );


  xor
  g888
  (
    n921,
    n735,
    n598,
    n750,
    n638
  );


  and
  g889
  (
    n869,
    n747,
    n704,
    n752,
    n762
  );


  xor
  g890
  (
    KeyWire_0_5,
    n752,
    n669,
    n599,
    n624
  );


  xor
  g891
  (
    n915,
    n604,
    n642,
    n708,
    n739
  );


  nand
  g892
  (
    n873,
    n610,
    n662,
    n678,
    n732
  );


  xor
  g893
  (
    n928,
    n720,
    n722,
    n693,
    n727
  );


  nand
  g894
  (
    n865,
    n748,
    n742,
    n668,
    n672
  );


  and
  g895
  (
    KeyWire_0_50,
    n739,
    n716,
    n751,
    n610
  );


  or
  g896
  (
    n874,
    n638,
    n692,
    n677,
    n623
  );


  nor
  g897
  (
    n890,
    n658,
    n651,
    n624,
    n732
  );


  nor
  g898
  (
    n904,
    n619,
    n714,
    n626,
    n675
  );


  xnor
  g899
  (
    n923,
    n673,
    n669,
    n635,
    n634
  );


  nand
  g900
  (
    n889,
    n646,
    n747,
    n756,
    n686
  );


  xnor
  g901
  (
    n929,
    n764,
    n742,
    n677,
    n736
  );


  xnor
  g902
  (
    n926,
    n637,
    n752,
    n760,
    n751
  );


  xnor
  g903
  (
    n892,
    n753,
    n758,
    n652
  );


  and
  g904
  (
    n942,
    n889,
    n821,
    n767,
    n909
  );


  nor
  g905
  (
    n951,
    n789,
    n814,
    n850,
    n842
  );


  xnor
  g906
  (
    n969,
    n810,
    n852,
    n801,
    n796
  );


  and
  g907
  (
    n977,
    n854,
    n824,
    n774,
    n771
  );


  or
  g908
  (
    n979,
    n864,
    n776,
    n799,
    n788
  );


  nand
  g909
  (
    n947,
    n813,
    n779,
    n882,
    n799
  );


  nor
  g910
  (
    n952,
    n821,
    n796,
    n786
  );


  nand
  g911
  (
    n1007,
    n782,
    n819,
    n816,
    n779
  );


  or
  g912
  (
    n959,
    n841,
    n823,
    n822,
    n781
  );


  xor
  g913
  (
    n970,
    n800,
    n765,
    n792,
    n868
  );


  xnor
  g914
  (
    n944,
    n791,
    n767,
    n788,
    n806
  );


  xnor
  g915
  (
    n997,
    n819,
    n766,
    n775,
    n804
  );


  nand
  g916
  (
    n992,
    n811,
    n782,
    n824,
    n818
  );


  xnor
  g917
  (
    n990,
    n861,
    n813,
    n810,
    n798
  );


  or
  g918
  (
    n975,
    n801,
    n800,
    n870,
    n846
  );


  xnor
  g919
  (
    n1001,
    n784,
    n782,
    n773,
    n875
  );


  and
  g920
  (
    n957,
    n802,
    n803,
    n888,
    n778
  );


  xnor
  g921
  (
    n966,
    n859,
    n781,
    n787,
    n885
  );


  xor
  g922
  (
    n986,
    n783,
    n791,
    n810,
    n865
  );


  nand
  g923
  (
    n981,
    n777,
    n770,
    n791,
    n805
  );


  xnor
  g924
  (
    n1004,
    n780,
    n847,
    n787,
    n803
  );


  and
  g925
  (
    n943,
    n775,
    n797,
    n902,
    n802
  );


  xnor
  g926
  (
    n996,
    n768,
    n824,
    n860,
    n783
  );


  xor
  g927
  (
    n955,
    n814,
    n891,
    n895,
    n881
  );


  nand
  g928
  (
    KeyWire_0_36,
    n856,
    n883,
    n790,
    n795
  );


  nor
  g929
  (
    n982,
    n818,
    n777,
    n820,
    n772
  );


  nand
  g930
  (
    n998,
    n822,
    n774,
    n773,
    n770
  );


  nand
  g931
  (
    n991,
    n869,
    n866,
    n809
  );


  nor
  g932
  (
    n993,
    n848,
    n793,
    n805,
    n804
  );


  or
  g933
  (
    n989,
    n800,
    n804,
    n778,
    n862
  );


  and
  g934
  (
    n958,
    n785,
    n803,
    n793,
    n774
  );


  or
  g935
  (
    n987,
    n787,
    n901,
    n867,
    n853
  );


  xor
  g936
  (
    n931,
    n820,
    n813,
    n872,
    n810
  );


  nand
  g937
  (
    n937,
    n817,
    n785,
    n780,
    n767
  );


  xnor
  g938
  (
    n936,
    n766,
    n804,
    n822,
    n788
  );


  and
  g939
  (
    n988,
    n816,
    n912,
    n814,
    n824
  );


  or
  g940
  (
    n948,
    n771,
    n792,
    n806,
    n887
  );


  nor
  g941
  (
    n963,
    n821,
    n779,
    n802,
    n904
  );


  nand
  g942
  (
    n980,
    n820,
    n812,
    n798,
    n838
  );


  xnor
  g943
  (
    n935,
    n815,
    n817,
    n789,
    n790
  );


  or
  g944
  (
    n953,
    n808,
    n781,
    n836,
    n855
  );


  or
  g945
  (
    n964,
    n843,
    n823,
    n898,
    n809
  );


  nand
  g946
  (
    n961,
    n799,
    n805,
    n798,
    n780
  );


  and
  g947
  (
    n940,
    n833,
    n821,
    n905,
    n894
  );


  and
  g948
  (
    n995,
    n793,
    n899,
    n771,
    n787
  );


  xor
  g949
  (
    n1002,
    n811,
    n858,
    n806,
    n782
  );


  nand
  g950
  (
    n983,
    n911,
    n822,
    n815,
    n784
  );


  nor
  g951
  (
    n939,
    n769,
    n813,
    n789,
    n771
  );


  and
  g952
  (
    n965,
    n817,
    n785,
    n812,
    n801
  );


  and
  g953
  (
    n1006,
    n908,
    n816,
    n835,
    n766
  );


  nor
  g954
  (
    n968,
    n793,
    n820,
    n768,
    n797
  );


  or
  g955
  (
    n973,
    n880,
    n783,
    n792,
    n808
  );


  xnor
  g956
  (
    n967,
    n834,
    n781,
    n910,
    n795
  );


  or
  g957
  (
    n960,
    n849,
    n785,
    n819,
    n788
  );


  or
  g958
  (
    n1003,
    n778,
    n844,
    n790,
    n772
  );


  or
  g959
  (
    n1000,
    n773,
    n797,
    n811,
    n784
  );


  or
  g960
  (
    n984,
    n768,
    n773,
    n794,
    n863
  );


  or
  g961
  (
    n938,
    n840,
    n775,
    n777,
    n776
  );


  xor
  g962
  (
    n978,
    n839,
    n805,
    n769,
    n900
  );


  xnor
  g963
  (
    n1009,
    n807,
    n818,
    n786,
    n851
  );


  nor
  g964
  (
    KeyWire_0_38,
    n775,
    n774,
    n806,
    n765
  );


  xnor
  g965
  (
    n945,
    n765,
    n769,
    n823,
    n837
  );


  xnor
  g966
  (
    n972,
    n799,
    n818,
    n795,
    n800
  );


  or
  g967
  (
    n933,
    n802,
    n797,
    n770,
    n816
  );


  nor
  g968
  (
    n930,
    n789,
    n906,
    n798,
    n876
  );


  or
  g969
  (
    n932,
    n809,
    n807,
    n768,
    n803
  );


  and
  g970
  (
    n950,
    n808,
    n791,
    n886,
    n874
  );


  xnor
  g971
  (
    n971,
    n873,
    n878,
    n770,
    n794
  );


  or
  g972
  (
    n956,
    n893,
    n786,
    n780,
    n815
  );


  xor
  g973
  (
    n946,
    n794,
    n884,
    n786,
    n814
  );


  and
  g974
  (
    n934,
    n896,
    n857,
    n815,
    n776
  );


  xor
  g975
  (
    n941,
    n792,
    n871,
    n877,
    n879
  );


  nand
  g976
  (
    n949,
    n783,
    n823,
    n772,
    n765
  );


  or
  g977
  (
    n1005,
    n779,
    n777,
    n812,
    n808
  );


  xnor
  g978
  (
    n974,
    n769,
    n903,
    n794,
    n845
  );


  xnor
  g979
  (
    n1008,
    n776,
    n892,
    n778,
    n772
  );


  xnor
  g980
  (
    n954,
    n796,
    n817,
    n784,
    n907
  );


  and
  g981
  (
    n985,
    n766,
    n811,
    n807,
    n790
  );


  xor
  g982
  (
    n976,
    n795,
    n890,
    n767,
    n897
  );


  xnor
  g983
  (
    n994,
    n801,
    n812,
    n807,
    n819
  );


  buf
  g984
  (
    KeyWire_0_4,
    n927
  );


  buf
  g985
  (
    n1028,
    n505
  );


  not
  g986
  (
    n1041,
    n982
  );


  buf
  g987
  (
    KeyWire_0_6,
    n984
  );


  not
  g988
  (
    n1045,
    n979
  );


  not
  g989
  (
    n1062,
    n942
  );


  not
  g990
  (
    KeyWire_0_21,
    n926
  );


  buf
  g991
  (
    n1026,
    n925
  );


  buf
  g992
  (
    n1051,
    n507
  );


  not
  g993
  (
    n1070,
    n507
  );


  not
  g994
  (
    n1039,
    n976
  );


  buf
  g995
  (
    n1012,
    n960
  );


  buf
  g996
  (
    n1064,
    n939
  );


  buf
  g997
  (
    n1054,
    n995
  );


  buf
  g998
  (
    n1018,
    n938
  );


  buf
  g999
  (
    n1015,
    n438
  );


  buf
  g1000
  (
    n1052,
    n940
  );


  not
  g1001
  (
    n1067,
    n972
  );


  not
  g1002
  (
    n1013,
    n950
  );


  buf
  g1003
  (
    n1027,
    n956
  );


  buf
  g1004
  (
    n1044,
    n439
  );


  buf
  g1005
  (
    n1072,
    n967
  );


  buf
  g1006
  (
    n1063,
    n929
  );


  buf
  g1007
  (
    n1048,
    n506
  );


  buf
  g1008
  (
    n1010,
    n981
  );


  not
  g1009
  (
    n1043,
    n964
  );


  buf
  g1010
  (
    n1038,
    n918
  );


  not
  g1011
  (
    n1053,
    n954
  );


  not
  g1012
  (
    n1031,
    n936
  );


  buf
  g1013
  (
    n1040,
    n955
  );


  buf
  g1014
  (
    n1058,
    n945
  );


  not
  g1015
  (
    n1023,
    n439
  );


  buf
  g1016
  (
    n1060,
    n916
  );


  not
  g1017
  (
    n1017,
    n952
  );


  not
  g1018
  (
    n1022,
    n963
  );


  not
  g1019
  (
    n1065,
    n506
  );


  buf
  g1020
  (
    n1021,
    n915
  );


  not
  g1021
  (
    n1011,
    n948
  );


  not
  g1022
  (
    KeyWire_0_29,
    n947
  );


  not
  g1023
  (
    n1049,
    n924
  );


  not
  g1024
  (
    n1025,
    n914
  );


  buf
  g1025
  (
    n1024,
    n951
  );


  not
  g1026
  (
    n1035,
    n994
  );


  buf
  g1027
  (
    n1032,
    n966
  );


  not
  g1028
  (
    n1014,
    n988
  );


  buf
  g1029
  (
    n1036,
    n1000
  );


  not
  g1030
  (
    n1046,
    n438
  );


  buf
  g1031
  (
    n1029,
    n941
  );


  buf
  g1032
  (
    n1019,
    n996
  );


  not
  g1033
  (
    n1047,
    n999
  );


  buf
  g1034
  (
    n1016,
    n25
  );


  nand
  g1035
  (
    n1020,
    n923,
    n978,
    n957,
    n971
  );


  or
  g1036
  (
    n1042,
    n969,
    n438,
    n993,
    n997
  );


  nor
  g1037
  (
    n1050,
    n937,
    n507,
    n989,
    n974
  );


  xnor
  g1038
  (
    n1071,
    n507,
    n983,
    n973,
    n968
  );


  nor
  g1039
  (
    n1069,
    n986,
    n985,
    n943,
    n917
  );


  and
  g1040
  (
    n1061,
    n919,
    n953,
    n987,
    n991
  );


  nand
  g1041
  (
    n1034,
    n980,
    n958,
    n992,
    n949
  );


  and
  g1042
  (
    n1066,
    n913,
    n439,
    n921,
    n505
  );


  xor
  g1043
  (
    n1059,
    n920,
    n998,
    n962,
    n506
  );


  xor
  g1044
  (
    n1057,
    n506,
    n990,
    n961,
    n922
  );


  nand
  g1045
  (
    n1055,
    n970,
    n928,
    n965,
    n977
  );


  or
  g1046
  (
    n1033,
    n959,
    n944,
    n946,
    n975
  );


  xor
  g1047
  (
    n1073,
    n1006,
    n1036,
    n1024,
    n1010
  );


  xnor
  g1048
  (
    n1084,
    n1064,
    n1054,
    n1065,
    n1025
  );


  or
  g1049
  (
    n1082,
    n1026,
    n1044,
    n1012,
    n1049
  );


  xnor
  g1050
  (
    n1087,
    n1003,
    n1027,
    n1066,
    n1054
  );


  and
  g1051
  (
    n1096,
    n1009,
    n1038,
    n1013,
    n1050
  );


  xor
  g1052
  (
    n1091,
    n1052,
    n1063,
    n1045,
    n1005
  );


  nand
  g1053
  (
    n1095,
    n1042,
    n1049,
    n1001,
    n1063
  );


  nor
  g1054
  (
    n1076,
    n1018,
    n1016,
    n1017,
    n1057
  );


  xor
  g1055
  (
    n1086,
    n1043,
    n1037,
    n1015,
    n1055
  );


  nand
  g1056
  (
    n1085,
    n1060,
    n1045,
    n1056,
    n1062
  );


  and
  g1057
  (
    n1094,
    n1014,
    n1035,
    n1068,
    n1031
  );


  xnor
  g1058
  (
    n1074,
    n1040,
    n1062,
    n1051,
    n1052
  );


  and
  g1059
  (
    n1081,
    n1048,
    n1060,
    n1047,
    n1033
  );


  xnor
  g1060
  (
    n1080,
    n1029,
    n1055,
    n1043,
    n1020
  );


  or
  g1061
  (
    n1092,
    n1050,
    n1041,
    n1040,
    n1032
  );


  nor
  g1062
  (
    n1090,
    n1066,
    n1053,
    n1002,
    n1059
  );


  or
  g1063
  (
    n1093,
    n1021,
    n1004,
    n1048,
    n1065
  );


  or
  g1064
  (
    n1089,
    n1057,
    n1067,
    n1059,
    n1064
  );


  or
  g1065
  (
    n1075,
    n1007,
    n1061,
    n1034,
    n1030
  );


  nor
  g1066
  (
    n1077,
    n1039,
    n1053,
    n1019,
    n1042
  );


  or
  g1067
  (
    n1088,
    n1056,
    n1046,
    n1058,
    n1023
  );


  xor
  g1068
  (
    n1078,
    n1008,
    n1046,
    n1028,
    n1047
  );


  xnor
  g1069
  (
    n1079,
    n1058,
    n1051,
    n1061,
    n1011
  );


  or
  g1070
  (
    n1083,
    n1044,
    n1067,
    n1041,
    n1022
  );


  xnor
  g1071
  (
    n1099,
    n1088,
    n1083,
    n1072,
    n1068
  );


  xor
  g1072
  (
    n1098,
    n1070,
    n1069,
    n1084,
    n1071
  );


  xnor
  g1073
  (
    n1100,
    n1081,
    n1082,
    n1070,
    n1085
  );


  and
  g1074
  (
    KeyWire_0_56,
    n1069,
    n1087,
    n1071,
    n1086
  );


  nand
  g1075
  (
    n1102,
    n1092,
    n1099,
    n1089,
    n1093
  );


  nand
  g1076
  (
    n1101,
    n1091,
    n1100,
    n1094,
    n1090
  );


  xnor
  g1077
  (
    n1103,
    n826,
    n1101,
    n1102
  );


  xnor
  g1078
  (
    n1105,
    n827,
    n826,
    n1102,
    n825
  );


  or
  g1079
  (
    n1104,
    n734,
    n733,
    n825,
    n1096
  );


  xor
  g1080
  (
    n1107,
    n827,
    n1072,
    n1102,
    n1095
  );


  or
  g1081
  (
    KeyWire_0_28,
    n826,
    n734,
    n827,
    n825
  );


  or
  g1082
  (
    n1106,
    n1101,
    n826,
    n733,
    n825
  );


  xnor
  g1083
  (
    n1114,
    n829,
    n828,
    n832,
    n827
  );


  xnor
  g1084
  (
    n1111,
    n1108,
    n828,
    n831,
    n830
  );


  nand
  g1085
  (
    n1112,
    n830,
    n1104,
    n829,
    n1106
  );


  nor
  g1086
  (
    KeyWire_0_52,
    n830,
    n1103,
    n828,
    n831
  );


  or
  g1087
  (
    n1115,
    n832,
    n1107,
    n830,
    n831
  );


  xnor
  g1088
  (
    n1113,
    n831,
    n1108,
    n829,
    n828
  );


  xor
  g1089
  (
    n1110,
    n832,
    n832,
    n1105,
    n829
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n99,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n558,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n700,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n137,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1030,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n848,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n1068,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n593,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n914,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n337,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n279,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n195,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n341,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n289,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n85,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n841,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n463,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n311,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n604,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n148,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n519,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1056,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n56,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n737,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n145,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n640,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n854,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n867,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1108,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1037,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n236,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n250,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n827,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n347,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n778,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n400,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n962,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n536,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n999,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n465,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n47,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n266,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n880,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n149,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n430,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n749,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n557,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n622,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n795,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n274,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n898,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n787,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n1109,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n316,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n439,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n881,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n1097,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n282,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n294,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n175,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n469,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n129,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n644,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n58,
    KeyNOTWire_0_63
  );


endmodule


