

module Stat_3000_431
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1816,
  n1831,
  n1858,
  n1875,
  n1876,
  n1873,
  n1871,
  n1877,
  n1872,
  n1870,
  n3018,
  n3013,
  n3028,
  n3022,
  n3020,
  n3012,
  n3015,
  n3019,
  n3021,
  n3016,
  n3011,
  n3023,
  n3026,
  n3024,
  n3025,
  n3030,
  n3027,
  n3029,
  n3031,
  n3032,
  n3017,
  n3014
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1816;output n1831;output n1858;output n1875;output n1876;output n1873;output n1871;output n1877;output n1872;output n1870;output n3018;output n3013;output n3028;output n3022;output n3020;output n3012;output n3015;output n3019;output n3021;output n3016;output n3011;output n3023;output n3026;output n3024;output n3025;output n3030;output n3027;output n3029;output n3031;output n3032;output n3017;output n3014;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1874;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;

  buf
  g0
  (
    n74,
    n14
  );


  buf
  g1
  (
    n109,
    n6
  );


  not
  g2
  (
    n134,
    n21
  );


  not
  g3
  (
    n41,
    n18
  );


  not
  g4
  (
    n39,
    n28
  );


  buf
  g5
  (
    n95,
    n31
  );


  not
  g6
  (
    n55,
    n17
  );


  not
  g7
  (
    n113,
    n13
  );


  not
  g8
  (
    n105,
    n31
  );


  buf
  g9
  (
    n121,
    n32
  );


  buf
  g10
  (
    n129,
    n15
  );


  not
  g11
  (
    n85,
    n4
  );


  buf
  g12
  (
    n125,
    n10
  );


  not
  g13
  (
    n112,
    n26
  );


  not
  g14
  (
    n103,
    n2
  );


  buf
  g15
  (
    n159,
    n13
  );


  buf
  g16
  (
    n50,
    n24
  );


  buf
  g17
  (
    n80,
    n16
  );


  not
  g18
  (
    n92,
    n7
  );


  not
  g19
  (
    n140,
    n8
  );


  not
  g20
  (
    n139,
    n18
  );


  not
  g21
  (
    n114,
    n21
  );


  not
  g22
  (
    n37,
    n30
  );


  buf
  g23
  (
    n34,
    n9
  );


  not
  g24
  (
    n47,
    n8
  );


  buf
  g25
  (
    n43,
    n21
  );


  not
  g26
  (
    n108,
    n31
  );


  buf
  g27
  (
    n77,
    n10
  );


  not
  g28
  (
    n144,
    n20
  );


  not
  g29
  (
    n59,
    n4
  );


  not
  g30
  (
    n54,
    n3
  );


  buf
  g31
  (
    n82,
    n22
  );


  buf
  g32
  (
    n87,
    n15
  );


  buf
  g33
  (
    n84,
    n10
  );


  not
  g34
  (
    n143,
    n12
  );


  not
  g35
  (
    n83,
    n9
  );


  buf
  g36
  (
    n68,
    n16
  );


  not
  g37
  (
    n124,
    n14
  );


  not
  g38
  (
    n40,
    n2
  );


  not
  g39
  (
    n130,
    n22
  );


  buf
  g40
  (
    KeyWire_0_24,
    n30
  );


  buf
  g41
  (
    n67,
    n1
  );


  not
  g42
  (
    n71,
    n27
  );


  not
  g43
  (
    n93,
    n13
  );


  not
  g44
  (
    n151,
    n14
  );


  buf
  g45
  (
    n127,
    n20
  );


  buf
  g46
  (
    n51,
    n7
  );


  buf
  g47
  (
    n153,
    n16
  );


  buf
  g48
  (
    n49,
    n25
  );


  buf
  g49
  (
    n88,
    n22
  );


  not
  g50
  (
    n102,
    n29
  );


  buf
  g51
  (
    n138,
    n20
  );


  buf
  g52
  (
    n106,
    n2
  );


  not
  g53
  (
    n133,
    n21
  );


  buf
  g54
  (
    n44,
    n30
  );


  buf
  g55
  (
    n91,
    n18
  );


  not
  g56
  (
    n148,
    n23
  );


  not
  g57
  (
    n119,
    n23
  );


  buf
  g58
  (
    n137,
    n32
  );


  buf
  g59
  (
    n117,
    n27
  );


  not
  g60
  (
    n66,
    n1
  );


  buf
  g61
  (
    n128,
    n14
  );


  buf
  g62
  (
    n57,
    n29
  );


  buf
  g63
  (
    n58,
    n12
  );


  not
  g64
  (
    n156,
    n3
  );


  buf
  g65
  (
    n135,
    n31
  );


  buf
  g66
  (
    n104,
    n15
  );


  buf
  g67
  (
    n81,
    n4
  );


  buf
  g68
  (
    n147,
    n19
  );


  not
  g69
  (
    n86,
    n25
  );


  not
  g70
  (
    n100,
    n9
  );


  not
  g71
  (
    n155,
    n24
  );


  buf
  g72
  (
    n110,
    n30
  );


  not
  g73
  (
    n158,
    n28
  );


  buf
  g74
  (
    n116,
    n22
  );


  not
  g75
  (
    n126,
    n19
  );


  buf
  g76
  (
    n99,
    n7
  );


  buf
  g77
  (
    n78,
    n18
  );


  not
  g78
  (
    n52,
    n13
  );


  not
  g79
  (
    n38,
    n32
  );


  buf
  g80
  (
    n136,
    n29
  );


  buf
  g81
  (
    n96,
    n1
  );


  not
  g82
  (
    n157,
    n27
  );


  not
  g83
  (
    n48,
    n10
  );


  not
  g84
  (
    n98,
    n6
  );


  buf
  g85
  (
    n70,
    n5
  );


  buf
  g86
  (
    n101,
    n3
  );


  buf
  g87
  (
    n33,
    n6
  );


  not
  g88
  (
    n42,
    n19
  );


  not
  g89
  (
    n149,
    n8
  );


  buf
  g90
  (
    n36,
    n27
  );


  buf
  g91
  (
    n90,
    n15
  );


  not
  g92
  (
    n61,
    n23
  );


  not
  g93
  (
    n56,
    n17
  );


  not
  g94
  (
    n160,
    n26
  );


  not
  g95
  (
    n46,
    n26
  );


  not
  g96
  (
    n141,
    n7
  );


  not
  g97
  (
    n152,
    n3
  );


  not
  g98
  (
    n60,
    n29
  );


  buf
  g99
  (
    n97,
    n5
  );


  buf
  g100
  (
    n65,
    n24
  );


  buf
  g101
  (
    n154,
    n20
  );


  buf
  g102
  (
    n94,
    n11
  );


  not
  g103
  (
    n123,
    n16
  );


  buf
  g104
  (
    n69,
    n25
  );


  not
  g105
  (
    n122,
    n17
  );


  not
  g106
  (
    n111,
    n12
  );


  buf
  g107
  (
    n150,
    n11
  );


  not
  g108
  (
    n63,
    n17
  );


  not
  g109
  (
    n89,
    n9
  );


  buf
  g110
  (
    n107,
    n12
  );


  not
  g111
  (
    n62,
    n11
  );


  buf
  g112
  (
    n45,
    n25
  );


  not
  g113
  (
    n72,
    n5
  );


  buf
  g114
  (
    n35,
    n24
  );


  buf
  g115
  (
    n73,
    n23
  );


  not
  g116
  (
    n115,
    n28
  );


  not
  g117
  (
    n131,
    n28
  );


  buf
  g118
  (
    n118,
    n6
  );


  not
  g119
  (
    n53,
    n2
  );


  not
  g120
  (
    n79,
    n26
  );


  buf
  g121
  (
    n120,
    n4
  );


  buf
  g122
  (
    n146,
    n11
  );


  buf
  g123
  (
    n75,
    n19
  );


  buf
  g124
  (
    n145,
    n5
  );


  buf
  g125
  (
    n76,
    n1
  );


  buf
  g126
  (
    n132,
    n32
  );


  buf
  g127
  (
    n142,
    n8
  );


  buf
  g128
  (
    n241,
    n76
  );


  buf
  g129
  (
    n635,
    n119
  );


  not
  g130
  (
    n397,
    n142
  );


  buf
  g131
  (
    KeyWire_0_11,
    n156
  );


  not
  g132
  (
    n345,
    n155
  );


  not
  g133
  (
    n504,
    n39
  );


  not
  g134
  (
    n205,
    n68
  );


  not
  g135
  (
    n204,
    n145
  );


  buf
  g136
  (
    n442,
    n73
  );


  not
  g137
  (
    n415,
    n157
  );


  not
  g138
  (
    n477,
    n100
  );


  buf
  g139
  (
    n422,
    n87
  );


  not
  g140
  (
    n474,
    n85
  );


  not
  g141
  (
    n171,
    n109
  );


  buf
  g142
  (
    n470,
    n152
  );


  buf
  g143
  (
    n520,
    n66
  );


  not
  g144
  (
    n627,
    n50
  );


  not
  g145
  (
    n375,
    n91
  );


  not
  g146
  (
    n272,
    n105
  );


  buf
  g147
  (
    n495,
    n39
  );


  buf
  g148
  (
    n651,
    n115
  );


  not
  g149
  (
    n349,
    n130
  );


  not
  g150
  (
    n215,
    n100
  );


  not
  g151
  (
    n178,
    n53
  );


  not
  g152
  (
    n254,
    n89
  );


  not
  g153
  (
    n589,
    n35
  );


  buf
  g154
  (
    n578,
    n158
  );


  not
  g155
  (
    n328,
    n46
  );


  buf
  g156
  (
    n311,
    n102
  );


  not
  g157
  (
    n505,
    n92
  );


  buf
  g158
  (
    n445,
    n58
  );


  not
  g159
  (
    n316,
    n113
  );


  buf
  g160
  (
    n219,
    n33
  );


  buf
  g161
  (
    n224,
    n107
  );


  not
  g162
  (
    n248,
    n65
  );


  buf
  g163
  (
    n469,
    n154
  );


  not
  g164
  (
    n304,
    n131
  );


  not
  g165
  (
    n420,
    n158
  );


  buf
  g166
  (
    n308,
    n112
  );


  not
  g167
  (
    n541,
    n152
  );


  buf
  g168
  (
    n533,
    n109
  );


  not
  g169
  (
    n337,
    n142
  );


  buf
  g170
  (
    n534,
    n47
  );


  buf
  g171
  (
    n388,
    n49
  );


  not
  g172
  (
    n623,
    n51
  );


  not
  g173
  (
    n535,
    n160
  );


  buf
  g174
  (
    n581,
    n141
  );


  buf
  g175
  (
    n602,
    n129
  );


  not
  g176
  (
    n334,
    n133
  );


  not
  g177
  (
    n658,
    n53
  );


  buf
  g178
  (
    n645,
    n53
  );


  not
  g179
  (
    n382,
    n69
  );


  buf
  g180
  (
    n634,
    n157
  );


  buf
  g181
  (
    n212,
    n59
  );


  buf
  g182
  (
    n582,
    n112
  );


  buf
  g183
  (
    n661,
    n86
  );


  buf
  g184
  (
    n267,
    n127
  );


  not
  g185
  (
    n360,
    n61
  );


  buf
  g186
  (
    n188,
    n113
  );


  buf
  g187
  (
    n406,
    n132
  );


  buf
  g188
  (
    n419,
    n42
  );


  buf
  g189
  (
    n438,
    n136
  );


  buf
  g190
  (
    n357,
    n62
  );


  buf
  g191
  (
    n618,
    n74
  );


  buf
  g192
  (
    n487,
    n55
  );


  not
  g193
  (
    n412,
    n46
  );


  not
  g194
  (
    n288,
    n45
  );


  not
  g195
  (
    n408,
    n102
  );


  not
  g196
  (
    n301,
    n54
  );


  not
  g197
  (
    n358,
    n58
  );


  not
  g198
  (
    n302,
    n60
  );


  buf
  g199
  (
    n362,
    n139
  );


  buf
  g200
  (
    n164,
    n43
  );


  buf
  g201
  (
    n237,
    n128
  );


  buf
  g202
  (
    n417,
    n111
  );


  buf
  g203
  (
    n299,
    n77
  );


  buf
  g204
  (
    KeyWire_0_57,
    n104
  );


  not
  g205
  (
    n173,
    n125
  );


  not
  g206
  (
    n401,
    n122
  );


  not
  g207
  (
    n343,
    n95
  );


  buf
  g208
  (
    n481,
    n64
  );


  not
  g209
  (
    n614,
    n58
  );


  not
  g210
  (
    n161,
    n94
  );


  not
  g211
  (
    n172,
    n131
  );


  not
  g212
  (
    n560,
    n67
  );


  buf
  g213
  (
    n361,
    n67
  );


  not
  g214
  (
    n571,
    n143
  );


  buf
  g215
  (
    n210,
    n44
  );


  not
  g216
  (
    n223,
    n88
  );


  not
  g217
  (
    n539,
    n157
  );


  buf
  g218
  (
    n368,
    n115
  );


  not
  g219
  (
    n255,
    n141
  );


  not
  g220
  (
    n273,
    n78
  );


  not
  g221
  (
    n377,
    n127
  );


  not
  g222
  (
    n271,
    n58
  );


  buf
  g223
  (
    n181,
    n60
  );


  buf
  g224
  (
    n190,
    n134
  );


  buf
  g225
  (
    n573,
    n116
  );


  not
  g226
  (
    n276,
    n70
  );


  buf
  g227
  (
    n296,
    n140
  );


  buf
  g228
  (
    n467,
    n160
  );


  not
  g229
  (
    n314,
    n83
  );


  buf
  g230
  (
    n546,
    n158
  );


  buf
  g231
  (
    n440,
    n139
  );


  buf
  g232
  (
    n496,
    n77
  );


  buf
  g233
  (
    n234,
    n92
  );


  buf
  g234
  (
    n568,
    n144
  );


  buf
  g235
  (
    n251,
    n95
  );


  not
  g236
  (
    n616,
    n87
  );


  not
  g237
  (
    n473,
    n59
  );


  buf
  g238
  (
    n354,
    n149
  );


  not
  g239
  (
    n335,
    n90
  );


  not
  g240
  (
    n291,
    n110
  );


  buf
  g241
  (
    n203,
    n50
  );


  buf
  g242
  (
    n229,
    n146
  );


  not
  g243
  (
    n405,
    n121
  );


  buf
  g244
  (
    n425,
    n115
  );


  not
  g245
  (
    n642,
    n49
  );


  buf
  g246
  (
    n545,
    n39
  );


  buf
  g247
  (
    n213,
    n44
  );


  buf
  g248
  (
    n170,
    n55
  );


  not
  g249
  (
    n333,
    n114
  );


  not
  g250
  (
    n421,
    n79
  );


  not
  g251
  (
    n284,
    n36
  );


  not
  g252
  (
    n565,
    n118
  );


  buf
  g253
  (
    n310,
    n79
  );


  buf
  g254
  (
    n399,
    n129
  );


  not
  g255
  (
    n322,
    n132
  );


  not
  g256
  (
    n242,
    n98
  );


  buf
  g257
  (
    n208,
    n157
  );


  not
  g258
  (
    n305,
    n132
  );


  not
  g259
  (
    n669,
    n122
  );


  buf
  g260
  (
    n256,
    n114
  );


  buf
  g261
  (
    n436,
    n91
  );


  buf
  g262
  (
    n657,
    n94
  );


  not
  g263
  (
    n189,
    n85
  );


  buf
  g264
  (
    n264,
    n57
  );


  not
  g265
  (
    n591,
    n71
  );


  not
  g266
  (
    n655,
    n72
  );


  not
  g267
  (
    n523,
    n95
  );


  not
  g268
  (
    n636,
    n88
  );


  not
  g269
  (
    n516,
    n43
  );


  buf
  g270
  (
    n387,
    n92
  );


  buf
  g271
  (
    n430,
    n70
  );


  buf
  g272
  (
    n601,
    n155
  );


  buf
  g273
  (
    n640,
    n40
  );


  buf
  g274
  (
    n629,
    n112
  );


  not
  g275
  (
    n447,
    n146
  );


  buf
  g276
  (
    n403,
    n48
  );


  not
  g277
  (
    n502,
    n127
  );


  not
  g278
  (
    n659,
    n115
  );


  buf
  g279
  (
    n286,
    n44
  );


  buf
  g280
  (
    n289,
    n39
  );


  buf
  g281
  (
    n610,
    n40
  );


  not
  g282
  (
    n197,
    n83
  );


  not
  g283
  (
    n390,
    n107
  );


  not
  g284
  (
    n320,
    n89
  );


  not
  g285
  (
    n348,
    n110
  );


  buf
  g286
  (
    n385,
    n85
  );


  not
  g287
  (
    n341,
    n113
  );


  buf
  g288
  (
    n169,
    n105
  );


  not
  g289
  (
    n567,
    n72
  );


  not
  g290
  (
    KeyWire_0_60,
    n47
  );


  not
  g291
  (
    n638,
    n139
  );


  not
  g292
  (
    n444,
    n101
  );


  buf
  g293
  (
    n558,
    n99
  );


  buf
  g294
  (
    n186,
    n97
  );


  buf
  g295
  (
    n446,
    n101
  );


  not
  g296
  (
    n239,
    n73
  );


  buf
  g297
  (
    n262,
    n72
  );


  buf
  g298
  (
    n471,
    n136
  );


  buf
  g299
  (
    n632,
    n82
  );


  not
  g300
  (
    n435,
    n116
  );


  buf
  g301
  (
    n265,
    n52
  );


  buf
  g302
  (
    KeyWire_0_22,
    n52
  );


  buf
  g303
  (
    n392,
    n144
  );


  not
  g304
  (
    n586,
    n117
  );


  not
  g305
  (
    n370,
    n86
  );


  buf
  g306
  (
    n268,
    n75
  );


  buf
  g307
  (
    n187,
    n127
  );


  not
  g308
  (
    n500,
    n113
  );


  buf
  g309
  (
    n269,
    n35
  );


  not
  g310
  (
    n460,
    n38
  );


  buf
  g311
  (
    n247,
    n100
  );


  buf
  g312
  (
    n259,
    n103
  );


  buf
  g313
  (
    n592,
    n105
  );


  buf
  g314
  (
    n300,
    n57
  );


  buf
  g315
  (
    n526,
    n79
  );


  not
  g316
  (
    n410,
    n138
  );


  not
  g317
  (
    n315,
    n89
  );


  buf
  g318
  (
    n654,
    n62
  );


  buf
  g319
  (
    n437,
    n136
  );


  buf
  g320
  (
    n249,
    n148
  );


  buf
  g321
  (
    n631,
    n118
  );


  not
  g322
  (
    n620,
    n142
  );


  buf
  g323
  (
    n585,
    n151
  );


  buf
  g324
  (
    n510,
    n104
  );


  not
  g325
  (
    n466,
    n117
  );


  buf
  g326
  (
    n409,
    n53
  );


  buf
  g327
  (
    n297,
    n93
  );


  not
  g328
  (
    n441,
    n91
  );


  not
  g329
  (
    n434,
    n130
  );


  not
  g330
  (
    n365,
    n60
  );


  not
  g331
  (
    n536,
    n101
  );


  not
  g332
  (
    n230,
    n47
  );


  not
  g333
  (
    n407,
    n43
  );


  buf
  g334
  (
    n646,
    n120
  );


  not
  g335
  (
    n509,
    n150
  );


  not
  g336
  (
    n217,
    n80
  );


  not
  g337
  (
    n404,
    n76
  );


  not
  g338
  (
    n569,
    n78
  );


  buf
  g339
  (
    n518,
    n63
  );


  buf
  g340
  (
    n483,
    n51
  );


  buf
  g341
  (
    n462,
    n138
  );


  buf
  g342
  (
    n461,
    n110
  );


  buf
  g343
  (
    KeyWire_0_9,
    n153
  );


  buf
  g344
  (
    n598,
    n111
  );


  not
  g345
  (
    n615,
    n82
  );


  not
  g346
  (
    n400,
    n120
  );


  not
  g347
  (
    n416,
    n71
  );


  not
  g348
  (
    n605,
    n67
  );


  not
  g349
  (
    n459,
    n38
  );


  not
  g350
  (
    n611,
    n75
  );


  not
  g351
  (
    n670,
    n33
  );


  buf
  g352
  (
    n346,
    n73
  );


  not
  g353
  (
    n531,
    n126
  );


  not
  g354
  (
    n630,
    n70
  );


  buf
  g355
  (
    n374,
    n141
  );


  not
  g356
  (
    n662,
    n93
  );


  buf
  g357
  (
    n488,
    n106
  );


  buf
  g358
  (
    n290,
    n160
  );


  not
  g359
  (
    n594,
    n52
  );


  not
  g360
  (
    n456,
    n106
  );


  buf
  g361
  (
    n564,
    n104
  );


  buf
  g362
  (
    n261,
    n137
  );


  buf
  g363
  (
    n206,
    n64
  );


  not
  g364
  (
    n307,
    n97
  );


  not
  g365
  (
    n625,
    n49
  );


  not
  g366
  (
    n547,
    n129
  );


  buf
  g367
  (
    n321,
    n154
  );


  not
  g368
  (
    n306,
    n72
  );


  buf
  g369
  (
    n191,
    n137
  );


  buf
  g370
  (
    n572,
    n117
  );


  not
  g371
  (
    n537,
    n88
  );


  buf
  g372
  (
    n340,
    n96
  );


  buf
  g373
  (
    n274,
    n150
  );


  buf
  g374
  (
    n463,
    n65
  );


  not
  g375
  (
    n218,
    n57
  );


  not
  g376
  (
    n559,
    n128
  );


  not
  g377
  (
    n168,
    n62
  );


  not
  g378
  (
    n257,
    n122
  );


  not
  g379
  (
    n476,
    n38
  );


  buf
  g380
  (
    n398,
    n132
  );


  not
  g381
  (
    n448,
    n69
  );


  buf
  g382
  (
    n336,
    n148
  );


  not
  g383
  (
    n599,
    n149
  );


  buf
  g384
  (
    n433,
    n91
  );


  not
  g385
  (
    n165,
    n52
  );


  buf
  g386
  (
    n351,
    n75
  );


  buf
  g387
  (
    n402,
    n90
  );


  not
  g388
  (
    n543,
    n121
  );


  buf
  g389
  (
    n293,
    n45
  );


  not
  g390
  (
    n540,
    n118
  );


  not
  g391
  (
    n450,
    n66
  );


  buf
  g392
  (
    n175,
    n81
  );


  buf
  g393
  (
    n182,
    n92
  );


  buf
  g394
  (
    n176,
    n145
  );


  not
  g395
  (
    n622,
    n99
  );


  not
  g396
  (
    n281,
    n46
  );


  buf
  g397
  (
    n295,
    n154
  );


  not
  g398
  (
    n637,
    n94
  );


  not
  g399
  (
    n619,
    n74
  );


  buf
  g400
  (
    n647,
    n149
  );


  buf
  g401
  (
    n489,
    n40
  );


  buf
  g402
  (
    n371,
    n133
  );


  not
  g403
  (
    n226,
    n158
  );


  not
  g404
  (
    n431,
    n80
  );


  not
  g405
  (
    n294,
    n135
  );


  not
  g406
  (
    n485,
    n148
  );


  buf
  g407
  (
    n277,
    n64
  );


  not
  g408
  (
    n644,
    n61
  );


  not
  g409
  (
    n613,
    n41
  );


  buf
  g410
  (
    n452,
    n67
  );


  not
  g411
  (
    n235,
    n107
  );


  buf
  g412
  (
    n575,
    n120
  );


  not
  g413
  (
    n606,
    n150
  );


  not
  g414
  (
    n593,
    n81
  );


  not
  g415
  (
    n517,
    n68
  );


  buf
  g416
  (
    n220,
    n159
  );


  buf
  g417
  (
    n350,
    n160
  );


  buf
  g418
  (
    n270,
    n56
  );


  not
  g419
  (
    n379,
    n84
  );


  buf
  g420
  (
    n184,
    n108
  );


  not
  g421
  (
    n183,
    n51
  );


  not
  g422
  (
    n660,
    n142
  );


  not
  g423
  (
    n648,
    n123
  );


  buf
  g424
  (
    n292,
    n153
  );


  buf
  g425
  (
    n426,
    n135
  );


  not
  g426
  (
    n458,
    n48
  );


  not
  g427
  (
    n475,
    n74
  );


  not
  g428
  (
    n185,
    n108
  );


  not
  g429
  (
    n424,
    n45
  );


  buf
  g430
  (
    n484,
    n124
  );


  buf
  g431
  (
    n652,
    n95
  );


  not
  g432
  (
    n278,
    n59
  );


  not
  g433
  (
    n525,
    n86
  );


  not
  g434
  (
    n221,
    n64
  );


  not
  g435
  (
    n391,
    n80
  );


  not
  g436
  (
    n228,
    n81
  );


  buf
  g437
  (
    n667,
    n71
  );


  not
  g438
  (
    n508,
    n152
  );


  buf
  g439
  (
    n665,
    n119
  );


  buf
  g440
  (
    n250,
    n41
  );


  buf
  g441
  (
    n554,
    n35
  );


  buf
  g442
  (
    n174,
    n147
  );


  buf
  g443
  (
    n275,
    n123
  );


  buf
  g444
  (
    n465,
    n101
  );


  buf
  g445
  (
    n364,
    n54
  );


  buf
  g446
  (
    n542,
    n123
  );


  buf
  g447
  (
    n472,
    n51
  );


  not
  g448
  (
    n209,
    n124
  );


  buf
  g449
  (
    n493,
    n74
  );


  buf
  g450
  (
    n561,
    n143
  );


  buf
  g451
  (
    n563,
    n138
  );


  buf
  g452
  (
    n427,
    n48
  );


  not
  g453
  (
    n522,
    n34
  );


  not
  g454
  (
    n544,
    n145
  );


  buf
  g455
  (
    n604,
    n96
  );


  not
  g456
  (
    n245,
    n159
  );


  buf
  g457
  (
    n232,
    n86
  );


  buf
  g458
  (
    n411,
    n128
  );


  buf
  g459
  (
    n672,
    n77
  );


  not
  g460
  (
    n222,
    n82
  );


  buf
  g461
  (
    n201,
    n65
  );


  not
  g462
  (
    n280,
    n90
  );


  buf
  g463
  (
    n179,
    n84
  );


  buf
  g464
  (
    KeyWire_0_37,
    n146
  );


  not
  g465
  (
    n464,
    n34
  );


  not
  g466
  (
    n524,
    n103
  );


  not
  g467
  (
    n347,
    n54
  );


  buf
  g468
  (
    n194,
    n125
  );


  not
  g469
  (
    n199,
    n138
  );


  buf
  g470
  (
    n538,
    n109
  );


  not
  g471
  (
    n303,
    n126
  );


  not
  g472
  (
    n590,
    n156
  );


  not
  g473
  (
    n244,
    n83
  );


  not
  g474
  (
    n468,
    n159
  );


  not
  g475
  (
    n584,
    n68
  );


  buf
  g476
  (
    n389,
    n116
  );


  not
  g477
  (
    n653,
    n59
  );


  not
  g478
  (
    n507,
    n118
  );


  not
  g479
  (
    n668,
    n37
  );


  buf
  g480
  (
    n650,
    n78
  );


  buf
  g481
  (
    n353,
    n62
  );


  buf
  g482
  (
    n608,
    n121
  );


  buf
  g483
  (
    n566,
    n153
  );


  not
  g484
  (
    n530,
    n126
  );


  not
  g485
  (
    n574,
    n98
  );


  not
  g486
  (
    n514,
    n37
  );


  not
  g487
  (
    n167,
    n70
  );


  buf
  g488
  (
    n359,
    n36
  );


  not
  g489
  (
    n423,
    n84
  );


  not
  g490
  (
    n587,
    n123
  );


  buf
  g491
  (
    n552,
    n119
  );


  buf
  g492
  (
    n455,
    n143
  );


  not
  g493
  (
    n319,
    n144
  );


  not
  g494
  (
    n532,
    n56
  );


  not
  g495
  (
    KeyWire_0_10,
    n45
  );


  not
  g496
  (
    n246,
    n97
  );


  not
  g497
  (
    n490,
    n35
  );


  buf
  g498
  (
    n352,
    n136
  );


  not
  g499
  (
    n621,
    n99
  );


  buf
  g500
  (
    n562,
    n154
  );


  not
  g501
  (
    n386,
    n146
  );


  buf
  g502
  (
    n317,
    n99
  );


  buf
  g503
  (
    n521,
    n75
  );


  not
  g504
  (
    n331,
    n120
  );


  not
  g505
  (
    n482,
    n38
  );


  not
  g506
  (
    n624,
    n143
  );


  not
  g507
  (
    n366,
    n102
  );


  not
  g508
  (
    n479,
    n148
  );


  not
  g509
  (
    n330,
    n96
  );


  not
  g510
  (
    n555,
    n106
  );


  buf
  g511
  (
    n383,
    n93
  );


  not
  g512
  (
    n513,
    n33
  );


  not
  g513
  (
    n193,
    n85
  );


  not
  g514
  (
    n609,
    n68
  );


  not
  g515
  (
    n633,
    n66
  );


  buf
  g516
  (
    n231,
    n133
  );


  not
  g517
  (
    n283,
    n135
  );


  not
  g518
  (
    n439,
    n110
  );


  not
  g519
  (
    n596,
    n144
  );


  not
  g520
  (
    n553,
    n116
  );


  not
  g521
  (
    n363,
    n122
  );


  not
  g522
  (
    n580,
    n103
  );


  buf
  g523
  (
    n163,
    n93
  );


  buf
  g524
  (
    n282,
    n129
  );


  not
  g525
  (
    n211,
    n133
  );


  not
  g526
  (
    n480,
    n63
  );


  not
  g527
  (
    n356,
    n48
  );


  buf
  g528
  (
    n233,
    n139
  );


  not
  g529
  (
    n326,
    n141
  );


  buf
  g530
  (
    n612,
    n134
  );


  buf
  g531
  (
    n327,
    n140
  );


  not
  g532
  (
    n339,
    n76
  );


  buf
  g533
  (
    n196,
    n124
  );


  buf
  g534
  (
    n641,
    n130
  );


  buf
  g535
  (
    n236,
    n151
  );


  not
  g536
  (
    n324,
    n112
  );


  not
  g537
  (
    n429,
    n153
  );


  buf
  g538
  (
    n414,
    n37
  );


  buf
  g539
  (
    n557,
    n135
  );


  not
  g540
  (
    n177,
    n140
  );


  buf
  g541
  (
    n603,
    n104
  );


  buf
  g542
  (
    KeyWire_0_39,
    n103
  );


  buf
  g543
  (
    n309,
    n100
  );


  not
  g544
  (
    n252,
    n76
  );


  not
  g545
  (
    n225,
    n119
  );


  buf
  g546
  (
    n227,
    n151
  );


  buf
  g547
  (
    n486,
    n130
  );


  buf
  g548
  (
    n548,
    n150
  );


  buf
  g549
  (
    n550,
    n73
  );


  not
  g550
  (
    n549,
    n134
  );


  buf
  g551
  (
    n373,
    n121
  );


  buf
  g552
  (
    n376,
    n156
  );


  buf
  g553
  (
    n279,
    n63
  );


  buf
  g554
  (
    n381,
    n149
  );


  buf
  g555
  (
    n266,
    n137
  );


  not
  g556
  (
    n499,
    n46
  );


  buf
  g557
  (
    n260,
    n125
  );


  not
  g558
  (
    n323,
    n82
  );


  buf
  g559
  (
    n192,
    n56
  );


  not
  g560
  (
    n639,
    n106
  );


  buf
  g561
  (
    n577,
    n50
  );


  not
  g562
  (
    n626,
    n105
  );


  not
  g563
  (
    n258,
    n87
  );


  buf
  g564
  (
    n576,
    n41
  );


  buf
  g565
  (
    n428,
    n63
  );


  not
  g566
  (
    n200,
    n117
  );


  not
  g567
  (
    n529,
    n87
  );


  not
  g568
  (
    n432,
    n42
  );


  not
  g569
  (
    n418,
    n151
  );


  not
  g570
  (
    n372,
    n36
  );


  not
  g571
  (
    n378,
    n42
  );


  buf
  g572
  (
    n551,
    n108
  );


  not
  g573
  (
    n367,
    n47
  );


  buf
  g574
  (
    n344,
    n81
  );


  buf
  g575
  (
    n443,
    n90
  );


  buf
  g576
  (
    n583,
    n44
  );


  not
  g577
  (
    n318,
    n107
  );


  buf
  g578
  (
    n457,
    n71
  );


  not
  g579
  (
    n202,
    n80
  );


  buf
  g580
  (
    n588,
    n88
  );


  not
  g581
  (
    n325,
    n145
  );


  buf
  g582
  (
    n656,
    n69
  );


  not
  g583
  (
    n579,
    n147
  );


  not
  g584
  (
    n395,
    n147
  );


  not
  g585
  (
    n285,
    n125
  );


  not
  g586
  (
    n449,
    n98
  );


  buf
  g587
  (
    n369,
    n128
  );


  buf
  g588
  (
    n332,
    n54
  );


  buf
  g589
  (
    n491,
    n94
  );


  buf
  g590
  (
    n453,
    n102
  );


  buf
  g591
  (
    n454,
    n147
  );


  buf
  g592
  (
    n240,
    n42
  );


  not
  g593
  (
    n503,
    n77
  );


  buf
  g594
  (
    n597,
    n131
  );


  not
  g595
  (
    n497,
    n114
  );


  not
  g596
  (
    n512,
    n37
  );


  buf
  g597
  (
    n556,
    n61
  );


  buf
  g598
  (
    KeyWire_0_8,
    n111
  );


  not
  g599
  (
    n355,
    n40
  );


  buf
  g600
  (
    n511,
    n60
  );


  not
  g601
  (
    n643,
    n34
  );


  not
  g602
  (
    n214,
    n140
  );


  not
  g603
  (
    n671,
    n66
  );


  not
  g604
  (
    n298,
    n50
  );


  buf
  g605
  (
    n384,
    n61
  );


  buf
  g606
  (
    n663,
    n69
  );


  not
  g607
  (
    n393,
    n114
  );


  not
  g608
  (
    n329,
    n56
  );


  not
  g609
  (
    n396,
    n33
  );


  not
  g610
  (
    n195,
    n126
  );


  not
  g611
  (
    n253,
    n84
  );


  buf
  g612
  (
    n570,
    n159
  );


  not
  g613
  (
    n664,
    n152
  );


  buf
  g614
  (
    n207,
    n79
  );


  buf
  g615
  (
    n243,
    n49
  );


  buf
  g616
  (
    n649,
    n156
  );


  not
  g617
  (
    n494,
    n83
  );


  buf
  g618
  (
    n394,
    n111
  );


  buf
  g619
  (
    n413,
    n43
  );


  not
  g620
  (
    n451,
    n57
  );


  buf
  g621
  (
    n478,
    n41
  );


  buf
  g622
  (
    n528,
    n34
  );


  not
  g623
  (
    n313,
    n96
  );


  buf
  g624
  (
    n519,
    n36
  );


  buf
  g625
  (
    n628,
    n134
  );


  buf
  g626
  (
    n607,
    n124
  );


  buf
  g627
  (
    n595,
    n155
  );


  not
  g628
  (
    n166,
    n131
  );


  not
  g629
  (
    n180,
    n155
  );


  not
  g630
  (
    KeyWire_0_1,
    n89
  );


  buf
  g631
  (
    n501,
    n137
  );


  buf
  g632
  (
    n380,
    n108
  );


  not
  g633
  (
    n287,
    n65
  );


  buf
  g634
  (
    n342,
    n55
  );


  not
  g635
  (
    n506,
    n109
  );


  not
  g636
  (
    n492,
    n98
  );


  not
  g637
  (
    KeyWire_0_30,
    n97
  );


  not
  g638
  (
    n162,
    n55
  );


  not
  g639
  (
    n263,
    n78
  );


  not
  g640
  (
    n1558,
    n212
  );


  buf
  g641
  (
    n746,
    n388
  );


  not
  g642
  (
    n1271,
    n227
  );


  not
  g643
  (
    n1594,
    n338
  );


  not
  g644
  (
    n1331,
    n288
  );


  not
  g645
  (
    n1650,
    n309
  );


  not
  g646
  (
    n1023,
    n410
  );


  buf
  g647
  (
    n1196,
    n300
  );


  buf
  g648
  (
    n900,
    n254
  );


  buf
  g649
  (
    n1007,
    n268
  );


  buf
  g650
  (
    n1349,
    n233
  );


  buf
  g651
  (
    n1153,
    n318
  );


  not
  g652
  (
    n679,
    n187
  );


  buf
  g653
  (
    n1458,
    n307
  );


  buf
  g654
  (
    n1629,
    n330
  );


  not
  g655
  (
    n1108,
    n204
  );


  not
  g656
  (
    n932,
    n372
  );


  not
  g657
  (
    KeyWire_0_61,
    n402
  );


  not
  g658
  (
    n1563,
    n307
  );


  not
  g659
  (
    n1200,
    n281
  );


  not
  g660
  (
    n1026,
    n354
  );


  not
  g661
  (
    n1692,
    n324
  );


  buf
  g662
  (
    n1649,
    n310
  );


  buf
  g663
  (
    n1336,
    n295
  );


  buf
  g664
  (
    n1579,
    n390
  );


  not
  g665
  (
    n818,
    n289
  );


  not
  g666
  (
    n1374,
    n285
  );


  buf
  g667
  (
    n1542,
    n218
  );


  buf
  g668
  (
    n720,
    n388
  );


  not
  g669
  (
    n774,
    n204
  );


  not
  g670
  (
    n1651,
    n199
  );


  not
  g671
  (
    n1203,
    n214
  );


  not
  g672
  (
    n1410,
    n219
  );


  not
  g673
  (
    n1597,
    n416
  );


  not
  g674
  (
    n993,
    n347
  );


  not
  g675
  (
    n842,
    n390
  );


  not
  g676
  (
    n896,
    n321
  );


  not
  g677
  (
    n1378,
    n186
  );


  buf
  g678
  (
    n1300,
    n232
  );


  not
  g679
  (
    n1494,
    n217
  );


  buf
  g680
  (
    n1146,
    n311
  );


  buf
  g681
  (
    n1113,
    n318
  );


  buf
  g682
  (
    n937,
    n303
  );


  not
  g683
  (
    n817,
    n238
  );


  buf
  g684
  (
    n870,
    n216
  );


  buf
  g685
  (
    n1583,
    n343
  );


  buf
  g686
  (
    n1325,
    n400
  );


  buf
  g687
  (
    n1642,
    n327
  );


  buf
  g688
  (
    n813,
    n392
  );


  buf
  g689
  (
    n1001,
    n337
  );


  not
  g690
  (
    n934,
    n406
  );


  buf
  g691
  (
    n1136,
    n298
  );


  buf
  g692
  (
    n749,
    n385
  );


  not
  g693
  (
    n1469,
    n272
  );


  buf
  g694
  (
    n907,
    n260
  );


  not
  g695
  (
    n897,
    n360
  );


  not
  g696
  (
    n841,
    n332
  );


  buf
  g697
  (
    n918,
    n267
  );


  not
  g698
  (
    n1332,
    n329
  );


  buf
  g699
  (
    n1387,
    n297
  );


  buf
  g700
  (
    n1189,
    n373
  );


  buf
  g701
  (
    n1131,
    n180
  );


  buf
  g702
  (
    n827,
    n343
  );


  not
  g703
  (
    n1490,
    n385
  );


  not
  g704
  (
    n1018,
    n220
  );


  buf
  g705
  (
    n1264,
    n391
  );


  not
  g706
  (
    n1037,
    n294
  );


  not
  g707
  (
    n1057,
    n179
  );


  buf
  g708
  (
    n951,
    n205
  );


  buf
  g709
  (
    n799,
    n399
  );


  buf
  g710
  (
    n703,
    n364
  );


  buf
  g711
  (
    n1339,
    n357
  );


  buf
  g712
  (
    n1260,
    n377
  );


  not
  g713
  (
    n862,
    n271
  );


  buf
  g714
  (
    n1307,
    n334
  );


  not
  g715
  (
    n1086,
    n240
  );


  buf
  g716
  (
    n1219,
    n262
  );


  buf
  g717
  (
    n1110,
    n323
  );


  buf
  g718
  (
    n973,
    n223
  );


  buf
  g719
  (
    n1237,
    n294
  );


  buf
  g720
  (
    n1148,
    n348
  );


  not
  g721
  (
    n1523,
    n364
  );


  buf
  g722
  (
    n1002,
    n292
  );


  not
  g723
  (
    n1027,
    n352
  );


  not
  g724
  (
    n984,
    n310
  );


  not
  g725
  (
    n686,
    n172
  );


  buf
  g726
  (
    n944,
    n330
  );


  not
  g727
  (
    n1350,
    n258
  );


  buf
  g728
  (
    n1071,
    n311
  );


  not
  g729
  (
    n964,
    n389
  );


  not
  g730
  (
    n1353,
    n277
  );


  not
  g731
  (
    n1637,
    n383
  );


  buf
  g732
  (
    n1658,
    n304
  );


  buf
  g733
  (
    n1564,
    n242
  );


  buf
  g734
  (
    n1524,
    n362
  );


  not
  g735
  (
    n874,
    n193
  );


  not
  g736
  (
    n1643,
    n360
  );


  not
  g737
  (
    KeyWire_0_31,
    n198
  );


  not
  g738
  (
    n1068,
    n197
  );


  buf
  g739
  (
    n901,
    n287
  );


  not
  g740
  (
    n1638,
    n361
  );


  not
  g741
  (
    n1596,
    n343
  );


  buf
  g742
  (
    n1489,
    n245
  );


  not
  g743
  (
    n747,
    n164
  );


  not
  g744
  (
    n877,
    n249
  );


  not
  g745
  (
    n1212,
    n204
  );


  not
  g746
  (
    n821,
    n245
  );


  buf
  g747
  (
    n927,
    n161
  );


  buf
  g748
  (
    n1053,
    n349
  );


  buf
  g749
  (
    n926,
    n340
  );


  buf
  g750
  (
    n681,
    n281
  );


  buf
  g751
  (
    n911,
    n320
  );


  not
  g752
  (
    n1622,
    n282
  );


  buf
  g753
  (
    n1101,
    n164
  );


  buf
  g754
  (
    n1299,
    n193
  );


  buf
  g755
  (
    n1459,
    n267
  );


  not
  g756
  (
    n1653,
    n363
  );


  buf
  g757
  (
    n775,
    n304
  );


  not
  g758
  (
    n1566,
    n348
  );


  buf
  g759
  (
    n1565,
    n201
  );


  buf
  g760
  (
    n715,
    n168
  );


  buf
  g761
  (
    n733,
    n384
  );


  not
  g762
  (
    n1655,
    n416
  );


  buf
  g763
  (
    n1497,
    n327
  );


  not
  g764
  (
    n816,
    n397
  );


  not
  g765
  (
    KeyWire_0_0,
    n187
  );


  buf
  g766
  (
    n1054,
    n272
  );


  not
  g767
  (
    n963,
    n170
  );


  buf
  g768
  (
    n737,
    n412
  );


  not
  g769
  (
    n903,
    n300
  );


  not
  g770
  (
    n1083,
    n276
  );


  not
  g771
  (
    n1283,
    n395
  );


  not
  g772
  (
    n1115,
    n287
  );


  not
  g773
  (
    n975,
    n223
  );


  not
  g774
  (
    n1373,
    n236
  );


  not
  g775
  (
    n1150,
    n254
  );


  not
  g776
  (
    n1227,
    n253
  );


  not
  g777
  (
    n1217,
    n295
  );


  buf
  g778
  (
    n754,
    n339
  );


  not
  g779
  (
    n1248,
    n285
  );


  not
  g780
  (
    n1278,
    n208
  );


  not
  g781
  (
    n1509,
    n382
  );


  not
  g782
  (
    n1379,
    n172
  );


  not
  g783
  (
    n1134,
    n415
  );


  buf
  g784
  (
    n1298,
    n282
  );


  buf
  g785
  (
    n924,
    n265
  );


  buf
  g786
  (
    n1333,
    n305
  );


  not
  g787
  (
    n1439,
    n172
  );


  buf
  g788
  (
    n1364,
    n256
  );


  buf
  g789
  (
    n1614,
    n385
  );


  not
  g790
  (
    n1032,
    n406
  );


  buf
  g791
  (
    n717,
    n163
  );


  buf
  g792
  (
    n1309,
    n179
  );


  not
  g793
  (
    n688,
    n225
  );


  not
  g794
  (
    n1234,
    n346
  );


  buf
  g795
  (
    n1289,
    n210
  );


  buf
  g796
  (
    KeyWire_0_14,
    n381
  );


  buf
  g797
  (
    n1537,
    n239
  );


  buf
  g798
  (
    n1178,
    n398
  );


  not
  g799
  (
    n930,
    n279
  );


  not
  g800
  (
    n844,
    n350
  );


  buf
  g801
  (
    n750,
    n274
  );


  buf
  g802
  (
    n1475,
    n335
  );


  buf
  g803
  (
    n1423,
    n290
  );


  not
  g804
  (
    n1409,
    n368
  );


  not
  g805
  (
    n1449,
    n261
  );


  not
  g806
  (
    n795,
    n167
  );


  buf
  g807
  (
    n706,
    n361
  );


  not
  g808
  (
    n1345,
    n308
  );


  buf
  g809
  (
    n719,
    n284
  );


  not
  g810
  (
    n753,
    n363
  );


  buf
  g811
  (
    n1641,
    n241
  );


  not
  g812
  (
    n1140,
    n222
  );


  not
  g813
  (
    n758,
    n325
  );


  not
  g814
  (
    n1620,
    n257
  );


  buf
  g815
  (
    n1615,
    n199
  );


  not
  g816
  (
    n728,
    n312
  );


  not
  g817
  (
    n1100,
    n286
  );


  buf
  g818
  (
    KeyWire_0_21,
    n418
  );


  not
  g819
  (
    n804,
    n270
  );


  not
  g820
  (
    n1102,
    n340
  );


  not
  g821
  (
    n1575,
    n229
  );


  buf
  g822
  (
    n1647,
    n319
  );


  buf
  g823
  (
    n1005,
    n386
  );


  not
  g824
  (
    n1043,
    n338
  );


  buf
  g825
  (
    n1452,
    n368
  );


  buf
  g826
  (
    n755,
    n409
  );


  buf
  g827
  (
    n1367,
    n194
  );


  buf
  g828
  (
    n1482,
    n336
  );


  not
  g829
  (
    n1492,
    n303
  );


  buf
  g830
  (
    n1078,
    n204
  );


  buf
  g831
  (
    n1394,
    n281
  );


  buf
  g832
  (
    n1171,
    n279
  );


  not
  g833
  (
    n1224,
    n222
  );


  buf
  g834
  (
    n789,
    n324
  );


  buf
  g835
  (
    n676,
    n278
  );


  buf
  g836
  (
    n1540,
    n294
  );


  not
  g837
  (
    n1662,
    n218
  );


  not
  g838
  (
    n791,
    n215
  );


  buf
  g839
  (
    n731,
    n401
  );


  buf
  g840
  (
    n1044,
    n276
  );


  not
  g841
  (
    n947,
    n169
  );


  buf
  g842
  (
    n1699,
    n191
  );


  not
  g843
  (
    n887,
    n191
  );


  not
  g844
  (
    KeyWire_0_13,
    n376
  );


  not
  g845
  (
    n806,
    n183
  );


  not
  g846
  (
    n1022,
    n349
  );


  not
  g847
  (
    n1518,
    n397
  );


  buf
  g848
  (
    KeyWire_0_51,
    n327
  );


  buf
  g849
  (
    n914,
    n406
  );


  not
  g850
  (
    n1166,
    n293
  );


  buf
  g851
  (
    n1275,
    n202
  );


  buf
  g852
  (
    n1012,
    n209
  );


  buf
  g853
  (
    n1014,
    n229
  );


  buf
  g854
  (
    n1609,
    n350
  );


  not
  g855
  (
    n1436,
    n335
  );


  not
  g856
  (
    n1607,
    n205
  );


  not
  g857
  (
    n942,
    n333
  );


  buf
  g858
  (
    n761,
    n383
  );


  buf
  g859
  (
    n1125,
    n168
  );


  buf
  g860
  (
    n1446,
    n404
  );


  not
  g861
  (
    n1689,
    n369
  );


  not
  g862
  (
    n1210,
    n270
  );


  not
  g863
  (
    n1390,
    n192
  );


  not
  g864
  (
    n1198,
    n400
  );


  buf
  g865
  (
    n1317,
    n284
  );


  buf
  g866
  (
    n931,
    n205
  );


  buf
  g867
  (
    n982,
    n377
  );


  buf
  g868
  (
    n985,
    n283
  );


  buf
  g869
  (
    n690,
    n278
  );


  not
  g870
  (
    n1344,
    n277
  );


  buf
  g871
  (
    n1553,
    n406
  );


  buf
  g872
  (
    n1585,
    n206
  );


  buf
  g873
  (
    n1222,
    n242
  );


  not
  g874
  (
    n1672,
    n354
  );


  buf
  g875
  (
    n1130,
    n399
  );


  not
  g876
  (
    n1516,
    n418
  );


  buf
  g877
  (
    KeyWire_0_17,
    n407
  );


  buf
  g878
  (
    n809,
    n258
  );


  buf
  g879
  (
    n1049,
    n184
  );


  not
  g880
  (
    n1546,
    n208
  );


  not
  g881
  (
    n1569,
    n214
  );


  buf
  g882
  (
    n702,
    n273
  );


  not
  g883
  (
    KeyWire_0_56,
    n196
  );


  buf
  g884
  (
    n1371,
    n313
  );


  not
  g885
  (
    n990,
    n166
  );


  buf
  g886
  (
    n952,
    n397
  );


  buf
  g887
  (
    n1004,
    n323
  );


  buf
  g888
  (
    n1059,
    n273
  );


  buf
  g889
  (
    n1411,
    n197
  );


  buf
  g890
  (
    n1177,
    n312
  );


  not
  g891
  (
    n1408,
    n336
  );


  buf
  g892
  (
    n945,
    n395
  );


  not
  g893
  (
    n704,
    n356
  );


  buf
  g894
  (
    n936,
    n186
  );


  buf
  g895
  (
    n1074,
    n190
  );


  buf
  g896
  (
    n689,
    n286
  );


  not
  g897
  (
    n1500,
    n412
  );


  not
  g898
  (
    n958,
    n316
  );


  buf
  g899
  (
    n977,
    n329
  );


  buf
  g900
  (
    n859,
    n182
  );


  buf
  g901
  (
    n1605,
    n171
  );


  buf
  g902
  (
    n1046,
    n230
  );


  not
  g903
  (
    n1461,
    n246
  );


  not
  g904
  (
    n692,
    n212
  );


  not
  g905
  (
    n1175,
    n345
  );


  buf
  g906
  (
    n819,
    n170
  );


  not
  g907
  (
    n1556,
    n237
  );


  buf
  g908
  (
    n1104,
    n378
  );


  buf
  g909
  (
    n863,
    n184
  );


  not
  g910
  (
    n1360,
    n377
  );


  not
  g911
  (
    n710,
    n275
  );


  not
  g912
  (
    n796,
    n169
  );


  not
  g913
  (
    n1380,
    n401
  );


  buf
  g914
  (
    n741,
    n242
  );


  buf
  g915
  (
    n1242,
    n213
  );


  buf
  g916
  (
    n1486,
    n203
  );


  not
  g917
  (
    n768,
    n246
  );


  not
  g918
  (
    n1584,
    n399
  );


  not
  g919
  (
    n1343,
    n337
  );


  buf
  g920
  (
    KeyWire_0_44,
    n405
  );


  not
  g921
  (
    n1174,
    n387
  );


  buf
  g922
  (
    n997,
    n331
  );


  buf
  g923
  (
    n1589,
    n290
  );


  not
  g924
  (
    n868,
    n370
  );


  not
  g925
  (
    n1623,
    n403
  );


  not
  g926
  (
    KeyWire_0_41,
    n330
  );


  not
  g927
  (
    n1414,
    n171
  );


  buf
  g928
  (
    n1590,
    n209
  );


  buf
  g929
  (
    n1539,
    n312
  );


  not
  g930
  (
    n1286,
    n237
  );


  buf
  g931
  (
    n1520,
    n188
  );


  not
  g932
  (
    n1159,
    n302
  );


  buf
  g933
  (
    n1297,
    n278
  );


  buf
  g934
  (
    n1082,
    n357
  );


  buf
  g935
  (
    n1268,
    n316
  );


  not
  g936
  (
    n1006,
    n236
  );


  buf
  g937
  (
    n1478,
    n240
  );


  not
  g938
  (
    n1031,
    n176
  );


  buf
  g939
  (
    n1481,
    n395
  );


  buf
  g940
  (
    n1127,
    n227
  );


  buf
  g941
  (
    n1690,
    n250
  );


  buf
  g942
  (
    n743,
    n214
  );


  not
  g943
  (
    n826,
    n333
  );


  buf
  g944
  (
    n1443,
    n404
  );


  buf
  g945
  (
    n941,
    n315
  );


  buf
  g946
  (
    n1639,
    n295
  );


  buf
  g947
  (
    n851,
    n165
  );


  not
  g948
  (
    n1093,
    n416
  );


  not
  g949
  (
    n965,
    n223
  );


  buf
  g950
  (
    n1058,
    n314
  );


  buf
  g951
  (
    n849,
    n170
  );


  buf
  g952
  (
    n1693,
    n321
  );


  not
  g953
  (
    n1599,
    n344
  );


  not
  g954
  (
    n1199,
    n282
  );


  buf
  g955
  (
    n1337,
    n408
  );


  buf
  g956
  (
    n968,
    n198
  );


  not
  g957
  (
    n1571,
    n244
  );


  buf
  g958
  (
    n1259,
    n219
  );


  not
  g959
  (
    n1517,
    n329
  );


  not
  g960
  (
    n1499,
    n217
  );


  not
  g961
  (
    n1285,
    n201
  );


  buf
  g962
  (
    n1691,
    n297
  );


  not
  g963
  (
    n1510,
    n338
  );


  buf
  g964
  (
    n1657,
    n370
  );


  buf
  g965
  (
    n1531,
    n347
  );


  buf
  g966
  (
    n1602,
    n249
  );


  not
  g967
  (
    n736,
    n192
  );


  buf
  g968
  (
    n954,
    n180
  );


  buf
  g969
  (
    n1147,
    n188
  );


  buf
  g970
  (
    n1488,
    n234
  );


  not
  g971
  (
    n1515,
    n252
  );


  buf
  g972
  (
    n1149,
    n318
  );


  buf
  g973
  (
    n1274,
    n414
  );


  not
  g974
  (
    n1095,
    n390
  );


  buf
  g975
  (
    n788,
    n371
  );


  buf
  g976
  (
    n1273,
    n350
  );


  buf
  g977
  (
    n732,
    n221
  );


  buf
  g978
  (
    n1696,
    n215
  );


  not
  g979
  (
    n1342,
    n325
  );


  buf
  g980
  (
    n1467,
    n199
  );


  buf
  g981
  (
    n1055,
    n394
  );


  buf
  g982
  (
    n1105,
    n341
  );


  buf
  g983
  (
    n1120,
    n380
  );


  not
  g984
  (
    n1167,
    n349
  );


  not
  g985
  (
    n1070,
    n247
  );


  not
  g986
  (
    n684,
    n263
  );


  not
  g987
  (
    n1106,
    n251
  );


  buf
  g988
  (
    n1163,
    n413
  );


  buf
  g989
  (
    n1207,
    n324
  );


  not
  g990
  (
    n1256,
    n316
  );


  buf
  g991
  (
    n1107,
    n210
  );


  not
  g992
  (
    n1081,
    n414
  );


  buf
  g993
  (
    n1625,
    n217
  );


  not
  g994
  (
    KeyWire_0_50,
    n273
  );


  buf
  g995
  (
    n1326,
    n419
  );


  not
  g996
  (
    n1228,
    n192
  );


  not
  g997
  (
    n961,
    n361
  );


  not
  g998
  (
    n999,
    n164
  );


  not
  g999
  (
    n894,
    n309
  );


  not
  g1000
  (
    n1576,
    n394
  );


  buf
  g1001
  (
    n802,
    n270
  );


  not
  g1002
  (
    n835,
    n306
  );


  not
  g1003
  (
    n1635,
    n253
  );


  buf
  g1004
  (
    n673,
    n301
  );


  not
  g1005
  (
    n1533,
    n210
  );


  buf
  g1006
  (
    n1035,
    n309
  );


  not
  g1007
  (
    n880,
    n384
  );


  not
  g1008
  (
    n1385,
    n351
  );


  buf
  g1009
  (
    n1122,
    n198
  );


  buf
  g1010
  (
    n694,
    n233
  );


  buf
  g1011
  (
    n1347,
    n407
  );


  not
  g1012
  (
    KeyWire_0_47,
    n253
  );


  not
  g1013
  (
    n843,
    n254
  );


  not
  g1014
  (
    n1279,
    n188
  );


  buf
  g1015
  (
    n1440,
    n355
  );


  buf
  g1016
  (
    n1677,
    n293
  );


  not
  g1017
  (
    n986,
    n381
  );


  buf
  g1018
  (
    n1369,
    n371
  );


  buf
  g1019
  (
    n1588,
    n264
  );


  not
  g1020
  (
    n1169,
    n265
  );


  buf
  g1021
  (
    n1039,
    n236
  );


  not
  g1022
  (
    n1646,
    n367
  );


  not
  g1023
  (
    n1477,
    n166
  );


  buf
  g1024
  (
    n1389,
    n305
  );


  not
  g1025
  (
    n1016,
    n180
  );


  buf
  g1026
  (
    n1645,
    n286
  );


  buf
  g1027
  (
    n1214,
    n376
  );


  not
  g1028
  (
    n1435,
    n229
  );


  not
  g1029
  (
    n1610,
    n325
  );


  not
  g1030
  (
    n723,
    n370
  );


  not
  g1031
  (
    n861,
    n268
  );


  buf
  g1032
  (
    n1463,
    n263
  );


  not
  g1033
  (
    n1335,
    n212
  );


  not
  g1034
  (
    n1644,
    n187
  );


  buf
  g1035
  (
    n1664,
    n304
  );


  not
  g1036
  (
    n966,
    n346
  );


  buf
  g1037
  (
    n1617,
    n353
  );


  not
  g1038
  (
    n1474,
    n215
  );


  not
  g1039
  (
    n707,
    n417
  );


  buf
  g1040
  (
    n1399,
    n326
  );


  buf
  g1041
  (
    n693,
    n265
  );


  buf
  g1042
  (
    KeyWire_0_32,
    n287
  );


  not
  g1043
  (
    n832,
    n418
  );


  buf
  g1044
  (
    n815,
    n248
  );


  not
  g1045
  (
    n1258,
    n319
  );


  buf
  g1046
  (
    n829,
    n236
  );


  buf
  g1047
  (
    n722,
    n391
  );


  not
  g1048
  (
    n1666,
    n193
  );


  not
  g1049
  (
    n1253,
    n256
  );


  buf
  g1050
  (
    n1096,
    n315
  );


  not
  g1051
  (
    n1464,
    n369
  );


  buf
  g1052
  (
    n1315,
    n363
  );


  not
  g1053
  (
    n1397,
    n197
  );


  buf
  g1054
  (
    n1314,
    n298
  );


  not
  g1055
  (
    n1493,
    n206
  );


  not
  g1056
  (
    n883,
    n296
  );


  not
  g1057
  (
    n1451,
    n310
  );


  buf
  g1058
  (
    n1063,
    n216
  );


  not
  g1059
  (
    n701,
    n337
  );


  buf
  g1060
  (
    n1444,
    n319
  );


  not
  g1061
  (
    n1305,
    n372
  );


  not
  g1062
  (
    n1679,
    n374
  );


  buf
  g1063
  (
    n1158,
    n276
  );


  buf
  g1064
  (
    n1424,
    n386
  );


  not
  g1065
  (
    n996,
    n213
  );


  buf
  g1066
  (
    n1247,
    n227
  );


  buf
  g1067
  (
    n1176,
    n173
  );


  buf
  g1068
  (
    n1181,
    n230
  );


  buf
  g1069
  (
    n1422,
    n167
  );


  buf
  g1070
  (
    n1220,
    n311
  );


  buf
  g1071
  (
    n1073,
    n165
  );


  not
  g1072
  (
    n1302,
    n225
  );


  not
  g1073
  (
    n910,
    n412
  );


  buf
  g1074
  (
    n836,
    n258
  );


  buf
  g1075
  (
    n1631,
    n394
  );


  not
  g1076
  (
    n1077,
    n218
  );


  not
  g1077
  (
    n1321,
    n203
  );


  not
  g1078
  (
    n1580,
    n374
  );


  buf
  g1079
  (
    n1051,
    n246
  );


  not
  g1080
  (
    n1328,
    n181
  );


  not
  g1081
  (
    n1396,
    n407
  );


  not
  g1082
  (
    n846,
    n279
  );


  buf
  g1083
  (
    n797,
    n290
  );


  not
  g1084
  (
    n678,
    n299
  );


  buf
  g1085
  (
    n1097,
    n163
  );


  not
  g1086
  (
    n1544,
    n305
  );


  buf
  g1087
  (
    n675,
    n228
  );


  not
  g1088
  (
    n1240,
    n380
  );


  buf
  g1089
  (
    n1080,
    n175
  );


  buf
  g1090
  (
    n1138,
    n401
  );


  not
  g1091
  (
    n1067,
    n225
  );


  not
  g1092
  (
    n1455,
    n194
  );


  buf
  g1093
  (
    n691,
    n343
  );


  buf
  g1094
  (
    n1291,
    n174
  );


  not
  g1095
  (
    n1266,
    n368
  );


  not
  g1096
  (
    n1334,
    n178
  );


  buf
  g1097
  (
    n1126,
    n412
  );


  not
  g1098
  (
    n1479,
    n235
  );


  buf
  g1099
  (
    n935,
    n371
  );


  not
  g1100
  (
    n1124,
    n289
  );


  buf
  g1101
  (
    n1603,
    n258
  );


  buf
  g1102
  (
    n1604,
    n195
  );


  buf
  g1103
  (
    KeyWire_0_16,
    n411
  );


  not
  g1104
  (
    n1245,
    n391
  );


  not
  g1105
  (
    n1504,
    n298
  );


  not
  g1106
  (
    n1249,
    n171
  );


  not
  g1107
  (
    n784,
    n322
  );


  buf
  g1108
  (
    n1034,
    n177
  );


  not
  g1109
  (
    n1064,
    n269
  );


  not
  g1110
  (
    n948,
    n161
  );


  not
  g1111
  (
    n1182,
    n232
  );


  not
  g1112
  (
    n1398,
    n244
  );


  buf
  g1113
  (
    n1688,
    n303
  );


  buf
  g1114
  (
    n1574,
    n206
  );


  not
  g1115
  (
    n726,
    n373
  );


  buf
  g1116
  (
    n909,
    n241
  );


  buf
  g1117
  (
    n1506,
    n408
  );


  not
  g1118
  (
    n1392,
    n171
  );


  buf
  g1119
  (
    n946,
    n355
  );


  buf
  g1120
  (
    n866,
    n256
  );


  not
  g1121
  (
    n916,
    n170
  );


  not
  g1122
  (
    n1634,
    n331
  );


  not
  g1123
  (
    n1184,
    n416
  );


  buf
  g1124
  (
    n1372,
    n306
  );


  not
  g1125
  (
    n923,
    n414
  );


  buf
  g1126
  (
    n1238,
    n313
  );


  buf
  g1127
  (
    n1473,
    n317
  );


  buf
  g1128
  (
    n1521,
    n391
  );


  not
  g1129
  (
    n1484,
    n228
  );


  not
  g1130
  (
    n1303,
    n333
  );


  buf
  g1131
  (
    n1251,
    n271
  );


  not
  g1132
  (
    n987,
    n248
  );


  buf
  g1133
  (
    n1438,
    n261
  );


  buf
  g1134
  (
    n1572,
    n238
  );


  not
  g1135
  (
    n1562,
    n189
  );


  not
  g1136
  (
    n1340,
    n174
  );


  not
  g1137
  (
    n1262,
    n292
  );


  not
  g1138
  (
    n820,
    n244
  );


  not
  g1139
  (
    n962,
    n285
  );


  buf
  g1140
  (
    n1040,
    n286
  );


  not
  g1141
  (
    n721,
    n385
  );


  buf
  g1142
  (
    n1447,
    n247
  );


  buf
  g1143
  (
    n1694,
    n181
  );


  not
  g1144
  (
    n1555,
    n167
  );


  not
  g1145
  (
    n1412,
    n226
  );


  buf
  g1146
  (
    n756,
    n299
  );


  not
  g1147
  (
    n1141,
    n342
  );


  not
  g1148
  (
    n1038,
    n352
  );


  not
  g1149
  (
    n839,
    n235
  );


  not
  g1150
  (
    n1429,
    n267
  );


  not
  g1151
  (
    n830,
    n331
  );


  buf
  g1152
  (
    n1684,
    n313
  );


  not
  g1153
  (
    n1172,
    n285
  );


  buf
  g1154
  (
    n831,
    n302
  );


  buf
  g1155
  (
    n724,
    n210
  );


  buf
  g1156
  (
    n853,
    n315
  );


  buf
  g1157
  (
    n1388,
    n162
  );


  buf
  g1158
  (
    n1324,
    n243
  );


  buf
  g1159
  (
    n1570,
    n252
  );


  buf
  g1160
  (
    n1202,
    n381
  );


  buf
  g1161
  (
    n1025,
    n220
  );


  not
  g1162
  (
    n1045,
    n243
  );


  not
  g1163
  (
    n1468,
    n280
  );


  buf
  g1164
  (
    n1129,
    n208
  );


  not
  g1165
  (
    n1033,
    n282
  );


  not
  g1166
  (
    n1621,
    n183
  );


  not
  g1167
  (
    n698,
    n201
  );


  buf
  g1168
  (
    KeyWire_0_53,
    n297
  );


  not
  g1169
  (
    n1180,
    n226
  );


  not
  g1170
  (
    n995,
    n200
  );


  buf
  g1171
  (
    n1470,
    n319
  );


  buf
  g1172
  (
    n1652,
    n393
  );


  not
  g1173
  (
    n1527,
    n270
  );


  buf
  g1174
  (
    n848,
    n186
  );


  buf
  g1175
  (
    n889,
    n362
  );


  not
  g1176
  (
    n805,
    n226
  );


  not
  g1177
  (
    n1287,
    n320
  );


  not
  g1178
  (
    n1352,
    n173
  );


  buf
  g1179
  (
    n807,
    n356
  );


  not
  g1180
  (
    n1462,
    n268
  );


  buf
  g1181
  (
    n840,
    n313
  );


  buf
  g1182
  (
    n1195,
    n311
  );


  buf
  g1183
  (
    n769,
    n201
  );


  buf
  g1184
  (
    n1229,
    n195
  );


  buf
  g1185
  (
    n1111,
    n383
  );


  not
  g1186
  (
    n1281,
    n198
  );


  not
  g1187
  (
    n1151,
    n251
  );


  buf
  g1188
  (
    n1681,
    n275
  );


  not
  g1189
  (
    n1183,
    n405
  );


  buf
  g1190
  (
    n1362,
    n413
  );


  buf
  g1191
  (
    n1296,
    n202
  );


  not
  g1192
  (
    KeyWire_0_45,
    n305
  );


  not
  g1193
  (
    n1512,
    n402
  );


  not
  g1194
  (
    n781,
    n389
  );


  buf
  g1195
  (
    n1030,
    n255
  );


  not
  g1196
  (
    n1072,
    n178
  );


  buf
  g1197
  (
    n1319,
    n358
  );


  buf
  g1198
  (
    n1327,
    n302
  );


  not
  g1199
  (
    n1232,
    n336
  );


  not
  g1200
  (
    n1630,
    n341
  );


  buf
  g1201
  (
    n847,
    n410
  );


  not
  g1202
  (
    n1508,
    n228
  );


  not
  g1203
  (
    n1257,
    n367
  );


  buf
  g1204
  (
    n759,
    n173
  );


  not
  g1205
  (
    n1656,
    n189
  );


  not
  g1206
  (
    n1277,
    n253
  );


  buf
  g1207
  (
    n1263,
    n351
  );


  not
  g1208
  (
    n825,
    n316
  );


  buf
  g1209
  (
    n950,
    n211
  );


  not
  g1210
  (
    n1441,
    n252
  );


  buf
  g1211
  (
    n1526,
    n267
  );


  not
  g1212
  (
    n1329,
    n323
  );


  not
  g1213
  (
    n1087,
    n308
  );


  buf
  g1214
  (
    n1310,
    n168
  );


  not
  g1215
  (
    n1156,
    n366
  );


  buf
  g1216
  (
    n1164,
    n217
  );


  buf
  g1217
  (
    n1582,
    n339
  );


  not
  g1218
  (
    n705,
    n289
  );


  buf
  g1219
  (
    n748,
    n173
  );


  not
  g1220
  (
    n1206,
    n339
  );


  buf
  g1221
  (
    n1193,
    n380
  );


  not
  g1222
  (
    n1428,
    n353
  );


  buf
  g1223
  (
    n1123,
    n231
  );


  not
  g1224
  (
    n1304,
    n303
  );


  buf
  g1225
  (
    n763,
    n273
  );


  buf
  g1226
  (
    n886,
    n200
  );


  buf
  g1227
  (
    n687,
    n300
  );


  not
  g1228
  (
    n760,
    n209
  );


  buf
  g1229
  (
    n1507,
    n396
  );


  not
  g1230
  (
    n872,
    n363
  );


  buf
  g1231
  (
    n1483,
    n404
  );


  buf
  g1232
  (
    n1092,
    n255
  );


  not
  g1233
  (
    n885,
    n278
  );


  buf
  g1234
  (
    KeyWire_0_48,
    n384
  );


  buf
  g1235
  (
    n1368,
    n411
  );


  not
  g1236
  (
    n915,
    n301
  );


  not
  g1237
  (
    n766,
    n317
  );


  buf
  g1238
  (
    n1254,
    n259
  );


  not
  g1239
  (
    n1323,
    n378
  );


  not
  g1240
  (
    n682,
    n194
  );


  not
  g1241
  (
    n879,
    n237
  );


  not
  g1242
  (
    n1320,
    n231
  );


  buf
  g1243
  (
    n1534,
    n181
  );


  not
  g1244
  (
    n1290,
    n400
  );


  not
  g1245
  (
    n1405,
    n335
  );


  not
  g1246
  (
    n884,
    n393
  );


  not
  g1247
  (
    n983,
    n224
  );


  not
  g1248
  (
    n899,
    n387
  );


  buf
  g1249
  (
    n1205,
    n274
  );


  not
  g1250
  (
    n1230,
    n219
  );


  buf
  g1251
  (
    n1495,
    n354
  );


  buf
  g1252
  (
    n1015,
    n191
  );


  buf
  g1253
  (
    n1491,
    n359
  );


  buf
  g1254
  (
    n1209,
    n324
  );


  not
  g1255
  (
    n1686,
    n195
  );


  not
  g1256
  (
    n1119,
    n381
  );


  buf
  g1257
  (
    n740,
    n317
  );


  buf
  g1258
  (
    n920,
    n280
  );


  buf
  g1259
  (
    n1395,
    n373
  );


  not
  g1260
  (
    n1619,
    n299
  );


  buf
  g1261
  (
    n860,
    n329
  );


  not
  g1262
  (
    n1308,
    n250
  );


  buf
  g1263
  (
    n898,
    n228
  );


  not
  g1264
  (
    n1384,
    n256
  );


  not
  g1265
  (
    n857,
    n203
  );


  buf
  g1266
  (
    n1383,
    n186
  );


  buf
  g1267
  (
    n1019,
    n238
  );


  buf
  g1268
  (
    n867,
    n252
  );


  buf
  g1269
  (
    n782,
    n283
  );


  buf
  g1270
  (
    n1062,
    n220
  );


  buf
  g1271
  (
    n1680,
    n320
  );


  buf
  g1272
  (
    n1060,
    n350
  );


  not
  g1273
  (
    n1514,
    n379
  );


  buf
  g1274
  (
    n989,
    n207
  );


  buf
  g1275
  (
    n1370,
    n331
  );


  buf
  g1276
  (
    n1415,
    n362
  );


  buf
  g1277
  (
    n1437,
    n272
  );


  buf
  g1278
  (
    n785,
    n208
  );


  buf
  g1279
  (
    n1687,
    n238
  );


  not
  g1280
  (
    n978,
    n266
  );


  buf
  g1281
  (
    n837,
    n178
  );


  not
  g1282
  (
    n751,
    n221
  );


  not
  g1283
  (
    n1400,
    n321
  );


  buf
  g1284
  (
    n1363,
    n369
  );


  buf
  g1285
  (
    n893,
    n375
  );


  not
  g1286
  (
    n716,
    n232
  );


  buf
  g1287
  (
    n1204,
    n235
  );


  not
  g1288
  (
    n1215,
    n202
  );


  buf
  g1289
  (
    n1450,
    n178
  );


  not
  g1290
  (
    n1048,
    n396
  );


  buf
  g1291
  (
    n711,
    n359
  );


  buf
  g1292
  (
    n1085,
    n352
  );


  buf
  g1293
  (
    n1535,
    n280
  );


  not
  g1294
  (
    n1135,
    n176
  );


  buf
  g1295
  (
    n1543,
    n239
  );


  not
  g1296
  (
    n1503,
    n293
  );


  not
  g1297
  (
    n957,
    n284
  );


  not
  g1298
  (
    n1261,
    n189
  );


  not
  g1299
  (
    n1354,
    n335
  );


  buf
  g1300
  (
    n1118,
    n410
  );


  buf
  g1301
  (
    n959,
    n167
  );


  buf
  g1302
  (
    n677,
    n200
  );


  not
  g1303
  (
    n876,
    n408
  );


  not
  g1304
  (
    n1557,
    n207
  );


  not
  g1305
  (
    n773,
    n332
  );


  not
  g1306
  (
    n1190,
    n417
  );


  buf
  g1307
  (
    n730,
    n405
  );


  buf
  g1308
  (
    n981,
    n366
  );


  not
  g1309
  (
    n1616,
    n243
  );


  not
  g1310
  (
    n787,
    n288
  );


  not
  g1311
  (
    n1430,
    n372
  );


  buf
  g1312
  (
    n1338,
    n386
  );


  not
  g1313
  (
    n1365,
    n247
  );


  buf
  g1314
  (
    n1377,
    n322
  );


  buf
  g1315
  (
    n1269,
    n354
  );


  buf
  g1316
  (
    n1084,
    n241
  );


  buf
  g1317
  (
    n1675,
    n231
  );


  not
  g1318
  (
    n764,
    n264
  );


  buf
  g1319
  (
    n1201,
    n292
  );


  buf
  g1320
  (
    n1221,
    n291
  );


  not
  g1321
  (
    n1236,
    n211
  );


  not
  g1322
  (
    n905,
    n359
  );


  buf
  g1323
  (
    n1216,
    n366
  );


  not
  g1324
  (
    n939,
    n263
  );


  buf
  g1325
  (
    n1393,
    n260
  );


  buf
  g1326
  (
    n967,
    n195
  );


  buf
  g1327
  (
    n1416,
    n246
  );


  buf
  g1328
  (
    n882,
    n360
  );


  not
  g1329
  (
    KeyWire_0_28,
    n361
  );


  buf
  g1330
  (
    n1160,
    n182
  );


  not
  g1331
  (
    n772,
    n239
  );


  not
  g1332
  (
    n1671,
    n224
  );


  not
  g1333
  (
    n1313,
    n392
  );


  buf
  g1334
  (
    n1663,
    n374
  );


  not
  g1335
  (
    n1050,
    n365
  );


  not
  g1336
  (
    n891,
    n257
  );


  not
  g1337
  (
    n943,
    n388
  );


  buf
  g1338
  (
    n1358,
    n339
  );


  buf
  g1339
  (
    n1255,
    n320
  );


  buf
  g1340
  (
    n1420,
    n200
  );


  buf
  g1341
  (
    n1480,
    n418
  );


  not
  g1342
  (
    n1357,
    n325
  );


  not
  g1343
  (
    KeyWire_0_19,
    n269
  );


  buf
  g1344
  (
    n1079,
    n211
  );


  not
  g1345
  (
    n1295,
    n261
  );


  not
  g1346
  (
    n890,
    n269
  );


  not
  g1347
  (
    n1528,
    n353
  );


  not
  g1348
  (
    n744,
    n344
  );


  buf
  g1349
  (
    n1626,
    n372
  );


  not
  g1350
  (
    n683,
    n352
  );


  not
  g1351
  (
    n680,
    n315
  );


  not
  g1352
  (
    n956,
    n362
  );


  buf
  g1353
  (
    n994,
    n399
  );


  not
  g1354
  (
    n738,
    n410
  );


  not
  g1355
  (
    n1186,
    n375
  );


  buf
  g1356
  (
    n1292,
    n341
  );


  buf
  g1357
  (
    n971,
    n379
  );


  buf
  g1358
  (
    n786,
    n259
  );


  not
  g1359
  (
    n1114,
    n300
  );


  not
  g1360
  (
    n955,
    n185
  );


  buf
  g1361
  (
    n906,
    n265
  );


  buf
  g1362
  (
    n1453,
    n390
  );


  not
  g1363
  (
    n1601,
    n192
  );


  not
  g1364
  (
    n992,
    n414
  );


  not
  g1365
  (
    n1538,
    n301
  );


  not
  g1366
  (
    n892,
    n386
  );


  buf
  g1367
  (
    n1432,
    n179
  );


  buf
  g1368
  (
    n1211,
    n308
  );


  not
  g1369
  (
    n1021,
    n207
  );


  not
  g1370
  (
    n1144,
    n358
  );


  not
  g1371
  (
    n792,
    n234
  );


  not
  g1372
  (
    n1382,
    n326
  );


  not
  g1373
  (
    n1628,
    n254
  );


  not
  g1374
  (
    n970,
    n262
  );


  not
  g1375
  (
    n1525,
    n403
  );


  buf
  g1376
  (
    n1433,
    n378
  );


  buf
  g1377
  (
    n1573,
    n244
  );


  buf
  g1378
  (
    n928,
    n342
  );


  buf
  g1379
  (
    n1636,
    n177
  );


  not
  g1380
  (
    n980,
    n185
  );


  buf
  g1381
  (
    n1244,
    n250
  );


  buf
  g1382
  (
    n800,
    n345
  );


  buf
  g1383
  (
    n1587,
    n407
  );


  buf
  g1384
  (
    n976,
    n298
  );


  not
  g1385
  (
    n1121,
    n367
  );


  not
  g1386
  (
    n912,
    n279
  );


  buf
  g1387
  (
    n1356,
    n358
  );


  buf
  g1388
  (
    n1042,
    n213
  );


  buf
  g1389
  (
    n1471,
    n255
  );


  buf
  g1390
  (
    n1185,
    n232
  );


  not
  g1391
  (
    n1154,
    n388
  );


  not
  g1392
  (
    n1676,
    n190
  );


  not
  g1393
  (
    n1683,
    n405
  );


  buf
  g1394
  (
    n1640,
    n408
  );


  buf
  g1395
  (
    n734,
    n411
  );


  not
  g1396
  (
    n1179,
    n393
  );


  not
  g1397
  (
    n1066,
    n373
  );


  buf
  g1398
  (
    n1530,
    n397
  );


  not
  g1399
  (
    n812,
    n347
  );


  buf
  g1400
  (
    n855,
    n249
  );


  buf
  g1401
  (
    n1595,
    n176
  );


  buf
  g1402
  (
    n1674,
    n337
  );


  buf
  g1403
  (
    n865,
    n274
  );


  not
  g1404
  (
    n938,
    n289
  );


  not
  g1405
  (
    n1028,
    n392
  );


  buf
  g1406
  (
    n1466,
    n377
  );


  not
  g1407
  (
    n1191,
    n375
  );


  buf
  g1408
  (
    n1445,
    n306
  );


  not
  g1409
  (
    n771,
    n392
  );


  buf
  g1410
  (
    n1427,
    n277
  );


  buf
  g1411
  (
    n824,
    n280
  );


  not
  g1412
  (
    n1608,
    n206
  );


  not
  g1413
  (
    n922,
    n355
  );


  buf
  g1414
  (
    n1413,
    n288
  );


  not
  g1415
  (
    n1402,
    n249
  );


  not
  g1416
  (
    n1442,
    n174
  );


  buf
  g1417
  (
    n1376,
    n226
  );


  not
  g1418
  (
    n1280,
    n168
  );


  not
  g1419
  (
    n1270,
    n342
  );


  not
  g1420
  (
    n794,
    n230
  );


  not
  g1421
  (
    n940,
    n338
  );


  buf
  g1422
  (
    n739,
    n376
  );


  not
  g1423
  (
    n869,
    n411
  );


  not
  g1424
  (
    n1697,
    n398
  );


  not
  g1425
  (
    n921,
    n351
  );


  not
  g1426
  (
    n1454,
    n216
  );


  buf
  g1427
  (
    n725,
    n389
  );


  buf
  g1428
  (
    n823,
    n312
  );


  not
  g1429
  (
    n1417,
    n330
  );


  buf
  g1430
  (
    n972,
    n413
  );


  not
  g1431
  (
    n1348,
    n239
  );


  buf
  g1432
  (
    n1618,
    n359
  );


  not
  g1433
  (
    n697,
    n235
  );


  buf
  g1434
  (
    n1076,
    n251
  );


  buf
  g1435
  (
    KeyWire_0_49,
    n292
  );


  buf
  g1436
  (
    n979,
    n283
  );


  buf
  g1437
  (
    n783,
    n205
  );


  buf
  g1438
  (
    n714,
    n348
  );


  buf
  g1439
  (
    n988,
    n290
  );


  not
  g1440
  (
    n1276,
    n389
  );


  not
  g1441
  (
    n713,
    n177
  );


  buf
  g1442
  (
    n1460,
    n229
  );


  buf
  g1443
  (
    n814,
    n328
  );


  not
  g1444
  (
    n974,
    n169
  );


  buf
  g1445
  (
    n1243,
    n387
  );


  buf
  g1446
  (
    n1381,
    n272
  );


  buf
  g1447
  (
    n1103,
    n189
  );


  not
  g1448
  (
    n1003,
    n263
  );


  not
  g1449
  (
    n960,
    n233
  );


  buf
  g1450
  (
    n1099,
    n220
  );


  not
  g1451
  (
    n1226,
    n398
  );


  buf
  g1452
  (
    n1231,
    n364
  );


  not
  g1453
  (
    n1559,
    n380
  );


  not
  g1454
  (
    KeyWire_0_7,
    n417
  );


  not
  g1455
  (
    n1404,
    n225
  );


  buf
  g1456
  (
    n1668,
    n349
  );


  not
  g1457
  (
    n902,
    n415
  );


  not
  g1458
  (
    n1513,
    n175
  );


  buf
  g1459
  (
    n904,
    n396
  );


  buf
  g1460
  (
    n875,
    n409
  );


  buf
  g1461
  (
    n1366,
    n370
  );


  buf
  g1462
  (
    n709,
    n304
  );


  not
  g1463
  (
    n1548,
    n175
  );


  not
  g1464
  (
    n1591,
    n284
  );


  not
  g1465
  (
    n1611,
    n181
  );


  not
  g1466
  (
    n1047,
    n196
  );


  buf
  g1467
  (
    n727,
    n199
  );


  buf
  g1468
  (
    n1187,
    n291
  );


  buf
  g1469
  (
    n1541,
    n287
  );


  not
  g1470
  (
    n1567,
    n308
  );


  not
  g1471
  (
    n1132,
    n214
  );


  not
  g1472
  (
    n1252,
    n271
  );


  buf
  g1473
  (
    n1250,
    n327
  );


  buf
  g1474
  (
    n1406,
    n332
  );


  not
  g1475
  (
    n1017,
    n187
  );


  buf
  g1476
  (
    n1165,
    n224
  );


  buf
  g1477
  (
    n779,
    n326
  );


  not
  g1478
  (
    n1293,
    n375
  );


  buf
  g1479
  (
    n998,
    n353
  );


  buf
  g1480
  (
    n1008,
    n185
  );


  not
  g1481
  (
    n1288,
    n231
  );


  not
  g1482
  (
    n1316,
    n296
  );


  buf
  g1483
  (
    n1109,
    n271
  );


  buf
  g1484
  (
    n1485,
    n334
  );


  not
  g1485
  (
    n803,
    n400
  );


  buf
  g1486
  (
    n834,
    n322
  );


  not
  g1487
  (
    n1143,
    n345
  );


  not
  g1488
  (
    n838,
    n365
  );


  buf
  g1489
  (
    n1197,
    n347
  );


  buf
  g1490
  (
    n1218,
    n241
  );


  not
  g1491
  (
    n1192,
    n257
  );


  not
  g1492
  (
    n852,
    n245
  );


  not
  g1493
  (
    n953,
    n409
  );


  buf
  g1494
  (
    n913,
    n302
  );


  buf
  g1495
  (
    n1670,
    n251
  );


  buf
  g1496
  (
    n765,
    n328
  );


  not
  g1497
  (
    n757,
    n366
  );


  buf
  g1498
  (
    n1698,
    n415
  );


  not
  g1499
  (
    n1000,
    n401
  );


  buf
  g1500
  (
    n1600,
    n340
  );


  not
  g1501
  (
    n1695,
    n215
  );


  buf
  g1502
  (
    n1052,
    n291
  );


  buf
  g1503
  (
    n1568,
    n223
  );


  buf
  g1504
  (
    n1465,
    n250
  );


  not
  g1505
  (
    n1375,
    n334
  );


  buf
  g1506
  (
    n1024,
    n179
  );


  not
  g1507
  (
    n745,
    n184
  );


  buf
  g1508
  (
    n1547,
    n248
  );


  buf
  g1509
  (
    n1487,
    n237
  );


  buf
  g1510
  (
    n919,
    n395
  );


  not
  g1511
  (
    n718,
    n216
  );


  buf
  g1512
  (
    n856,
    n261
  );


  buf
  g1513
  (
    n1550,
    n417
  );


  not
  g1514
  (
    n790,
    n166
  );


  buf
  g1515
  (
    n699,
    n219
  );


  not
  g1516
  (
    n778,
    n358
  );


  not
  g1517
  (
    n1665,
    n172
  );


  buf
  g1518
  (
    n1029,
    n222
  );


  buf
  g1519
  (
    n1142,
    n209
  );


  not
  g1520
  (
    n1661,
    n277
  );


  buf
  g1521
  (
    n808,
    n196
  );


  buf
  g1522
  (
    n1267,
    n264
  );


  not
  g1523
  (
    n929,
    n174
  );


  buf
  g1524
  (
    n708,
    n188
  );


  not
  g1525
  (
    n770,
    n297
  );


  not
  g1526
  (
    n850,
    n274
  );


  not
  g1527
  (
    n1065,
    n314
  );


  not
  g1528
  (
    n1246,
    n344
  );


  buf
  g1529
  (
    n1624,
    n369
  );


  not
  g1530
  (
    n1041,
    n266
  );


  buf
  g1531
  (
    n1318,
    n415
  );


  not
  g1532
  (
    n1501,
    n196
  );


  buf
  g1533
  (
    n1457,
    n357
  );


  buf
  g1534
  (
    n1419,
    n177
  );


  buf
  g1535
  (
    n1551,
    n262
  );


  not
  g1536
  (
    n1386,
    n374
  );


  buf
  g1537
  (
    n949,
    n288
  );


  not
  g1538
  (
    n1311,
    n182
  );


  not
  g1539
  (
    n1239,
    n404
  );


  buf
  g1540
  (
    n1152,
    n379
  );


  not
  g1541
  (
    n1225,
    n403
  );


  not
  g1542
  (
    n685,
    n368
  );


  buf
  g1543
  (
    n1294,
    n230
  );


  buf
  g1544
  (
    n1592,
    n248
  );


  buf
  g1545
  (
    n1194,
    n306
  );


  buf
  g1546
  (
    n833,
    n364
  );


  buf
  g1547
  (
    n1351,
    n348
  );


  not
  g1548
  (
    n1633,
    n269
  );


  buf
  g1549
  (
    n1545,
    n224
  );


  buf
  g1550
  (
    n1272,
    n382
  );


  not
  g1551
  (
    n1112,
    n266
  );


  buf
  g1552
  (
    n798,
    n376
  );


  buf
  g1553
  (
    n1673,
    n175
  );


  buf
  g1554
  (
    n801,
    n323
  );


  not
  g1555
  (
    n752,
    n221
  );


  buf
  g1556
  (
    n1161,
    n328
  );


  buf
  g1557
  (
    n1128,
    n334
  );


  buf
  g1558
  (
    n1069,
    n281
  );


  not
  g1559
  (
    n1654,
    n240
  );


  buf
  g1560
  (
    n811,
    n413
  );


  buf
  g1561
  (
    n1312,
    n227
  );


  not
  g1562
  (
    n1346,
    n183
  );


  buf
  g1563
  (
    n933,
    n351
  );


  buf
  g1564
  (
    n1532,
    n318
  );


  buf
  g1565
  (
    n881,
    n165
  );


  not
  g1566
  (
    KeyWire_0_3,
    n197
  );


  not
  g1567
  (
    n1418,
    n262
  );


  not
  g1568
  (
    n1188,
    n299
  );


  not
  g1569
  (
    n1529,
    n333
  );


  not
  g1570
  (
    n1010,
    n378
  );


  buf
  g1571
  (
    n1170,
    n314
  );


  not
  g1572
  (
    n1456,
    n247
  );


  buf
  g1573
  (
    n1322,
    n234
  );


  not
  g1574
  (
    n1301,
    n393
  );


  not
  g1575
  (
    n925,
    n268
  );


  buf
  g1576
  (
    n1448,
    n387
  );


  not
  g1577
  (
    n1075,
    n382
  );


  not
  g1578
  (
    n1613,
    n341
  );


  buf
  g1579
  (
    n1137,
    n365
  );


  not
  g1580
  (
    n1173,
    n264
  );


  buf
  g1581
  (
    KeyWire_0_54,
    n169
  );


  not
  g1582
  (
    n1359,
    n283
  );


  buf
  g1583
  (
    n767,
    n296
  );


  buf
  g1584
  (
    n1088,
    n259
  );


  buf
  g1585
  (
    n712,
    n293
  );


  not
  g1586
  (
    n1426,
    n242
  );


  not
  g1587
  (
    n1593,
    n301
  );


  buf
  g1588
  (
    KeyWire_0_40,
    n185
  );


  not
  g1589
  (
    n969,
    n211
  );


  not
  g1590
  (
    n1667,
    n233
  );


  buf
  g1591
  (
    n1606,
    n260
  );


  buf
  g1592
  (
    n1586,
    n328
  );


  not
  g1593
  (
    n991,
    n182
  );


  not
  g1594
  (
    n1117,
    n166
  );


  not
  g1595
  (
    n1011,
    n344
  );


  not
  g1596
  (
    n1598,
    n346
  );


  buf
  g1597
  (
    n1094,
    n243
  );


  not
  g1598
  (
    n793,
    n402
  );


  buf
  g1599
  (
    n1213,
    n218
  );


  buf
  g1600
  (
    KeyWire_0_36,
    n162
  );


  not
  g1601
  (
    n888,
    n245
  );


  buf
  g1602
  (
    n1577,
    n213
  );


  not
  g1603
  (
    n864,
    n207
  );


  buf
  g1604
  (
    n810,
    n240
  );


  not
  g1605
  (
    n845,
    n355
  );


  buf
  g1606
  (
    n908,
    n336
  );


  not
  g1607
  (
    n1009,
    n403
  );


  buf
  g1608
  (
    n695,
    n321
  );


  not
  g1609
  (
    n895,
    n294
  );


  not
  g1610
  (
    n1361,
    n402
  );


  buf
  g1611
  (
    n1265,
    n190
  );


  buf
  g1612
  (
    n917,
    n255
  );


  not
  g1613
  (
    n1013,
    n176
  );


  buf
  g1614
  (
    n1578,
    n367
  );


  buf
  g1615
  (
    n1560,
    n190
  );


  not
  g1616
  (
    n1612,
    n165
  );


  not
  g1617
  (
    n1284,
    n379
  );


  not
  g1618
  (
    n1682,
    n221
  );


  not
  g1619
  (
    n1519,
    n180
  );


  buf
  g1620
  (
    n1554,
    n317
  );


  buf
  g1621
  (
    KeyWire_0_12,
    n309
  );


  not
  g1622
  (
    n1056,
    n296
  );


  buf
  g1623
  (
    n822,
    n357
  );


  not
  g1624
  (
    n700,
    n275
  );


  buf
  g1625
  (
    n1061,
    n183
  );


  not
  g1626
  (
    n1235,
    n259
  );


  not
  g1627
  (
    n1552,
    n184
  );


  buf
  g1628
  (
    KeyWire_0_25,
    n371
  );


  not
  g1629
  (
    n1020,
    n212
  );


  not
  g1630
  (
    n1223,
    n222
  );


  not
  g1631
  (
    n735,
    n383
  );


  not
  g1632
  (
    n1403,
    n202
  );


  buf
  g1633
  (
    n1241,
    n384
  );


  buf
  g1634
  (
    n1036,
    n307
  );


  not
  g1635
  (
    n696,
    n419
  );


  buf
  g1636
  (
    n1669,
    n322
  );


  buf
  g1637
  (
    n1090,
    n345
  );


  buf
  g1638
  (
    n1162,
    n307
  );


  not
  g1639
  (
    n1659,
    n314
  );


  buf
  g1640
  (
    n1678,
    n396
  );


  not
  g1641
  (
    n1341,
    n275
  );


  buf
  g1642
  (
    n873,
    n398
  );


  buf
  g1643
  (
    n1098,
    n409
  );


  buf
  g1644
  (
    n1561,
    n365
  );


  buf
  g1645
  (
    n1476,
    n332
  );


  buf
  g1646
  (
    n1401,
    n191
  );


  not
  g1647
  (
    n828,
    n326
  );


  not
  g1648
  (
    n1133,
    n260
  );


  not
  g1649
  (
    n1407,
    n394
  );


  buf
  g1650
  (
    n1496,
    n356
  );


  not
  g1651
  (
    n1330,
    n203
  );


  buf
  g1652
  (
    n729,
    n310
  );


  buf
  g1653
  (
    n1627,
    n346
  );


  not
  g1654
  (
    n878,
    n342
  );


  not
  g1655
  (
    n1648,
    n382
  );


  buf
  g1656
  (
    n742,
    n193
  );


  buf
  g1657
  (
    n1632,
    n360
  );


  buf
  g1658
  (
    n1434,
    n257
  );


  not
  g1659
  (
    n871,
    n340
  );


  buf
  g1660
  (
    n1431,
    n291
  );


  not
  g1661
  (
    n1155,
    n295
  );


  not
  g1662
  (
    n858,
    n266
  );


  buf
  g1663
  (
    n1168,
    n276
  );


  not
  g1664
  (
    n1091,
    n356
  );


  not
  g1665
  (
    n674,
    n234
  );


  not
  g1666
  (
    n1089,
    n194
  );


  not
  g1667
  (
    n1722,
    n692
  );


  buf
  g1668
  (
    n1702,
    n696
  );


  buf
  g1669
  (
    n1725,
    n697
  );


  buf
  g1670
  (
    n1711,
    n680
  );


  not
  g1671
  (
    n1700,
    n679
  );


  not
  g1672
  (
    n1706,
    n682
  );


  not
  g1673
  (
    n1717,
    n677
  );


  buf
  g1674
  (
    n1715,
    n700
  );


  not
  g1675
  (
    n1708,
    n698
  );


  buf
  g1676
  (
    n1707,
    n691
  );


  buf
  g1677
  (
    n1723,
    n685
  );


  buf
  g1678
  (
    n1710,
    n688
  );


  not
  g1679
  (
    n1718,
    n694
  );


  buf
  g1680
  (
    n1726,
    n699
  );


  not
  g1681
  (
    n1701,
    n687
  );


  not
  g1682
  (
    n1724,
    n675
  );


  buf
  g1683
  (
    n1716,
    n681
  );


  not
  g1684
  (
    n1721,
    n690
  );


  buf
  g1685
  (
    n1703,
    n695
  );


  not
  g1686
  (
    n1719,
    n673
  );


  buf
  g1687
  (
    n1714,
    n689
  );


  buf
  g1688
  (
    n1720,
    n674
  );


  buf
  g1689
  (
    n1705,
    n678
  );


  buf
  g1690
  (
    n1727,
    n686
  );


  buf
  g1691
  (
    n1712,
    n683
  );


  buf
  g1692
  (
    n1709,
    n676
  );


  buf
  g1693
  (
    n1713,
    n693
  );


  not
  g1694
  (
    n1704,
    n684
  );


  nand
  g1695
  (
    n1732,
    n722,
    n720,
    n705,
    n1700
  );


  xor
  g1696
  (
    n1731,
    n1708,
    n1703,
    n1704,
    n1705
  );


  nor
  g1697
  (
    n1728,
    n715,
    n718,
    n701,
    n723
  );


  xnor
  g1698
  (
    n1734,
    n703,
    n710,
    n708,
    n1707
  );


  or
  g1699
  (
    n1730,
    n702,
    n711,
    n704,
    n727
  );


  xnor
  g1700
  (
    n1729,
    n714,
    n707,
    n709,
    n725
  );


  xnor
  g1701
  (
    n1736,
    n712,
    n1702,
    n716,
    n726
  );


  nor
  g1702
  (
    n1735,
    n706,
    n713,
    n1701,
    n724
  );


  or
  g1703
  (
    n1733,
    n719,
    n717,
    n1706,
    n721
  );


  xor
  g1704
  (
    n1738,
    n735,
    n748,
    n1735,
    n753
  );


  nand
  g1705
  (
    n1743,
    n739,
    n749,
    n747,
    n1734
  );


  nor
  g1706
  (
    n1737,
    n741,
    n740,
    n751,
    n737
  );


  xor
  g1707
  (
    n1739,
    n750,
    n1733,
    n729,
    n730
  );


  nor
  g1708
  (
    n1741,
    n744,
    n754,
    n743,
    n752
  );


  and
  g1709
  (
    n1740,
    n742,
    n1730,
    n1729,
    n733
  );


  nand
  g1710
  (
    n1745,
    n1728,
    n738,
    n1732,
    n1731
  );


  xor
  g1711
  (
    n1744,
    n728,
    n732,
    n745,
    n731
  );


  xnor
  g1712
  (
    n1742,
    n734,
    n736,
    n746,
    n1736
  );


  nor
  g1713
  (
    n1751,
    n755,
    n1742,
    n1745,
    n1740
  );


  nand
  g1714
  (
    n1749,
    n1716,
    n1743,
    n1714,
    n763
  );


  nor
  g1715
  (
    n1748,
    n762,
    n1714,
    n1710,
    n1744
  );


  nor
  g1716
  (
    n1755,
    n765,
    n1713,
    n1737,
    n1745
  );


  nand
  g1717
  (
    n1750,
    n757,
    n1718,
    n1709,
    n1710
  );


  xor
  g1718
  (
    n1754,
    n1738,
    n1711,
    n756
  );


  xnor
  g1719
  (
    n1752,
    n1718,
    n1739,
    n1717,
    n1712
  );


  or
  g1720
  (
    n1747,
    n1712,
    n758,
    n1713,
    n761
  );


  nand
  g1721
  (
    n1753,
    n1717,
    n764,
    n1741,
    n1715
  );


  or
  g1722
  (
    n1746,
    n760,
    n759,
    n1716,
    n1715
  );


  xor
  g1723
  (
    n1759,
    n766,
    n1746
  );


  xnor
  g1724
  (
    n1764,
    n768,
    n1748
  );


  xnor
  g1725
  (
    n1758,
    n1725,
    n1721,
    n1724,
    n769
  );


  nor
  g1726
  (
    n1756,
    n1721,
    n770,
    n1719,
    n1722
  );


  or
  g1727
  (
    n1762,
    n774,
    n1723,
    n1726
  );


  xnor
  g1728
  (
    n1760,
    n1754,
    n1719,
    n772,
    n1750
  );


  and
  g1729
  (
    n1765,
    n1720,
    n1726,
    n1753,
    n1725
  );


  and
  g1730
  (
    n1761,
    n767,
    n1720,
    n1727,
    n773
  );


  or
  g1731
  (
    n1757,
    n1751,
    n1747,
    n1722,
    n771
  );


  xor
  g1732
  (
    n1763,
    n1755,
    n1749,
    n1724,
    n1752
  );


  not
  g1733
  (
    n1774,
    n1765
  );


  buf
  g1734
  (
    n1777,
    n1758
  );


  not
  g1735
  (
    n1784,
    n1764
  );


  buf
  g1736
  (
    n1768,
    n1764
  );


  buf
  g1737
  (
    n1782,
    n1763
  );


  buf
  g1738
  (
    n1776,
    n1756
  );


  buf
  g1739
  (
    n1770,
    n1765
  );


  not
  g1740
  (
    n1767,
    n1765
  );


  not
  g1741
  (
    n1771,
    n1756
  );


  buf
  g1742
  (
    n1772,
    n1758
  );


  not
  g1743
  (
    n1785,
    n1762
  );


  not
  g1744
  (
    n1788,
    n775
  );


  buf
  g1745
  (
    n1786,
    n1759
  );


  buf
  g1746
  (
    n1780,
    n1759
  );


  buf
  g1747
  (
    n1775,
    n1760
  );


  buf
  g1748
  (
    n1783,
    n1765
  );


  buf
  g1749
  (
    n1787,
    n1761
  );


  buf
  g1750
  (
    n1766,
    n1763
  );


  buf
  g1751
  (
    n1779,
    n1762
  );


  not
  g1752
  (
    n1789,
    n1757
  );


  buf
  g1753
  (
    n1781,
    n1761
  );


  not
  g1754
  (
    n1773,
    n1757
  );


  not
  g1755
  (
    n1769,
    n1764
  );


  or
  g1756
  (
    n1778,
    n1760,
    n1764
  );


  not
  g1757
  (
    n1790,
    n1769
  );


  buf
  g1758
  (
    n1793,
    n1768
  );


  not
  g1759
  (
    n1798,
    n1772
  );


  buf
  g1760
  (
    n1796,
    n776
  );


  and
  g1761
  (
    n1794,
    n779,
    n1774
  );


  and
  g1762
  (
    n1792,
    n781,
    n782,
    n1774,
    n1767
  );


  and
  g1763
  (
    n1795,
    n1773,
    n1770,
    n1766,
    n1771
  );


  xnor
  g1764
  (
    n1799,
    n1766,
    n1767,
    n1770,
    n1775
  );


  or
  g1765
  (
    n1797,
    n1773,
    n780,
    n1771,
    n1769
  );


  xnor
  g1766
  (
    n1791,
    n1768,
    n778,
    n777,
    n1772
  );


  not
  g1767
  (
    n1805,
    n794
  );


  buf
  g1768
  (
    n1802,
    n1792
  );


  not
  g1769
  (
    n1809,
    n789
  );


  buf
  g1770
  (
    n1807,
    n785
  );


  not
  g1771
  (
    n1803,
    n791
  );


  buf
  g1772
  (
    n1806,
    n786
  );


  or
  g1773
  (
    n1800,
    n1796,
    n1791,
    n784
  );


  xor
  g1774
  (
    n1801,
    n1799,
    n1790,
    n790,
    n788
  );


  nor
  g1775
  (
    n1810,
    n793,
    n1799,
    n787,
    n1795
  );


  nand
  g1776
  (
    n1808,
    n1797,
    n792,
    n783,
    n1798
  );


  xor
  g1777
  (
    n1804,
    n795,
    n1793,
    n1775,
    n1794
  );


  nand
  g1778
  (
    n1812,
    n1802,
    n1778,
    n1776,
    n1784
  );


  xnor
  g1779
  (
    n1817,
    n1777,
    n1781,
    n1801,
    n1782
  );


  xnor
  g1780
  (
    n1815,
    n1785,
    n1779,
    n1807,
    n1800
  );


  nand
  g1781
  (
    n1818,
    n1783,
    n1779,
    n1781,
    n1805
  );


  nand
  g1782
  (
    n1813,
    n1777,
    n1787,
    n1780,
    n1776
  );


  xor
  g1783
  (
    n1816,
    n1785,
    n1783,
    n1804,
    n1803
  );


  xnor
  g1784
  (
    n1814,
    n1784,
    n1780,
    n1808,
    n1782
  );


  or
  g1785
  (
    n1811,
    n1806,
    n1786,
    n1778
  );


  not
  g1786
  (
    n1824,
    n1816
  );


  buf
  g1787
  (
    n1819,
    n796
  );


  buf
  g1788
  (
    n1820,
    n1815
  );


  buf
  g1789
  (
    n1823,
    n1814
  );


  and
  g1790
  (
    n1822,
    n1788,
    n1788,
    n1787,
    n797
  );


  nand
  g1791
  (
    n1821,
    n798,
    n1817,
    n1813,
    n1812
  );


  xnor
  g1792
  (
    n1827,
    n1820,
    n1824,
    n800,
    n1818
  );


  xor
  g1793
  (
    n1826,
    n1823,
    n1821,
    n1822,
    n1789
  );


  nor
  g1794
  (
    n1825,
    n1819,
    n799,
    n1809,
    n1789
  );


  not
  g1795
  (
    n1829,
    n1825
  );


  buf
  g1796
  (
    n1828,
    n1826
  );


  buf
  g1797
  (
    n1830,
    n1828
  );


  buf
  g1798
  (
    n1831,
    n1830
  );


  not
  g1799
  (
    n1832,
    n1830
  );


  and
  g1800
  (
    n1833,
    n1832,
    n1829
  );


  not
  g1801
  (
    n1835,
    n1833
  );


  not
  g1802
  (
    n1834,
    n1833
  );


  buf
  g1803
  (
    n1836,
    n1835
  );


  not
  g1804
  (
    n1837,
    n1834
  );


  not
  g1805
  (
    n1844,
    n1836
  );


  buf
  g1806
  (
    n1842,
    n1837
  );


  buf
  g1807
  (
    n1838,
    n1836
  );


  buf
  g1808
  (
    n1843,
    n1836
  );


  buf
  g1809
  (
    n1845,
    n1837
  );


  not
  g1810
  (
    n1841,
    n1837
  );


  not
  g1811
  (
    n1839,
    n1836
  );


  buf
  g1812
  (
    n1840,
    n1837
  );


  not
  g1813
  (
    n1846,
    n1838
  );


  buf
  g1814
  (
    n1847,
    n1838
  );


  buf
  g1815
  (
    n1850,
    n1846
  );


  not
  g1816
  (
    n1849,
    n1846
  );


  buf
  g1817
  (
    n1848,
    n1847
  );


  not
  g1818
  (
    n1851,
    n1847
  );


  not
  g1819
  (
    n1852,
    n1848
  );


  buf
  g1820
  (
    n1853,
    n1848
  );


  buf
  g1821
  (
    n1855,
    n1853
  );


  not
  g1822
  (
    n1854,
    n1853
  );


  buf
  g1823
  (
    n1857,
    n1852
  );


  buf
  g1824
  (
    n1856,
    n1853
  );


  xor
  g1825
  (
    n1858,
    n1850,
    n1849,
    n1854
  );


  and
  g1826
  (
    n1859,
    n801,
    n1849,
    n1854
  );


  buf
  g1827
  (
    n1860,
    n1859
  );


  buf
  g1828
  (
    n1863,
    n1860
  );


  buf
  g1829
  (
    n1862,
    n1855
  );


  xor
  g1830
  (
    n1861,
    n1856,
    n1856,
    n1855,
    n1860
  );


  and
  g1831
  (
    n1864,
    n1853,
    n1857,
    n1860
  );


  buf
  g1832
  (
    n1869,
    n1861
  );


  not
  g1833
  (
    n1867,
    n1861
  );


  not
  g1834
  (
    n1865,
    n1862
  );


  not
  g1835
  (
    n1868,
    n1862
  );


  buf
  g1836
  (
    n1866,
    n1862
  );


  nor
  g1837
  (
    n1871,
    n1864,
    n1865,
    n1868
  );


  and
  g1838
  (
    n1875,
    n1866,
    n1867
  );


  nand
  g1839
  (
    n1877,
    n1847,
    n1868,
    n1863
  );


  nor
  g1840
  (
    n1874,
    n1850,
    n1863,
    n803
  );


  nand
  g1841
  (
    n1870,
    n1850,
    n1839,
    n1863,
    n1857
  );


  and
  g1842
  (
    n1876,
    n1866,
    n1865,
    n1839,
    n1847
  );


  xnor
  g1843
  (
    n1873,
    n1865,
    n1866
  );


  nand
  g1844
  (
    n1872,
    n802,
    n1864,
    n1862,
    n1867
  );


  not
  g1845
  (
    n1878,
    n1877
  );


  buf
  g1846
  (
    n1879,
    n1878
  );


  not
  g1847
  (
    n1880,
    n1878
  );


  xnor
  g1848
  (
    n1881,
    n1851,
    n1880
  );


  and
  g1849
  (
    n1885,
    n1864,
    n1880
  );


  xnor
  g1850
  (
    n1882,
    n1851,
    n1810
  );


  nor
  g1851
  (
    n1884,
    n1869,
    n1864
  );


  and
  g1852
  (
    n1883,
    n1851,
    n1869
  );


  and
  g1853
  (
    n1887,
    n1880,
    n1879,
    n1857
  );


  xnor
  g1854
  (
    n1888,
    n1850,
    n1880,
    n1879
  );


  xor
  g1855
  (
    n1886,
    n1851,
    n1869,
    n1789
  );


  nand
  g1856
  (
    n1889,
    n1882,
    n1881
  );


  not
  g1857
  (
    n1890,
    n1889
  );


  buf
  g1858
  (
    n1892,
    n1890
  );


  buf
  g1859
  (
    n1891,
    n1890
  );


  and
  g1860
  (
    n1893,
    n1727,
    n1886
  );


  and
  g1861
  (
    KeyWire_0_5,
    n1886,
    n1892
  );


  nand
  g1862
  (
    n1896,
    n1891,
    n1884
  );


  nand
  g1863
  (
    n1900,
    n1840,
    n1891
  );


  xnor
  g1864
  (
    n1894,
    n1883,
    n1892
  );


  and
  g1865
  (
    n1895,
    n1892,
    n1887,
    n1827
  );


  or
  g1866
  (
    n1898,
    n1885,
    n1885,
    n1892,
    n1884
  );


  xnor
  g1867
  (
    n1899,
    n1887,
    n1891,
    n1883
  );


  not
  g1868
  (
    n1908,
    n1895
  );


  buf
  g1869
  (
    n1929,
    n1888
  );


  not
  g1870
  (
    n1923,
    n1893
  );


  not
  g1871
  (
    n1902,
    n1899
  );


  buf
  g1872
  (
    n1932,
    n1843
  );


  not
  g1873
  (
    n1930,
    n1893
  );


  not
  g1874
  (
    n1924,
    n1894
  );


  buf
  g1875
  (
    n1926,
    n1842
  );


  not
  g1876
  (
    n1925,
    n1842
  );


  not
  g1877
  (
    n1917,
    n1899
  );


  not
  g1878
  (
    n1904,
    n1895
  );


  not
  g1879
  (
    n1918,
    n1900
  );


  not
  g1880
  (
    n1931,
    n1896
  );


  not
  g1881
  (
    n1916,
    n1896
  );


  buf
  g1882
  (
    n1913,
    n1900
  );


  buf
  g1883
  (
    n1906,
    n1893
  );


  buf
  g1884
  (
    n1914,
    n1895
  );


  buf
  g1885
  (
    n1911,
    n1842
  );


  not
  g1886
  (
    n1909,
    n1898
  );


  not
  g1887
  (
    n1907,
    n1898
  );


  buf
  g1888
  (
    n1912,
    n1840
  );


  not
  g1889
  (
    n1922,
    n1898
  );


  not
  g1890
  (
    n1903,
    n1843
  );


  buf
  g1891
  (
    n1919,
    n1899
  );


  not
  g1892
  (
    n1910,
    n1890
  );


  buf
  g1893
  (
    n1928,
    n1899
  );


  not
  g1894
  (
    n1920,
    n1841
  );


  not
  g1895
  (
    n1915,
    n1900
  );


  nand
  g1896
  (
    n1901,
    n1895,
    n1896,
    n1888
  );


  nor
  g1897
  (
    n1921,
    n1841,
    n1893,
    n1900,
    n1890
  );


  and
  g1898
  (
    n1927,
    n1894,
    n1897
  );


  and
  g1899
  (
    n1905,
    n1894,
    n1897,
    n1898
  );


  buf
  g1900
  (
    n1994,
    n1917
  );


  not
  g1901
  (
    n2017,
    n1906
  );


  not
  g1902
  (
    n1959,
    n1926
  );


  buf
  g1903
  (
    n1958,
    n1920
  );


  buf
  g1904
  (
    n1966,
    n1924
  );


  not
  g1905
  (
    n1940,
    n1927
  );


  buf
  g1906
  (
    n1984,
    n1912
  );


  buf
  g1907
  (
    n1950,
    n1923
  );


  buf
  g1908
  (
    n2008,
    n1906
  );


  not
  g1909
  (
    n1991,
    n1916
  );


  buf
  g1910
  (
    n1953,
    n1906
  );


  buf
  g1911
  (
    n2023,
    n1922
  );


  not
  g1912
  (
    n2038,
    n1931
  );


  not
  g1913
  (
    n1947,
    n1914
  );


  buf
  g1914
  (
    n2016,
    n1921
  );


  not
  g1915
  (
    n1937,
    n1932
  );


  buf
  g1916
  (
    n2033,
    n1919
  );


  not
  g1917
  (
    KeyWire_0_27,
    n1912
  );


  not
  g1918
  (
    n1964,
    n1918
  );


  not
  g1919
  (
    n2001,
    n1911
  );


  buf
  g1920
  (
    n2041,
    n1905
  );


  not
  g1921
  (
    n2056,
    n1905
  );


  buf
  g1922
  (
    n1939,
    n1909
  );


  buf
  g1923
  (
    n1946,
    n1918
  );


  buf
  g1924
  (
    n2011,
    n1911
  );


  buf
  g1925
  (
    n1981,
    n1922
  );


  not
  g1926
  (
    n1979,
    n1908
  );


  not
  g1927
  (
    n2000,
    n1907
  );


  buf
  g1928
  (
    n2044,
    n1909
  );


  not
  g1929
  (
    n2021,
    n1910
  );


  buf
  g1930
  (
    n1955,
    n1921
  );


  buf
  g1931
  (
    n1935,
    n1924
  );


  buf
  g1932
  (
    n2019,
    n1912
  );


  buf
  g1933
  (
    n1962,
    n1906
  );


  buf
  g1934
  (
    n1978,
    n1911
  );


  not
  g1935
  (
    n2010,
    n1925
  );


  not
  g1936
  (
    n1993,
    n1917
  );


  not
  g1937
  (
    n1965,
    n1923
  );


  not
  g1938
  (
    n1956,
    n1925
  );


  not
  g1939
  (
    n1995,
    n1927
  );


  buf
  g1940
  (
    n1948,
    n1916
  );


  not
  g1941
  (
    n2050,
    n1903
  );


  buf
  g1942
  (
    n2025,
    n1920
  );


  buf
  g1943
  (
    n1992,
    n1926
  );


  buf
  g1944
  (
    n1996,
    n1924
  );


  buf
  g1945
  (
    n2032,
    n1912
  );


  not
  g1946
  (
    n2018,
    n1917
  );


  not
  g1947
  (
    n1943,
    n1913
  );


  buf
  g1948
  (
    n2049,
    n1911
  );


  not
  g1949
  (
    n2035,
    n1922
  );


  buf
  g1950
  (
    n2043,
    n1913
  );


  buf
  g1951
  (
    n2048,
    n1910
  );


  not
  g1952
  (
    n1949,
    n1901
  );


  not
  g1953
  (
    n2036,
    n1928
  );


  buf
  g1954
  (
    n2022,
    n1932
  );


  buf
  g1955
  (
    n2060,
    n1909
  );


  not
  g1956
  (
    n2042,
    n1843
  );


  not
  g1957
  (
    n2058,
    n1927
  );


  buf
  g1958
  (
    KeyWire_0_35,
    n1908
  );


  buf
  g1959
  (
    n1988,
    n1925
  );


  buf
  g1960
  (
    n2045,
    n1930
  );


  not
  g1961
  (
    n2047,
    n1921
  );


  buf
  g1962
  (
    n1967,
    n1905
  );


  buf
  g1963
  (
    n2002,
    n1901
  );


  buf
  g1964
  (
    n1933,
    n1922
  );


  not
  g1965
  (
    n2007,
    n1931
  );


  buf
  g1966
  (
    n2029,
    n1915
  );


  not
  g1967
  (
    n2028,
    n1929
  );


  not
  g1968
  (
    n1942,
    n1909
  );


  not
  g1969
  (
    n2057,
    n1920
  );


  buf
  g1970
  (
    n2006,
    n1914
  );


  buf
  g1971
  (
    n1980,
    n1904
  );


  buf
  g1972
  (
    n2055,
    n1903
  );


  buf
  g1973
  (
    n2009,
    n1930
  );


  not
  g1974
  (
    n2059,
    n1916
  );


  buf
  g1975
  (
    n1974,
    n1907
  );


  buf
  g1976
  (
    n1998,
    n1910
  );


  not
  g1977
  (
    n2024,
    n1905
  );


  buf
  g1978
  (
    n2039,
    n1928
  );


  buf
  g1979
  (
    n1945,
    n1928
  );


  not
  g1980
  (
    n2014,
    n1903
  );


  not
  g1981
  (
    n2027,
    n1904
  );


  not
  g1982
  (
    n2012,
    n1914
  );


  buf
  g1983
  (
    n1936,
    n1916
  );


  not
  g1984
  (
    n2003,
    n1901
  );


  not
  g1985
  (
    n2034,
    n1923
  );


  buf
  g1986
  (
    n1944,
    n1928
  );


  buf
  g1987
  (
    n1982,
    n1924
  );


  not
  g1988
  (
    n1951,
    n1915
  );


  not
  g1989
  (
    n1983,
    n1921
  );


  buf
  g1990
  (
    n1986,
    n1930
  );


  not
  g1991
  (
    n2015,
    n1926
  );


  buf
  g1992
  (
    n1985,
    n1914
  );


  not
  g1993
  (
    n2005,
    n1904
  );


  not
  g1994
  (
    n1990,
    n1908
  );


  buf
  g1995
  (
    n2053,
    n1915
  );


  not
  g1996
  (
    n2004,
    n1918
  );


  not
  g1997
  (
    n1941,
    n1919
  );


  not
  g1998
  (
    n2026,
    n1932
  );


  not
  g1999
  (
    n1963,
    n1931
  );


  buf
  g2000
  (
    n2040,
    n1925
  );


  not
  g2001
  (
    n1999,
    n1917
  );


  not
  g2002
  (
    n2052,
    n1903
  );


  not
  g2003
  (
    n1961,
    n1918
  );


  buf
  g2004
  (
    n1971,
    n1920
  );


  not
  g2005
  (
    n2051,
    n1908
  );


  buf
  g2006
  (
    n1938,
    n1930
  );


  not
  g2007
  (
    n1934,
    n1932
  );


  not
  g2008
  (
    n1989,
    n1902
  );


  not
  g2009
  (
    n2030,
    n1931
  );


  not
  g2010
  (
    n2020,
    n1913
  );


  buf
  g2011
  (
    n1968,
    n1923
  );


  not
  g2012
  (
    n1975,
    n1910
  );


  not
  g2013
  (
    n1952,
    n1915
  );


  buf
  g2014
  (
    n1969,
    n1919
  );


  not
  g2015
  (
    KeyWire_0_59,
    n1929
  );


  buf
  g2016
  (
    n1987,
    n1902
  );


  not
  g2017
  (
    n2031,
    n1902
  );


  not
  g2018
  (
    n1970,
    n1904
  );


  buf
  g2019
  (
    n1972,
    n1929
  );


  not
  g2020
  (
    KeyWire_0_33,
    n1913
  );


  not
  g2021
  (
    n2037,
    n1929
  );


  not
  g2022
  (
    n1997,
    n1927
  );


  not
  g2023
  (
    n2046,
    n1901
  );


  buf
  g2024
  (
    n1960,
    n1907
  );


  not
  g2025
  (
    n1954,
    n1907
  );


  buf
  g2026
  (
    n1977,
    n1919
  );


  xnor
  g2027
  (
    n1976,
    n1902,
    n1926
  );


  not
  g2028
  (
    n2061,
    n2032
  );


  buf
  g2029
  (
    n2410,
    n588
  );


  not
  g2030
  (
    n2362,
    n436
  );


  buf
  g2031
  (
    n2213,
    n509
  );


  not
  g2032
  (
    n2569,
    n2030
  );


  not
  g2033
  (
    n2090,
    n660
  );


  buf
  g2034
  (
    n2337,
    n1998
  );


  buf
  g2035
  (
    n2561,
    n647
  );


  not
  g2036
  (
    n2212,
    n555
  );


  not
  g2037
  (
    n2448,
    n2032
  );


  not
  g2038
  (
    n2388,
    n470
  );


  buf
  g2039
  (
    n2524,
    n550
  );


  not
  g2040
  (
    n2485,
    n428
  );


  buf
  g2041
  (
    n2472,
    n598
  );


  buf
  g2042
  (
    n2255,
    n529
  );


  not
  g2043
  (
    n2404,
    n454
  );


  not
  g2044
  (
    n2505,
    n1990
  );


  buf
  g2045
  (
    n2133,
    n512
  );


  buf
  g2046
  (
    n2370,
    n1940
  );


  buf
  g2047
  (
    n2308,
    n550
  );


  buf
  g2048
  (
    n2446,
    n617
  );


  not
  g2049
  (
    n2180,
    n2020
  );


  buf
  g2050
  (
    n2250,
    n557
  );


  not
  g2051
  (
    n2269,
    n552
  );


  not
  g2052
  (
    n2164,
    n1945
  );


  not
  g2053
  (
    n2307,
    n2055
  );


  buf
  g2054
  (
    n2390,
    n514
  );


  not
  g2055
  (
    n2491,
    n485
  );


  not
  g2056
  (
    n2270,
    n626
  );


  not
  g2057
  (
    n2525,
    n2040
  );


  not
  g2058
  (
    n2199,
    n2014
  );


  not
  g2059
  (
    n2365,
    n548
  );


  buf
  g2060
  (
    n2267,
    n623
  );


  buf
  g2061
  (
    n2293,
    n2023
  );


  not
  g2062
  (
    n2193,
    n1978
  );


  buf
  g2063
  (
    n2175,
    n1844
  );


  buf
  g2064
  (
    n2568,
    n2056
  );


  not
  g2065
  (
    n2427,
    n1971
  );


  not
  g2066
  (
    n2473,
    n641
  );


  buf
  g2067
  (
    n2477,
    n2008
  );


  not
  g2068
  (
    n2204,
    n2036
  );


  not
  g2069
  (
    n2351,
    n2042
  );


  not
  g2070
  (
    n2431,
    n2028
  );


  buf
  g2071
  (
    n2219,
    n619
  );


  buf
  g2072
  (
    n2095,
    n573
  );


  buf
  g2073
  (
    n2252,
    n1948
  );


  not
  g2074
  (
    n2274,
    n629
  );


  buf
  g2075
  (
    n2126,
    n427
  );


  buf
  g2076
  (
    n2342,
    n671
  );


  not
  g2077
  (
    n2552,
    n566
  );


  not
  g2078
  (
    n2153,
    n589
  );


  buf
  g2079
  (
    n2397,
    n524
  );


  not
  g2080
  (
    n2504,
    n464
  );


  buf
  g2081
  (
    n2438,
    n1988
  );


  buf
  g2082
  (
    n2484,
    n659
  );


  buf
  g2083
  (
    n2369,
    n516
  );


  not
  g2084
  (
    n2110,
    n557
  );


  not
  g2085
  (
    n2523,
    n1964
  );


  buf
  g2086
  (
    n2348,
    n633
  );


  buf
  g2087
  (
    n2242,
    n2053
  );


  buf
  g2088
  (
    n2558,
    n486
  );


  buf
  g2089
  (
    n2393,
    n606
  );


  buf
  g2090
  (
    n2177,
    n638
  );


  not
  g2091
  (
    n2236,
    n483
  );


  not
  g2092
  (
    n2124,
    n1987
  );


  not
  g2093
  (
    n2194,
    n1997
  );


  not
  g2094
  (
    n2435,
    n1957
  );


  not
  g2095
  (
    n2486,
    n1990
  );


  not
  g2096
  (
    n2453,
    n1981
  );


  not
  g2097
  (
    n2184,
    n1986
  );


  not
  g2098
  (
    n2380,
    n466
  );


  not
  g2099
  (
    n2157,
    n1959
  );


  not
  g2100
  (
    n2066,
    n580
  );


  buf
  g2101
  (
    n2544,
    n2018
  );


  buf
  g2102
  (
    KeyWire_0_4,
    n445
  );


  buf
  g2103
  (
    n2235,
    n600
  );


  not
  g2104
  (
    n2521,
    n453
  );


  not
  g2105
  (
    n2187,
    n636
  );


  not
  g2106
  (
    n2230,
    n636
  );


  not
  g2107
  (
    n2560,
    n558
  );


  buf
  g2108
  (
    n2254,
    n523
  );


  not
  g2109
  (
    n2289,
    n1980
  );


  not
  g2110
  (
    n2433,
    n568
  );


  not
  g2111
  (
    n2275,
    n631
  );


  buf
  g2112
  (
    n2502,
    n452
  );


  buf
  g2113
  (
    n2172,
    n2059
  );


  buf
  g2114
  (
    n2559,
    n663
  );


  not
  g2115
  (
    n2530,
    n485
  );


  not
  g2116
  (
    n2081,
    n2045
  );


  not
  g2117
  (
    n2413,
    n463
  );


  buf
  g2118
  (
    n2454,
    n2017
  );


  buf
  g2119
  (
    n2548,
    n1981
  );


  buf
  g2120
  (
    n2398,
    n442
  );


  buf
  g2121
  (
    n2449,
    n569
  );


  buf
  g2122
  (
    n2459,
    n1994
  );


  buf
  g2123
  (
    n2387,
    n1936
  );


  not
  g2124
  (
    n2517,
    n422
  );


  not
  g2125
  (
    n2541,
    n507
  );


  not
  g2126
  (
    n2445,
    n652
  );


  not
  g2127
  (
    n2266,
    n1941
  );


  buf
  g2128
  (
    n2518,
    n473
  );


  not
  g2129
  (
    n2374,
    n585
  );


  buf
  g2130
  (
    n2241,
    n668
  );


  buf
  g2131
  (
    n2245,
    n426
  );


  buf
  g2132
  (
    n2354,
    n448
  );


  buf
  g2133
  (
    n2174,
    n535
  );


  not
  g2134
  (
    n2511,
    n1944
  );


  not
  g2135
  (
    n2371,
    n584
  );


  buf
  g2136
  (
    n2494,
    n492
  );


  buf
  g2137
  (
    n2476,
    n645
  );


  not
  g2138
  (
    n2443,
    n539
  );


  not
  g2139
  (
    n2196,
    n577
  );


  buf
  g2140
  (
    n2392,
    n624
  );


  buf
  g2141
  (
    n2149,
    n611
  );


  buf
  g2142
  (
    n2528,
    n535
  );


  not
  g2143
  (
    n2161,
    n550
  );


  buf
  g2144
  (
    KeyWire_0_52,
    n588
  );


  buf
  g2145
  (
    KeyWire_0_58,
    n2013
  );


  buf
  g2146
  (
    n2515,
    n1988
  );


  buf
  g2147
  (
    n2223,
    n2055
  );


  not
  g2148
  (
    n2304,
    n497
  );


  buf
  g2149
  (
    n2253,
    n522
  );


  not
  g2150
  (
    n2455,
    n536
  );


  not
  g2151
  (
    n2132,
    n1989
  );


  buf
  g2152
  (
    n2144,
    n1959
  );


  not
  g2153
  (
    n2221,
    n478
  );


  buf
  g2154
  (
    n2423,
    n646
  );


  buf
  g2155
  (
    n2323,
    n544
  );


  not
  g2156
  (
    n2186,
    n2004
  );


  not
  g2157
  (
    KeyWire_0_55,
    n504
  );


  not
  g2158
  (
    n2279,
    n1954
  );


  buf
  g2159
  (
    n2137,
    n454
  );


  buf
  g2160
  (
    n2556,
    n2021
  );


  buf
  g2161
  (
    n2408,
    n565
  );


  not
  g2162
  (
    n2539,
    n1975
  );


  buf
  g2163
  (
    n2417,
    n1845
  );


  buf
  g2164
  (
    n2496,
    n2058
  );


  buf
  g2165
  (
    n2118,
    n471
  );


  buf
  g2166
  (
    n2412,
    n1987
  );


  not
  g2167
  (
    n2229,
    n593
  );


  not
  g2168
  (
    n2233,
    n2037
  );


  not
  g2169
  (
    n2310,
    n468
  );


  buf
  g2170
  (
    n2129,
    n499
  );


  not
  g2171
  (
    n2216,
    n1950
  );


  not
  g2172
  (
    n2563,
    n439
  );


  not
  g2173
  (
    n2069,
    n467
  );


  buf
  g2174
  (
    n2116,
    n1963
  );


  not
  g2175
  (
    n2495,
    n602
  );


  buf
  g2176
  (
    n2469,
    n2046
  );


  not
  g2177
  (
    n2214,
    n490
  );


  buf
  g2178
  (
    n2281,
    n640
  );


  not
  g2179
  (
    n2322,
    n2028
  );


  not
  g2180
  (
    n2509,
    n2022
  );


  buf
  g2181
  (
    n2460,
    n451
  );


  not
  g2182
  (
    n2420,
    n2038
  );


  buf
  g2183
  (
    n2158,
    n1933
  );


  not
  g2184
  (
    n2403,
    n618
  );


  buf
  g2185
  (
    n2508,
    n550
  );


  not
  g2186
  (
    n2462,
    n431
  );


  not
  g2187
  (
    n2309,
    n1962
  );


  not
  g2188
  (
    n2067,
    n1977
  );


  buf
  g2189
  (
    n2226,
    n479
  );


  not
  g2190
  (
    n2538,
    n1956
  );


  not
  g2191
  (
    n2077,
    n1957
  );


  not
  g2192
  (
    n2074,
    n592
  );


  buf
  g2193
  (
    n2426,
    n635
  );


  buf
  g2194
  (
    n2381,
    n555
  );


  buf
  g2195
  (
    n2104,
    n1959
  );


  buf
  g2196
  (
    n2114,
    n476
  );


  or
  g2197
  (
    n2303,
    n543,
    n2015,
    n428,
    n470
  );


  nor
  g2198
  (
    n2470,
    n480,
    n506,
    n604,
    n642
  );


  xnor
  g2199
  (
    n2150,
    n436,
    n559,
    n1966,
    n558
  );


  xnor
  g2200
  (
    n2335,
    n567,
    n600,
    n548,
    n457
  );


  xnor
  g2201
  (
    n2185,
    n516,
    n434,
    n1969,
    n589
  );


  xnor
  g2202
  (
    n2551,
    n542,
    n1938,
    n566,
    n440
  );


  xor
  g2203
  (
    n2346,
    n545,
    n597,
    n486,
    n476
  );


  or
  g2204
  (
    n2471,
    n2054,
    n573,
    n2000,
    n439
  );


  xnor
  g2205
  (
    KeyWire_0_20,
    n2017,
    n451,
    n575,
    n569
  );


  nand
  g2206
  (
    n2195,
    n468,
    n450,
    n1942,
    n1965
  );


  xnor
  g2207
  (
    n2357,
    n651,
    n1978,
    n1988,
    n1943
  );


  nor
  g2208
  (
    n2097,
    n1966,
    n1945,
    n530,
    n2038
  );


  and
  g2209
  (
    n2297,
    n537,
    n446,
    n460,
    n668
  );


  xnor
  g2210
  (
    n2360,
    n527,
    n2036,
    n670,
    n444
  );


  xnor
  g2211
  (
    n2405,
    n430,
    n436,
    n651,
    n581
  );


  and
  g2212
  (
    n2501,
    n610,
    n1948,
    n2013,
    n2027
  );


  nand
  g2213
  (
    n2188,
    n1967,
    n543,
    n1958,
    n455
  );


  nand
  g2214
  (
    n2166,
    n445,
    n2006,
    n1965,
    n525
  );


  xor
  g2215
  (
    n2414,
    n421,
    n2042,
    n447,
    n1954
  );


  and
  g2216
  (
    n2456,
    n549,
    n491,
    n490,
    n585
  );


  xnor
  g2217
  (
    n2447,
    n478,
    n2023,
    n672,
    n434
  );


  nor
  g2218
  (
    n2497,
    n1960,
    n515,
    n2046,
    n449
  );


  nand
  g2219
  (
    n2567,
    n630,
    n470,
    n447,
    n637
  );


  xnor
  g2220
  (
    n2131,
    n440,
    n473,
    n521,
    n443
  );


  nand
  g2221
  (
    n2465,
    n660,
    n523,
    n649,
    n482
  );


  nor
  g2222
  (
    n2436,
    n596,
    n518,
    n1989,
    n517
  );


  nand
  g2223
  (
    n2105,
    n581,
    n2021,
    n1844,
    n646
  );


  and
  g2224
  (
    n2458,
    n1998,
    n590,
    n1953,
    n504
  );


  or
  g2225
  (
    n2315,
    n459,
    n515,
    n2049,
    n1992
  );


  xnor
  g2226
  (
    n2243,
    n535,
    n1960,
    n2038,
    n544
  );


  xor
  g2227
  (
    n2064,
    n2034,
    n492,
    n572,
    n658
  );


  or
  g2228
  (
    n2467,
    n615,
    n438,
    n2035,
    n672
  );


  xor
  g2229
  (
    n2557,
    n599,
    n2007,
    n532,
    n2043
  );


  or
  g2230
  (
    n2209,
    n1942,
    n503,
    n567,
    n424
  );


  or
  g2231
  (
    n2092,
    n484,
    n479,
    n542,
    n606
  );


  xor
  g2232
  (
    KeyWire_0_38,
    n546,
    n2033,
    n518,
    n507
  );


  xnor
  g2233
  (
    n2094,
    n431,
    n647,
    n435,
    n640
  );


  or
  g2234
  (
    n2356,
    n448,
    n461,
    n578,
    n1994
  );


  nor
  g2235
  (
    n2262,
    n637,
    n1941,
    n609,
    n487
  );


  xor
  g2236
  (
    n2280,
    n662,
    n616,
    n2053,
    n1962
  );


  and
  g2237
  (
    n2522,
    n2002,
    n521,
    n586,
    n2048
  );


  or
  g2238
  (
    n2318,
    n2049,
    n1963,
    n438,
    n2060
  );


  nand
  g2239
  (
    n2244,
    n441,
    n1977,
    n458,
    n477
  );


  and
  g2240
  (
    n2181,
    n2003,
    n428,
    n2030,
    n656
  );


  nor
  g2241
  (
    n2202,
    n2019,
    n1943,
    n632,
    n495
  );


  or
  g2242
  (
    n2119,
    n560,
    n602,
    n1951,
    n1949
  );


  and
  g2243
  (
    n2160,
    n517,
    n474,
    n635,
    n2055
  );


  nand
  g2244
  (
    n2500,
    n651,
    n627,
    n464,
    n1952
  );


  xnor
  g2245
  (
    n2531,
    n1953,
    n652,
    n1973,
    n636
  );


  nand
  g2246
  (
    n2514,
    n451,
    n2009,
    n467,
    n463
  );


  or
  g2247
  (
    n2134,
    n466,
    n1955,
    n591,
    n2003
  );


  and
  g2248
  (
    n2364,
    n587,
    n1988,
    n516,
    n607
  );


  nand
  g2249
  (
    n2278,
    n520,
    n593,
    n2001,
    n488
  );


  and
  g2250
  (
    n2396,
    n2027,
    n652,
    n1940,
    n653
  );


  or
  g2251
  (
    n2481,
    n461,
    n1964,
    n495,
    n615
  );


  nand
  g2252
  (
    n2384,
    n2021,
    n424,
    n2017,
    n557
  );


  nor
  g2253
  (
    n2386,
    n482,
    n540,
    n435,
    n556
  );


  and
  g2254
  (
    n2378,
    n502,
    n628,
    n2050,
    n429
  );


  nand
  g2255
  (
    n2321,
    n563,
    n502,
    n2056,
    n1943
  );


  nand
  g2256
  (
    KeyWire_0_29,
    n2041,
    n657,
    n665,
    n2052
  );


  nor
  g2257
  (
    n2546,
    n603,
    n1977,
    n2051,
    n453
  );


  and
  g2258
  (
    n2419,
    n632,
    n512,
    n560,
    n430
  );


  and
  g2259
  (
    n2492,
    n541,
    n588,
    n606,
    n570
  );


  or
  g2260
  (
    n2200,
    n522,
    n493,
    n1948,
    n611
  );


  nor
  g2261
  (
    n2325,
    n562,
    n1958,
    n2003,
    n1946
  );


  nand
  g2262
  (
    n2121,
    n483,
    n1980,
    n670,
    n630
  );


  nand
  g2263
  (
    n2217,
    n533,
    n627,
    n630,
    n1975
  );


  or
  g2264
  (
    n2237,
    n658,
    n497,
    n1974,
    n638
  );


  xor
  g2265
  (
    n2120,
    n2053,
    n525,
    n559,
    n531
  );


  nor
  g2266
  (
    n2442,
    n544,
    n2005,
    n465,
    n577
  );


  or
  g2267
  (
    n2532,
    n1968,
    n528,
    n669,
    n646
  );


  nand
  g2268
  (
    n2550,
    n1939,
    n1970,
    n2031,
    n481
  );


  or
  g2269
  (
    n2088,
    n420,
    n519,
    n1961,
    n572
  );


  and
  g2270
  (
    n2345,
    n2015,
    n2043,
    n1961,
    n638
  );


  or
  g2271
  (
    n2276,
    n664,
    n2034,
    n437,
    n2031
  );


  nor
  g2272
  (
    n2135,
    n1995,
    n2041,
    n604,
    n519
  );


  nand
  g2273
  (
    n2545,
    n515,
    n636,
    n558,
    n645
  );


  xnor
  g2274
  (
    n2268,
    n509,
    n504,
    n647,
    n1947
  );


  xnor
  g2275
  (
    n2128,
    n2010,
    n578,
    n453,
    n421
  );


  nor
  g2276
  (
    n2344,
    n1934,
    n1960,
    n626,
    n523
  );


  and
  g2277
  (
    n2296,
    n588,
    n2026,
    n2012,
    n513
  );


  nand
  g2278
  (
    n2355,
    n640,
    n632,
    n489,
    n479
  );


  nor
  g2279
  (
    n2434,
    n2047,
    n1938,
    n614,
    n654
  );


  nor
  g2280
  (
    n2316,
    n664,
    n1967,
    n1979,
    n594
  );


  nor
  g2281
  (
    n2367,
    n2037,
    n643,
    n667,
    n489
  );


  nand
  g2282
  (
    n2340,
    n623,
    n2021,
    n1963,
    n477
  );


  or
  g2283
  (
    n2277,
    n605,
    n483,
    n624,
    n542
  );


  xor
  g2284
  (
    n2075,
    n567,
    n597,
    n666,
    n491
  );


  xnor
  g2285
  (
    n2080,
    n427,
    n597,
    n2035,
    n1987
  );


  xnor
  g2286
  (
    n2457,
    n446,
    n2044,
    n592,
    n667
  );


  and
  g2287
  (
    n2425,
    n565,
    n462,
    n2036,
    n463
  );


  nor
  g2288
  (
    n2339,
    n534,
    n670,
    n2023,
    n480
  );


  or
  g2289
  (
    n2102,
    n542,
    n2011,
    n1982,
    n625
  );


  nor
  g2290
  (
    n2488,
    n505,
    n1969,
    n658,
    n534
  );


  xor
  g2291
  (
    n2093,
    n496,
    n561,
    n2002,
    n656
  );


  nand
  g2292
  (
    n2444,
    n526,
    n451,
    n622,
    n2043
  );


  nor
  g2293
  (
    n2421,
    n669,
    n1945,
    n574,
    n434
  );


  nand
  g2294
  (
    n2302,
    n2023,
    n2001,
    n564,
    n670
  );


  or
  g2295
  (
    n2320,
    n528,
    n425,
    n1979,
    n556
  );


  xor
  g2296
  (
    n2299,
    n618,
    n613,
    n552,
    n522
  );


  nor
  g2297
  (
    n2111,
    n1978,
    n601,
    n620,
    n2015
  );


  or
  g2298
  (
    n2273,
    n1968,
    n505,
    n480,
    n1971
  );


  xnor
  g2299
  (
    n2100,
    n584,
    n430,
    n614,
    n468
  );


  xnor
  g2300
  (
    n2076,
    n549,
    n546,
    n2008,
    n604
  );


  nor
  g2301
  (
    n2570,
    n1984,
    n568,
    n447,
    n2001
  );


  nor
  g2302
  (
    n2096,
    n621,
    n547,
    n486,
    n506
  );


  nor
  g2303
  (
    n2562,
    n667,
    n654,
    n452,
    n2005
  );


  and
  g2304
  (
    n2107,
    n671,
    n541,
    n1939,
    n572
  );


  nor
  g2305
  (
    n2331,
    n1990,
    n2060,
    n578,
    n463
  );


  nand
  g2306
  (
    n2228,
    n1976,
    n1962,
    n478,
    n533
  );


  nand
  g2307
  (
    n2429,
    n2057,
    n2012,
    n492,
    n468
  );


  xor
  g2308
  (
    n2101,
    n497,
    n427,
    n571,
    n2014
  );


  and
  g2309
  (
    n2191,
    n471,
    n2010,
    n1938,
    n664
  );


  xnor
  g2310
  (
    n2542,
    n553,
    n459,
    n628,
    n612
  );


  xnor
  g2311
  (
    n2327,
    n513,
    n529,
    n455,
    n1935
  );


  xor
  g2312
  (
    n2537,
    n2027,
    n595,
    n2029,
    n2025
  );


  nor
  g2313
  (
    n2383,
    n1993,
    n1946,
    n538,
    n640
  );


  nand
  g2314
  (
    n2227,
    n629,
    n1963,
    n510,
    n499
  );


  and
  g2315
  (
    n2084,
    n422,
    n649,
    n1984,
    n657
  );


  xnor
  g2316
  (
    n2475,
    n583,
    n497,
    n1961,
    n566
  );


  nand
  g2317
  (
    n2073,
    n437,
    n2011,
    n554,
    n657
  );


  and
  g2318
  (
    n2198,
    n642,
    n654,
    n518,
    n2032
  );


  xnor
  g2319
  (
    n2334,
    n538,
    n1936,
    n605,
    n1952
  );


  or
  g2320
  (
    n2437,
    n539,
    n442,
    n1942,
    n650
  );


  and
  g2321
  (
    n2317,
    n456,
    n563,
    n2052,
    n634
  );


  xnor
  g2322
  (
    n2463,
    n528,
    n487,
    n2054,
    n662
  );


  nor
  g2323
  (
    n2468,
    n553,
    n1949,
    n523,
    n540
  );


  and
  g2324
  (
    n2527,
    n620,
    n2004,
    n629,
    n2052
  );


  or
  g2325
  (
    n2203,
    n617,
    n2032,
    n603,
    n464
  );


  xor
  g2326
  (
    n2535,
    n425,
    n665,
    n431,
    n1994
  );


  and
  g2327
  (
    n2106,
    n526,
    n557,
    n532,
    n617
  );


  nor
  g2328
  (
    n2192,
    n561,
    n641,
    n611,
    n2048
  );


  xor
  g2329
  (
    n2117,
    n2045,
    n2002,
    n548,
    n420
  );


  or
  g2330
  (
    n2113,
    n596,
    n1972,
    n469,
    n614
  );


  xnor
  g2331
  (
    n2341,
    n594,
    n643,
    n517,
    n1991
  );


  and
  g2332
  (
    n2513,
    n648,
    n481,
    n2047,
    n619
  );


  xnor
  g2333
  (
    n2347,
    n611,
    n476,
    n653,
    n579
  );


  nand
  g2334
  (
    n2248,
    n511,
    n650,
    n607,
    n608
  );


  nor
  g2335
  (
    n2130,
    n612,
    n481,
    n2004,
    n651
  );


  and
  g2336
  (
    n2206,
    n607,
    n444,
    n631,
    n500
  );


  nor
  g2337
  (
    n2072,
    n662,
    n1844,
    n459,
    n637
  );


  nand
  g2338
  (
    n2543,
    n624,
    n543,
    n661,
    n2018
  );


  nand
  g2339
  (
    n2264,
    n1961,
    n530,
    n571,
    n526
  );


  xor
  g2340
  (
    n2263,
    n630,
    n583,
    n528,
    n491
  );


  and
  g2341
  (
    n2312,
    n481,
    n1953,
    n2040,
    n1964
  );


  nor
  g2342
  (
    n2176,
    n467,
    n1982,
    n2007,
    n450
  );


  or
  g2343
  (
    n2285,
    n1944,
    n1955,
    n660,
    n612
  );


  xor
  g2344
  (
    n2526,
    n2028,
    n465,
    n1993,
    n572
  );


  xor
  g2345
  (
    n2328,
    n2051,
    n650,
    n645,
    n599
  );


  and
  g2346
  (
    n2483,
    n2006,
    n1996,
    n582,
    n1946
  );


  nand
  g2347
  (
    n2127,
    n538,
    n1977,
    n655,
    n639
  );


  xor
  g2348
  (
    n2490,
    n514,
    n473,
    n432,
    n2020
  );


  nor
  g2349
  (
    n2138,
    n437,
    n621,
    n456,
    n2015
  );


  nor
  g2350
  (
    n2498,
    n456,
    n433,
    n632,
    n591
  );


  nand
  g2351
  (
    n2284,
    n593,
    n1989,
    n482,
    n493
  );


  or
  g2352
  (
    n2089,
    n475,
    n462,
    n2025,
    n1999
  );


  and
  g2353
  (
    n2155,
    n2007,
    n456,
    n602,
    n426
  );


  and
  g2354
  (
    n2489,
    n564,
    n495,
    n1955,
    n2046
  );


  nand
  g2355
  (
    n2142,
    n527,
    n2006,
    n2057,
    n1956
  );


  xnor
  g2356
  (
    n2288,
    n1972,
    n1933,
    n420,
    n520
  );


  nor
  g2357
  (
    n2210,
    n1993,
    n579,
    n1996,
    n1985
  );


  nor
  g2358
  (
    n2358,
    n635,
    n2051,
    n472,
    n622
  );


  xor
  g2359
  (
    n2140,
    n443,
    n1986,
    n516,
    n498
  );


  nand
  g2360
  (
    n2156,
    n505,
    n624,
    n461,
    n1998
  );


  xnor
  g2361
  (
    n2529,
    n625,
    n634,
    n562,
    n2046
  );


  nor
  g2362
  (
    n2178,
    n603,
    n1998,
    n583,
    n425
  );


  or
  g2363
  (
    n2154,
    n562,
    n1950,
    n457,
    n498
  );


  nor
  g2364
  (
    n2238,
    n556,
    n484,
    n1976,
    n580
  );


  nor
  g2365
  (
    n2087,
    n548,
    n482,
    n655,
    n615
  );


  or
  g2366
  (
    n2549,
    n1995,
    n1962,
    n1996,
    n454
  );


  nor
  g2367
  (
    n2062,
    n484,
    n444,
    n555,
    n582
  );


  or
  g2368
  (
    n2218,
    n494,
    n587,
    n609,
    n2035
  );


  or
  g2369
  (
    n2510,
    n2025,
    n1937,
    n487,
    n574
  );


  nand
  g2370
  (
    n2294,
    n2026,
    n563,
    n609,
    n494
  );


  nor
  g2371
  (
    n2363,
    n580,
    n586,
    n591,
    n454
  );


  or
  g2372
  (
    n2295,
    n500,
    n614,
    n668,
    n2011
  );


  or
  g2373
  (
    n2222,
    n423,
    n2057,
    n615,
    n657
  );


  nor
  g2374
  (
    n2389,
    n655,
    n602,
    n558,
    n1949
  );


  and
  g2375
  (
    n2205,
    n527,
    n455,
    n1991,
    n2000
  );


  xnor
  g2376
  (
    n2163,
    n1937,
    n530,
    n1843,
    n2005
  );


  or
  g2377
  (
    n2197,
    n627,
    n460,
    n506,
    n503
  );


  xnor
  g2378
  (
    n2234,
    n1964,
    n534,
    n1992,
    n2018
  );


  xor
  g2379
  (
    n2068,
    n2022,
    n568,
    n644,
    n2059
  );


  xor
  g2380
  (
    n2499,
    n639,
    n1990,
    n2016,
    n625
  );


  or
  g2381
  (
    n2298,
    n537,
    n2014,
    n434,
    n2049
  );


  nand
  g2382
  (
    n2082,
    n1845,
    n601,
    n1991,
    n498
  );


  or
  g2383
  (
    n2324,
    n474,
    n472,
    n2042,
    n532
  );


  and
  g2384
  (
    n2141,
    n639,
    n1993,
    n1957,
    n2030
  );


  or
  g2385
  (
    n2461,
    n587,
    n543,
    n1934,
    n2017
  );


  xor
  g2386
  (
    n2091,
    n522,
    n531,
    n503,
    n470
  );


  and
  g2387
  (
    n2146,
    n2016,
    n612,
    n2000,
    n462
  );


  xor
  g2388
  (
    n2151,
    n671,
    n475,
    n565,
    n666
  );


  and
  g2389
  (
    n2313,
    n566,
    n592,
    n518,
    n499
  );


  or
  g2390
  (
    n2411,
    n1997,
    n510,
    n1999,
    n487
  );


  and
  g2391
  (
    n2215,
    n647,
    n422,
    n2060,
    n525
  );


  xnor
  g2392
  (
    n2260,
    n1982,
    n1972,
    n2059,
    n505
  );


  and
  g2393
  (
    n2441,
    n1985,
    n608,
    n442,
    n2009
  );


  and
  g2394
  (
    n2173,
    n524,
    n1952,
    n654,
    n1997
  );


  nor
  g2395
  (
    n2272,
    n457,
    n1937,
    n551,
    n666
  );


  or
  g2396
  (
    n2338,
    n598,
    n554,
    n575,
    n1983
  );


  xor
  g2397
  (
    n2231,
    n2053,
    n474,
    n2024,
    n2036
  );


  nand
  g2398
  (
    n2319,
    n627,
    n671,
    n424,
    n2056
  );


  or
  g2399
  (
    n2136,
    n1845,
    n2047,
    n619,
    n2012
  );


  nand
  g2400
  (
    n2145,
    n656,
    n452,
    n529,
    n1970
  );


  nand
  g2401
  (
    n2554,
    n422,
    n573,
    n549,
    n585
  );


  nor
  g2402
  (
    KeyWire_0_26,
    n1940,
    n521,
    n493,
    n2039
  );


  nor
  g2403
  (
    n2286,
    n2034,
    n617,
    n449,
    n440
  );


  xnor
  g2404
  (
    n2306,
    n621,
    n580,
    n537,
    n1939
  );


  nand
  g2405
  (
    n2249,
    n649,
    n2008,
    n1973,
    n605
  );


  and
  g2406
  (
    n2391,
    n475,
    n582,
    n1985,
    n2058
  );


  xnor
  g2407
  (
    n2329,
    n577,
    n653,
    n431,
    n576
  );


  xor
  g2408
  (
    KeyWire_0_34,
    n641,
    n438,
    n634,
    n478
  );


  or
  g2409
  (
    n2534,
    n619,
    n643,
    n476,
    n1947
  );


  and
  g2410
  (
    n2394,
    n510,
    n2044,
    n429,
    n642
  );


  nand
  g2411
  (
    n2125,
    n2060,
    n1970,
    n633,
    n2019
  );


  xnor
  g2412
  (
    n2109,
    n639,
    n2005,
    n1976,
    n2002
  );


  xor
  g2413
  (
    n2208,
    n423,
    n2047,
    n536,
    n501
  );


  xnor
  g2414
  (
    n2070,
    n667,
    n509,
    n610,
    n586
  );


  xnor
  g2415
  (
    n2512,
    n2058,
    n537,
    n622,
    n1994
  );


  nor
  g2416
  (
    n2333,
    n2058,
    n429,
    n2059,
    n1934
  );


  or
  g2417
  (
    n2406,
    n638,
    n618,
    n1951,
    n546
  );


  and
  g2418
  (
    n2373,
    n540,
    n472,
    n466,
    n589
  );


  nor
  g2419
  (
    n2375,
    n2013,
    n661,
    n545,
    n604
  );


  nand
  g2420
  (
    n2452,
    n662,
    n2043,
    n1945,
    n583
  );


  or
  g2421
  (
    n2372,
    n2035,
    n1983,
    n477,
    n559
  );


  xnor
  g2422
  (
    n2225,
    n587,
    n1845,
    n469,
    n633
  );


  nand
  g2423
  (
    n2079,
    n461,
    n626,
    n2013,
    n608
  );


  and
  g2424
  (
    n2122,
    n620,
    n546,
    n2007,
    n489
  );


  xor
  g2425
  (
    n2301,
    n1999,
    n601,
    n547,
    n2019
  );


  nand
  g2426
  (
    n2379,
    n1979,
    n460,
    n2056,
    n472
  );


  and
  g2427
  (
    n2399,
    n477,
    n489,
    n471,
    n509
  );


  and
  g2428
  (
    n2416,
    n502,
    n535,
    n435,
    n669
  );


  nor
  g2429
  (
    n2083,
    n2039,
    n466,
    n508,
    n526
  );


  xor
  g2430
  (
    n2170,
    n496,
    n2024,
    n1956,
    n1971
  );


  nand
  g2431
  (
    n2439,
    n1984,
    n1936,
    n554,
    n625
  );


  xnor
  g2432
  (
    n2479,
    n519,
    n2000,
    n2042,
    n2044
  );


  nor
  g2433
  (
    n2359,
    n1971,
    n608,
    n2051,
    n479
  );


  xor
  g2434
  (
    n2401,
    n573,
    n500,
    n2037,
    n628
  );


  xor
  g2435
  (
    n2430,
    n419,
    n480,
    n2057,
    n2001
  );


  xnor
  g2436
  (
    n2123,
    n570,
    n610,
    n565,
    n527
  );


  xnor
  g2437
  (
    n2466,
    n1983,
    n2050,
    n551,
    n2040
  );


  nor
  g2438
  (
    n2366,
    n540,
    n530,
    n1973,
    n661
  );


  xnor
  g2439
  (
    n2332,
    n592,
    n465,
    n1989,
    n1951
  );


  xor
  g2440
  (
    n2400,
    n616,
    n547,
    n1943,
    n1941
  );


  or
  g2441
  (
    n2232,
    n485,
    n2029,
    n665,
    n672
  );


  nor
  g2442
  (
    n2519,
    n658,
    n490,
    n659,
    n586
  );


  nor
  g2443
  (
    n2395,
    n2044,
    n433,
    n539,
    n1935
  );


  and
  g2444
  (
    n2553,
    n605,
    n425,
    n469,
    n643
  );


  nor
  g2445
  (
    n2086,
    n1942,
    n634,
    n423,
    n620
  );


  xnor
  g2446
  (
    n2326,
    n520,
    n635,
    n426,
    n2038
  );


  or
  g2447
  (
    n2224,
    n1986,
    n607,
    n506,
    n533
  );


  xnor
  g2448
  (
    n2239,
    n444,
    n2022,
    n1967,
    n569
  );


  and
  g2449
  (
    n2065,
    n2016,
    n595,
    n1980,
    n613
  );


  xnor
  g2450
  (
    n2516,
    n432,
    n512,
    n1960,
    n581
  );


  and
  g2451
  (
    n2314,
    n579,
    n435,
    n515,
    n2031
  );


  xor
  g2452
  (
    n2482,
    n517,
    n502,
    n486,
    n567
  );


  and
  g2453
  (
    n2402,
    n1999,
    n1997,
    n508,
    n1973
  );


  and
  g2454
  (
    n2183,
    n561,
    n1995,
    n648,
    n578
  );


  xnor
  g2455
  (
    n2071,
    n594,
    n563,
    n1946,
    n1992
  );


  xor
  g2456
  (
    n2143,
    n1957,
    n1935,
    n539,
    n2048
  );


  and
  g2457
  (
    n2247,
    n2003,
    n1954,
    n672,
    n488
  );


  or
  g2458
  (
    n2415,
    n1944,
    n494,
    n1983,
    n590
  );


  xor
  g2459
  (
    n2487,
    n568,
    n1986,
    n484,
    n570
  );


  and
  g2460
  (
    n2385,
    n483,
    n513,
    n641,
    n1948
  );


  or
  g2461
  (
    n2211,
    n621,
    n436,
    n584,
    n2045
  );


  and
  g2462
  (
    n2451,
    n663,
    n551,
    n595,
    n2020
  );


  and
  g2463
  (
    n2507,
    n2028,
    n553,
    n1966,
    n576
  );


  xor
  g2464
  (
    n2162,
    n1970,
    n2052,
    n459,
    n1940
  );


  nand
  g2465
  (
    n2063,
    n597,
    n458,
    n1978,
    n623
  );


  xor
  g2466
  (
    n2493,
    n469,
    n1980,
    n1995,
    n613
  );


  xor
  g2467
  (
    n2103,
    n1958,
    n575,
    n493,
    n498
  );


  nor
  g2468
  (
    n2422,
    n1975,
    n598,
    n652,
    n495
  );


  and
  g2469
  (
    n2418,
    n2055,
    n488,
    n448,
    n508
  );


  xnor
  g2470
  (
    n2353,
    n2039,
    n599,
    n610,
    n595
  );


  nand
  g2471
  (
    n2207,
    n1935,
    n655,
    n1949,
    n1941
  );


  and
  g2472
  (
    n2382,
    n613,
    n446,
    n1965,
    n2037
  );


  xnor
  g2473
  (
    n2165,
    n622,
    n2054,
    n554,
    n560
  );


  nor
  g2474
  (
    n2478,
    n541,
    n2009,
    n2006,
    n1967
  );


  and
  g2475
  (
    n2566,
    n553,
    n510,
    n1955,
    n2041
  );


  nand
  g2476
  (
    n2361,
    n1952,
    n519,
    n1976,
    n445
  );


  xnor
  g2477
  (
    n2533,
    n458,
    n2039,
    n449,
    n1958
  );


  xor
  g2478
  (
    n2098,
    n564,
    n534,
    n644,
    n2024
  );


  nand
  g2479
  (
    n2139,
    n507,
    n508,
    n458,
    n564
  );


  and
  g2480
  (
    n2112,
    n2033,
    n511,
    n2045,
    n433
  );


  nand
  g2481
  (
    n2287,
    n1844,
    n545,
    n442,
    n1974
  );


  and
  g2482
  (
    n2290,
    n1974,
    n2004,
    n2033,
    n666
  );


  xor
  g2483
  (
    n2108,
    n576,
    n2012,
    n552,
    n663
  );


  or
  g2484
  (
    n2377,
    n520,
    n2009,
    n547,
    n437
  );


  and
  g2485
  (
    n2171,
    n660,
    n603,
    n421,
    n2048
  );


  or
  g2486
  (
    n2506,
    n631,
    n465,
    n2026,
    n496
  );


  and
  g2487
  (
    n2336,
    n514,
    n2050,
    n494,
    n511
  );


  xnor
  g2488
  (
    n2300,
    n501,
    n492,
    n428,
    n429
  );


  xnor
  g2489
  (
    n2189,
    n650,
    n2033,
    n561,
    n584
  );


  and
  g2490
  (
    n2190,
    n447,
    n594,
    n2026,
    n2040
  );


  and
  g2491
  (
    n2330,
    n421,
    n656,
    n1965,
    n541
  );


  nand
  g2492
  (
    n2503,
    n432,
    n1947,
    n1966,
    n2024
  );


  xnor
  g2493
  (
    n2565,
    n659,
    n648,
    n560,
    n2054
  );


  xor
  g2494
  (
    n2376,
    n504,
    n623,
    n1982,
    n441
  );


  or
  g2495
  (
    n2169,
    n445,
    n665,
    n2019,
    n2027
  );


  nor
  g2496
  (
    n2085,
    n2011,
    n606,
    n661,
    n562
  );


  and
  g2497
  (
    n2179,
    n1985,
    n438,
    n448,
    n1996
  );


  or
  g2498
  (
    n2368,
    n574,
    n574,
    n649,
    n533
  );


  nor
  g2499
  (
    KeyWire_0_2,
    n590,
    n1953,
    n600,
    n500
  );


  or
  g2500
  (
    n2152,
    n513,
    n2014,
    n424,
    n432
  );


  xor
  g2501
  (
    n2182,
    n598,
    n1950,
    n2008,
    n430
  );


  xor
  g2502
  (
    n2282,
    n2010,
    n1956,
    n2020,
    n423
  );


  or
  g2503
  (
    n2099,
    n646,
    n571,
    n575,
    n441
  );


  or
  g2504
  (
    n2291,
    n524,
    n2018,
    n471,
    n644
  );


  nand
  g2505
  (
    n2305,
    n1944,
    n1969,
    n452,
    n1992
  );


  or
  g2506
  (
    n2564,
    n439,
    n1968,
    n669,
    n593
  );


  xnor
  g2507
  (
    n2464,
    n488,
    n633,
    n485,
    n532
  );


  xor
  g2508
  (
    n2147,
    n1951,
    n1950,
    n474,
    n464
  );


  or
  g2509
  (
    n2078,
    n551,
    n569,
    n1954,
    n457
  );


  or
  g2510
  (
    n2167,
    n644,
    n659,
    n473,
    n577
  );


  xnor
  g2511
  (
    n2246,
    n552,
    n1984,
    n491,
    n475
  );


  xnor
  g2512
  (
    n2424,
    n443,
    n2029,
    n507,
    n579
  );


  nand
  g2513
  (
    n2350,
    n1939,
    n549,
    n1981,
    n1991
  );


  and
  g2514
  (
    n2265,
    n599,
    n2010,
    n499,
    n1969
  );


  xnor
  g2515
  (
    n2258,
    n426,
    n2031,
    n536,
    n576
  );


  xor
  g2516
  (
    n2407,
    n596,
    n531,
    n653,
    n524
  );


  xor
  g2517
  (
    n2343,
    n496,
    n589,
    n525,
    n443
  );


  nor
  g2518
  (
    n2271,
    n2034,
    n420,
    n1947,
    n642
  );


  nor
  g2519
  (
    n2240,
    n601,
    n616,
    n631,
    n600
  );


  xnor
  g2520
  (
    n2251,
    n2041,
    n446,
    n490,
    n1974
  );


  and
  g2521
  (
    n2283,
    n545,
    n2025,
    n453,
    n529
  );


  or
  g2522
  (
    n2555,
    n591,
    n531,
    n585,
    n582
  );


  nand
  g2523
  (
    n2480,
    n1975,
    n1981,
    n512,
    n1938
  );


  xnor
  g2524
  (
    n2540,
    n663,
    n439,
    n664,
    n668
  );


  nor
  g2525
  (
    n2201,
    n648,
    n1937,
    n449,
    n511
  );


  or
  g2526
  (
    n2148,
    n514,
    n616,
    n2029,
    n460
  );


  or
  g2527
  (
    n2159,
    n462,
    n544,
    n538,
    n450
  );


  and
  g2528
  (
    n2450,
    n581,
    n1987,
    n419,
    n467
  );


  and
  g2529
  (
    n2259,
    n596,
    n501,
    n521,
    n555
  );


  xor
  g2530
  (
    n2428,
    n2050,
    n556,
    n629,
    n1968
  );


  or
  g2531
  (
    n2409,
    n645,
    n536,
    n637,
    n441
  );


  xor
  g2532
  (
    n2474,
    n2049,
    n570,
    n559,
    n450
  );


  nor
  g2533
  (
    n2220,
    n609,
    n628,
    n503,
    n1959
  );


  and
  g2534
  (
    n2257,
    n455,
    n2030,
    n2022,
    n1936
  );


  xnor
  g2535
  (
    KeyWire_0_15,
    n440,
    n618,
    n2016,
    n1934
  );


  or
  g2536
  (
    n2311,
    n1979,
    n590,
    n1972,
    n571
  );


  nor
  g2537
  (
    n2115,
    n427,
    n501,
    n433,
    n626
  );


  nor
  g2538
  (
    n2605,
    n1185,
    n865,
    n1320
  );


  xor
  g2539
  (
    n2907,
    n1536,
    n1078,
    n1379
  );


  xnor
  g2540
  (
    n2660,
    n1243,
    n2245,
    n2344,
    n1034
  );


  xnor
  g2541
  (
    n2587,
    n1281,
    n1637,
    n2459,
    n2364
  );


  and
  g2542
  (
    n2879,
    n1383,
    n991,
    n921,
    n1474
  );


  and
  g2543
  (
    n2653,
    n912,
    n1464,
    n1250,
    n1343
  );


  or
  g2544
  (
    n2727,
    n828,
    n1602,
    n1068,
    n2117
  );


  and
  g2545
  (
    n2844,
    n2500,
    n2360,
    n1192,
    n2385
  );


  nor
  g2546
  (
    n2690,
    n2552,
    n2299,
    n1666,
    n1214
  );


  and
  g2547
  (
    n2886,
    n1187,
    n2278,
    n2132,
    n2323
  );


  and
  g2548
  (
    n2883,
    n1642,
    n978,
    n2486,
    n1172
  );


  nand
  g2549
  (
    n2662,
    n1404,
    n881,
    n2448,
    n1420
  );


  or
  g2550
  (
    n2623,
    n2116,
    n1455,
    n2509,
    n2414
  );


  or
  g2551
  (
    n2843,
    n1401,
    n1213,
    n1410,
    n2186
  );


  xor
  g2552
  (
    n2700,
    n886,
    n1591,
    n1378,
    n2562
  );


  xor
  g2553
  (
    n2830,
    n2149,
    n836,
    n1441,
    n1162
  );


  xnor
  g2554
  (
    n2762,
    n1066,
    n1305,
    n903,
    n2553
  );


  and
  g2555
  (
    n2701,
    n2438,
    n955,
    n877,
    n929
  );


  and
  g2556
  (
    n2910,
    n939,
    n1044,
    n2536,
    n2103
  );


  nand
  g2557
  (
    n2868,
    n1201,
    n1451,
    n1030,
    n1291
  );


  xor
  g2558
  (
    n2905,
    n2260,
    n888,
    n1104,
    n2119
  );


  xor
  g2559
  (
    n2884,
    n2286,
    n853,
    n879,
    n1503
  );


  xnor
  g2560
  (
    n2691,
    n2238,
    n1399,
    n1296,
    n2558
  );


  xnor
  g2561
  (
    n2800,
    n838,
    n1691,
    n1309,
    n1101
  );


  xor
  g2562
  (
    n2812,
    n2387,
    n1613,
    n1431,
    n2475
  );


  or
  g2563
  (
    n2659,
    n924,
    n1335,
    n2519,
    n1042
  );


  xnor
  g2564
  (
    n2854,
    n2546,
    n1587,
    n1136,
    n1247
  );


  nand
  g2565
  (
    n2889,
    n1523,
    n874,
    n1607,
    n938
  );


  nor
  g2566
  (
    n2842,
    n2392,
    n2322,
    n2432,
    n2240
  );


  nor
  g2567
  (
    n2644,
    n1585,
    n1499,
    n1472,
    n910
  );


  nand
  g2568
  (
    n2719,
    n968,
    n894,
    n919,
    n1077
  );


  nor
  g2569
  (
    n2922,
    n2568,
    n2489,
    n2504,
    n2391
  );


  and
  g2570
  (
    n2867,
    n1069,
    n963,
    n855,
    n2168
  );


  xnor
  g2571
  (
    n2602,
    n1462,
    n2404,
    n1609,
    n2137
  );


  and
  g2572
  (
    n2792,
    n844,
    n2461,
    n1385,
    n2095
  );


  nand
  g2573
  (
    n2829,
    n1649,
    n2274,
    n1052,
    n2456
  );


  nand
  g2574
  (
    n2920,
    n2211,
    n1220,
    n1498,
    n923
  );


  and
  g2575
  (
    n2598,
    n933,
    n1696,
    n1382,
    n2347
  );


  and
  g2576
  (
    n2861,
    n920,
    n825,
    n2268,
    n2452
  );


  xnor
  g2577
  (
    n2752,
    n1210,
    n1226,
    n2405,
    n1260
  );


  and
  g2578
  (
    n2797,
    n926,
    n1515,
    n2317,
    n1606
  );


  xnor
  g2579
  (
    n2694,
    n845,
    n1135,
    n2421,
    n2166
  );


  or
  g2580
  (
    n2864,
    n1456,
    n2273,
    n2130,
    n2141
  );


  or
  g2581
  (
    n2919,
    n1163,
    n1510,
    n2378,
    n1211
  );


  nor
  g2582
  (
    n2651,
    n1173,
    n1149,
    n2363,
    n870
  );


  or
  g2583
  (
    n2876,
    n1507,
    n1482,
    n1511,
    n2366
  );


  xnor
  g2584
  (
    n2833,
    n2239,
    n1393,
    n1589,
    n1153
  );


  xor
  g2585
  (
    n2898,
    n2189,
    n1065,
    n1660,
    n1158
  );


  nor
  g2586
  (
    n2869,
    n1533,
    n2181,
    n2261,
    n2557
  );


  nor
  g2587
  (
    n2607,
    n1692,
    n1395,
    n1408,
    n1359
  );


  nand
  g2588
  (
    n2579,
    n2297,
    n1377,
    n1661,
    n1390
  );


  xor
  g2589
  (
    n2768,
    n2267,
    n2092,
    n2534,
    n1290
  );


  or
  g2590
  (
    n2726,
    n1471,
    n1543,
    n954,
    n2518
  );


  nand
  g2591
  (
    n2865,
    n2341,
    n1484,
    n2225,
    n1434
  );


  nand
  g2592
  (
    n2737,
    n2449,
    n1415,
    n1470,
    n1570
  );


  xnor
  g2593
  (
    n2652,
    n1346,
    n2316,
    n1341,
    n1009
  );


  xor
  g2594
  (
    n2738,
    n832,
    n2336,
    n1119,
    n2259
  );


  nand
  g2595
  (
    n2717,
    n2511,
    n1165,
    n1270,
    n2532
  );


  or
  g2596
  (
    n2755,
    n1697,
    n1063,
    n1411,
    n1224
  );


  xor
  g2597
  (
    n2610,
    n1204,
    n2516,
    n2473,
    n1433
  );


  xor
  g2598
  (
    n2591,
    n2277,
    n1110,
    n858,
    n2453
  );


  and
  g2599
  (
    n2803,
    n1081,
    n2515,
    n2174,
    n1171
  );


  nor
  g2600
  (
    n2704,
    n1271,
    n981,
    n1632,
    n2325
  );


  nand
  g2601
  (
    n2714,
    n1500,
    n2228,
    n2235,
    n2544
  );


  or
  g2602
  (
    n2645,
    n1221,
    n1245,
    n1612,
    n1690
  );


  or
  g2603
  (
    n2697,
    n1155,
    n1116,
    n1300,
    n1641
  );


  xnor
  g2604
  (
    n2713,
    n937,
    n931,
    n2476,
    n1579
  );


  nor
  g2605
  (
    n2784,
    n2150,
    n1048,
    n1313,
    n1447
  );


  xnor
  g2606
  (
    n2724,
    n2255,
    n1495,
    n1358,
    n1046
  );


  xor
  g2607
  (
    n2888,
    n1349,
    n2410,
    n2066,
    n1516
  );


  xnor
  g2608
  (
    n2706,
    n1005,
    n1638,
    n2242,
    n1053
  );


  xor
  g2609
  (
    n2841,
    n1361,
    n2159,
    n1647,
    n2298
  );


  and
  g2610
  (
    n2725,
    n2388,
    n1563,
    n1107,
    n1483
  );


  or
  g2611
  (
    n2680,
    n2447,
    n2418,
    n1592,
    n2063
  );


  nor
  g2612
  (
    n2572,
    n2281,
    n2241,
    n1279,
    n1113
  );


  xor
  g2613
  (
    n2915,
    n1397,
    n2280,
    n917,
    n2350
  );


  and
  g2614
  (
    n2821,
    n804,
    n2236,
    n1079,
    n909
  );


  or
  g2615
  (
    n2685,
    n1036,
    n1012,
    n2146,
    n2199
  );


  and
  g2616
  (
    n2676,
    n2482,
    n1272,
    n1630,
    n1038
  );


  and
  g2617
  (
    n2743,
    n959,
    n1685,
    n1025,
    n1453
  );


  nor
  g2618
  (
    n2663,
    n2098,
    n1405,
    n2570,
    n2138
  );


  or
  g2619
  (
    n2614,
    n2389,
    n1476,
    n1645,
    n1098
  );


  or
  g2620
  (
    n2838,
    n1248,
    n1253,
    n990,
    n2072
  );


  xnor
  g2621
  (
    n2748,
    n2480,
    n1229,
    n2287,
    n884
  );


  xor
  g2622
  (
    n2603,
    n1575,
    n1049,
    n2233,
    n1094
  );


  xor
  g2623
  (
    n2739,
    n1156,
    n1132,
    n2365,
    n2151
  );


  xnor
  g2624
  (
    n2809,
    n1352,
    n1635,
    n2219,
    n1479
  );


  and
  g2625
  (
    n2871,
    n1103,
    n2229,
    n1108,
    n810
  );


  xnor
  g2626
  (
    n2798,
    n1159,
    n1586,
    n833,
    n2324
  );


  and
  g2627
  (
    n2604,
    n2538,
    n2210,
    n1651,
    n1659
  );


  xnor
  g2628
  (
    n2708,
    n1519,
    n987,
    n1086,
    n1062
  );


  and
  g2629
  (
    n2613,
    n1106,
    n1488,
    n1329,
    n1478
  );


  and
  g2630
  (
    n2649,
    n2481,
    n984,
    n1561,
    n1633
  );


  xnor
  g2631
  (
    n2799,
    n2145,
    n2428,
    n2442,
    n1573
  );


  nand
  g2632
  (
    n2575,
    n2477,
    n1562,
    n2069,
    n2462
  );


  xnor
  g2633
  (
    n2832,
    n1332,
    n1384,
    n2490,
    n1282
  );


  and
  g2634
  (
    n2790,
    n2083,
    n1386,
    n1508,
    n1091
  );


  nor
  g2635
  (
    n2763,
    n1540,
    n2468,
    n2315,
    n1344
  );


  and
  g2636
  (
    n2847,
    n902,
    n2252,
    n988,
    n1342
  );


  or
  g2637
  (
    n2771,
    n2133,
    n2180,
    n2437,
    n1620
  );


  nor
  g2638
  (
    n2880,
    n940,
    n2431,
    n1608,
    n2422
  );


  and
  g2639
  (
    n2596,
    n2455,
    n1437,
    n1436,
    n2182
  );


  xor
  g2640
  (
    n2816,
    n1125,
    n2470,
    n2310,
    n1581
  );


  nor
  g2641
  (
    n2577,
    n1460,
    n964,
    n1310,
    n2177
  );


  xor
  g2642
  (
    n2734,
    n2091,
    n1000,
    n2533,
    n1502
  );


  or
  g2643
  (
    n2901,
    n1152,
    n878,
    n1016,
    n899
  );


  nand
  g2644
  (
    n2695,
    n1301,
    n1463,
    n882,
    n1539
  );


  xnor
  g2645
  (
    n2828,
    n1675,
    n2358,
    n2296,
    n1365
  );


  or
  g2646
  (
    n2622,
    n1655,
    n2156,
    n1496,
    n2107
  );


  nand
  g2647
  (
    n2722,
    n970,
    n1597,
    n1501,
    n1619
  );


  and
  g2648
  (
    n2894,
    n1514,
    n1676,
    n1409,
    n1139
  );


  xnor
  g2649
  (
    n2887,
    n1681,
    n2309,
    n1285,
    n2346
  );


  nor
  g2650
  (
    n2658,
    n2231,
    n2221,
    n1075,
    n2303
  );


  nand
  g2651
  (
    n2896,
    n934,
    n1233,
    n1636,
    n2213
  );


  or
  g2652
  (
    n2785,
    n2564,
    n1055,
    n1373,
    n1089
  );


  and
  g2653
  (
    n2656,
    n1008,
    n2335,
    n1461,
    n1193
  );


  nand
  g2654
  (
    n2692,
    n2232,
    n1672,
    n1297,
    n1096
  );


  or
  g2655
  (
    n2912,
    n2301,
    n1467,
    n2294,
    n1526
  );


  or
  g2656
  (
    n2606,
    n2248,
    n1311,
    n2528,
    n1258
  );


  or
  g2657
  (
    n2666,
    n1150,
    n2202,
    n1123,
    n1531
  );


  xor
  g2658
  (
    n2782,
    n1569,
    n2305,
    n830,
    n2373
  );


  xnor
  g2659
  (
    n2599,
    n1648,
    n1120,
    n1051,
    n2089
  );


  and
  g2660
  (
    n2845,
    n1217,
    n1288,
    n2204,
    n1315
  );


  or
  g2661
  (
    n2628,
    n1164,
    n1554,
    n2176,
    n818
  );


  and
  g2662
  (
    n2720,
    n928,
    n2357,
    n2311,
    n1186
  );


  and
  g2663
  (
    n2787,
    n860,
    n1137,
    n2099,
    n2464
  );


  and
  g2664
  (
    n2916,
    n1095,
    n2173,
    n898,
    n2474
  );


  nor
  g2665
  (
    n2616,
    n2065,
    n1306,
    n1177,
    n2551
  );


  and
  g2666
  (
    n2627,
    n1190,
    n2527,
    n1583,
    n1392
  );


  nand
  g2667
  (
    n2902,
    n1147,
    n1218,
    n2412,
    n2400
  );


  and
  g2668
  (
    n2822,
    n2487,
    n1355,
    n2188,
    n1255
  );


  and
  g2669
  (
    n2683,
    n890,
    n1584,
    n2348,
    n1076
  );


  and
  g2670
  (
    n2730,
    n1422,
    n1225,
    n861,
    n2131
  );


  and
  g2671
  (
    n2840,
    n1574,
    n1695,
    n2326,
    n1356
  );


  and
  g2672
  (
    n2594,
    n1231,
    n1154,
    n1559,
    n1535
  );


  or
  g2673
  (
    n2857,
    n1146,
    n2381,
    n1654,
    n2403
  );


  nand
  g2674
  (
    n2633,
    n1209,
    n2193,
    n2520,
    n1580
  );


  xor
  g2675
  (
    n2735,
    n2494,
    n2114,
    n1195,
    n1273
  );


  nand
  g2676
  (
    KeyWire_0_46,
    n1351,
    n1235,
    n1459,
    n2469
  );


  xor
  g2677
  (
    n2674,
    n911,
    n2435,
    n2081,
    n2155
  );


  nand
  g2678
  (
    n2754,
    n1544,
    n2147,
    n1438,
    n958
  );


  nor
  g2679
  (
    n2654,
    n2275,
    n1194,
    n1576,
    n1184
  );


  nand
  g2680
  (
    KeyWire_0_23,
    n1133,
    n1617,
    n1307,
    n1400
  );


  and
  g2681
  (
    n2705,
    n2407,
    n1521,
    n2415,
    n1480
  );


  xor
  g2682
  (
    n2612,
    n2064,
    n2471,
    n2258,
    n1264
  );


  xnor
  g2683
  (
    n2764,
    n2256,
    n2111,
    n2550,
    n2554
  );


  xnor
  g2684
  (
    n2657,
    n1566,
    n1330,
    n1360,
    n992
  );


  and
  g2685
  (
    n2686,
    n2169,
    n1284,
    n1109,
    n2368
  );


  xnor
  g2686
  (
    n2573,
    n2224,
    n2370,
    n1067,
    n852
  );


  xnor
  g2687
  (
    n2583,
    n1114,
    n2078,
    n1624,
    n1338
  );


  nor
  g2688
  (
    n2778,
    n2152,
    n2093,
    n1277,
    n2445
  );


  or
  g2689
  (
    n2890,
    n1669,
    n1170,
    n1045,
    n1457
  );


  nand
  g2690
  (
    n2665,
    n966,
    n1318,
    n895,
    n1299
  );


  nor
  g2691
  (
    n2624,
    n1442,
    n1212,
    n2406,
    n2086
  );


  or
  g2692
  (
    n2702,
    n824,
    n1626,
    n1428,
    n1683
  );


  or
  g2693
  (
    n2766,
    n805,
    n1370,
    n2343,
    n2122
  );


  or
  g2694
  (
    n2873,
    n2506,
    n2222,
    n1550,
    n875
  );


  nand
  g2695
  (
    n2729,
    n2136,
    n1203,
    n2230,
    n2067
  );


  nor
  g2696
  (
    n2750,
    n2104,
    n2144,
    n2270,
    n1407
  );


  xor
  g2697
  (
    n2740,
    n2444,
    n862,
    n2250,
    n1694
  );


  and
  g2698
  (
    n2848,
    n1429,
    n1682,
    n1601,
    n1047
  );


  xor
  g2699
  (
    n2742,
    n2411,
    n2153,
    n2307,
    n2206
  );


  and
  g2700
  (
    n2813,
    n1032,
    n2143,
    n1375,
    n2109
  );


  nor
  g2701
  (
    n2851,
    n2427,
    n1517,
    n975,
    n2382
  );


  and
  g2702
  (
    n2595,
    n2543,
    n1037,
    n2423,
    n2510
  );


  xor
  g2703
  (
    n2780,
    n1611,
    n1327,
    n1105,
    n974
  );


  nor
  g2704
  (
    n2642,
    n1458,
    n2499,
    n943,
    n1181
  );


  xnor
  g2705
  (
    n2904,
    n1525,
    n2154,
    n1532,
    n1430
  );


  or
  g2706
  (
    n2588,
    n1662,
    n905,
    n1031,
    n1621
  );


  and
  g2707
  (
    n2736,
    n1207,
    n2361,
    n2417,
    n1371
  );


  and
  g2708
  (
    n2849,
    n1673,
    n977,
    n998,
    n872
  );


  or
  g2709
  (
    n2921,
    n1588,
    n1593,
    n2096,
    n1357
  );


  and
  g2710
  (
    n2707,
    n2483,
    n843,
    n1222,
    n2450
  );


  nand
  g2711
  (
    n2574,
    n1674,
    n2430,
    n2115,
    n821
  );


  xor
  g2712
  (
    n2671,
    n1481,
    n969,
    n2522,
    n871
  );


  nand
  g2713
  (
    n2639,
    n957,
    n965,
    n819,
    n1653
  );


  and
  g2714
  (
    n2796,
    n2314,
    n834,
    n1506,
    n2306
  );


  or
  g2715
  (
    n2757,
    n2371,
    n935,
    n985,
    n1168
  );


  xnor
  g2716
  (
    n2804,
    n1688,
    n889,
    n2243,
    n945
  );


  xnor
  g2717
  (
    n2877,
    n807,
    n1174,
    n2272,
    n2380
  );


  and
  g2718
  (
    n2721,
    n2257,
    n1557,
    n2165,
    n1530
  );


  nor
  g2719
  (
    n2571,
    n2175,
    n1259,
    n1265,
    n1080
  );


  and
  g2720
  (
    n2918,
    n1440,
    n1236,
    n1041,
    n1021
  );


  xor
  g2721
  (
    n2677,
    n1492,
    n1452,
    n2201,
    n941
  );


  xnor
  g2722
  (
    n2900,
    n1274,
    n1398,
    n2279,
    n1443
  );


  xnor
  g2723
  (
    n2745,
    n1287,
    n1126,
    n1064,
    n1509
  );


  and
  g2724
  (
    n2856,
    n1219,
    n2217,
    n1180,
    n864
  );


  nor
  g2725
  (
    n2731,
    n980,
    n2539,
    n1088,
    n1416
  );


  nand
  g2726
  (
    n2789,
    n1317,
    n1486,
    n1616,
    n1276
  );


  xor
  g2727
  (
    n2909,
    n1699,
    n2349,
    n2192,
    n1527
  );


  nor
  g2728
  (
    n2818,
    n1027,
    n820,
    n1680,
    n2134
  );


  xor
  g2729
  (
    n2621,
    n2401,
    n953,
    n1169,
    n1551
  );


  nor
  g2730
  (
    n2749,
    n1679,
    n2187,
    n2071,
    n1205
  );


  nand
  g2731
  (
    n2668,
    n1175,
    n2501,
    n1505,
    n2079
  );


  xor
  g2732
  (
    n2814,
    n1176,
    n1019,
    n2327,
    n2458
  );


  nor
  g2733
  (
    n2715,
    n2395,
    n1197,
    n1667,
    n2090
  );


  nor
  g2734
  (
    n2853,
    n2399,
    n896,
    n1454,
    n2249
  );


  nand
  g2735
  (
    KeyWire_0_6,
    n1534,
    n2386,
    n1689,
    n1129
  );


  xnor
  g2736
  (
    n2664,
    n2285,
    n2283,
    n1002,
    n1614
  );


  xnor
  g2737
  (
    n2824,
    n1246,
    n2355,
    n1128,
    n851
  );


  nand
  g2738
  (
    n2881,
    n1202,
    n2185,
    n837,
    n863
  );


  xor
  g2739
  (
    n2815,
    n1326,
    n1541,
    n2123,
    n2214
  );


  or
  g2740
  (
    n2772,
    n1389,
    n999,
    n2140,
    n2263
  );


  and
  g2741
  (
    n2576,
    n2313,
    n2318,
    n841,
    n1678
  );


  nand
  g2742
  (
    n2646,
    n839,
    n812,
    n2508,
    n2319
  );


  xor
  g2743
  (
    n2913,
    n859,
    n2408,
    n1157,
    n868
  );


  nor
  g2744
  (
    n2744,
    n1639,
    n2342,
    n2124,
    n1435
  );


  nor
  g2745
  (
    n2801,
    n1206,
    n916,
    n1605,
    n1191
  );


  xnor
  g2746
  (
    n2600,
    n848,
    n993,
    n907,
    n854
  );


  and
  g2747
  (
    n2643,
    n1652,
    n2495,
    n2436,
    n1387
  );


  xor
  g2748
  (
    n2672,
    n1671,
    n1060,
    n2209,
    n2524
  );


  and
  g2749
  (
    n2834,
    n1421,
    n2565,
    n2247,
    n2352
  );


  and
  g2750
  (
    n2673,
    n1006,
    n1090,
    n1424,
    n2561
  );


  nand
  g2751
  (
    n2629,
    n892,
    n2178,
    n1553,
    n2547
  );


  and
  g2752
  (
    n2781,
    n983,
    n1085,
    n1198,
    n1578
  );


  nor
  g2753
  (
    n2753,
    n1278,
    n1350,
    n1518,
    n2376
  );


  and
  g2754
  (
    n2874,
    n2284,
    n2172,
    n1059,
    n960
  );


  xnor
  g2755
  (
    n2878,
    n2216,
    n1369,
    n1599,
    n2463
  );


  and
  g2756
  (
    n2589,
    n1241,
    n1595,
    n1334,
    n2205
  );


  xor
  g2757
  (
    n2765,
    n1449,
    n2502,
    n2197,
    n2251
  );


  xnor
  g2758
  (
    n2866,
    n2540,
    n2208,
    n1010,
    n1650
  );


  xor
  g2759
  (
    n2641,
    n2340,
    n906,
    n1121,
    n1057
  );


  and
  g2760
  (
    n2593,
    n2491,
    n1418,
    n1323,
    n1670
  );


  xor
  g2761
  (
    n2609,
    n2374,
    n1473,
    n1485,
    n2488
  );


  or
  g2762
  (
    n2584,
    n1555,
    n2293,
    n995,
    n2409
  );


  nor
  g2763
  (
    n2728,
    n2466,
    n1232,
    n835,
    n1004
  );


  nor
  g2764
  (
    n2590,
    n2457,
    n2443,
    n846,
    n1141
  );


  xor
  g2765
  (
    n2783,
    n1618,
    n2290,
    n2333,
    n1412
  );


  nand
  g2766
  (
    n2827,
    n1083,
    n2157,
    n2525,
    n1199
  );


  xnor
  g2767
  (
    n2647,
    n1266,
    n1353,
    n2126,
    n2521
  );


  or
  g2768
  (
    n2819,
    n1182,
    n2429,
    n2158,
    n2383
  );


  nor
  g2769
  (
    n2870,
    n2215,
    n1015,
    n2198,
    n891
  );


  xnor
  g2770
  (
    n2689,
    n814,
    n811,
    n2531,
    n1227
  );


  nor
  g2771
  (
    n2774,
    n1646,
    n869,
    n2332,
    n2454
  );


  or
  g2772
  (
    n2863,
    n815,
    n1366,
    n1560,
    n2075
  );


  or
  g2773
  (
    n2794,
    n1596,
    n936,
    n1376,
    n1140
  );


  nor
  g2774
  (
    n2831,
    n1093,
    n949,
    n1568,
    n866
  );


  and
  g2775
  (
    n2620,
    n2128,
    n1631,
    n1547,
    n1124
  );


  and
  g2776
  (
    n2746,
    n856,
    n2396,
    n2331,
    n1295
  );


  and
  g2777
  (
    n2626,
    n2367,
    n1286,
    n2328,
    n2397
  );


  nor
  g2778
  (
    n2899,
    n1465,
    n1657,
    n1644,
    n831
  );


  xnor
  g2779
  (
    n2773,
    n1693,
    n994,
    n1368,
    n1043
  );


  nor
  g2780
  (
    n2760,
    n2460,
    n1267,
    n2339,
    n1138
  );


  xor
  g2781
  (
    n2895,
    n2496,
    n1028,
    n2330,
    n1257
  );


  xor
  g2782
  (
    n2650,
    n2203,
    n1268,
    n2375,
    n1477
  );


  or
  g2783
  (
    n2710,
    n2424,
    n971,
    n1374,
    n1558
  );


  nand
  g2784
  (
    n2810,
    n2513,
    n2142,
    n1396,
    n1223
  );


  xnor
  g2785
  (
    n2679,
    n2195,
    n913,
    n2194,
    n2127
  );


  xor
  g2786
  (
    n2769,
    n1594,
    n2353,
    n883,
    n1289
  );


  or
  g2787
  (
    n2817,
    n1622,
    n873,
    n1242,
    n2291
  );


  and
  g2788
  (
    n2891,
    n897,
    n2087,
    n2262,
    n1237
  );


  nand
  g2789
  (
    n2682,
    n2304,
    n2207,
    n1444,
    n2077
  );


  xnor
  g2790
  (
    n2608,
    n1339,
    n1234,
    n806,
    n2246
  );


  xor
  g2791
  (
    n2655,
    n813,
    n2377,
    n979,
    n1337
  );


  xor
  g2792
  (
    n2823,
    n1115,
    n1074,
    n1325,
    n2440
  );


  xor
  g2793
  (
    n2578,
    n967,
    n2541,
    n1196,
    n847
  );


  or
  g2794
  (
    n2807,
    n956,
    n1322,
    n1308,
    n2183
  );


  xor
  g2795
  (
    n2592,
    n2276,
    n876,
    n1469,
    n2108
  );


  and
  g2796
  (
    n2625,
    n1698,
    n1112,
    n2321,
    n2535
  );


  xnor
  g2797
  (
    n2835,
    n1564,
    n927,
    n2295,
    n2161
  );


  xnor
  g2798
  (
    n2723,
    n901,
    n2073,
    n1072,
    n1665
  );


  nor
  g2799
  (
    n2636,
    n2441,
    n1298,
    n2110,
    n1406
  );


  nand
  g2800
  (
    n2759,
    n2264,
    n1336,
    n1130,
    n2200
  );


  nor
  g2801
  (
    n2758,
    n1634,
    n1663,
    n1493,
    n1014
  );


  xnor
  g2802
  (
    n2640,
    n1269,
    n1134,
    n1572,
    n1304
  );


  nor
  g2803
  (
    n2786,
    n1439,
    n1629,
    n2244,
    n1380
  );


  nor
  g2804
  (
    n2638,
    n1546,
    n840,
    n2372,
    n1643
  );


  xnor
  g2805
  (
    n2777,
    n1446,
    n2129,
    n1528,
    n885
  );


  nand
  g2806
  (
    KeyWire_0_62,
    n2390,
    n1494,
    n2416,
    n1216
  );


  or
  g2807
  (
    n2805,
    n1677,
    n1003,
    n2308,
    n1228
  );


  and
  g2808
  (
    n2836,
    n986,
    n1127,
    n2556,
    n2162
  );


  nand
  g2809
  (
    n2917,
    n1627,
    n1050,
    n822,
    n2451
  );


  xor
  g2810
  (
    n2687,
    n1280,
    n1362,
    n1188,
    n1314
  );


  nor
  g2811
  (
    n2820,
    n1520,
    n1565,
    n1333,
    n2478
  );


  xor
  g2812
  (
    n2688,
    n2292,
    n2523,
    n1615,
    n2567
  );


  nor
  g2813
  (
    n2775,
    n1118,
    n942,
    n1249,
    n972
  );


  nor
  g2814
  (
    n2839,
    n2542,
    n1178,
    n1251,
    n1381
  );


  or
  g2815
  (
    n2825,
    n1087,
    n2384,
    n2529,
    n1364
  );


  xnor
  g2816
  (
    n2632,
    n1487,
    n1522,
    n2507,
    n946
  );


  nand
  g2817
  (
    n2767,
    n2102,
    n1039,
    n2479,
    n2492
  );


  xnor
  g2818
  (
    n2699,
    n1413,
    n817,
    n961,
    n925
  );


  nand
  g2819
  (
    n2908,
    n1256,
    n1099,
    n857,
    n1179
  );


  xnor
  g2820
  (
    n2914,
    n1208,
    n2517,
    n2503,
    n2085
  );


  nand
  g2821
  (
    n2872,
    n1345,
    n2467,
    n1402,
    n816
  );


  or
  g2822
  (
    n2911,
    n1261,
    n1161,
    n1388,
    n1166
  );


  nand
  g2823
  (
    n2601,
    n2334,
    n1061,
    n2288,
    n1425
  );


  or
  g2824
  (
    n2846,
    n1018,
    n1183,
    n2135,
    n2312
  );


  nor
  g2825
  (
    n2788,
    n2439,
    n1600,
    n944,
    n2184
  );


  xor
  g2826
  (
    n2850,
    n1347,
    n2266,
    n1026,
    n2106
  );


  nand
  g2827
  (
    n2855,
    n1497,
    n2549,
    n2300,
    n1142
  );


  and
  g2828
  (
    n2862,
    n1252,
    n1552,
    n2118,
    n1513
  );


  xnor
  g2829
  (
    n2903,
    n915,
    n1070,
    n1468,
    n2434
  );


  nor
  g2830
  (
    n2897,
    n2062,
    n2337,
    n1417,
    n1466
  );


  xor
  g2831
  (
    n2858,
    n930,
    n1604,
    n1263,
    n2359
  );


  xor
  g2832
  (
    n2808,
    n2101,
    n1567,
    n2354,
    n1590
  );


  nand
  g2833
  (
    n2859,
    n2271,
    n1512,
    n2393,
    n2530
  );


  nor
  g2834
  (
    n2661,
    n1538,
    n2097,
    n2514,
    n2080
  );


  or
  g2835
  (
    n2693,
    n1024,
    n1097,
    n1548,
    n2125
  );


  xor
  g2836
  (
    n2795,
    n948,
    n1504,
    n2394,
    n1448
  );


  nor
  g2837
  (
    n2718,
    n1160,
    n1189,
    n1029,
    n1293
  );


  nor
  g2838
  (
    n2875,
    n2419,
    n2234,
    n1537,
    n1603
  );


  nand
  g2839
  (
    n2670,
    n1001,
    n989,
    n1571,
    n2112
  );


  and
  g2840
  (
    n2826,
    n1324,
    n2560,
    n1040,
    n2148
  );


  and
  g2841
  (
    n2585,
    n2379,
    n829,
    n1151,
    n1423
  );


  nand
  g2842
  (
    n2634,
    n2269,
    n1372,
    n1023,
    n1215
  );


  or
  g2843
  (
    n2681,
    n2068,
    n1549,
    n918,
    n908
  );


  and
  g2844
  (
    n2906,
    n2465,
    n1239,
    n2171,
    n2512
  );


  xor
  g2845
  (
    n2580,
    n1056,
    n1007,
    n2170,
    n2402
  );


  nor
  g2846
  (
    KeyWire_0_43,
    n1610,
    n2191,
    n1426,
    n2074
  );


  nand
  g2847
  (
    n2779,
    n1623,
    n2493,
    n2105,
    n2220
  );


  or
  g2848
  (
    n2882,
    n2223,
    n914,
    n2070,
    n1524
  );


  or
  g2849
  (
    n2860,
    n1490,
    n1033,
    n1687,
    n887
  );


  nor
  g2850
  (
    n2635,
    n2555,
    n2100,
    n2320,
    n2413
  );


  xnor
  g2851
  (
    n2716,
    n1011,
    n951,
    n2563,
    n1529
  );


  nor
  g2852
  (
    n2582,
    n1254,
    n2433,
    n1668,
    n1082
  );


  nor
  g2853
  (
    n2885,
    n1391,
    n1122,
    n2362,
    n1131
  );


  nor
  g2854
  (
    n2711,
    n1664,
    n1419,
    n1319,
    n1686
  );


  nor
  g2855
  (
    n2837,
    n976,
    n1167,
    n808,
    n1363
  );


  or
  g2856
  (
    n2893,
    n950,
    n2338,
    n904,
    n962
  );


  xnor
  g2857
  (
    n2791,
    n1598,
    n1432,
    n1354,
    n1625
  );


  nand
  g2858
  (
    n2747,
    n2212,
    n2082,
    n2559,
    n1144
  );


  nor
  g2859
  (
    n2703,
    n2254,
    n952,
    n2472,
    n1328
  );


  xor
  g2860
  (
    n2761,
    n2426,
    n2227,
    n2218,
    n1013
  );


  or
  g2861
  (
    n2741,
    n1450,
    n842,
    n809,
    n2113
  );


  xnor
  g2862
  (
    n2630,
    n1321,
    n2484,
    n1340,
    n1545
  );


  nor
  g2863
  (
    n2597,
    n2545,
    n1582,
    n1445,
    n2167
  );


  nand
  g2864
  (
    n2770,
    n2190,
    n1017,
    n1275,
    n2282
  );


  xnor
  g2865
  (
    n2617,
    n1020,
    n2084,
    n1200,
    n2226
  );


  and
  g2866
  (
    n2811,
    n1491,
    n1348,
    n922,
    n826
  );


  xor
  g2867
  (
    n2619,
    n827,
    n850,
    n1117,
    n1262
  );


  nor
  g2868
  (
    n2684,
    n2329,
    n2497,
    n1316,
    n1628
  );


  xnor
  g2869
  (
    n2675,
    n2351,
    n2160,
    n1092,
    n2446
  );


  and
  g2870
  (
    n2696,
    n1100,
    n1084,
    n1238,
    n2253
  );


  or
  g2871
  (
    n2712,
    n2061,
    n1058,
    n1427,
    n1302
  );


  xor
  g2872
  (
    n2678,
    n2088,
    n1294,
    n1303,
    n1230
  );


  nand
  g2873
  (
    n2776,
    n1283,
    n2425,
    n2265,
    n1102
  );


  nand
  g2874
  (
    n2637,
    n1542,
    n1022,
    n1111,
    n2526
  );


  and
  g2875
  (
    n2618,
    n2094,
    n2120,
    n1073,
    n2237
  );


  nand
  g2876
  (
    n2586,
    n2505,
    n2369,
    n1394,
    n2076
  );


  nor
  g2877
  (
    n2733,
    n2566,
    n973,
    n1489,
    n1475
  );


  xnor
  g2878
  (
    n2669,
    n2163,
    n1240,
    n1656,
    n1312
  );


  xnor
  g2879
  (
    n2709,
    n1148,
    n2420,
    n2302,
    n893
  );


  xor
  g2880
  (
    n2581,
    n1292,
    n1035,
    n2121,
    n849
  );


  nor
  g2881
  (
    n2698,
    n2345,
    n947,
    n2398,
    n1143
  );


  xor
  g2882
  (
    n2806,
    n982,
    n1556,
    n2485,
    n1658
  );


  nand
  g2883
  (
    n2667,
    n2164,
    n1145,
    n2537,
    n1414
  );


  xnor
  g2884
  (
    n2631,
    n823,
    n932,
    n2289,
    n2196
  );


  and
  g2885
  (
    n2892,
    n996,
    n867,
    n1403,
    n2569
  );


  and
  g2886
  (
    n2756,
    n900,
    n1367,
    n1684,
    n997
  );


  xor
  g2887
  (
    n2802,
    n2179,
    n2498,
    n1244,
    n1071
  );


  nand
  g2888
  (
    n2793,
    n1640,
    n2356,
    n1577,
    n2548
  );


  xor
  g2889
  (
    n2852,
    n880,
    n2139,
    n1331,
    n1054
  );


  or
  g2890
  (
    n2993,
    n2818,
    n2820,
    n2608,
    n2641
  );


  nand
  g2891
  (
    n3000,
    n2634,
    n2711,
    n2830,
    n2823
  );


  nand
  g2892
  (
    n2940,
    n2601,
    n2784,
    n2579,
    n2593
  );


  and
  g2893
  (
    n2958,
    n2875,
    n2620,
    n2745,
    n2714
  );


  or
  g2894
  (
    n2994,
    n2598,
    n2886,
    n2746,
    n2873
  );


  nand
  g2895
  (
    n2995,
    n2864,
    n2572,
    n2616,
    n2670
  );


  xnor
  g2896
  (
    n3009,
    n2907,
    n2898,
    n2910,
    n2644
  );


  and
  g2897
  (
    n2968,
    n2607,
    n2840,
    n2815,
    n2887
  );


  nor
  g2898
  (
    n2972,
    n2787,
    n2854,
    n2643,
    n2869
  );


  nor
  g2899
  (
    n2946,
    n2624,
    n2770,
    n2871,
    n2651
  );


  xor
  g2900
  (
    n2929,
    n2668,
    n2636,
    n2577,
    n2780
  );


  and
  g2901
  (
    n2979,
    n2621,
    n2847,
    n2719,
    n2680
  );


  xor
  g2902
  (
    n2983,
    n2759,
    n2891,
    n2747,
    n2656
  );


  xnor
  g2903
  (
    n2988,
    n2908,
    n2816,
    n2631,
    n2900
  );


  xnor
  g2904
  (
    n2938,
    n2799,
    n2674,
    n2715,
    n2896
  );


  or
  g2905
  (
    n3003,
    n2622,
    n2742,
    n2732,
    n2739
  );


  or
  g2906
  (
    n2975,
    n2673,
    n2612,
    n2657,
    n2812
  );


  xor
  g2907
  (
    n3004,
    n2689,
    n2748,
    n2588,
    n2669
  );


  and
  g2908
  (
    n2931,
    n2790,
    n2626,
    n2755,
    n2913
  );


  nand
  g2909
  (
    n2982,
    n2623,
    n2785,
    n2709,
    n2817
  );


  nand
  g2910
  (
    n2943,
    n2663,
    n2632,
    n2629,
    n2918
  );


  xnor
  g2911
  (
    n2973,
    n2686,
    n2852,
    n2591,
    n2822
  );


  xnor
  g2912
  (
    n2930,
    n2850,
    n2844,
    n2602,
    n2861
  );


  nor
  g2913
  (
    n2996,
    n2839,
    n2633,
    n2849,
    n2723
  );


  or
  g2914
  (
    n2962,
    n2700,
    n2571,
    n2863,
    n2718
  );


  xor
  g2915
  (
    n2927,
    n2792,
    n2738,
    n2888,
    n2605
  );


  and
  g2916
  (
    n2992,
    n2772,
    n2776,
    n2862,
    n2685
  );


  xor
  g2917
  (
    n2936,
    n2843,
    n2660,
    n2574,
    n2857
  );


  nor
  g2918
  (
    n2990,
    n2791,
    n2826,
    n2800,
    n2694
  );


  nor
  g2919
  (
    n2956,
    n2858,
    n2824,
    n2777,
    n2675
  );


  or
  g2920
  (
    n3007,
    n2740,
    n2583,
    n2582,
    n2892
  );


  nor
  g2921
  (
    n2977,
    n2690,
    n2769,
    n2684,
    n2754
  );


  nor
  g2922
  (
    n2937,
    n2774,
    n2614,
    n2771,
    n2665
  );


  nand
  g2923
  (
    n3002,
    n2894,
    n2883,
    n2695,
    n2609
  );


  xnor
  g2924
  (
    n2967,
    n2735,
    n2828,
    n2835,
    n2842
  );


  nand
  g2925
  (
    n2966,
    n2794,
    n2726,
    n2576,
    n2806
  );


  nand
  g2926
  (
    n2953,
    n2678,
    n2751,
    n2646,
    n2741
  );


  and
  g2927
  (
    n2997,
    n2731,
    n2595,
    n2859,
    n2586
  );


  and
  g2928
  (
    n2941,
    n2724,
    n2833,
    n2692,
    n2615
  );


  xor
  g2929
  (
    KeyWire_0_42,
    n2763,
    n2821,
    n2807,
    n2637
  );


  and
  g2930
  (
    n2924,
    n2855,
    n2902,
    n2672,
    n2808
  );


  nand
  g2931
  (
    n2999,
    n2903,
    n2736,
    n2650,
    n2853
  );


  and
  g2932
  (
    n2978,
    n2762,
    n2728,
    n2878,
    n2897
  );


  or
  g2933
  (
    n3006,
    n2676,
    n2890,
    n2638,
    n2645
  );


  or
  g2934
  (
    n2942,
    n2640,
    n2720,
    n2885,
    n2836
  );


  or
  g2935
  (
    n2964,
    n2596,
    n2677,
    n2846,
    n2912
  );


  nand
  g2936
  (
    n2926,
    n2805,
    n2617,
    n2721,
    n2834
  );


  and
  g2937
  (
    n2947,
    n2659,
    n2837,
    n2851,
    n2716
  );


  xnor
  g2938
  (
    n2969,
    n2838,
    n2809,
    n2793,
    n2813
  );


  and
  g2939
  (
    n2985,
    n2671,
    n2703,
    n2693,
    n2688
  );


  nor
  g2940
  (
    n2952,
    n2635,
    n2639,
    n2810,
    n2647
  );


  or
  g2941
  (
    n2981,
    n2662,
    n2919,
    n2604,
    n2893
  );


  xor
  g2942
  (
    n2976,
    n2752,
    n2722,
    n2921,
    n2750
  );


  xor
  g2943
  (
    n2948,
    n2687,
    n2845,
    n2712,
    n2882
  );


  nand
  g2944
  (
    n2934,
    n2920,
    n2814,
    n2899,
    n2917
  );


  nand
  g2945
  (
    n2971,
    n2867,
    n2655,
    n2827,
    n2679
  );


  or
  g2946
  (
    n2974,
    n2743,
    n2877,
    n2901,
    n2915
  );


  and
  g2947
  (
    n2932,
    n2765,
    n2611,
    n2707,
    n2653
  );


  nand
  g2948
  (
    n2957,
    n2613,
    n2879,
    n2801,
    n2603
  );


  or
  g2949
  (
    n2987,
    n2737,
    n2768,
    n2708,
    n2578
  );


  xnor
  g2950
  (
    n2980,
    n2592,
    n2895,
    n2832,
    n2804
  );


  nor
  g2951
  (
    n2954,
    n2764,
    n2666,
    n2581,
    n2597
  );


  and
  g2952
  (
    n2961,
    n2701,
    n2865,
    n2795,
    n2696
  );


  or
  g2953
  (
    n2950,
    n2773,
    n2905,
    n2627,
    n2819
  );


  nand
  g2954
  (
    n2949,
    n2756,
    n2649,
    n2587,
    n2642
  );


  or
  g2955
  (
    n2963,
    n2757,
    n2667,
    n2691,
    n2734
  );


  xor
  g2956
  (
    n2944,
    n2625,
    n2652,
    n2802,
    n2786
  );


  nand
  g2957
  (
    n2991,
    n2749,
    n2585,
    n2904,
    n2580
  );


  or
  g2958
  (
    n2955,
    n2761,
    n2658,
    n2648,
    n2848
  );


  xnor
  g2959
  (
    KeyWire_0_18,
    n2775,
    n2906,
    n2767,
    n2758
  );


  or
  g2960
  (
    n3008,
    n2618,
    n2872,
    n2706,
    n2841
  );


  xor
  g2961
  (
    n2951,
    n2781,
    n2916,
    n2699,
    n2702
  );


  and
  g2962
  (
    n3005,
    n2874,
    n2600,
    n2884,
    n2876
  );


  and
  g2963
  (
    n3001,
    n2911,
    n2778,
    n2594,
    n2914
  );


  nand
  g2964
  (
    n2923,
    n2730,
    n2766,
    n2881,
    n2796
  );


  or
  g2965
  (
    n2933,
    n2681,
    n2573,
    n2798,
    n2630
  );


  or
  g2966
  (
    n2989,
    n2661,
    n2783,
    n2704,
    n2705
  );


  or
  g2967
  (
    n2925,
    n2788,
    n2825,
    n2599,
    n2698
  );


  or
  g2968
  (
    n2960,
    n2683,
    n2831,
    n2811,
    n2619
  );


  nor
  g2969
  (
    n2984,
    n2589,
    n2779,
    n2654,
    n2880
  );


  or
  g2970
  (
    n2928,
    n2789,
    n2610,
    n2664,
    n2729
  );


  xnor
  g2971
  (
    n2965,
    n2803,
    n2725,
    n2797,
    n2713
  );


  nand
  g2972
  (
    n2986,
    n2860,
    n2760,
    n2866,
    n2682
  );


  xor
  g2973
  (
    n2939,
    n2889,
    n2829,
    n2717,
    n2606
  );


  and
  g2974
  (
    n2998,
    n2782,
    n2744,
    n2590,
    n2870
  );


  xnor
  g2975
  (
    n2945,
    n2733,
    n2575,
    n2727,
    n2710
  );


  nor
  g2976
  (
    n2959,
    n2697,
    n2868,
    n2856,
    n2584
  );


  and
  g2977
  (
    n3010,
    n2628,
    n2922,
    n2753,
    n2909
  );


  xor
  g2978
  (
    n3025,
    n2959,
    n2943,
    n2991,
    n2987
  );


  or
  g2979
  (
    n3028,
    n2923,
    n2955,
    n2990,
    n2979
  );


  nand
  g2980
  (
    n3031,
    n2984,
    n2958,
    n3001,
    n2933
  );


  nand
  g2981
  (
    n3027,
    n2983,
    n2946,
    n3002,
    n2945
  );


  or
  g2982
  (
    n3019,
    n2978,
    n2992,
    n2981,
    n2962
  );


  nor
  g2983
  (
    n3018,
    n2932,
    n2977,
    n2973,
    n2942
  );


  nand
  g2984
  (
    n3017,
    n2956,
    n2985,
    n2976,
    n2940
  );


  or
  g2985
  (
    n3021,
    n2998,
    n2937,
    n3008,
    n2952
  );


  and
  g2986
  (
    n3023,
    n2927,
    n3004,
    n2989,
    n2953
  );


  xor
  g2987
  (
    n3032,
    n2938,
    n2997,
    n2965,
    n2934
  );


  nor
  g2988
  (
    n3030,
    n2960,
    n3003,
    n2986,
    n2929
  );


  nor
  g2989
  (
    n3022,
    n2924,
    n2926,
    n3009,
    n3000
  );


  nand
  g2990
  (
    n3029,
    n2925,
    n3010,
    n2974,
    n2963
  );


  nor
  g2991
  (
    n3016,
    n2948,
    n2950,
    n2996,
    n3006
  );


  xnor
  g2992
  (
    n3015,
    n2964,
    n2951,
    n2954,
    n2930
  );


  xnor
  g2993
  (
    n3012,
    n2972,
    n2971,
    n2936,
    n3007
  );


  nand
  g2994
  (
    n3020,
    n3005,
    n2939,
    n2999,
    n2995
  );


  xor
  g2995
  (
    n3014,
    n2988,
    n2928,
    n2931,
    n2957
  );


  xnor
  g2996
  (
    n3024,
    n2980,
    n2993,
    n2994,
    n2947
  );


  nand
  g2997
  (
    n3013,
    n2935,
    n2969,
    n2982,
    n2968
  );


  xor
  g2998
  (
    KeyWire_0_63,
    n2970,
    n2961,
    n2966,
    n2967
  );


  xor
  g2999
  (
    n3011,
    n2944,
    n2949,
    n2975,
    n2941
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1157,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n312,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n2261,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1660,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n2168,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1897,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n2648,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1282,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n238,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n216,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n617,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n515,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1536,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1116,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1139,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n2547,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1511,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1355,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n2970,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1425,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n2352,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1581,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n527,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n2611,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n64,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n1145,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n2536,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1957,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1498,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n2432,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n600,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n762,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n780,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n2013,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n2349,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n2054,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n1522,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n198,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n2440,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n338,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n777,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n1685,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n2935,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n2615,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n1391,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n854,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n2751,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n1549,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1421,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n1306,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n1233,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n1502,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n2256,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1505,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n1208,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n2520,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n776,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n498,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n2292,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n1973,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n666,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n1472,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n2732,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n3026,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


