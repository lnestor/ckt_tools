

module Stat_1000_104
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n731,
  n623,
  n637,
  n649,
  n677,
  n718,
  n675,
  n616,
  n668,
  n707,
  n643,
  n626,
  n701,
  n625,
  n735,
  n681,
  n627,
  n1022,
  n1020,
  n1019,
  n1031,
  n1026,
  n1029,
  n1023,
  n1021,
  n1024,
  n1025,
  n1027,
  n1030,
  n1028,
  n1018,
  n1032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n731;
  output n623;
  output n637;
  output n649;
  output n677;
  output n718;
  output n675;
  output n616;
  output n668;
  output n707;
  output n643;
  output n626;
  output n701;
  output n625;
  output n735;
  output n681;
  output n627;
  output n1022;
  output n1020;
  output n1019;
  output n1031;
  output n1026;
  output n1029;
  output n1023;
  output n1021;
  output n1024;
  output n1025;
  output n1027;
  output n1030;
  output n1028;
  output n1018;
  output n1032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n624;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n676;
  wire n678;
  wire n679;
  wire n680;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n732;
  wire n733;
  wire n734;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n158,
    n30
  );


  not
  g1
  (
    n71,
    n16
  );


  buf
  g2
  (
    n147,
    n11
  );


  buf
  g3
  (
    n101,
    n22
  );


  not
  g4
  (
    n96,
    n22
  );


  not
  g5
  (
    KeyWire_0_2,
    n29
  );


  buf
  g6
  (
    n159,
    n27
  );


  buf
  g7
  (
    n37,
    n10
  );


  buf
  g8
  (
    n126,
    n10
  );


  buf
  g9
  (
    KeyWire_0_56,
    n4
  );


  not
  g10
  (
    n120,
    n27
  );


  buf
  g11
  (
    n152,
    n32
  );


  not
  g12
  (
    n47,
    n23
  );


  not
  g13
  (
    n41,
    n8
  );


  buf
  g14
  (
    n110,
    n24
  );


  not
  g15
  (
    n90,
    n13
  );


  buf
  g16
  (
    n72,
    n5
  );


  buf
  g17
  (
    n99,
    n1
  );


  not
  g18
  (
    n69,
    n25
  );


  not
  g19
  (
    n145,
    n26
  );


  buf
  g20
  (
    KeyWire_0_35,
    n1
  );


  buf
  g21
  (
    n98,
    n25
  );


  not
  g22
  (
    n60,
    n6
  );


  not
  g23
  (
    n116,
    n3
  );


  buf
  g24
  (
    n92,
    n18
  );


  buf
  g25
  (
    n82,
    n28
  );


  not
  g26
  (
    KeyWire_0_58,
    n8
  );


  buf
  g27
  (
    n49,
    n12
  );


  buf
  g28
  (
    n61,
    n15
  );


  buf
  g29
  (
    n132,
    n14
  );


  not
  g30
  (
    n58,
    n16
  );


  buf
  g31
  (
    n67,
    n21
  );


  buf
  g32
  (
    n106,
    n21
  );


  buf
  g33
  (
    KeyWire_0_3,
    n6
  );


  not
  g34
  (
    n140,
    n15
  );


  buf
  g35
  (
    n93,
    n19
  );


  not
  g36
  (
    n121,
    n17
  );


  not
  g37
  (
    n64,
    n13
  );


  not
  g38
  (
    n115,
    n18
  );


  not
  g39
  (
    n130,
    n20
  );


  buf
  g40
  (
    n112,
    n5
  );


  buf
  g41
  (
    n76,
    n28
  );


  not
  g42
  (
    n156,
    n7
  );


  buf
  g43
  (
    n89,
    n26
  );


  buf
  g44
  (
    n87,
    n7
  );


  buf
  g45
  (
    n46,
    n26
  );


  buf
  g46
  (
    n77,
    n4
  );


  buf
  g47
  (
    n33,
    n14
  );


  buf
  g48
  (
    n80,
    n18
  );


  not
  g49
  (
    n151,
    n32
  );


  buf
  g50
  (
    n108,
    n31
  );


  buf
  g51
  (
    n52,
    n11
  );


  not
  g52
  (
    n48,
    n17
  );


  not
  g53
  (
    n36,
    n26
  );


  buf
  g54
  (
    n128,
    n12
  );


  not
  g55
  (
    n65,
    n20
  );


  not
  g56
  (
    n119,
    n15
  );


  buf
  g57
  (
    n102,
    n7
  );


  buf
  g58
  (
    n153,
    n12
  );


  buf
  g59
  (
    n134,
    n2
  );


  not
  g60
  (
    n114,
    n7
  );


  buf
  g61
  (
    n40,
    n1
  );


  buf
  g62
  (
    n94,
    n20
  );


  buf
  g63
  (
    n74,
    n19
  );


  buf
  g64
  (
    n63,
    n24
  );


  not
  g65
  (
    n154,
    n31
  );


  buf
  g66
  (
    n38,
    n25
  );


  buf
  g67
  (
    n43,
    n15
  );


  not
  g68
  (
    KeyWire_0_19,
    n11
  );


  not
  g69
  (
    n113,
    n22
  );


  not
  g70
  (
    n42,
    n21
  );


  buf
  g71
  (
    n44,
    n10
  );


  not
  g72
  (
    n133,
    n8
  );


  not
  g73
  (
    n143,
    n30
  );


  buf
  g74
  (
    n85,
    n31
  );


  not
  g75
  (
    n45,
    n27
  );


  buf
  g76
  (
    n81,
    n16
  );


  buf
  g77
  (
    n57,
    n3
  );


  not
  g78
  (
    n104,
    n4
  );


  buf
  g79
  (
    n111,
    n24
  );


  not
  g80
  (
    n95,
    n14
  );


  buf
  g81
  (
    n68,
    n19
  );


  buf
  g82
  (
    n124,
    n30
  );


  buf
  g83
  (
    n34,
    n17
  );


  buf
  g84
  (
    n100,
    n9
  );


  not
  g85
  (
    n105,
    n28
  );


  not
  g86
  (
    n123,
    n29
  );


  not
  g87
  (
    n53,
    n29
  );


  buf
  g88
  (
    n39,
    n23
  );


  buf
  g89
  (
    n139,
    n1
  );


  buf
  g90
  (
    n125,
    n13
  );


  buf
  g91
  (
    n160,
    n3
  );


  not
  g92
  (
    n131,
    n21
  );


  buf
  g93
  (
    n97,
    n22
  );


  buf
  g94
  (
    n122,
    n4
  );


  buf
  g95
  (
    n138,
    n32
  );


  not
  g96
  (
    n127,
    n23
  );


  buf
  g97
  (
    n84,
    n14
  );


  buf
  g98
  (
    n51,
    n27
  );


  buf
  g99
  (
    n117,
    n3
  );


  not
  g100
  (
    n146,
    n6
  );


  buf
  g101
  (
    n149,
    n5
  );


  buf
  g102
  (
    n141,
    n2
  );


  buf
  g103
  (
    n135,
    n10
  );


  buf
  g104
  (
    n83,
    n20
  );


  buf
  g105
  (
    n142,
    n9
  );


  buf
  g106
  (
    n78,
    n28
  );


  buf
  g107
  (
    n75,
    n12
  );


  not
  g108
  (
    n88,
    n16
  );


  buf
  g109
  (
    n54,
    n29
  );


  not
  g110
  (
    n109,
    n31
  );


  not
  g111
  (
    n155,
    n2
  );


  buf
  g112
  (
    n148,
    n9
  );


  not
  g113
  (
    n86,
    n8
  );


  buf
  g114
  (
    n66,
    n11
  );


  buf
  g115
  (
    n118,
    n19
  );


  buf
  g116
  (
    n137,
    n18
  );


  not
  g117
  (
    n91,
    n9
  );


  not
  g118
  (
    n103,
    n17
  );


  buf
  g119
  (
    n70,
    n5
  );


  not
  g120
  (
    n129,
    n32
  );


  not
  g121
  (
    n56,
    n23
  );


  buf
  g122
  (
    n107,
    n2
  );


  not
  g123
  (
    n62,
    n13
  );


  buf
  g124
  (
    n79,
    n30
  );


  not
  g125
  (
    KeyWire_0_33,
    n24
  );


  buf
  g126
  (
    n50,
    n25
  );


  not
  g127
  (
    KeyWire_0_14,
    n6
  );


  xor
  g128
  (
    n273,
    n112,
    n82
  );


  xor
  g129
  (
    n274,
    n115,
    n33
  );


  and
  g130
  (
    n300,
    n83,
    n112
  );


  nor
  g131
  (
    n180,
    n99,
    n41
  );


  or
  g132
  (
    n250,
    n52,
    n38
  );


  nand
  g133
  (
    n181,
    n80,
    n77
  );


  nand
  g134
  (
    n230,
    n46,
    n114
  );


  and
  g135
  (
    n276,
    n52,
    n90
  );


  xnor
  g136
  (
    n196,
    n62,
    n94
  );


  or
  g137
  (
    n182,
    n56,
    n62
  );


  and
  g138
  (
    n167,
    n84,
    n91
  );


  and
  g139
  (
    n322,
    n60,
    n56
  );


  and
  g140
  (
    n177,
    n82,
    n47
  );


  nand
  g141
  (
    n261,
    n122,
    n98
  );


  xor
  g142
  (
    n166,
    n63,
    n50
  );


  or
  g143
  (
    n169,
    n124,
    n115
  );


  xor
  g144
  (
    n236,
    n87,
    n111
  );


  nand
  g145
  (
    n282,
    n100,
    n77
  );


  nand
  g146
  (
    n279,
    n33,
    n106
  );


  and
  g147
  (
    n227,
    n60,
    n52
  );


  or
  g148
  (
    n268,
    n44,
    n106
  );


  and
  g149
  (
    n319,
    n65,
    n104
  );


  xnor
  g150
  (
    n259,
    n126,
    n46
  );


  nor
  g151
  (
    n294,
    n81,
    n55
  );


  nor
  g152
  (
    n246,
    n57,
    n118
  );


  xor
  g153
  (
    n321,
    n86,
    n65
  );


  and
  g154
  (
    n216,
    n35,
    n67
  );


  nor
  g155
  (
    n314,
    n43,
    n58
  );


  nor
  g156
  (
    n299,
    n71,
    n103
  );


  and
  g157
  (
    n239,
    n70,
    n117
  );


  or
  g158
  (
    n281,
    n72,
    n94
  );


  and
  g159
  (
    n188,
    n89,
    n94
  );


  xnor
  g160
  (
    n211,
    n47,
    n41
  );


  nand
  g161
  (
    n218,
    n71,
    n74
  );


  and
  g162
  (
    n286,
    n87,
    n69
  );


  xnor
  g163
  (
    n215,
    n86,
    n57
  );


  nand
  g164
  (
    n290,
    n104,
    n46
  );


  or
  g165
  (
    n317,
    n39,
    n93
  );


  nor
  g166
  (
    KeyWire_0_24,
    n108,
    n81
  );


  nand
  g167
  (
    n219,
    n107,
    n44
  );


  and
  g168
  (
    n187,
    n39,
    n91
  );


  nand
  g169
  (
    n285,
    n61,
    n92
  );


  or
  g170
  (
    n217,
    n105,
    n107
  );


  and
  g171
  (
    n208,
    n117,
    n44
  );


  nand
  g172
  (
    n309,
    n86,
    n97
  );


  or
  g173
  (
    n170,
    n85,
    n114
  );


  or
  g174
  (
    n249,
    n92,
    n45
  );


  xor
  g175
  (
    n207,
    n48,
    n106
  );


  xnor
  g176
  (
    n256,
    n73,
    n60
  );


  nand
  g177
  (
    n210,
    n122,
    n40
  );


  nand
  g178
  (
    KeyWire_0_44,
    n75,
    n123
  );


  or
  g179
  (
    KeyWire_0_21,
    n68,
    n85
  );


  xor
  g180
  (
    n292,
    n37,
    n80
  );


  xor
  g181
  (
    n265,
    n117,
    n85
  );


  xor
  g182
  (
    n229,
    n73,
    n113
  );


  nand
  g183
  (
    n185,
    n96,
    n121
  );


  or
  g184
  (
    n209,
    n63,
    n114
  );


  and
  g185
  (
    n260,
    n45,
    n102
  );


  xor
  g186
  (
    n289,
    n93,
    n111
  );


  xnor
  g187
  (
    n320,
    n110,
    n72
  );


  xnor
  g188
  (
    n164,
    n72,
    n71
  );


  xnor
  g189
  (
    n168,
    n88,
    n89
  );


  xnor
  g190
  (
    n172,
    n110,
    n34
  );


  nand
  g191
  (
    n226,
    n72,
    n52
  );


  and
  g192
  (
    n306,
    n78,
    n67
  );


  nor
  g193
  (
    n315,
    n42,
    n113
  );


  xnor
  g194
  (
    n271,
    n42,
    n57
  );


  nand
  g195
  (
    n162,
    n101,
    n125
  );


  or
  g196
  (
    KeyWire_0_40,
    n119,
    n122
  );


  or
  g197
  (
    n225,
    n63,
    n100
  );


  xor
  g198
  (
    n310,
    n83,
    n89
  );


  xnor
  g199
  (
    n194,
    n109,
    n83
  );


  nand
  g200
  (
    n221,
    n62,
    n86
  );


  xor
  g201
  (
    n288,
    n74,
    n63
  );


  or
  g202
  (
    n308,
    n88,
    n110
  );


  xor
  g203
  (
    n203,
    n34,
    n67
  );


  xnor
  g204
  (
    n272,
    n61,
    n59
  );


  and
  g205
  (
    n243,
    n121,
    n119
  );


  and
  g206
  (
    n312,
    n36,
    n74
  );


  and
  g207
  (
    n264,
    n123,
    n57
  );


  xor
  g208
  (
    n206,
    n68,
    n116
  );


  or
  g209
  (
    n298,
    n76,
    n98
  );


  xnor
  g210
  (
    n220,
    n101,
    n118
  );


  and
  g211
  (
    KeyWire_0_60,
    n45,
    n41
  );


  and
  g212
  (
    n176,
    n125,
    n45
  );


  xor
  g213
  (
    n174,
    n40,
    n125
  );


  and
  g214
  (
    n305,
    n46,
    n98
  );


  xor
  g215
  (
    n235,
    n40,
    n64
  );


  nor
  g216
  (
    n200,
    n53,
    n66
  );


  xor
  g217
  (
    n269,
    n58,
    n109
  );


  nand
  g218
  (
    n171,
    n38,
    n74
  );


  or
  g219
  (
    n297,
    n82,
    n33
  );


  and
  g220
  (
    n247,
    n102,
    n69
  );


  and
  g221
  (
    n237,
    n107,
    n34
  );


  xor
  g222
  (
    n313,
    n95,
    n55
  );


  and
  g223
  (
    n301,
    n61,
    n38
  );


  nor
  g224
  (
    KeyWire_0_10,
    n96,
    n61
  );


  nand
  g225
  (
    n280,
    n59,
    n44
  );


  and
  g226
  (
    n202,
    n66,
    n64
  );


  xnor
  g227
  (
    n253,
    n114,
    n65
  );


  nor
  g228
  (
    n192,
    n39,
    n43
  );


  and
  g229
  (
    n223,
    n37,
    n64
  );


  and
  g230
  (
    n296,
    n104,
    n91
  );


  xor
  g231
  (
    n233,
    n49,
    n108
  );


  xnor
  g232
  (
    n284,
    n73,
    n106
  );


  xnor
  g233
  (
    n163,
    n35,
    n78
  );


  nor
  g234
  (
    n267,
    n59,
    n81
  );


  xor
  g235
  (
    n193,
    n101,
    n113
  );


  nand
  g236
  (
    n303,
    n121,
    n105
  );


  xor
  g237
  (
    n183,
    n84,
    n108
  );


  xnor
  g238
  (
    n266,
    n124,
    n66
  );


  and
  g239
  (
    n302,
    n68,
    n54
  );


  or
  g240
  (
    n191,
    n89,
    n95
  );


  nor
  g241
  (
    n198,
    n53,
    n40
  );


  xnor
  g242
  (
    n224,
    n116,
    n124
  );


  and
  g243
  (
    KeyWire_0_63,
    n69,
    n97
  );


  and
  g244
  (
    n287,
    n48,
    n92
  );


  nor
  g245
  (
    n242,
    n112,
    n75
  );


  nand
  g246
  (
    KeyWire_0_17,
    n85,
    n33
  );


  nand
  g247
  (
    n254,
    n79,
    n120
  );


  xor
  g248
  (
    n234,
    n87,
    n35
  );


  and
  g249
  (
    n190,
    n119,
    n51
  );


  xor
  g250
  (
    n318,
    n94,
    n104
  );


  nand
  g251
  (
    n255,
    n93,
    n109
  );


  or
  g252
  (
    KeyWire_0_47,
    n103,
    n49
  );


  xor
  g253
  (
    n197,
    n43,
    n41
  );


  or
  g254
  (
    n204,
    n116,
    n69
  );


  nand
  g255
  (
    n252,
    n111,
    n48
  );


  or
  g256
  (
    KeyWire_0_25,
    n77,
    n103
  );


  and
  g257
  (
    n304,
    n53,
    n97
  );


  and
  g258
  (
    KeyWire_0_23,
    n36,
    n120
  );


  nor
  g259
  (
    n195,
    n120,
    n77
  );


  and
  g260
  (
    n175,
    n98,
    n67
  );


  nor
  g261
  (
    n248,
    n96,
    n124
  );


  xor
  g262
  (
    n283,
    n60,
    n113
  );


  xnor
  g263
  (
    n173,
    n62,
    n50
  );


  and
  g264
  (
    n311,
    n56,
    n108
  );


  nor
  g265
  (
    n228,
    n64,
    n51
  );


  xor
  g266
  (
    n245,
    n95,
    n37
  );


  or
  g267
  (
    n258,
    n120,
    n88
  );


  nor
  g268
  (
    n324,
    n102,
    n79
  );


  xor
  g269
  (
    n232,
    n42,
    n107,
    n80
  );


  xnor
  g270
  (
    n275,
    n58,
    n122,
    n79,
    n84
  );


  nand
  g271
  (
    n295,
    n118,
    n79,
    n73,
    n65
  );


  xnor
  g272
  (
    n244,
    n84,
    n78,
    n93,
    n54
  );


  nor
  g273
  (
    n316,
    n123,
    n119,
    n95,
    n101
  );


  xnor
  g274
  (
    n205,
    n103,
    n97,
    n105,
    n70
  );


  xor
  g275
  (
    n186,
    n111,
    n88,
    n109,
    n55
  );


  nor
  g276
  (
    n291,
    n49,
    n58,
    n75,
    n71
  );


  and
  g277
  (
    n257,
    n48,
    n91,
    n110,
    n121
  );


  and
  g278
  (
    KeyWire_0_8,
    n70,
    n117,
    n99,
    n76
  );


  or
  g279
  (
    n213,
    n80,
    n116,
    n87,
    n105
  );


  xor
  g280
  (
    n212,
    n100,
    n54,
    n112,
    n102
  );


  nor
  g281
  (
    n278,
    n56,
    n82,
    n38,
    n118
  );


  xnor
  g282
  (
    n323,
    n90,
    n99,
    n34,
    n75
  );


  xnor
  g283
  (
    n231,
    n83,
    n37,
    n81,
    n59
  );


  and
  g284
  (
    n165,
    n96,
    n70,
    n76,
    n55
  );


  xnor
  g285
  (
    n222,
    n68,
    n125,
    n76,
    n54
  );


  and
  g286
  (
    n178,
    n50,
    n115,
    n123,
    n92
  );


  nand
  g287
  (
    n270,
    n47,
    n42,
    n39,
    n90
  );


  nand
  g288
  (
    n161,
    n90,
    n49,
    n66,
    n36
  );


  or
  g289
  (
    n184,
    n36,
    n115,
    n43,
    n99
  );


  or
  g290
  (
    n251,
    n47,
    n78,
    n51,
    n100
  );


  and
  g291
  (
    n263,
    n35,
    n50,
    n53,
    n51
  );


  not
  g292
  (
    n378,
    n273
  );


  not
  g293
  (
    n463,
    n191
  );


  buf
  g294
  (
    n487,
    n296
  );


  buf
  g295
  (
    n349,
    n224
  );


  not
  g296
  (
    n453,
    n240
  );


  not
  g297
  (
    n383,
    n201
  );


  buf
  g298
  (
    n471,
    n182
  );


  not
  g299
  (
    n454,
    n209
  );


  not
  g300
  (
    n413,
    n278
  );


  not
  g301
  (
    n426,
    n181
  );


  not
  g302
  (
    n470,
    n288
  );


  not
  g303
  (
    n412,
    n264
  );


  buf
  g304
  (
    n386,
    n258
  );


  buf
  g305
  (
    n358,
    n301
  );


  buf
  g306
  (
    n340,
    n284
  );


  not
  g307
  (
    n385,
    n288
  );


  buf
  g308
  (
    n356,
    n244
  );


  nor
  g309
  (
    n394,
    n255,
    n251
  );


  nand
  g310
  (
    n434,
    n269,
    n248,
    n196,
    n216
  );


  and
  g311
  (
    n488,
    n279,
    n269,
    n271,
    n130
  );


  and
  g312
  (
    n457,
    n280,
    n210,
    n282,
    n135
  );


  or
  g313
  (
    n384,
    n225,
    n218,
    n242,
    n164
  );


  xor
  g314
  (
    n351,
    n260,
    n278,
    n205
  );


  nor
  g315
  (
    n360,
    n185,
    n130,
    n303,
    n180
  );


  xor
  g316
  (
    n331,
    n258,
    n228,
    n131,
    n213
  );


  or
  g317
  (
    n490,
    n247,
    n166,
    n274,
    n199
  );


  xnor
  g318
  (
    n414,
    n275,
    n289,
    n204,
    n128
  );


  xnor
  g319
  (
    n461,
    n255,
    n166,
    n215,
    n201
  );


  xnor
  g320
  (
    n456,
    n283,
    n289,
    n245,
    n187
  );


  xor
  g321
  (
    n432,
    n205,
    n273,
    n202,
    n210
  );


  nor
  g322
  (
    KeyWire_0_41,
    n287,
    n236,
    n127,
    n231
  );


  xor
  g323
  (
    n410,
    n176,
    n180,
    n262,
    n302
  );


  nor
  g324
  (
    n326,
    n133,
    n194,
    n192,
    n280
  );


  nor
  g325
  (
    n425,
    n169,
    n236,
    n244,
    n276
  );


  nand
  g326
  (
    n407,
    n260,
    n183,
    n217
  );


  xor
  g327
  (
    n485,
    n229,
    n199,
    n261,
    n162
  );


  nand
  g328
  (
    KeyWire_0_4,
    n179,
    n168,
    n250,
    n212
  );


  or
  g329
  (
    n439,
    n194,
    n294,
    n127,
    n201
  );


  xnor
  g330
  (
    n477,
    n272,
    n254,
    n245,
    n191
  );


  xor
  g331
  (
    n372,
    n163,
    n251,
    n190,
    n184
  );


  or
  g332
  (
    n436,
    n280,
    n246,
    n216,
    n263
  );


  nand
  g333
  (
    n376,
    n255,
    n189,
    n168,
    n266
  );


  xnor
  g334
  (
    n474,
    n232,
    n248,
    n161,
    n164
  );


  xor
  g335
  (
    n341,
    n135,
    n185,
    n178,
    n212
  );


  nand
  g336
  (
    n330,
    n294,
    n255,
    n170,
    n285
  );


  nand
  g337
  (
    n466,
    n221,
    n238,
    n271,
    n136
  );


  nor
  g338
  (
    n444,
    n299,
    n166,
    n195,
    n256
  );


  or
  g339
  (
    n449,
    n192,
    n207,
    n238,
    n128
  );


  xor
  g340
  (
    n409,
    n275,
    n228,
    n206,
    n291
  );


  xnor
  g341
  (
    n482,
    n173,
    n130,
    n259,
    n186
  );


  nand
  g342
  (
    n411,
    n276,
    n233,
    n249
  );


  and
  g343
  (
    n357,
    n269,
    n167,
    n211,
    n196
  );


  or
  g344
  (
    n421,
    n239,
    n232,
    n198,
    n191
  );


  nor
  g345
  (
    n334,
    n266,
    n194,
    n133,
    n275
  );


  xor
  g346
  (
    n364,
    n136,
    n252,
    n267,
    n246
  );


  nand
  g347
  (
    n390,
    n135,
    n240,
    n248,
    n188
  );


  xor
  g348
  (
    n445,
    n301,
    n184,
    n203,
    n226
  );


  xor
  g349
  (
    n489,
    n177,
    n247,
    n281,
    n165
  );


  or
  g350
  (
    n345,
    n182,
    n216,
    n208,
    n244
  );


  nand
  g351
  (
    n325,
    n194,
    n253,
    n201,
    n273
  );


  xnor
  g352
  (
    n440,
    n132,
    n185,
    n218,
    n281
  );


  xor
  g353
  (
    n458,
    n263,
    n298,
    n294,
    n174
  );


  xnor
  g354
  (
    n481,
    n244,
    n282,
    n227,
    n195
  );


  or
  g355
  (
    n479,
    n293,
    n189,
    n130,
    n268
  );


  xor
  g356
  (
    n393,
    n243,
    n253,
    n248,
    n167
  );


  nand
  g357
  (
    KeyWire_0_55,
    n284,
    n241,
    n256,
    n212
  );


  xnor
  g358
  (
    n455,
    n246,
    n265,
    n254,
    n172
  );


  and
  g359
  (
    n374,
    n173,
    n241,
    n131,
    n285
  );


  and
  g360
  (
    n430,
    n263,
    n203,
    n235,
    n282
  );


  xor
  g361
  (
    n438,
    n219,
    n290,
    n198,
    n170
  );


  and
  g362
  (
    KeyWire_0_15,
    n174,
    n169,
    n286,
    n186
  );


  nand
  g363
  (
    n329,
    n213,
    n126,
    n250,
    n303
  );


  or
  g364
  (
    n348,
    n209,
    n275,
    n261,
    n163
  );


  nor
  g365
  (
    n381,
    n175,
    n219,
    n167,
    n231
  );


  nor
  g366
  (
    n361,
    n227,
    n242,
    n204,
    n129
  );


  and
  g367
  (
    n443,
    n134,
    n240,
    n221,
    n237
  );


  nand
  g368
  (
    n366,
    n258,
    n279,
    n226,
    n289
  );


  nor
  g369
  (
    n469,
    n272,
    n300,
    n190,
    n269
  );


  nor
  g370
  (
    n419,
    n210,
    n178,
    n177,
    n252
  );


  xor
  g371
  (
    n408,
    n220,
    n268,
    n128,
    n242
  );


  xnor
  g372
  (
    n406,
    n170,
    n276,
    n213,
    n172
  );


  nor
  g373
  (
    n465,
    n224,
    n281,
    n285,
    n193
  );


  xnor
  g374
  (
    n459,
    n227,
    n170,
    n206,
    n203
  );


  nor
  g375
  (
    n328,
    n165,
    n210,
    n173,
    n181
  );


  xnor
  g376
  (
    n452,
    n250,
    n220,
    n134,
    n200
  );


  xor
  g377
  (
    n427,
    n291,
    n270,
    n245,
    n274
  );


  or
  g378
  (
    n442,
    n193,
    n172,
    n195
  );


  or
  g379
  (
    n446,
    n222,
    n292,
    n188,
    n168
  );


  nor
  g380
  (
    KeyWire_0_18,
    n181,
    n293,
    n162,
    n183
  );


  nand
  g381
  (
    n415,
    n126,
    n287,
    n161,
    n192
  );


  xor
  g382
  (
    n342,
    n223,
    n207,
    n175,
    n229
  );


  xor
  g383
  (
    n335,
    n225,
    n249,
    n287,
    n265
  );


  or
  g384
  (
    n365,
    n128,
    n230,
    n182,
    n129
  );


  nand
  g385
  (
    n354,
    n229,
    n257,
    n301,
    n175
  );


  xnor
  g386
  (
    n382,
    n176,
    n214,
    n204,
    n233
  );


  xnor
  g387
  (
    n373,
    n277,
    n230,
    n208,
    n184
  );


  or
  g388
  (
    n450,
    n260,
    n188,
    n258,
    n223
  );


  nand
  g389
  (
    n472,
    n228,
    n278,
    n217,
    n259
  );


  nand
  g390
  (
    n387,
    n203,
    n234,
    n214,
    n131
  );


  xor
  g391
  (
    n460,
    n230,
    n239,
    n232,
    n133
  );


  nand
  g392
  (
    n424,
    n192,
    n266,
    n298,
    n129
  );


  nand
  g393
  (
    n401,
    n302,
    n250,
    n221,
    n256
  );


  nand
  g394
  (
    n433,
    n205,
    n190,
    n171,
    n289
  );


  nor
  g395
  (
    n346,
    n178,
    n207,
    n165,
    n209
  );


  xnor
  g396
  (
    n375,
    n300,
    n221,
    n284,
    n297
  );


  nor
  g397
  (
    n431,
    n131,
    n199,
    n240,
    n161
  );


  or
  g398
  (
    n350,
    n232,
    n126,
    n268,
    n237
  );


  or
  g399
  (
    n429,
    n259,
    n164,
    n222,
    n162
  );


  or
  g400
  (
    n362,
    n223,
    n202,
    n283,
    n264
  );


  and
  g401
  (
    n396,
    n288,
    n163,
    n286,
    n291
  );


  and
  g402
  (
    n451,
    n197,
    n296,
    n283,
    n247
  );


  and
  g403
  (
    n403,
    n127,
    n174,
    n290,
    n206
  );


  nand
  g404
  (
    n391,
    n241,
    n134,
    n185,
    n299
  );


  or
  g405
  (
    n435,
    n177,
    n271,
    n163
  );


  or
  g406
  (
    n473,
    n292,
    n231,
    n219,
    n272
  );


  or
  g407
  (
    n347,
    n169,
    n245,
    n277,
    n179
  );


  xor
  g408
  (
    KeyWire_0_34,
    n287,
    n279,
    n295,
    n189
  );


  nand
  g409
  (
    n344,
    n263,
    n206,
    n300,
    n261
  );


  nor
  g410
  (
    n417,
    n262,
    n186,
    n236,
    n195
  );


  nand
  g411
  (
    n416,
    n251,
    n173,
    n270,
    n252
  );


  nor
  g412
  (
    n448,
    n297,
    n183,
    n268,
    n257
  );


  nor
  g413
  (
    n486,
    n270,
    n225,
    n175,
    n299
  );


  nand
  g414
  (
    n395,
    n267,
    n292,
    n181,
    n246
  );


  xor
  g415
  (
    n338,
    n187,
    n234,
    n238,
    n243
  );


  nand
  g416
  (
    n462,
    n298,
    n276,
    n217,
    n171
  );


  and
  g417
  (
    n389,
    n134,
    n262,
    n197,
    n238
  );


  nor
  g418
  (
    n353,
    n215,
    n296,
    n171,
    n252
  );


  or
  g419
  (
    n336,
    n233,
    n296,
    n298,
    n236
  );


  nand
  g420
  (
    n428,
    n212,
    n198,
    n174,
    n264
  );


  or
  g421
  (
    KeyWire_0_26,
    n167,
    n234,
    n282,
    n227
  );


  nand
  g422
  (
    n355,
    n189,
    n202,
    n237,
    n253
  );


  nor
  g423
  (
    n467,
    n253,
    n229,
    n198,
    n215
  );


  xor
  g424
  (
    n370,
    n135,
    n292,
    n274,
    n171
  );


  and
  g425
  (
    n369,
    n211,
    n211,
    n224,
    n294
  );


  xnor
  g426
  (
    n398,
    n290,
    n265,
    n165,
    n247
  );


  and
  g427
  (
    n468,
    n168,
    n286,
    n205,
    n235
  );


  or
  g428
  (
    n483,
    n211,
    n200,
    n295,
    n272
  );


  and
  g429
  (
    n359,
    n230,
    n196,
    n200
  );


  xor
  g430
  (
    n363,
    n132,
    n226,
    n166,
    n207
  );


  xnor
  g431
  (
    n402,
    n164,
    n184,
    n214,
    n179
  );


  nor
  g432
  (
    n423,
    n277,
    n213,
    n267,
    n182
  );


  xnor
  g433
  (
    n388,
    n243,
    n169,
    n235,
    n237
  );


  and
  g434
  (
    n405,
    n228,
    n266,
    n187,
    n265
  );


  and
  g435
  (
    n480,
    n133,
    n239,
    n204,
    n127
  );


  nand
  g436
  (
    n464,
    n302,
    n286,
    n279,
    n193
  );


  nand
  g437
  (
    n399,
    n257,
    n262,
    n270,
    n225
  );


  and
  g438
  (
    n484,
    n176,
    n220,
    n178,
    n186
  );


  xnor
  g439
  (
    n397,
    n299,
    n235,
    n233,
    n188
  );


  and
  g440
  (
    KeyWire_0_61,
    n297,
    n197,
    n301,
    n293
  );


  xnor
  g441
  (
    KeyWire_0_7,
    n177,
    n241,
    n231,
    n216
  );


  xor
  g442
  (
    n333,
    n256,
    n254,
    n234,
    n214
  );


  nor
  g443
  (
    n332,
    n226,
    n187,
    n239,
    n222
  );


  and
  g444
  (
    n441,
    n223,
    n191,
    n220,
    n260
  );


  nand
  g445
  (
    n379,
    n215,
    n293,
    n300,
    n190
  );


  nor
  g446
  (
    n371,
    n297,
    n281,
    n285,
    n257
  );


  xor
  g447
  (
    n420,
    n302,
    n199,
    n242,
    n295
  );


  xnor
  g448
  (
    n475,
    n129,
    n288,
    n208,
    n274
  );


  xnor
  g449
  (
    n367,
    n180,
    n180,
    n273,
    n219
  );


  nand
  g450
  (
    n400,
    n291,
    n222,
    n161,
    n218
  );


  and
  g451
  (
    n343,
    n283,
    n259,
    n208,
    n249
  );


  xor
  g452
  (
    n352,
    n218,
    n209,
    n132,
    n295
  );


  nand
  g453
  (
    n368,
    n290,
    n267,
    n132,
    n196
  );


  xor
  g454
  (
    n478,
    n197,
    n280,
    n251,
    n254
  );


  nor
  g455
  (
    n418,
    n179,
    n277,
    n261,
    n162
  );


  nand
  g456
  (
    n380,
    n264,
    n176,
    n284,
    n224
  );


  nor
  g457
  (
    n404,
    n243,
    n193,
    n202,
    n217
  );


  xnor
  g458
  (
    KeyWire_0_38,
    n330,
    n339,
    n336,
    n326
  );


  and
  g459
  (
    n504,
    n331,
    n339,
    n334,
    n328
  );


  xor
  g460
  (
    n501,
    n326,
    n327,
    n330,
    n332
  );


  xor
  g461
  (
    n493,
    n338,
    n331,
    n341,
    n333
  );


  and
  g462
  (
    n499,
    n332,
    n334,
    n331,
    n338
  );


  or
  g463
  (
    n505,
    n340,
    n329,
    n339
  );


  xor
  g464
  (
    n497,
    n336,
    n332,
    n333
  );


  or
  g465
  (
    n495,
    n333,
    n335,
    n340
  );


  xnor
  g466
  (
    KeyWire_0_52,
    n327,
    n341
  );


  or
  g467
  (
    KeyWire_0_9,
    n329,
    n326,
    n328,
    n337
  );


  nand
  g468
  (
    n500,
    n330,
    n334,
    n335,
    n331
  );


  nand
  g469
  (
    n492,
    n327,
    n340,
    n330,
    n337
  );


  and
  g470
  (
    n506,
    n337,
    n326,
    n338
  );


  xnor
  g471
  (
    n496,
    n329,
    n341,
    n339,
    n335
  );


  nor
  g472
  (
    n494,
    n334,
    n328,
    n337
  );


  nand
  g473
  (
    KeyWire_0_11,
    n340,
    n336,
    n332
  );


  buf
  g474
  (
    n509,
    n496
  );


  buf
  g475
  (
    n511,
    n501
  );


  buf
  g476
  (
    n515,
    n504
  );


  buf
  g477
  (
    n512,
    n497
  );


  buf
  g478
  (
    n528,
    n501
  );


  buf
  g479
  (
    n508,
    n506
  );


  buf
  g480
  (
    n524,
    n493
  );


  buf
  g481
  (
    n510,
    n503
  );


  not
  g482
  (
    KeyWire_0_54,
    n502
  );


  buf
  g483
  (
    n526,
    n506
  );


  not
  g484
  (
    n518,
    n505
  );


  not
  g485
  (
    n519,
    n504
  );


  not
  g486
  (
    n523,
    n500
  );


  not
  g487
  (
    n507,
    n491
  );


  buf
  g488
  (
    n527,
    n492
  );


  not
  g489
  (
    n522,
    n495
  );


  buf
  g490
  (
    n521,
    n499
  );


  buf
  g491
  (
    n516,
    n503
  );


  buf
  g492
  (
    n513,
    n502
  );


  buf
  g493
  (
    KeyWire_0_28,
    n505
  );


  not
  g494
  (
    n525,
    n494
  );


  not
  g495
  (
    n520,
    n498
  );


  nand
  g496
  (
    n539,
    n359,
    n384,
    n361,
    n377
  );


  xnor
  g497
  (
    n541,
    n366,
    n525,
    n516,
    n141
  );


  xnor
  g498
  (
    n578,
    n352,
    n364,
    n513,
    n142
  );


  nor
  g499
  (
    n604,
    n520,
    n350,
    n515,
    n347
  );


  or
  g500
  (
    n582,
    n523,
    n521,
    n364,
    n385
  );


  xor
  g501
  (
    n542,
    n382,
    n523,
    n365,
    n142
  );


  xnor
  g502
  (
    n581,
    n512,
    n140,
    n357,
    n511
  );


  or
  g503
  (
    n580,
    n143,
    n352,
    n521,
    n353
  );


  xor
  g504
  (
    n546,
    n356,
    n362,
    n345,
    n368
  );


  xnor
  g505
  (
    n571,
    n374,
    n381,
    n369,
    n520
  );


  or
  g506
  (
    n559,
    n368,
    n151,
    n376,
    n511
  );


  xnor
  g507
  (
    KeyWire_0_45,
    n526,
    n362,
    n146,
    n350
  );


  xor
  g508
  (
    n595,
    n377,
    n507,
    n140,
    n347
  );


  xor
  g509
  (
    KeyWire_0_30,
    n344,
    n524,
    n148,
    n510
  );


  nor
  g510
  (
    n566,
    n375,
    n508,
    n140,
    n520
  );


  xor
  g511
  (
    n588,
    n522,
    n383,
    n517,
    n142
  );


  or
  g512
  (
    n589,
    n136,
    n150,
    n382,
    n377
  );


  or
  g513
  (
    n548,
    n138,
    n146,
    n344,
    n515
  );


  xnor
  g514
  (
    n600,
    n375,
    n371,
    n342,
    n142
  );


  xnor
  g515
  (
    n573,
    n345,
    n374,
    n382,
    n358
  );


  nor
  g516
  (
    n596,
    n378,
    n373,
    n342,
    n374
  );


  or
  g517
  (
    n602,
    n525,
    n373,
    n511,
    n517
  );


  xor
  g518
  (
    KeyWire_0_13,
    n516,
    n346,
    n378,
    n141
  );


  xor
  g519
  (
    n556,
    n518,
    n526,
    n350,
    n381
  );


  xor
  g520
  (
    KeyWire_0_12,
    n372,
    n523,
    n347,
    n371
  );


  nor
  g521
  (
    n530,
    n360,
    n521,
    n371,
    n348
  );


  xor
  g522
  (
    KeyWire_0_62,
    n507,
    n150,
    n526,
    n370
  );


  and
  g523
  (
    n545,
    n527,
    n138,
    n139,
    n363
  );


  nand
  g524
  (
    n532,
    n349,
    n373,
    n375,
    n147
  );


  xor
  g525
  (
    n607,
    n383,
    n342,
    n139,
    n145
  );


  and
  g526
  (
    n586,
    n517,
    n510,
    n144,
    n379
  );


  nor
  g527
  (
    n585,
    n357,
    n379,
    n514,
    n360
  );


  xnor
  g528
  (
    n557,
    n149,
    n152,
    n145,
    n513
  );


  or
  g529
  (
    n553,
    n147,
    n362,
    n366,
    n376
  );


  xor
  g530
  (
    n584,
    n151,
    n380,
    n385,
    n508
  );


  nand
  g531
  (
    n533,
    n345,
    n357,
    n141,
    n368
  );


  xnor
  g532
  (
    n540,
    n513,
    n152,
    n144,
    n524
  );


  and
  g533
  (
    n558,
    n522,
    n522,
    n361,
    n360
  );


  nand
  g534
  (
    n565,
    n149,
    n514,
    n355,
    n508
  );


  and
  g535
  (
    n603,
    n380,
    n348,
    n346,
    n507
  );


  and
  g536
  (
    KeyWire_0_57,
    n521,
    n152,
    n355,
    n377
  );


  or
  g537
  (
    n583,
    n352,
    n526,
    n149,
    n358
  );


  xnor
  g538
  (
    n576,
    n520,
    n375,
    n356,
    n516
  );


  xnor
  g539
  (
    n606,
    n145,
    n363,
    n376,
    n349
  );


  nand
  g540
  (
    n592,
    n378,
    n510,
    n148,
    n508
  );


  or
  g541
  (
    n608,
    n347,
    n381,
    n518,
    n354
  );


  nor
  g542
  (
    n555,
    n380,
    n352,
    n145,
    n140
  );


  and
  g543
  (
    n579,
    n514,
    n137,
    n365,
    n362
  );


  or
  g544
  (
    KeyWire_0_32,
    n354,
    n371,
    n382,
    n343
  );


  xnor
  g545
  (
    n552,
    n370,
    n150,
    n512,
    n137
  );


  or
  g546
  (
    n550,
    n146,
    n374,
    n345,
    n381
  );


  xor
  g547
  (
    n609,
    n523,
    n512,
    n364,
    n148
  );


  and
  g548
  (
    n531,
    n525,
    n144,
    n346,
    n343
  );


  nor
  g549
  (
    n551,
    n141,
    n517,
    n363,
    n139
  );


  nor
  g550
  (
    n605,
    n385,
    n376,
    n379,
    n518
  );


  nor
  g551
  (
    n594,
    n510,
    n366,
    n351
  );


  nor
  g552
  (
    n599,
    n509,
    n369,
    n357,
    n519
  );


  and
  g553
  (
    n568,
    n370,
    n151,
    n384,
    n380
  );


  and
  g554
  (
    n601,
    n372,
    n370,
    n348,
    n358
  );


  nand
  g555
  (
    n554,
    n355,
    n136,
    n515,
    n361
  );


  xor
  g556
  (
    n543,
    n509,
    n348,
    n369,
    n356
  );


  and
  g557
  (
    n567,
    n353,
    n151,
    n378,
    n139
  );


  or
  g558
  (
    n538,
    n153,
    n137,
    n372,
    n356
  );


  or
  g559
  (
    n569,
    n519,
    n149,
    n351,
    n150
  );


  xnor
  g560
  (
    n570,
    n519,
    n346,
    n518,
    n359
  );


  or
  g561
  (
    n561,
    n509,
    n358,
    n351,
    n350
  );


  xor
  g562
  (
    n537,
    n367,
    n524,
    n355
  );


  or
  g563
  (
    n535,
    n379,
    n383,
    n367
  );


  xor
  g564
  (
    n597,
    n148,
    n384,
    n138,
    n519
  );


  xnor
  g565
  (
    n564,
    n147,
    n143,
    n361,
    n369
  );


  xor
  g566
  (
    n560,
    n513,
    n515,
    n509,
    n344
  );


  xor
  g567
  (
    n544,
    n516,
    n144,
    n368,
    n143
  );


  nor
  g568
  (
    n549,
    n365,
    n360,
    n364,
    n343
  );


  xor
  g569
  (
    KeyWire_0_42,
    n365,
    n359,
    n349,
    n512
  );


  xor
  g570
  (
    n587,
    n511,
    n351,
    n514,
    n138
  );


  or
  g571
  (
    n593,
    n147,
    n143,
    n525,
    n367
  );


  and
  g572
  (
    n563,
    n146,
    n137,
    n363,
    n385
  );


  and
  g573
  (
    n591,
    n367,
    n522,
    n353,
    n384
  );


  xor
  g574
  (
    KeyWire_0_39,
    n353,
    n372,
    n354,
    n507
  );


  nor
  g575
  (
    n575,
    n152,
    n342,
    n359,
    n349
  );


  nand
  g576
  (
    n534,
    n343,
    n344,
    n373,
    n354
  );


  not
  g577
  (
    n624,
    n574
  );


  buf
  g578
  (
    n636,
    n552
  );


  not
  g579
  (
    n685,
    n570
  );


  buf
  g580
  (
    n639,
    n533
  );


  buf
  g581
  (
    n680,
    n553
  );


  not
  g582
  (
    n659,
    n528
  );


  buf
  g583
  (
    n627,
    n311
  );


  not
  g584
  (
    n629,
    n420
  );


  or
  g585
  (
    KeyWire_0_20,
    n403,
    n562,
    n429,
    n425
  );


  xnor
  g586
  (
    n737,
    n576,
    n399,
    n557,
    n542
  );


  nand
  g587
  (
    n697,
    n571,
    n405,
    n569,
    n418
  );


  xor
  g588
  (
    n653,
    n423,
    n538,
    n561,
    n319
  );


  and
  g589
  (
    n692,
    n542,
    n319,
    n404,
    n153
  );


  and
  g590
  (
    n654,
    n541,
    n569,
    n316,
    n320
  );


  xor
  g591
  (
    KeyWire_0_36,
    n530,
    n427,
    n155,
    n408
  );


  or
  g592
  (
    n615,
    n406,
    n571,
    n155,
    n555
  );


  and
  g593
  (
    n704,
    n573,
    n157,
    n564,
    n558
  );


  xnor
  g594
  (
    KeyWire_0_51,
    n430,
    n321,
    n407
  );


  xnor
  g595
  (
    n610,
    n321,
    n533,
    n547,
    n426
  );


  xnor
  g596
  (
    n727,
    n578,
    n323,
    n572,
    n389
  );


  nand
  g597
  (
    n613,
    n569,
    n413,
    n540,
    n318
  );


  and
  g598
  (
    n709,
    n424,
    n552,
    n309,
    n417
  );


  or
  g599
  (
    n681,
    n154,
    n323,
    n420,
    n401
  );


  nand
  g600
  (
    n663,
    n318,
    n321,
    n315,
    n409
  );


  and
  g601
  (
    n725,
    n565,
    n417,
    n309,
    n429
  );


  xor
  g602
  (
    n626,
    n156,
    n414,
    n399,
    n548
  );


  and
  g603
  (
    n675,
    n540,
    n576,
    n553,
    n570
  );


  xnor
  g604
  (
    n733,
    n552,
    n393,
    n426,
    n391
  );


  and
  g605
  (
    n688,
    n567,
    n559,
    n532,
    n527
  );


  and
  g606
  (
    n694,
    n530,
    n427,
    n551,
    n418
  );


  xnor
  g607
  (
    n631,
    n546,
    n548,
    n306,
    n391
  );


  and
  g608
  (
    n635,
    n534,
    n306,
    n533,
    n550
  );


  and
  g609
  (
    n650,
    n547,
    n566,
    n306,
    n549
  );


  xnor
  g610
  (
    n705,
    n397,
    n566,
    n396,
    n569
  );


  xnor
  g611
  (
    n662,
    n316,
    n428,
    n580,
    n390
  );


  or
  g612
  (
    n655,
    n411,
    n532,
    n393,
    n539
  );


  nand
  g613
  (
    n721,
    n431,
    n529,
    n560,
    n538
  );


  and
  g614
  (
    n652,
    n397,
    n420,
    n419,
    n579
  );


  nor
  g615
  (
    n728,
    n554,
    n546,
    n529,
    n310
  );


  nor
  g616
  (
    n684,
    n578,
    n560,
    n535,
    n318
  );


  nand
  g617
  (
    n634,
    n578,
    n406,
    n537,
    n309
  );


  and
  g618
  (
    n637,
    n547,
    n571,
    n398,
    n317
  );


  nor
  g619
  (
    n646,
    n568,
    n531,
    n416,
    n408
  );


  and
  g620
  (
    n690,
    n403,
    n531,
    n555,
    n395
  );


  nand
  g621
  (
    KeyWire_0_59,
    n323,
    n415,
    n389,
    n423
  );


  xnor
  g622
  (
    n642,
    n410,
    n577,
    n430,
    n386
  );


  or
  g623
  (
    n656,
    n554,
    n403,
    n536,
    n424
  );


  nand
  g624
  (
    n730,
    n154,
    n407,
    n320,
    n315
  );


  nand
  g625
  (
    n630,
    n535,
    n426,
    n549,
    n539
  );


  nand
  g626
  (
    n643,
    n401,
    n541,
    n554,
    n422
  );


  or
  g627
  (
    n726,
    n574,
    n303,
    n539,
    n552
  );


  nor
  g628
  (
    n710,
    n556,
    n561,
    n306,
    n425
  );


  xnor
  g629
  (
    n625,
    n404,
    n565,
    n413,
    n392
  );


  or
  g630
  (
    n689,
    n422,
    n153,
    n429,
    n304
  );


  nor
  g631
  (
    n638,
    n545,
    n559,
    n412,
    n536
  );


  or
  g632
  (
    n683,
    n431,
    n407,
    n528,
    n413
  );


  or
  g633
  (
    n723,
    n315,
    n551,
    n402,
    n400
  );


  xnor
  g634
  (
    n648,
    n316,
    n540,
    n421,
    n533
  );


  and
  g635
  (
    n686,
    n402,
    n393,
    n430,
    n406
  );


  and
  g636
  (
    n735,
    n568,
    n421,
    n551,
    n317
  );


  and
  g637
  (
    n671,
    n410,
    n308,
    n419,
    n563
  );


  xnor
  g638
  (
    n701,
    n314,
    n576,
    n418,
    n313
  );


  and
  g639
  (
    n677,
    n544,
    n425,
    n570,
    n314
  );


  nand
  g640
  (
    n687,
    n546,
    n317,
    n388,
    n556
  );


  nand
  g641
  (
    n696,
    n537,
    n313,
    n156,
    n558
  );


  nand
  g642
  (
    n695,
    n398,
    n312,
    n402,
    n553
  );


  nand
  g643
  (
    n693,
    n153,
    n155,
    n577,
    n311
  );


  nand
  g644
  (
    n645,
    n547,
    n415,
    n538,
    n412
  );


  or
  g645
  (
    n706,
    n565,
    n568,
    n391,
    n555
  );


  nor
  g646
  (
    n738,
    n527,
    n409,
    n579,
    n570
  );


  xnor
  g647
  (
    n658,
    n428,
    n558,
    n539,
    n531
  );


  nor
  g648
  (
    n729,
    n541,
    n572,
    n558,
    n307
  );


  nor
  g649
  (
    n665,
    n549,
    n529,
    n577,
    n550
  );


  nand
  g650
  (
    KeyWire_0_53,
    n392,
    n412,
    n553,
    n556
  );


  nor
  g651
  (
    n703,
    n398,
    n554,
    n312,
    n424
  );


  xnor
  g652
  (
    n673,
    n394,
    n304,
    n534,
    n423
  );


  xnor
  g653
  (
    n647,
    n575,
    n408,
    n560,
    n534
  );


  nand
  g654
  (
    n660,
    n154,
    n308,
    n557,
    n420
  );


  and
  g655
  (
    n736,
    n305,
    n308,
    n312,
    n572
  );


  xnor
  g656
  (
    n708,
    n395,
    n317,
    n387,
    n562
  );


  or
  g657
  (
    n672,
    n398,
    n312,
    n561,
    n154
  );


  nor
  g658
  (
    n611,
    n536,
    n397,
    n405,
    n411
  );


  nor
  g659
  (
    n714,
    n563,
    n322,
    n562,
    n542
  );


  xnor
  g660
  (
    n612,
    n564,
    n572,
    n422,
    n313
  );


  xnor
  g661
  (
    n712,
    n396,
    n386,
    n417,
    n401
  );


  or
  g662
  (
    n640,
    n545,
    n548,
    n405,
    n426
  );


  nor
  g663
  (
    n702,
    n557,
    n573,
    n571,
    n544
  );


  or
  g664
  (
    KeyWire_0_6,
    n409,
    n425,
    n390,
    n305
  );


  and
  g665
  (
    n732,
    n549,
    n575,
    n528,
    n431
  );


  xnor
  g666
  (
    n682,
    n532,
    n156,
    n559,
    n556
  );


  xor
  g667
  (
    n657,
    n419,
    n565,
    n395,
    n403
  );


  nand
  g668
  (
    n678,
    n555,
    n411,
    n563,
    n416
  );


  and
  g669
  (
    n616,
    n307,
    n396,
    n427,
    n527
  );


  nor
  g670
  (
    n623,
    n545,
    n394,
    n577,
    n406
  );


  nand
  g671
  (
    n632,
    n396,
    n307,
    n575,
    n546
  );


  xor
  g672
  (
    n641,
    n416,
    n537,
    n566,
    n389
  );


  xor
  g673
  (
    n731,
    n395,
    n404,
    n580,
    n305
  );


  xnor
  g674
  (
    n699,
    n324,
    n568,
    n315,
    n532
  );


  or
  g675
  (
    n619,
    n562,
    n404,
    n388,
    n544
  );


  nor
  g676
  (
    n628,
    n400,
    n540,
    n544,
    n430
  );


  xor
  g677
  (
    n667,
    n543,
    n431,
    n576,
    n399
  );


  or
  g678
  (
    n633,
    n566,
    n538,
    n316,
    n402
  );


  or
  g679
  (
    n691,
    n543,
    n387,
    n559,
    n310
  );


  nand
  g680
  (
    n676,
    n414,
    n543,
    n567,
    n400
  );


  and
  g681
  (
    n666,
    n543,
    n407,
    n394,
    n542
  );


  xor
  g682
  (
    n649,
    n550,
    n564,
    n392,
    n531
  );


  xor
  g683
  (
    n614,
    n310,
    n319,
    n416,
    n389
  );


  xnor
  g684
  (
    n722,
    n567,
    n388,
    n390,
    n320
  );


  and
  g685
  (
    n720,
    n415,
    n412,
    n541,
    n319
  );


  and
  g686
  (
    KeyWire_0_27,
    n573,
    n564,
    n417,
    n308
  );


  xor
  g687
  (
    n661,
    n535,
    n423,
    n529,
    n307
  );


  nor
  g688
  (
    n734,
    n418,
    n422,
    n397,
    n563
  );


  nand
  g689
  (
    n664,
    n427,
    n311,
    n415,
    n303
  );


  xor
  g690
  (
    n668,
    n537,
    n155,
    n387,
    n424
  );


  nor
  g691
  (
    n711,
    n392,
    n414,
    n567
  );


  or
  g692
  (
    n715,
    n322,
    n386,
    n318,
    n388
  );


  nor
  g693
  (
    n724,
    n387,
    n400,
    n310,
    n530
  );


  and
  g694
  (
    n698,
    n530,
    n573,
    n386,
    n419
  );


  xor
  g695
  (
    n674,
    n534,
    n313,
    n579,
    n575
  );


  and
  g696
  (
    n620,
    n428,
    n560,
    n323,
    n535
  );


  nand
  g697
  (
    n713,
    n391,
    n401,
    n428,
    n390
  );


  xnor
  g698
  (
    n617,
    n304,
    n561,
    n410,
    n421
  );


  and
  g699
  (
    n618,
    n393,
    n574,
    n309,
    n408
  );


  xnor
  g700
  (
    n718,
    n304,
    n409,
    n413,
    n394
  );


  nand
  g701
  (
    n651,
    n156,
    n320,
    n574,
    n548
  );


  xor
  g702
  (
    n622,
    n314,
    n551,
    n536,
    n399
  );


  xor
  g703
  (
    n719,
    n305,
    n528,
    n579,
    n557
  );


  and
  g704
  (
    n739,
    n311,
    n322,
    n410,
    n578
  );


  xor
  g705
  (
    n669,
    n550,
    n421,
    n545,
    n411
  );


  xor
  g706
  (
    n717,
    n314,
    n405,
    n429,
    n322
  );


  nand
  g707
  (
    n784,
    n476,
    n717,
    n471,
    n599
  );


  and
  g708
  (
    n813,
    n658,
    n462,
    n736,
    n437
  );


  and
  g709
  (
    n824,
    n619,
    n478,
    n615,
    n584
  );


  nand
  g710
  (
    n956,
    n669,
    n604,
    n725,
    n629
  );


  xor
  g711
  (
    n918,
    n679,
    n159,
    n718,
    n651
  );


  nand
  g712
  (
    n752,
    n717,
    n693,
    n683,
    n684
  );


  and
  g713
  (
    n929,
    n586,
    n460,
    n665,
    n733
  );


  and
  g714
  (
    n838,
    n682,
    n646,
    n457,
    n664
  );


  and
  g715
  (
    n923,
    n600,
    n461,
    n724,
    n693
  );


  xnor
  g716
  (
    n879,
    n665,
    n444,
    n659,
    n607
  );


  and
  g717
  (
    n859,
    n650,
    n704,
    n456,
    n652
  );


  or
  g718
  (
    n753,
    n601,
    n675,
    n720,
    n725
  );


  and
  g719
  (
    n863,
    n721,
    n478,
    n581,
    n714
  );


  xor
  g720
  (
    n846,
    n620,
    n448,
    n724,
    n726
  );


  nand
  g721
  (
    n827,
    n450,
    n725,
    n625,
    n443
  );


  or
  g722
  (
    n869,
    n680,
    n477,
    n604,
    n489
  );


  and
  g723
  (
    n819,
    n721,
    n483,
    n607,
    n713
  );


  xnor
  g724
  (
    n772,
    n696,
    n667,
    n457,
    n676
  );


  or
  g725
  (
    n804,
    n728,
    n594,
    n709,
    n676
  );


  xnor
  g726
  (
    n886,
    n617,
    n702,
    n605,
    n634
  );


  or
  g727
  (
    n945,
    n655,
    n463,
    n476,
    n643
  );


  nor
  g728
  (
    n925,
    n617,
    n667,
    n588,
    n683
  );


  nor
  g729
  (
    n820,
    n485,
    n721,
    n690,
    n583
  );


  nand
  g730
  (
    n759,
    n695,
    n641,
    n642,
    n451
  );


  xor
  g731
  (
    n877,
    n606,
    n682,
    n635,
    n704
  );


  and
  g732
  (
    n816,
    n587,
    n592,
    n705,
    n619
  );


  xnor
  g733
  (
    n791,
    n593,
    n616,
    n454,
    n601
  );


  nor
  g734
  (
    n950,
    n435,
    n701,
    n641,
    n636
  );


  nand
  g735
  (
    n740,
    n597,
    n632,
    n662,
    n681
  );


  xor
  g736
  (
    KeyWire_0_48,
    n727,
    n608,
    n638,
    n702
  );


  and
  g737
  (
    n912,
    n657,
    n633,
    n732,
    n157
  );


  xnor
  g738
  (
    n774,
    n719,
    n447,
    n437,
    n470
  );


  and
  g739
  (
    n832,
    n722,
    n688,
    n643,
    n697
  );


  and
  g740
  (
    n953,
    n588,
    n697,
    n466,
    n660
  );


  or
  g741
  (
    n903,
    n631,
    n454,
    n666,
    n738
  );


  or
  g742
  (
    n823,
    n622,
    n720,
    n624,
    n672
  );


  or
  g743
  (
    n775,
    n475,
    n694,
    n686,
    n636
  );


  nand
  g744
  (
    n814,
    n690,
    n490,
    n446,
    n689
  );


  nand
  g745
  (
    n907,
    n451,
    n590,
    n719,
    n685
  );


  xnor
  g746
  (
    n882,
    n635,
    n432,
    n644,
    n734
  );


  xnor
  g747
  (
    n921,
    n677,
    n626,
    n600,
    n478
  );


  nor
  g748
  (
    n788,
    n471,
    n598,
    n490,
    n673
  );


  nor
  g749
  (
    n857,
    n604,
    n475,
    n631,
    n589
  );


  xor
  g750
  (
    n761,
    n588,
    n732,
    n451,
    n484
  );


  xor
  g751
  (
    n856,
    n645,
    n484,
    n728,
    n480
  );


  xnor
  g752
  (
    n942,
    n590,
    n620,
    n488,
    n443
  );


  xor
  g753
  (
    n811,
    n611,
    n623,
    n657,
    n690
  );


  or
  g754
  (
    n762,
    n653,
    n442,
    n463,
    n458
  );


  xor
  g755
  (
    n828,
    n692,
    n664,
    n643,
    n609
  );


  and
  g756
  (
    n826,
    n580,
    n662,
    n658,
    n617
  );


  nor
  g757
  (
    n890,
    n472,
    n731,
    n640,
    n614
  );


  xor
  g758
  (
    n944,
    n613,
    n433,
    n472,
    n597
  );


  or
  g759
  (
    n906,
    n699,
    n686,
    n587,
    n729
  );


  xor
  g760
  (
    KeyWire_0_50,
    n598,
    n730,
    n639,
    n695
  );


  nor
  g761
  (
    n795,
    n649,
    n665,
    n630,
    n706
  );


  and
  g762
  (
    n936,
    n463,
    n607,
    n731,
    n643
  );


  nor
  g763
  (
    n798,
    n618,
    n656,
    n446,
    n603
  );


  xnor
  g764
  (
    n924,
    n436,
    n735,
    n733,
    n585
  );


  or
  g765
  (
    n755,
    n699,
    n652,
    n472,
    n677
  );


  nand
  g766
  (
    n872,
    n698,
    n159,
    n662,
    n605
  );


  nor
  g767
  (
    n742,
    n631,
    n680,
    n661,
    n648
  );


  xnor
  g768
  (
    n931,
    n658,
    n622,
    n713,
    n451
  );


  nor
  g769
  (
    n844,
    n585,
    n669,
    n735,
    n639
  );


  xor
  g770
  (
    KeyWire_0_5,
    n458,
    n440,
    n645,
    n456
  );


  and
  g771
  (
    n951,
    n481,
    n690,
    n487,
    n594
  );


  nor
  g772
  (
    n747,
    n649,
    n630,
    n593,
    n638
  );


  nand
  g773
  (
    n852,
    n652,
    n473,
    n470,
    n589
  );


  xor
  g774
  (
    n881,
    n473,
    n723,
    n625,
    n734
  );


  nand
  g775
  (
    n917,
    n675,
    n660,
    n640,
    n635
  );


  xor
  g776
  (
    n947,
    n687,
    n739,
    n447,
    n621
  );


  xor
  g777
  (
    n938,
    n478,
    n629,
    n476,
    n461
  );


  nor
  g778
  (
    n803,
    n472,
    n648,
    n602
  );


  nand
  g779
  (
    n941,
    n482,
    n632,
    n437,
    n646
  );


  or
  g780
  (
    n901,
    n461,
    n465,
    n582,
    n659
  );


  xor
  g781
  (
    n770,
    n632,
    n455,
    n474,
    n623
  );


  xnor
  g782
  (
    n905,
    n461,
    n488,
    n730,
    n669
  );


  nor
  g783
  (
    n751,
    n474,
    n726,
    n711,
    n668
  );


  or
  g784
  (
    n922,
    n708,
    n710,
    n722,
    n467
  );


  xor
  g785
  (
    n842,
    n682,
    n468,
    n584,
    n712
  );


  nand
  g786
  (
    n861,
    n608,
    n678,
    n696,
    n433
  );


  and
  g787
  (
    n833,
    n701,
    n609,
    n466,
    n624
  );


  and
  g788
  (
    n900,
    n666,
    n444,
    n489,
    n160
  );


  nand
  g789
  (
    n948,
    n675,
    n606,
    n637,
    n670
  );


  nor
  g790
  (
    KeyWire_0_37,
    n678,
    n160,
    n674,
    n599
  );


  and
  g791
  (
    n949,
    n434,
    n696,
    n453,
    n645
  );


  xnor
  g792
  (
    n836,
    n732,
    n704,
    n734,
    n606
  );


  nand
  g793
  (
    n760,
    n716,
    n698,
    n679,
    n673
  );


  xor
  g794
  (
    n766,
    n452,
    n600,
    n691,
    n708
  );


  xnor
  g795
  (
    n800,
    n598,
    n700,
    n449,
    n738
  );


  nand
  g796
  (
    n779,
    n710,
    n586,
    n441,
    n696
  );


  and
  g797
  (
    n777,
    n455,
    n441,
    n629,
    n703
  );


  nand
  g798
  (
    n909,
    n585,
    n674,
    n490,
    n626
  );


  nand
  g799
  (
    n837,
    n160,
    n625,
    n483
  );


  nor
  g800
  (
    n904,
    n444,
    n439,
    n459,
    n638
  );


  nand
  g801
  (
    KeyWire_0_0,
    n464,
    n691,
    n723,
    n581
  );


  nand
  g802
  (
    KeyWire_0_43,
    n469,
    n605,
    n738,
    n636
  );


  xnor
  g803
  (
    n865,
    n477,
    n597,
    n709,
    n716
  );


  nor
  g804
  (
    n939,
    n708,
    n644,
    n669,
    n589
  );


  nor
  g805
  (
    n932,
    n718,
    n440,
    n714,
    n583
  );


  xnor
  g806
  (
    n785,
    n651,
    n449,
    n655,
    n694
  );


  nand
  g807
  (
    n749,
    n606,
    n432,
    n730,
    n677
  );


  and
  g808
  (
    n802,
    n710,
    n468,
    n707,
    n477
  );


  and
  g809
  (
    n822,
    n468,
    n456,
    n440,
    n641
  );


  and
  g810
  (
    n748,
    n703,
    n453,
    n434,
    n432
  );


  xnor
  g811
  (
    n843,
    n436,
    n450,
    n595,
    n712
  );


  or
  g812
  (
    n792,
    n627,
    n485,
    n452,
    n474
  );


  and
  g813
  (
    n817,
    n628,
    n726,
    n596,
    n729
  );


  nor
  g814
  (
    n758,
    n700,
    n158,
    n716,
    n602
  );


  nand
  g815
  (
    n873,
    n705,
    n434,
    n462,
    n654
  );


  or
  g816
  (
    n896,
    n444,
    n435,
    n436,
    n642
  );


  nor
  g817
  (
    n794,
    n637,
    n620,
    n724,
    n583
  );


  or
  g818
  (
    KeyWire_0_1,
    n706,
    n589,
    n692,
    n694
  );


  and
  g819
  (
    n864,
    n657,
    n682,
    n640,
    n590
  );


  nor
  g820
  (
    n831,
    n474,
    n439,
    n660,
    n647
  );


  and
  g821
  (
    n916,
    n450,
    n596,
    n672,
    n693
  );


  or
  g822
  (
    n850,
    n486,
    n720,
    n630,
    n469
  );


  xor
  g823
  (
    n952,
    n157,
    n728,
    n717,
    n442
  );


  and
  g824
  (
    n888,
    n442,
    n157,
    n699,
    n443
  );


  xnor
  g825
  (
    n889,
    n653,
    n678,
    n679,
    n623
  );


  xnor
  g826
  (
    n883,
    n477,
    n595,
    n715,
    n707
  );


  and
  g827
  (
    n809,
    n628,
    n702,
    n686,
    n637
  );


  xnor
  g828
  (
    n913,
    n603,
    n487,
    n612,
    n645
  );


  nand
  g829
  (
    n899,
    n698,
    n715,
    n473,
    n686
  );


  or
  g830
  (
    n845,
    n667,
    n455,
    n650,
    n711
  );


  nand
  g831
  (
    n744,
    n731,
    n612,
    n688,
    n448
  );


  and
  g832
  (
    n866,
    n593,
    n703,
    n483,
    n449
  );


  or
  g833
  (
    n765,
    n714,
    n619,
    n691,
    n471
  );


  xnor
  g834
  (
    n825,
    n588,
    n615,
    n159,
    n694
  );


  xnor
  g835
  (
    n767,
    n432,
    n666,
    n622,
    n445
  );


  nor
  g836
  (
    n935,
    n711,
    n621,
    n618,
    n446
  );


  xor
  g837
  (
    n875,
    n734,
    n460,
    n674,
    n727
  );


  nor
  g838
  (
    n781,
    n433,
    n722,
    n582,
    n616
  );


  xor
  g839
  (
    n847,
    n663,
    n739,
    n633,
    n490
  );


  nor
  g840
  (
    n898,
    n608,
    n688,
    n698,
    n596
  );


  xnor
  g841
  (
    n928,
    n158,
    n159,
    n678,
    n695
  );


  xor
  g842
  (
    n943,
    n603,
    n671,
    n475,
    n470
  );


  and
  g843
  (
    n926,
    n482,
    n624,
    n460,
    n715
  );


  nor
  g844
  (
    n764,
    n700,
    n464,
    n626,
    n673
  );


  and
  g845
  (
    n839,
    n658,
    n685,
    n707,
    n729
  );


  and
  g846
  (
    n745,
    n654,
    n158,
    n597,
    n467
  );


  nor
  g847
  (
    n884,
    n668,
    n656,
    n701,
    n726
  );


  and
  g848
  (
    n915,
    n458,
    n663,
    n709,
    n731
  );


  and
  g849
  (
    n750,
    n459,
    n466,
    n446,
    n644
  );


  nor
  g850
  (
    n920,
    n656,
    n609,
    n708,
    n685
  );


  xnor
  g851
  (
    n829,
    n445,
    n438,
    n621,
    n634
  );


  nand
  g852
  (
    n893,
    n651,
    n719,
    n725,
    n652
  );


  or
  g853
  (
    n927,
    n480,
    n691,
    n634,
    n668
  );


  xor
  g854
  (
    n911,
    n622,
    n706,
    n650,
    n671
  );


  or
  g855
  (
    n880,
    n604,
    n627,
    n633,
    n479
  );


  xnor
  g856
  (
    n937,
    n650,
    n685,
    n480,
    n590
  );


  and
  g857
  (
    n955,
    n466,
    n661,
    n687,
    n448
  );


  nand
  g858
  (
    KeyWire_0_31,
    n485,
    n671,
    n445,
    n627
  );


  xor
  g859
  (
    n854,
    n659,
    n733,
    n719,
    n594
  );


  xnor
  g860
  (
    n754,
    n489,
    n467,
    n628,
    n692
  );


  nand
  g861
  (
    n855,
    n602,
    n443,
    n692,
    n670
  );


  xor
  g862
  (
    n946,
    n587,
    n663,
    n601,
    n651
  );


  or
  g863
  (
    n768,
    n720,
    n448,
    n716,
    n687
  );


  xnor
  g864
  (
    n796,
    n469,
    n591,
    n624,
    n482
  );


  xor
  g865
  (
    n862,
    n664,
    n617,
    n614,
    n482
  );


  xnor
  g866
  (
    n786,
    n677,
    n647,
    n437,
    n735
  );


  nand
  g867
  (
    n806,
    n450,
    n459,
    n739,
    n586
  );


  or
  g868
  (
    n858,
    n592,
    n605,
    n632,
    n736
  );


  xnor
  g869
  (
    n835,
    n438,
    n736,
    n584,
    n681
  );


  xor
  g870
  (
    n940,
    n457,
    n465,
    n456,
    n712
  );


  nand
  g871
  (
    n776,
    n641,
    n637,
    n689,
    n681
  );


  xnor
  g872
  (
    n780,
    n683,
    n705,
    n663,
    n638
  );


  nor
  g873
  (
    KeyWire_0_22,
    n462,
    n598,
    n656,
    n438
  );


  xnor
  g874
  (
    n756,
    n486,
    n675,
    n697,
    n458
  );


  nand
  g875
  (
    n810,
    n667,
    n724,
    n647,
    n661
  );


  nand
  g876
  (
    n910,
    n654,
    n676,
    n439,
    n592
  );


  and
  g877
  (
    n801,
    n618,
    n581,
    n706,
    n653
  );


  xor
  g878
  (
    n746,
    n462,
    n486,
    n728,
    n680
  );


  xnor
  g879
  (
    n790,
    n619,
    n487,
    n479,
    n488
  );


  nand
  g880
  (
    n895,
    n730,
    n608,
    n160,
    n649
  );


  xnor
  g881
  (
    n773,
    n704,
    n665,
    n584,
    n657
  );


  xnor
  g882
  (
    n821,
    n441,
    n631,
    n599,
    n435
  );


  nand
  g883
  (
    n805,
    n666,
    n591,
    n627,
    n435
  );


  nor
  g884
  (
    n902,
    n648,
    n596,
    n447,
    n683
  );


  xnor
  g885
  (
    n763,
    n487,
    n693,
    n737,
    n646
  );


  and
  g886
  (
    n954,
    n712,
    n459,
    n463,
    n460
  );


  xnor
  g887
  (
    n757,
    n595,
    n684,
    n445,
    n473
  );


  or
  g888
  (
    n892,
    n626,
    n697,
    n469,
    n452
  );


  xnor
  g889
  (
    n818,
    n713,
    n736,
    n722,
    n738
  );


  xor
  g890
  (
    n897,
    n727,
    n486,
    n737,
    n464
  );


  nor
  g891
  (
    n885,
    n707,
    n436,
    n639,
    n479
  );


  and
  g892
  (
    n782,
    n587,
    n453,
    n684,
    n702
  );


  and
  g893
  (
    n769,
    n705,
    n684,
    n471,
    n653
  );


  and
  g894
  (
    n840,
    n628,
    n672,
    n709,
    n465
  );


  or
  g895
  (
    n812,
    n648,
    n636,
    n618,
    n735
  );


  and
  g896
  (
    n808,
    n452,
    n673,
    n635,
    n455
  );


  nand
  g897
  (
    n874,
    n732,
    n672,
    n642,
    n733
  );


  xnor
  g898
  (
    n807,
    n674,
    n454,
    n467,
    n687
  );


  and
  g899
  (
    n894,
    n639,
    n670,
    n601,
    n158
  );


  nor
  g900
  (
    n848,
    n689,
    n642,
    n620,
    n703
  );


  xor
  g901
  (
    n876,
    n649,
    n655,
    n454,
    n464
  );


  nand
  g902
  (
    n891,
    n668,
    n438,
    n442,
    n433
  );


  and
  g903
  (
    n741,
    n723,
    n583,
    n727,
    n591
  );


  nor
  g904
  (
    n834,
    n644,
    n646,
    n447,
    n481
  );


  xor
  g905
  (
    n934,
    n721,
    n713,
    n470,
    n623
  );


  and
  g906
  (
    n793,
    n457,
    n679,
    n489,
    n655
  );


  or
  g907
  (
    n860,
    n586,
    n465,
    n485,
    n661
  );


  and
  g908
  (
    n919,
    n441,
    n449,
    n599,
    n592
  );


  or
  g909
  (
    n783,
    n634,
    n481,
    n591,
    n711
  );


  or
  g910
  (
    n933,
    n585,
    n613,
    n654,
    n609
  );


  xnor
  g911
  (
    n830,
    n593,
    n700,
    n737,
    n600
  );


  xor
  g912
  (
    n957,
    n681,
    n710,
    n715,
    n714
  );


  xnor
  g913
  (
    n799,
    n660,
    n488,
    n671,
    n676
  );


  nor
  g914
  (
    n878,
    n737,
    n603,
    n607,
    n475
  );


  and
  g915
  (
    n771,
    n453,
    n699,
    n439,
    n484
  );


  nand
  g916
  (
    n797,
    n594,
    n580,
    n595,
    n582
  );


  and
  g917
  (
    n908,
    n689,
    n662,
    n659,
    n479
  );


  or
  g918
  (
    n789,
    n476,
    n633,
    n664,
    n581
  );


  xor
  g919
  (
    n870,
    n630,
    n480,
    n647,
    n688
  );


  xnor
  g920
  (
    n868,
    n670,
    n625,
    n629,
    n484
  );


  nand
  g921
  (
    n787,
    n640,
    n718,
    n717,
    n729
  );


  or
  g922
  (
    n841,
    n440,
    n701,
    n723,
    n621
  );


  and
  g923
  (
    n743,
    n468,
    n434,
    n718,
    n582
  );


  and
  g924
  (
    n914,
    n680,
    n739,
    n695,
    n481
  );


  and
  g925
  (
    n983,
    n824,
    n767,
    n928,
    n868
  );


  and
  g926
  (
    n979,
    n799,
    n895,
    n893,
    n952
  );


  xor
  g927
  (
    n973,
    n810,
    n942,
    n936,
    n919
  );


  or
  g928
  (
    n960,
    n842,
    n807,
    n778,
    n918
  );


  nor
  g929
  (
    n1013,
    n814,
    n782,
    n945,
    n948
  );


  nor
  g930
  (
    n964,
    n761,
    n836,
    n950,
    n941
  );


  or
  g931
  (
    n971,
    n780,
    n932,
    n917,
    n774
  );


  nor
  g932
  (
    n965,
    n783,
    n884,
    n921,
    n853
  );


  xor
  g933
  (
    n997,
    n852,
    n813,
    n869,
    n896
  );


  xor
  g934
  (
    n989,
    n792,
    n885,
    n907,
    n944
  );


  nor
  g935
  (
    n966,
    n832,
    n851,
    n950,
    n938
  );


  and
  g936
  (
    n975,
    n882,
    n881,
    n771,
    n891
  );


  nor
  g937
  (
    n990,
    n957,
    n759,
    n887,
    n827
  );


  nor
  g938
  (
    n995,
    n945,
    n826,
    n935,
    n812
  );


  xnor
  g939
  (
    n976,
    n776,
    n809,
    n946,
    n784
  );


  or
  g940
  (
    n1011,
    n841,
    n937,
    n769,
    n837
  );


  xor
  g941
  (
    n982,
    n954,
    n899,
    n839,
    n931
  );


  xnor
  g942
  (
    n1004,
    n788,
    n828,
    n930,
    n938
  );


  nand
  g943
  (
    n968,
    n875,
    n324,
    n956,
    n903
  );


  nor
  g944
  (
    n998,
    n858,
    n889,
    n805,
    n900
  );


  or
  g945
  (
    n980,
    n855,
    n872,
    n854,
    n905
  );


  xnor
  g946
  (
    n963,
    n946,
    n864,
    n949,
    n951
  );


  xor
  g947
  (
    n999,
    n927,
    n867,
    n877,
    n796
  );


  or
  g948
  (
    n1000,
    n838,
    n890,
    n932,
    n870
  );


  nor
  g949
  (
    KeyWire_0_49,
    n781,
    n791,
    n760,
    n808
  );


  or
  g950
  (
    n981,
    n862,
    n848,
    n786,
    n873
  );


  xnor
  g951
  (
    KeyWire_0_29,
    n821,
    n910,
    n806,
    n940
  );


  nand
  g952
  (
    n986,
    n772,
    n789,
    n757,
    n324
  );


  nor
  g953
  (
    n970,
    n888,
    n770,
    n795,
    n787
  );


  xor
  g954
  (
    n1002,
    n755,
    n897,
    n941,
    n947
  );


  nor
  g955
  (
    n969,
    n880,
    n871,
    n861,
    n804
  );


  xor
  g956
  (
    n988,
    n816,
    n773,
    n825,
    n785
  );


  xnor
  g957
  (
    n984,
    n798,
    n777,
    n878,
    n811
  );


  or
  g958
  (
    n978,
    n925,
    n765,
    n764,
    n833
  );


  and
  g959
  (
    n1015,
    n859,
    n819,
    n883,
    n803
  );


  xnor
  g960
  (
    n1008,
    n955,
    n956,
    n797,
    n834
  );


  nor
  g961
  (
    n961,
    n860,
    n914,
    n754,
    n953
  );


  xnor
  g962
  (
    n991,
    n840,
    n763,
    n911,
    n944
  );


  or
  g963
  (
    n972,
    n955,
    n902,
    n845,
    n324
  );


  or
  g964
  (
    n977,
    n779,
    n915,
    n904,
    n879
  );


  or
  g965
  (
    KeyWire_0_46,
    n857,
    n892,
    n898,
    n913
  );


  or
  g966
  (
    n1003,
    n933,
    n766,
    n849,
    n912
  );


  or
  g967
  (
    n974,
    n934,
    n802,
    n758,
    n943
  );


  nor
  g968
  (
    n1007,
    n909,
    n957,
    n906,
    n937
  );


  nand
  g969
  (
    n962,
    n936,
    n790,
    n843,
    n948
  );


  and
  g970
  (
    n993,
    n929,
    n924,
    n822,
    n947
  );


  xor
  g971
  (
    n959,
    n863,
    n876,
    n856,
    n866
  );


  nand
  g972
  (
    n958,
    n931,
    n927,
    n952,
    n916
  );


  nor
  g973
  (
    n1001,
    n957,
    n901,
    n933,
    n942
  );


  or
  g974
  (
    n985,
    n847,
    n823,
    n835,
    n886
  );


  xnor
  g975
  (
    KeyWire_0_16,
    n926,
    n844,
    n831,
    n928
  );


  nor
  g976
  (
    n1009,
    n939,
    n954,
    n850,
    n957
  );


  nand
  g977
  (
    n987,
    n930,
    n756,
    n951,
    n815
  );


  or
  g978
  (
    n1006,
    n768,
    n920,
    n940,
    n846
  );


  and
  g979
  (
    n992,
    n801,
    n953,
    n817,
    n820
  );


  nor
  g980
  (
    n1005,
    n934,
    n894,
    n818,
    n935
  );


  xor
  g981
  (
    n1016,
    n908,
    n794,
    n923,
    n874
  );


  nor
  g982
  (
    n1012,
    n929,
    n829,
    n800,
    n775
  );


  xor
  g983
  (
    n1014,
    n949,
    n830,
    n793,
    n922
  );


  and
  g984
  (
    n994,
    n865,
    n939,
    n943,
    n762
  );


  or
  g985
  (
    n1025,
    n1007,
    n1003,
    n981,
    n982
  );


  nand
  g986
  (
    n1028,
    n972,
    n1002,
    n975,
    n971
  );


  and
  g987
  (
    n1019,
    n979,
    n1006,
    n994,
    n985
  );


  nor
  g988
  (
    n1030,
    n1001,
    n1015,
    n1010,
    n966
  );


  xor
  g989
  (
    n1032,
    n973,
    n987,
    n1017,
    n1012
  );


  or
  g990
  (
    n1027,
    n963,
    n977,
    n1014,
    n978
  );


  xnor
  g991
  (
    n1023,
    n980,
    n1008,
    n961,
    n988
  );


  and
  g992
  (
    n1020,
    n960,
    n1004,
    n1005,
    n990
  );


  nand
  g993
  (
    n1024,
    n1016,
    n969,
    n995,
    n970
  );


  xnor
  g994
  (
    n1018,
    n1000,
    n984,
    n958,
    n967
  );


  nor
  g995
  (
    n1031,
    n1009,
    n976,
    n991,
    n999
  );


  nand
  g996
  (
    n1029,
    n992,
    n989,
    n983,
    n959
  );


  or
  g997
  (
    n1021,
    n965,
    n968,
    n996,
    n962
  );


  or
  g998
  (
    n1026,
    n986,
    n1013,
    n974,
    n997
  );


  xor
  g999
  (
    n1022,
    n964,
    n1011,
    n998,
    n993
  );


  xnor
  KeyGate_0_0
  (
    n867,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n887,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n157,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n144,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n422,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n778,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n716,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n392,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n240,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n498,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n214,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n503,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n562,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n547,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n150,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n337,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n1017,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n189,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n377,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n136,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n679,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n238,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n849,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n262,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n307,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n199,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n437,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n621,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n517,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n967,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n574,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n853,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n598,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n35,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n476,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n55,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n700,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n930,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n491,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n536,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n241,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n447,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n529,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n815,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n179,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n577,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n996,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n293,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n851,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n1010,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n871,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n670,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n502,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n707,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n514,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n327,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n73,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n590,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n59,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n644,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n201,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n339,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n572,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n277,
    KeyNOTWire_0_63
  );


endmodule

