// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_2749_29_1 written by SynthGen on 2021/06/15 15:06:09
module Stat_2749_29_1( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25,
 n2466, n2459, n2515, n2748, n2757, n2770, n2755, n2774,
 n2759, n2742, n2766, n2747, n2773, n2743, n2772, n2761,
 n2749, n2752, n2763, n2746, n2762, n2768, n2758, n2741,
 n2753, n2764, n2751, n2767, n2750, n2756, n2745, n2769,
 n2760, n2765, n2744, n2754, n2771);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25;

output n2466, n2459, n2515, n2748, n2757, n2770, n2755, n2774,
 n2759, n2742, n2766, n2747, n2773, n2743, n2772, n2761,
 n2749, n2752, n2763, n2746, n2762, n2768, n2758, n2741,
 n2753, n2764, n2751, n2767, n2750, n2756, n2745, n2769,
 n2760, n2765, n2744, n2754, n2771;

wire n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
 n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
 n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
 n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
 n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
 n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
 n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
 n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
 n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
 n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
 n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
 n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
 n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
 n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
 n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
 n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
 n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
 n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
 n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
 n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
 n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
 n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
 n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
 n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
 n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
 n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
 n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
 n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
 n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
 n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
 n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
 n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
 n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
 n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
 n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
 n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
 n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
 n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
 n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
 n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
 n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
 n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
 n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
 n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
 n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
 n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
 n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
 n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
 n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
 n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
 n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
 n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
 n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
 n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
 n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
 n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
 n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
 n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
 n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
 n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
 n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
 n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
 n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
 n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
 n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
 n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
 n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
 n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
 n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
 n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
 n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
 n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
 n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
 n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
 n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
 n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
 n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
 n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
 n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
 n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
 n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
 n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
 n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
 n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
 n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
 n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
 n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
 n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
 n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
 n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
 n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
 n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
 n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
 n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
 n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
 n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
 n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
 n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
 n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
 n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
 n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
 n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
 n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
 n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
 n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
 n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
 n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
 n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
 n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
 n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
 n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
 n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
 n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
 n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
 n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
 n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
 n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
 n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
 n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
 n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
 n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
 n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
 n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
 n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
 n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
 n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
 n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
 n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
 n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
 n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
 n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
 n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
 n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
 n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
 n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
 n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
 n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
 n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
 n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
 n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
 n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
 n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
 n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
 n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
 n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
 n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
 n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
 n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
 n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
 n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
 n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
 n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
 n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
 n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
 n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
 n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
 n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
 n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
 n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
 n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
 n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
 n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
 n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
 n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
 n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
 n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
 n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
 n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
 n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
 n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
 n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
 n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
 n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
 n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
 n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
 n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
 n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
 n2458, n2460, n2461, n2462, n2463, n2464, n2465, n2467,
 n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
 n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
 n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
 n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
 n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
 n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2516,
 n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
 n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
 n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
 n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
 n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556,
 n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
 n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
 n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
 n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
 n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596,
 n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
 n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
 n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
 n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
 n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
 n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
 n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
 n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
 n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
 n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
 n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
 n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
 n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
 n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
 n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
 n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
 n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
 n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740;

buf  g0 (n88, n12);
buf  g1 (n105, n9);
not  g2 (n90, n13);
buf  g3 (n106, n9);
buf  g4 (n92, n19);
buf  g5 (n63, n7);
not  g6 (n57, n13);
buf  g7 (n77, n5);
not  g8 (n66, n2);
not  g9 (n85, n6);
buf  g10 (n50, n16);
not  g11 (n47, n4);
buf  g12 (n40, n19);
not  g13 (n51, n4);
buf  g14 (n84, n15);
not  g15 (n37, n4);
not  g16 (n30, n5);
not  g17 (n73, n21);
not  g18 (n75, n19);
not  g19 (n97, n18);
buf  g20 (n98, n3);
buf  g21 (n76, n8);
buf  g22 (n48, n8);
buf  g23 (n46, n6);
buf  g24 (n29, n3);
buf  g25 (n100, n20);
not  g26 (n86, n13);
not  g27 (n42, n2);
buf  g28 (n59, n12);
not  g29 (n81, n17);
not  g30 (n104, n18);
buf  g31 (n55, n14);
buf  g32 (n53, n6);
buf  g33 (n83, n14);
not  g34 (n28, n20);
buf  g35 (n54, n14);
not  g36 (n101, n3);
buf  g37 (n33, n9);
not  g38 (n45, n7);
buf  g39 (n64, n5);
not  g40 (n102, n17);
not  g41 (n89, n2);
not  g42 (n44, n9);
not  g43 (n79, n15);
not  g44 (n68, n1);
not  g45 (n43, n10);
not  g46 (n74, n1);
not  g47 (n65, n18);
buf  g48 (n60, n16);
not  g49 (n26, n12);
buf  g50 (n34, n5);
buf  g51 (n35, n19);
buf  g52 (n52, n15);
buf  g53 (n78, n17);
buf  g54 (n71, n7);
buf  g55 (n31, n1);
not  g56 (n61, n17);
not  g57 (n36, n14);
buf  g58 (n38, n1);
buf  g59 (n87, n11);
not  g60 (n41, n12);
buf  g61 (n67, n11);
not  g62 (n70, n3);
not  g63 (n94, n10);
buf  g64 (n96, n4);
buf  g65 (n103, n18);
buf  g66 (n39, n16);
buf  g67 (n49, n11);
not  g68 (n32, n10);
not  g69 (n91, n16);
not  g70 (n93, n20);
not  g71 (n95, n13);
not  g72 (n99, n2);
not  g73 (n62, n7);
buf  g74 (n58, n11);
buf  g75 (n82, n20);
buf  g76 (n80, n8);
not  g77 (n69, n15);
buf  g78 (n72, n10);
buf  g79 (n56, n8);
buf  g80 (n27, n6);
buf  g81 (n330, n60);
not  g82 (n410, n32);
not  g83 (n411, n30);
buf  g84 (n159, n36);
not  g85 (n109, n81);
buf  g86 (n336, n92);
buf  g87 (n230, n36);
not  g88 (n279, n45);
buf  g89 (n254, n46);
buf  g90 (n396, n43);
buf  g91 (n133, n44);
not  g92 (n340, n96);
buf  g93 (n256, n90);
buf  g94 (n343, n102);
not  g95 (n223, n39);
not  g96 (n124, n101);
not  g97 (n320, n95);
buf  g98 (n354, n49);
buf  g99 (n355, n104);
not  g100 (n307, n37);
not  g101 (n260, n85);
not  g102 (n383, n80);
buf  g103 (n392, n104);
buf  g104 (n333, n46);
buf  g105 (n132, n94);
not  g106 (n121, n95);
buf  g107 (n128, n47);
buf  g108 (n202, n50);
buf  g109 (n306, n74);
buf  g110 (n193, n90);
not  g111 (n118, n47);
buf  g112 (n135, n44);
buf  g113 (n196, n99);
buf  g114 (n273, n46);
not  g115 (n235, n104);
not  g116 (n155, n76);
not  g117 (n368, n30);
buf  g118 (n374, n66);
not  g119 (n208, n40);
not  g120 (n263, n81);
not  g121 (n236, n86);
not  g122 (n324, n71);
buf  g123 (n421, n89);
buf  g124 (n394, n44);
not  g125 (n364, n43);
not  g126 (n420, n82);
buf  g127 (n348, n27);
buf  g128 (n220, n63);
buf  g129 (n422, n70);
not  g130 (n325, n52);
buf  g131 (n402, n77);
not  g132 (n321, n50);
buf  g133 (n184, n103);
buf  g134 (n219, n54);
not  g135 (n244, n56);
not  g136 (n268, n88);
buf  g137 (n391, n41);
not  g138 (n186, n99);
buf  g139 (n185, n35);
buf  g140 (n406, n79);
buf  g141 (n258, n58);
buf  g142 (n141, n99);
buf  g143 (n337, n78);
buf  g144 (n351, n52);
buf  g145 (n115, n64);
buf  g146 (n416, n42);
not  g147 (n366, n29);
buf  g148 (n281, n75);
buf  g149 (n180, n82);
buf  g150 (n187, n77);
not  g151 (n171, n89);
buf  g152 (n267, n101);
buf  g153 (n117, n70);
not  g154 (n203, n77);
not  g155 (n216, n80);
buf  g156 (n127, n75);
buf  g157 (n301, n49);
not  g158 (n151, n61);
buf  g159 (n309, n92);
buf  g160 (n123, n102);
buf  g161 (n249, n97);
not  g162 (n169, n96);
buf  g163 (n362, n86);
not  g164 (n125, n27);
not  g165 (n298, n72);
buf  g166 (n276, n67);
not  g167 (n190, n96);
not  g168 (n363, n66);
buf  g169 (n404, n62);
buf  g170 (n111, n63);
buf  g171 (n382, n63);
buf  g172 (n405, n92);
buf  g173 (n138, n26);
buf  g174 (n367, n53);
not  g175 (n308, n42);
not  g176 (n409, n87);
not  g177 (n142, n28);
buf  g178 (n126, n34);
buf  g179 (n418, n44);
buf  g180 (n311, n78);
not  g181 (n250, n67);
buf  g182 (n211, n47);
buf  g183 (n120, n59);
buf  g184 (n173, n104);
not  g185 (n417, n33);
buf  g186 (n357, n89);
not  g187 (n174, n42);
buf  g188 (n144, n31);
buf  g189 (n261, n51);
not  g190 (n122, n66);
buf  g191 (n361, n77);
buf  g192 (n365, n29);
buf  g193 (n304, n31);
not  g194 (n168, n48);
not  g195 (n302, n59);
not  g196 (n401, n76);
buf  g197 (n188, n49);
buf  g198 (n242, n37);
not  g199 (n269, n60);
buf  g200 (n257, n30);
buf  g201 (n136, n37);
not  g202 (n339, n38);
buf  g203 (n240, n50);
not  g204 (n214, n38);
buf  g205 (n295, n55);
buf  g206 (n114, n97);
not  g207 (n403, n55);
buf  g208 (n108, n64);
not  g209 (n386, n79);
not  g210 (n356, n86);
not  g211 (n318, n81);
buf  g212 (n177, n47);
not  g213 (n119, n65);
not  g214 (n413, n85);
not  g215 (n226, n88);
not  g216 (n253, n33);
buf  g217 (n369, n73);
buf  g218 (n234, n34);
buf  g219 (n229, n33);
buf  g220 (n389, n58);
buf  g221 (n313, n84);
not  g222 (n178, n90);
not  g223 (n210, n70);
buf  g224 (n205, n60);
buf  g225 (n310, n60);
buf  g226 (n189, n28);
buf  g227 (n238, n83);
not  g228 (n140, n76);
buf  g229 (n329, n98);
not  g230 (n378, n65);
buf  g231 (n291, n102);
buf  g232 (n283, n101);
buf  g233 (n160, n45);
not  g234 (n282, n29);
buf  g235 (n312, n49);
buf  g236 (n350, n32);
buf  g237 (n342, n91);
not  g238 (n262, n61);
buf  g239 (n370, n88);
buf  g240 (n259, n93);
buf  g241 (n194, n29);
not  g242 (n130, n62);
buf  g243 (n204, n68);
not  g244 (n266, n71);
not  g245 (n233, n41);
buf  g246 (n395, n68);
buf  g247 (n264, n69);
not  g248 (n148, n56);
not  g249 (n349, n69);
not  g250 (n317, n83);
buf  g251 (n110, n53);
not  g252 (n407, n74);
buf  g253 (n289, n69);
buf  g254 (n344, n64);
buf  g255 (n326, n80);
not  g256 (n284, n78);
buf  g257 (n373, n28);
not  g258 (n166, n32);
buf  g259 (n172, n35);
buf  g260 (n359, n68);
not  g261 (n247, n96);
not  g262 (n241, n57);
buf  g263 (n332, n83);
buf  g264 (n319, n64);
buf  g265 (n143, n55);
not  g266 (n314, n51);
buf  g267 (n360, n85);
buf  g268 (n248, n45);
buf  g269 (n182, n56);
buf  g270 (n290, n78);
buf  g271 (n346, n35);
not  g272 (n154, n54);
buf  g273 (n408, n94);
not  g274 (n165, n51);
not  g275 (n293, n65);
buf  g276 (n162, n98);
buf  g277 (n251, n98);
not  g278 (n224, n74);
buf  g279 (n137, n54);
not  g280 (n399, n100);
buf  g281 (n227, n84);
not  g282 (n419, n83);
buf  g283 (n222, n61);
not  g284 (n385, n70);
not  g285 (n153, n102);
not  g286 (n278, n100);
not  g287 (n334, n73);
buf  g288 (n287, n69);
buf  g289 (n305, n46);
not  g290 (n272, n36);
not  g291 (n371, n95);
buf  g292 (n175, n58);
not  g293 (n200, n90);
not  g294 (n397, n97);
buf  g295 (n294, n52);
buf  g296 (n280, n100);
not  g297 (n335, n45);
buf  g298 (n237, n42);
not  g299 (n163, n84);
buf  g300 (n331, n74);
not  g301 (n167, n99);
buf  g302 (n255, n38);
buf  g303 (n415, n39);
not  g304 (n164, n26);
buf  g305 (n183, n73);
not  g306 (n303, n27);
not  g307 (n381, n57);
not  g308 (n323, n65);
not  g309 (n379, n91);
buf  g310 (n412, n87);
buf  g311 (n400, n56);
buf  g312 (n372, n71);
buf  g313 (n129, n89);
not  g314 (n384, n75);
buf  g315 (n112, n35);
buf  g316 (n245, n75);
buf  g317 (n393, n63);
not  g318 (n116, n43);
buf  g319 (n288, n72);
not  g320 (n286, n91);
not  g321 (n158, n97);
buf  g322 (n156, n54);
buf  g323 (n265, n50);
not  g324 (n231, n36);
not  g325 (n145, n95);
buf  g326 (n358, n68);
not  g327 (n375, n103);
buf  g328 (n297, n28);
buf  g329 (n315, n48);
not  g330 (n414, n66);
buf  g331 (n218, n34);
not  g332 (n192, n85);
not  g333 (n191, n62);
not  g334 (n274, n93);
buf  g335 (n341, n87);
buf  g336 (n207, n94);
buf  g337 (n398, n61);
not  g338 (n387, n55);
not  g339 (n376, n38);
not  g340 (n328, n58);
buf  g341 (n139, n30);
not  g342 (n179, n48);
not  g343 (n345, n73);
buf  g344 (n292, n67);
not  g345 (n327, n98);
buf  g346 (n149, n81);
buf  g347 (n201, n59);
not  g348 (n161, n41);
not  g349 (n390, n51);
buf  g350 (n146, n82);
not  g351 (n107, n27);
buf  g352 (n195, n62);
not  g353 (n170, n79);
not  g354 (n181, n52);
not  g355 (n299, n37);
not  g356 (n388, n72);
buf  g357 (n232, n101);
buf  g358 (n296, n67);
buf  g359 (n217, n39);
buf  g360 (n277, n79);
buf  g361 (n197, n93);
buf  g362 (n199, n86);
not  g363 (n221, n41);
not  g364 (n252, n40);
not  g365 (n209, n92);
not  g366 (n338, n34);
not  g367 (n380, n57);
not  g368 (n131, n59);
buf  g369 (n134, n80);
not  g370 (n150, n103);
not  g371 (n215, n91);
not  g372 (n157, n31);
not  g373 (n147, n87);
not  g374 (n347, n53);
not  g375 (n352, n31);
not  g376 (n228, n100);
buf  g377 (n212, n43);
buf  g378 (n316, n40);
not  g379 (n243, n53);
not  g380 (n152, n76);
not  g381 (n246, n33);
not  g382 (n271, n88);
not  g383 (n300, n40);
not  g384 (n322, n82);
buf  g385 (n377, n94);
not  g386 (n225, n32);
buf  g387 (n113, n26);
not  g388 (n176, n93);
not  g389 (n353, n39);
buf  g390 (n239, n71);
not  g391 (n206, n72);
not  g392 (n275, n26);
not  g393 (n198, n84);
not  g394 (n270, n48);
not  g395 (n213, n57);
not  g396 (n285, n103);
not  g397 (n651, n303);
not  g398 (n1268, n407);
not  g399 (n1030, n240);
not  g400 (n886, n151);
not  g401 (n1204, n239);
buf  g402 (n1128, n374);
not  g403 (n1091, n174);
buf  g404 (n1545, n392);
buf  g405 (n798, n313);
not  g406 (n1044, n252);
not  g407 (n1616, n265);
buf  g408 (n1640, n362);
not  g409 (n1067, n404);
not  g410 (n496, n202);
not  g411 (n1312, n171);
not  g412 (n1353, n421);
not  g413 (n1038, n107);
buf  g414 (n581, n142);
not  g415 (n826, n238);
not  g416 (n1025, n331);
buf  g417 (n1114, n335);
not  g418 (n1408, n419);
not  g419 (n836, n383);
not  g420 (n915, n397);
buf  g421 (n674, n166);
not  g422 (n440, n414);
not  g423 (n1051, n218);
buf  g424 (n1306, n171);
not  g425 (n1130, n140);
not  g426 (n1646, n217);
buf  g427 (n1533, n321);
buf  g428 (n1496, n163);
buf  g429 (n788, n196);
buf  g430 (n525, n177);
not  g431 (n743, n253);
buf  g432 (n438, n346);
buf  g433 (n458, n333);
not  g434 (n775, n379);
not  g435 (n617, n294);
buf  g436 (n1278, n185);
not  g437 (n1056, n390);
not  g438 (n938, n337);
buf  g439 (n1052, n359);
buf  g440 (n570, n404);
not  g441 (n1347, n367);
not  g442 (n907, n348);
not  g443 (n1265, n161);
buf  g444 (n1614, n223);
buf  g445 (n999, n187);
buf  g446 (n1293, n157);
not  g447 (n1491, n220);
buf  g448 (n538, n211);
not  g449 (n585, n322);
buf  g450 (n903, n145);
buf  g451 (n1003, n351);
not  g452 (n1463, n277);
buf  g453 (n1097, n347);
buf  g454 (n856, n299);
not  g455 (n1156, n193);
buf  g456 (n1064, n410);
buf  g457 (n771, n184);
buf  g458 (n567, n228);
buf  g459 (n919, n395);
buf  g460 (n709, n255);
not  g461 (n1193, n280);
not  g462 (n1512, n284);
buf  g463 (n1477, n250);
not  g464 (n1604, n351);
not  g465 (n1664, n301);
not  g466 (n618, n355);
buf  g467 (n573, n170);
buf  g468 (n1569, n134);
buf  g469 (n1652, n310);
buf  g470 (n610, n170);
buf  g471 (n1279, n198);
buf  g472 (n1162, n197);
not  g473 (n1473, n316);
buf  g474 (n1682, n247);
buf  g475 (n833, n131);
not  g476 (n1553, n416);
buf  g477 (n1529, n225);
not  g478 (n435, n300);
buf  g479 (n1430, n380);
buf  g480 (n888, n384);
not  g481 (n948, n162);
buf  g482 (n757, n116);
buf  g483 (n582, n288);
buf  g484 (n1208, n386);
not  g485 (n443, n270);
not  g486 (n1191, n293);
buf  g487 (n656, n365);
not  g488 (n866, n173);
buf  g489 (n859, n267);
buf  g490 (n428, n123);
not  g491 (n1339, n360);
buf  g492 (n1543, n222);
not  g493 (n1550, n401);
not  g494 (n1078, n189);
buf  g495 (n1443, n261);
buf  g496 (n1133, n114);
buf  g497 (n801, n379);
buf  g498 (n532, n307);
not  g499 (n621, n376);
not  g500 (n1547, n185);
buf  g501 (n1615, n265);
not  g502 (n1027, n301);
buf  g503 (n1618, n282);
buf  g504 (n764, n143);
buf  g505 (n1358, n200);
not  g506 (n1561, n395);
buf  g507 (n624, n224);
not  g508 (n756, n241);
not  g509 (n1313, n378);
not  g510 (n1062, n124);
buf  g511 (n975, n164);
not  g512 (n639, n107);
not  g513 (n664, n279);
not  g514 (n1511, n258);
buf  g515 (n1404, n357);
buf  g516 (n1612, n160);
buf  g517 (n1518, n264);
not  g518 (n831, n209);
not  g519 (n569, n385);
not  g520 (n1623, n392);
buf  g521 (n1455, n325);
buf  g522 (n1231, n205);
not  g523 (n998, n268);
buf  g524 (n1548, n175);
not  g525 (n464, n314);
buf  g526 (n1377, n274);
not  g527 (n712, n371);
buf  g528 (n1402, n192);
buf  g529 (n1409, n252);
buf  g530 (n970, n307);
not  g531 (n901, n165);
buf  g532 (n1461, n202);
buf  g533 (n657, n308);
not  g534 (n462, n197);
buf  g535 (n916, n236);
not  g536 (n855, n286);
not  g537 (n439, n312);
not  g538 (n746, n248);
buf  g539 (n1144, n261);
buf  g540 (n1571, n333);
not  g541 (n729, n299);
not  g542 (n1656, n268);
buf  g543 (n549, n133);
not  g544 (n1609, n109);
buf  g545 (n1648, n229);
not  g546 (n1601, n239);
buf  g547 (n1307, n361);
not  g548 (n1223, n335);
not  g549 (n542, n269);
not  g550 (n1387, n288);
not  g551 (n739, n326);
buf  g552 (n981, n359);
buf  g553 (n1102, n317);
buf  g554 (n1633, n340);
not  g555 (n1600, n410);
buf  g556 (n1281, n416);
buf  g557 (n780, n224);
buf  g558 (n620, n417);
buf  g559 (n1292, n321);
not  g560 (n654, n421);
not  g561 (n1254, n374);
buf  g562 (n1126, n366);
buf  g563 (n1369, n117);
buf  g564 (n425, n283);
not  g565 (n1450, n181);
not  g566 (n1579, n374);
buf  g567 (n1636, n233);
not  g568 (n518, n405);
buf  g569 (n1673, n385);
buf  g570 (n666, n406);
buf  g571 (n744, n270);
not  g572 (n619, n125);
not  g573 (n544, n177);
not  g574 (n734, n248);
buf  g575 (n1232, n419);
not  g576 (n885, n227);
not  g577 (n1419, n164);
not  g578 (n467, n375);
not  g579 (n1457, n259);
not  g580 (n471, n114);
not  g581 (n973, n195);
buf  g582 (n1053, n128);
not  g583 (n1414, n300);
not  g584 (n1163, n378);
not  g585 (n1176, n293);
buf  g586 (n936, n348);
not  g587 (n1017, n208);
buf  g588 (n1494, n236);
buf  g589 (n1077, n240);
buf  g590 (n926, n108);
buf  g591 (n1207, n417);
buf  g592 (n632, n378);
buf  g593 (n784, n405);
buf  g594 (n1337, n210);
buf  g595 (n1345, n169);
buf  g596 (n1079, n201);
buf  g597 (n898, n275);
buf  g598 (n884, n207);
buf  g599 (n1523, n377);
buf  g600 (n495, n253);
buf  g601 (n956, n337);
buf  g602 (n1197, n176);
not  g603 (n1563, n339);
buf  g604 (n929, n163);
buf  g605 (n1214, n120);
not  g606 (n1624, n388);
buf  g607 (n1593, n365);
buf  g608 (n1532, n206);
buf  g609 (n676, n358);
not  g610 (n1297, n314);
not  g611 (n1684, n213);
buf  g612 (n672, n243);
buf  g613 (n1479, n308);
buf  g614 (n670, n344);
not  g615 (n1177, n377);
not  g616 (n1088, n246);
buf  g617 (n1249, n241);
not  g618 (n700, n133);
buf  g619 (n953, n389);
not  g620 (n993, n195);
not  g621 (n842, n277);
not  g622 (n485, n236);
buf  g623 (n810, n269);
not  g624 (n1354, n115);
not  g625 (n1334, n269);
not  g626 (n447, n258);
not  g627 (n1273, n282);
not  g628 (n1438, n232);
buf  g629 (n730, n136);
buf  g630 (n942, n110);
buf  g631 (n1662, n216);
buf  g632 (n694, n415);
not  g633 (n701, n310);
buf  g634 (n1350, n411);
buf  g635 (n851, n236);
not  g636 (n850, n247);
buf  g637 (n1597, n139);
not  g638 (n590, n365);
buf  g639 (n1186, n346);
buf  g640 (n649, n120);
buf  g641 (n1531, n407);
buf  g642 (n1021, n323);
not  g643 (n1008, n414);
not  g644 (n1653, n400);
buf  g645 (n655, n394);
buf  g646 (n1175, n353);
buf  g647 (n1514, n413);
not  g648 (n1014, n110);
not  g649 (n691, n112);
not  g650 (n605, n203);
not  g651 (n935, n204);
not  g652 (n1433, n118);
not  g653 (n738, n363);
not  g654 (n1449, n279);
not  g655 (n545, n180);
buf  g656 (n586, n353);
not  g657 (n1559, n158);
buf  g658 (n943, n284);
not  g659 (n1210, n146);
buf  g660 (n1356, n233);
buf  g661 (n1309, n320);
buf  g662 (n1539, n206);
buf  g663 (n1493, n372);
not  g664 (n494, n209);
buf  g665 (n1229, n364);
buf  g666 (n722, n131);
buf  g667 (n1431, n297);
not  g668 (n524, n110);
not  g669 (n1454, n317);
not  g670 (n949, n353);
buf  g671 (n865, n227);
not  g672 (n977, n276);
buf  g673 (n1280, n276);
not  g674 (n768, n179);
not  g675 (n1425, n201);
not  g676 (n1002, n134);
buf  g677 (n776, n235);
buf  g678 (n578, n221);
not  g679 (n1150, n237);
not  g680 (n1073, n378);
buf  g681 (n1226, n167);
not  g682 (n1271, n128);
not  g683 (n1023, n418);
buf  g684 (n767, n168);
not  g685 (n719, n156);
not  g686 (n832, n109);
buf  g687 (n520, n108);
not  g688 (n1360, n198);
not  g689 (n910, n335);
not  g690 (n614, n161);
not  g691 (n733, n362);
not  g692 (n1185, n286);
not  g693 (n1215, n111);
buf  g694 (n1372, n209);
not  g695 (n822, n237);
buf  g696 (n1534, n380);
buf  g697 (n1109, n406);
buf  g698 (n1098, n350);
buf  g699 (n1211, n290);
buf  g700 (n952, n366);
buf  g701 (n976, n370);
not  g702 (n1535, n259);
buf  g703 (n627, n143);
not  g704 (n1467, n319);
buf  g705 (n1040, n313);
buf  g706 (n1359, n112);
buf  g707 (n747, n387);
not  g708 (n1606, n163);
buf  g709 (n1300, n326);
buf  g710 (n1287, n258);
buf  g711 (n1391, n413);
not  g712 (n1244, n206);
not  g713 (n1024, n303);
not  g714 (n1448, n403);
buf  g715 (n1240, n251);
not  g716 (n1367, n205);
not  g717 (n553, n222);
buf  g718 (n516, n256);
buf  g719 (n1153, n252);
buf  g720 (n1355, n247);
not  g721 (n1295, n173);
buf  g722 (n482, n207);
buf  g723 (n1198, n373);
buf  g724 (n1217, n125);
not  g725 (n896, n308);
not  g726 (n491, n157);
not  g727 (n797, n255);
buf  g728 (n1299, n284);
buf  g729 (n772, n191);
buf  g730 (n1241, n249);
buf  g731 (n1131, n395);
not  g732 (n1421, n194);
not  g733 (n1000, n393);
buf  g734 (n880, n152);
not  g735 (n1283, n259);
buf  g736 (n1630, n382);
buf  g737 (n720, n330);
not  g738 (n668, n200);
buf  g739 (n1272, n415);
not  g740 (n870, n355);
not  g741 (n1092, n324);
buf  g742 (n1143, n389);
not  g743 (n1351, n204);
not  g744 (n450, n167);
not  g745 (n812, n172);
not  g746 (n761, n158);
buf  g747 (n459, n134);
not  g748 (n890, n145);
buf  g749 (n1440, n292);
not  g750 (n827, n272);
not  g751 (n1558, n213);
buf  g752 (n1298, n399);
not  g753 (n1034, n245);
not  g754 (n522, n114);
not  g755 (n579, n336);
not  g756 (n873, n262);
buf  g757 (n1598, n295);
not  g758 (n1196, n342);
not  g759 (n1517, n294);
buf  g760 (n1560, n261);
not  g761 (n457, n395);
buf  g762 (n882, n307);
not  g763 (n592, n317);
buf  g764 (n1666, n295);
not  g765 (n1058, n363);
not  g766 (n714, n380);
buf  g767 (n1480, n242);
buf  g768 (n741, n108);
buf  g769 (n1031, n140);
not  g770 (n1575, n192);
not  g771 (n692, n152);
buf  g772 (n1263, n408);
not  g773 (n785, n371);
buf  g774 (n1610, n256);
buf  g775 (n753, n413);
buf  g776 (n1371, n366);
buf  g777 (n779, n150);
not  g778 (n623, n285);
not  g779 (n951, n214);
not  g780 (n1202, n229);
not  g781 (n1234, n265);
buf  g782 (n1066, n142);
not  g783 (n642, n190);
buf  g784 (n1582, n153);
not  g785 (n807, n183);
not  g786 (n823, n198);
buf  g787 (n960, n119);
not  g788 (n511, n183);
not  g789 (n726, n352);
not  g790 (n1602, n306);
not  g791 (n1503, n186);
buf  g792 (n690, n138);
not  g793 (n905, n162);
not  g794 (n1645, n393);
buf  g795 (n1206, n401);
not  g796 (n737, n274);
not  g797 (n1256, n180);
not  g798 (n446, n316);
not  g799 (n1108, n157);
buf  g800 (n1568, n205);
buf  g801 (n1199, n110);
buf  g802 (n503, n296);
not  g803 (n1227, n314);
not  g804 (n631, n344);
not  g805 (n1070, n219);
not  g806 (n868, n147);
not  g807 (n1622, n353);
buf  g808 (n748, n396);
not  g809 (n510, n324);
buf  g810 (n1412, n359);
not  g811 (n1305, n329);
buf  g812 (n429, n266);
buf  g813 (n887, n152);
buf  g814 (n1389, n234);
not  g815 (n1237, n203);
buf  g816 (n1519, n122);
not  g817 (n628, n223);
buf  g818 (n895, n160);
buf  g819 (n1142, n199);
not  g820 (n1022, n364);
not  g821 (n1145, n373);
buf  g822 (n1410, n390);
buf  g823 (n1260, n244);
not  g824 (n892, n418);
buf  g825 (n878, n229);
not  g826 (n1498, n183);
buf  g827 (n1669, n419);
not  g828 (n616, n391);
buf  g829 (n505, n308);
not  g830 (n1190, n313);
not  g831 (n1269, n369);
buf  g832 (n922, n150);
buf  g833 (n1047, n309);
buf  g834 (n1469, n119);
buf  g835 (n1405, n126);
not  g836 (n436, n185);
buf  g837 (n1524, n277);
buf  g838 (n652, n318);
not  g839 (n1643, n334);
not  g840 (n609, n243);
not  g841 (n1546, n188);
not  g842 (n728, n259);
buf  g843 (n556, n216);
not  g844 (n736, n318);
buf  g845 (n1654, n220);
not  g846 (n1658, n412);
not  g847 (n663, n363);
not  g848 (n1119, n188);
buf  g849 (n1344, n398);
buf  g850 (n717, n396);
buf  g851 (n693, n165);
buf  g852 (n1382, n190);
buf  g853 (n897, n339);
buf  g854 (n466, n172);
not  g855 (n486, n257);
not  g856 (n562, n389);
not  g857 (n945, n107);
not  g858 (n531, n135);
buf  g859 (n1671, n372);
buf  g860 (n937, n177);
not  g861 (n724, n329);
not  g862 (n608, n412);
buf  g863 (n1608, n421);
buf  g864 (n647, n253);
buf  g865 (n997, n238);
not  g866 (n962, n407);
buf  g867 (n1581, n255);
buf  g868 (n644, n139);
buf  g869 (n790, n194);
not  g870 (n1333, n286);
not  g871 (n1500, n147);
buf  g872 (n1557, n180);
buf  g873 (n1054, n291);
not  g874 (n1378, n343);
not  g875 (n571, n168);
not  g876 (n643, n243);
buf  g877 (n584, n345);
not  g878 (n983, n169);
buf  g879 (n455, n319);
not  g880 (n1587, n138);
not  g881 (n1200, n220);
not  g882 (n704, n340);
buf  g883 (n1248, n328);
buf  g884 (n667, n176);
not  g885 (n1501, n211);
not  g886 (n1173, n350);
not  g887 (n982, n151);
not  g888 (n1046, n149);
buf  g889 (n665, n302);
buf  g890 (n1154, n372);
not  g891 (n1107, n175);
not  g892 (n1452, n398);
buf  g893 (n561, n154);
not  g894 (n1082, n210);
not  g895 (n1506, n300);
buf  g896 (n611, n121);
buf  g897 (n874, n333);
buf  g898 (n1386, n315);
buf  g899 (n474, n164);
not  g900 (n1168, n324);
buf  g901 (n1286, n276);
not  g902 (n1605, n323);
buf  g903 (n735, n210);
buf  g904 (n1444, n219);
buf  g905 (n1084, n119);
buf  g906 (n1507, n332);
buf  g907 (n1069, n418);
buf  g908 (n1617, n119);
not  g909 (n540, n303);
not  g910 (n1613, n351);
not  g911 (n1460, n296);
not  g912 (n1564, n306);
not  g913 (n1267, n154);
buf  g914 (n1028, n218);
not  g915 (n658, n144);
not  g916 (n526, n283);
buf  g917 (n671, n260);
buf  g918 (n1018, n265);
buf  g919 (n1399, n346);
not  g920 (n599, n137);
buf  g921 (n917, n143);
buf  g922 (n1415, n337);
not  g923 (n1158, n356);
buf  g924 (n669, n141);
buf  g925 (n819, n198);
buf  g926 (n1001, n127);
not  g927 (n1488, n144);
not  g928 (n751, n138);
not  g929 (n1549, n248);
not  g930 (n1160, n289);
not  g931 (n1187, n174);
not  g932 (n1422, n354);
not  g933 (n995, n148);
not  g934 (n933, n135);
not  g935 (n1129, n254);
not  g936 (n1179, n183);
not  g937 (n1426, n133);
buf  g938 (n1105, n123);
not  g939 (n899, n332);
buf  g940 (n1236, n270);
not  g941 (n488, n379);
not  g942 (n793, n212);
not  g943 (n845, n375);
buf  g944 (n876, n158);
not  g945 (n820, n264);
not  g946 (n1420, n297);
not  g947 (n1435, n397);
buf  g948 (n990, n294);
not  g949 (n1577, n281);
not  g950 (n1192, n381);
not  g951 (n843, n213);
buf  g952 (n1651, n384);
not  g953 (n1112, n368);
not  g954 (n430, n318);
buf  g955 (n706, n288);
buf  g956 (n1320, n200);
not  g957 (n1655, n239);
buf  g958 (n1036, n360);
not  g959 (n799, n345);
buf  g960 (n1282, n297);
not  g961 (n858, n381);
not  g962 (n760, n208);
not  g963 (n1570, n287);
not  g964 (n1417, n362);
not  g965 (n763, n332);
not  g966 (n1049, n367);
not  g967 (n1159, n120);
buf  g968 (n437, n234);
buf  g969 (n1311, n331);
buf  g970 (n992, n230);
not  g971 (n925, n412);
not  g972 (n1484, n398);
buf  g973 (n1619, n392);
not  g974 (n1060, n310);
not  g975 (n1352, n369);
not  g976 (n1537, n331);
buf  g977 (n1584, n382);
not  g978 (n1328, n342);
buf  g979 (n1376, n388);
not  g980 (n504, n360);
not  g981 (n1310, n271);
buf  g982 (n1665, n408);
not  g983 (n479, n270);
buf  g984 (n808, n152);
buf  g985 (n750, n126);
buf  g986 (n475, n153);
not  g987 (n1057, n279);
buf  g988 (n1111, n137);
not  g989 (n635, n250);
not  g990 (n1331, n386);
buf  g991 (n1674, n170);
buf  g992 (n835, n402);
not  g993 (n1627, n411);
buf  g994 (n1330, n316);
buf  g995 (n1657, n182);
buf  g996 (n1148, n364);
not  g997 (n1370, n333);
buf  g998 (n1125, n294);
buf  g999 (n955, n320);
buf  g1000 (n1416, n342);
not  g1001 (n1515, n289);
not  g1002 (n1221, n260);
not  g1003 (n1659, n189);
not  g1004 (n1045, n201);
buf  g1005 (n770, n317);
not  g1006 (n492, n370);
buf  g1007 (n782, n175);
not  g1008 (n1670, n121);
buf  g1009 (n521, n242);
buf  g1010 (n931, n376);
not  g1011 (n848, n387);
not  g1012 (n918, n153);
not  g1013 (n773, n136);
not  g1014 (n547, n131);
buf  g1015 (n580, n336);
not  g1016 (n791, n336);
not  g1017 (n424, n107);
not  g1018 (n591, n304);
not  g1019 (n978, n146);
not  g1020 (n991, n379);
not  g1021 (n685, n136);
not  g1022 (n1122, n338);
not  g1023 (n1458, n141);
not  g1024 (n431, n129);
buf  g1025 (n1242, n228);
buf  g1026 (n1124, n281);
not  g1027 (n1315, n272);
buf  g1028 (n1403, n229);
buf  g1029 (n1401, n394);
buf  g1030 (n1274, n320);
not  g1031 (n1135, n400);
buf  g1032 (n441, n422);
buf  g1033 (n1341, n288);
buf  g1034 (n1323, n128);
not  g1035 (n1629, n422);
not  g1036 (n984, n278);
not  g1037 (n857, n289);
not  g1038 (n1411, n122);
buf  g1039 (n576, n285);
not  g1040 (n564, n149);
not  g1041 (n725, n408);
not  g1042 (n423, n359);
not  g1043 (n877, n251);
buf  g1044 (n537, n367);
not  g1045 (n602, n178);
not  g1046 (n946, n358);
buf  g1047 (n678, n420);
buf  g1048 (n1261, n362);
not  g1049 (n909, n196);
buf  g1050 (n947, n118);
not  g1051 (n478, n140);
buf  g1052 (n731, n365);
buf  g1053 (n1428, n235);
buf  g1054 (n1540, n373);
not  g1055 (n1573, n227);
buf  g1056 (n834, n393);
buf  g1057 (n572, n117);
buf  g1058 (n565, n215);
buf  g1059 (n715, n357);
not  g1060 (n588, n178);
buf  g1061 (n1486, n138);
not  g1062 (n1294, n159);
not  g1063 (n1075, n351);
not  g1064 (n1121, n194);
buf  g1065 (n965, n202);
not  g1066 (n1184, n296);
buf  g1067 (n512, n340);
buf  g1068 (n762, n272);
not  g1069 (n1365, n214);
buf  g1070 (n939, n328);
buf  g1071 (n1120, n386);
not  g1072 (n1118, n151);
not  g1073 (n523, n160);
not  g1074 (n1620, n297);
buf  g1075 (n1576, n130);
not  g1076 (n852, n256);
buf  g1077 (n449, n208);
not  g1078 (n593, n403);
not  g1079 (n502, n154);
buf  g1080 (n489, n238);
buf  g1081 (n575, n415);
buf  g1082 (n1554, n295);
not  g1083 (n653, n146);
buf  g1084 (n944, n170);
not  g1085 (n1361, n277);
buf  g1086 (n769, n405);
not  g1087 (n1116, n272);
not  g1088 (n1117, n167);
buf  g1089 (n1157, n249);
buf  g1090 (n1522, n154);
buf  g1091 (n932, n280);
buf  g1092 (n1137, n211);
buf  g1093 (n1203, n349);
buf  g1094 (n1076, n337);
buf  g1095 (n1343, n253);
not  g1096 (n796, n327);
not  g1097 (n1141, n127);
not  g1098 (n988, n231);
buf  g1099 (n681, n230);
not  g1100 (n626, n305);
buf  g1101 (n1255, n231);
not  g1102 (n716, n191);
buf  g1103 (n1201, n373);
buf  g1104 (n454, n377);
not  g1105 (n968, n330);
not  g1106 (n1037, n123);
buf  g1107 (n920, n143);
buf  g1108 (n1134, n363);
not  g1109 (n1136, n244);
buf  g1110 (n1388, n151);
buf  g1111 (n660, n132);
buf  g1112 (n1209, n218);
buf  g1113 (n673, n262);
buf  g1114 (n1115, n196);
buf  g1115 (n814, n226);
not  g1116 (n598, n296);
buf  g1117 (n1383, n231);
buf  g1118 (n840, n402);
buf  g1119 (n1326, n161);
buf  g1120 (n587, n247);
buf  g1121 (n1374, n406);
not  g1122 (n1213, n394);
not  g1123 (n1680, n260);
buf  g1124 (n1181, n391);
not  g1125 (n1093, n135);
buf  g1126 (n1099, n109);
not  g1127 (n867, n417);
buf  g1128 (n1650, n184);
not  g1129 (n921, n371);
buf  g1130 (n1625, n241);
buf  g1131 (n1663, n245);
buf  g1132 (n615, n326);
buf  g1133 (n1423, n283);
not  g1134 (n994, n341);
buf  g1135 (n1565, n302);
not  g1136 (n996, n279);
buf  g1137 (n821, n216);
not  g1138 (n1316, n305);
buf  g1139 (n1147, n269);
buf  g1140 (n710, n356);
not  g1141 (n1170, n370);
buf  g1142 (n1649, n380);
not  g1143 (n1089, n202);
buf  g1144 (n1110, n290);
not  g1145 (n828, n148);
not  g1146 (n794, n117);
buf  g1147 (n815, n287);
not  g1148 (n594, n197);
not  g1149 (n680, n383);
not  g1150 (n755, n221);
not  g1151 (n847, n167);
buf  g1152 (n1586, n345);
not  g1153 (n1155, n157);
not  g1154 (n559, n315);
buf  g1155 (n574, n328);
not  g1156 (n1302, n358);
not  g1157 (n1063, n187);
not  g1158 (n1555, n148);
not  g1159 (n636, n116);
not  g1160 (n1011, n193);
buf  g1161 (n568, n181);
buf  g1162 (n1510, n133);
buf  g1163 (n1594, n364);
buf  g1164 (n1578, n292);
not  g1165 (n558, n121);
buf  g1166 (n1456, n261);
not  g1167 (n1020, n255);
not  g1168 (n456, n238);
buf  g1169 (n875, n372);
buf  g1170 (n830, n221);
buf  g1171 (n1478, n187);
buf  g1172 (n1074, n268);
not  g1173 (n1471, n340);
not  g1174 (n1591, n268);
not  g1175 (n1580, n182);
buf  g1176 (n1349, n278);
not  g1177 (n1485, n112);
not  g1178 (n1667, n123);
not  g1179 (n1676, n322);
buf  g1180 (n637, n230);
buf  g1181 (n1357, n118);
not  g1182 (n1585, n386);
not  g1183 (n902, n287);
not  g1184 (n971, n226);
not  g1185 (n811, n267);
not  g1186 (n1453, n169);
not  g1187 (n1483, n210);
buf  g1188 (n766, n285);
buf  g1189 (n472, n136);
buf  g1190 (n1475, n203);
buf  g1191 (n911, n168);
buf  g1192 (n445, n228);
not  g1193 (n924, n181);
buf  g1194 (n711, n338);
buf  g1195 (n1166, n334);
buf  g1196 (n1472, n356);
buf  g1197 (n809, n182);
not  g1198 (n707, n113);
not  g1199 (n646, n212);
buf  g1200 (n718, n252);
buf  g1201 (n1424, n114);
not  g1202 (n1288, n420);
buf  g1203 (n500, n233);
buf  g1204 (n1291, n262);
buf  g1205 (n1188, n274);
buf  g1206 (n595, n113);
buf  g1207 (n817, n313);
buf  g1208 (n1290, n311);
buf  g1209 (n1362, n382);
buf  g1210 (n684, n341);
buf  g1211 (n986, n299);
not  g1212 (n1441, n298);
buf  g1213 (n554, n118);
buf  g1214 (n589, n388);
buf  g1215 (n541, n312);
buf  g1216 (n1152, n121);
not  g1217 (n1032, n176);
buf  g1218 (n1238, n306);
not  g1219 (n1220, n207);
buf  g1220 (n1140, n127);
not  g1221 (n535, n391);
not  g1222 (n453, n222);
buf  g1223 (n1132, n239);
not  g1224 (n515, n327);
buf  g1225 (n778, n358);
not  g1226 (n1502, n323);
buf  g1227 (n1520, n287);
buf  g1228 (n703, n273);
not  g1229 (n806, n302);
buf  g1230 (n1660, n142);
buf  g1231 (n846, n181);
not  g1232 (n1631, n115);
buf  g1233 (n686, n350);
buf  g1234 (n539, n311);
buf  g1235 (n607, n367);
buf  g1236 (n1253, n127);
buf  g1237 (n513, n321);
buf  g1238 (n1041, n352);
buf  g1239 (n473, n195);
not  g1240 (n930, n376);
buf  g1241 (n1462, n400);
not  g1242 (n787, n284);
buf  g1243 (n1364, n162);
not  g1244 (n839, n266);
not  g1245 (n1638, n217);
not  g1246 (n816, n357);
not  g1247 (n1257, n344);
not  g1248 (n1308, n352);
buf  g1249 (n1637, n223);
buf  g1250 (n1167, n111);
not  g1251 (n1275, n295);
buf  g1252 (n1262, n275);
buf  g1253 (n1635, n187);
not  g1254 (n481, n403);
not  g1255 (n1218, n307);
not  g1256 (n1247, n124);
buf  g1257 (n563, n324);
not  g1258 (n950, n111);
buf  g1259 (n476, n189);
buf  g1260 (n1525, n159);
buf  g1261 (n1151, n149);
not  g1262 (n527, n328);
not  g1263 (n550, n305);
buf  g1264 (n854, n147);
buf  g1265 (n1492, n285);
not  g1266 (n783, n214);
not  g1267 (n1050, n186);
buf  g1268 (n1626, n360);
not  g1269 (n461, n235);
not  g1270 (n805, n155);
not  g1271 (n1174, n342);
buf  g1272 (n883, n414);
not  g1273 (n1149, n267);
not  g1274 (n777, n421);
buf  g1275 (n493, n137);
not  g1276 (n1055, n320);
not  g1277 (n1487, n184);
not  g1278 (n1392, n341);
buf  g1279 (n1029, n249);
buf  g1280 (n1068, n361);
buf  g1281 (n1385, n335);
not  g1282 (n1180, n186);
not  g1283 (n1544, n155);
not  g1284 (n872, n227);
buf  g1285 (n543, n300);
buf  g1286 (n792, n225);
buf  g1287 (n934, n402);
buf  g1288 (n1015, n401);
not  g1289 (n687, n179);
not  g1290 (n529, n172);
not  g1291 (n1225, n190);
buf  g1292 (n597, n153);
not  g1293 (n634, n146);
not  g1294 (n604, n311);
buf  g1295 (n1301, n366);
buf  g1296 (n1342, n390);
not  g1297 (n1489, n318);
not  g1298 (n1634, n322);
not  g1299 (n566, n248);
buf  g1300 (n941, n263);
not  g1301 (n1346, n245);
not  g1302 (n640, n332);
not  g1303 (n708, n398);
buf  g1304 (n1407, n212);
not  g1305 (n662, n412);
not  g1306 (n689, n256);
not  g1307 (n1406, n116);
not  g1308 (n683, n338);
not  g1309 (n699, n411);
not  g1310 (n1642, n302);
not  g1311 (n1442, n387);
not  g1312 (n1246, n411);
buf  g1313 (n596, n301);
buf  g1314 (n1672, n275);
not  g1315 (n1508, n273);
buf  g1316 (n603, n343);
buf  g1317 (n1516, n390);
buf  g1318 (n862, n219);
buf  g1319 (n1087, n173);
not  g1320 (n1285, n246);
not  g1321 (n914, n115);
not  g1322 (n1434, n354);
buf  g1323 (n818, n244);
not  g1324 (n1596, n204);
buf  g1325 (n1482, n267);
not  g1326 (n1497, n368);
buf  g1327 (n427, n301);
not  g1328 (n825, n278);
not  g1329 (n1012, n168);
buf  g1330 (n1284, n132);
buf  g1331 (n1427, n396);
buf  g1332 (n659, n289);
buf  g1333 (n752, n336);
not  g1334 (n1321, n165);
buf  g1335 (n1224, n193);
not  g1336 (n1080, n159);
not  g1337 (n1447, n420);
buf  g1338 (n448, n218);
buf  g1339 (n928, n266);
not  g1340 (n1526, n338);
buf  g1341 (n509, n281);
not  g1342 (n1465, n176);
buf  g1343 (n583, n185);
not  g1344 (n1567, n207);
not  g1345 (n1641, n334);
buf  g1346 (n1628, n190);
buf  g1347 (n1381, n124);
not  g1348 (n732, n254);
buf  g1349 (n1165, n303);
buf  g1350 (n1681, n175);
not  g1351 (n754, n375);
buf  g1352 (n721, n254);
not  g1353 (n802, n361);
buf  g1354 (n1235, n389);
buf  g1355 (n638, n397);
buf  g1356 (n470, n231);
buf  g1357 (n1325, n215);
not  g1358 (n844, n329);
buf  g1359 (n487, n132);
not  g1360 (n1446, n250);
not  g1361 (n1171, n262);
buf  g1362 (n954, n215);
buf  g1363 (n497, n315);
not  g1364 (n702, n208);
not  g1365 (n1026, n330);
buf  g1366 (n893, n221);
buf  g1367 (n1139, n339);
not  g1368 (n1138, n321);
buf  g1369 (n841, n326);
buf  g1370 (n1336, n179);
buf  g1371 (n1481, n293);
not  g1372 (n629, n383);
buf  g1373 (n891, n135);
not  g1374 (n499, n257);
buf  g1375 (n853, n130);
not  g1376 (n1019, n319);
not  g1377 (n1296, n309);
buf  g1378 (n795, n109);
not  g1379 (n1006, n194);
not  g1380 (n498, n420);
buf  g1381 (n1266, n243);
not  g1382 (n879, n249);
not  g1383 (n1205, n130);
buf  g1384 (n501, n155);
buf  g1385 (n1398, n266);
buf  g1386 (n1010, n149);
not  g1387 (n1400, n137);
buf  g1388 (n1566, n355);
not  g1389 (n1182, n246);
not  g1390 (n1332, n330);
not  g1391 (n1551, n258);
buf  g1392 (n432, n173);
buf  g1393 (n483, n383);
not  g1394 (n980, n226);
buf  g1395 (n1394, n271);
not  g1396 (n1086, n240);
buf  g1397 (n705, n352);
buf  g1398 (n1230, n327);
not  g1399 (n987, n199);
buf  g1400 (n1085, n376);
not  g1401 (n1521, n142);
buf  g1402 (n1590, n309);
buf  g1403 (n1380, n369);
buf  g1404 (n1081, n399);
buf  g1405 (n548, n331);
not  g1406 (n1340, n196);
not  g1407 (n477, n311);
buf  g1408 (n442, n148);
buf  g1409 (n1161, n164);
not  g1410 (n452, n263);
not  g1411 (n1219, n241);
not  g1412 (n861, n213);
not  g1413 (n800, n225);
buf  g1414 (n460, n354);
buf  g1415 (n959, n159);
not  g1416 (n1530, n348);
not  g1417 (n727, n371);
not  g1418 (n864, n325);
buf  g1419 (n742, n278);
not  g1420 (n1303, n286);
buf  g1421 (n1096, n323);
not  g1422 (n688, n242);
buf  g1423 (n967, n171);
not  g1424 (n426, n113);
not  g1425 (n1588, n128);
buf  g1426 (n1277, n280);
buf  g1427 (n1396, n179);
buf  g1428 (n940, n381);
not  g1429 (n894, n156);
not  g1430 (n1189, n339);
not  g1431 (n1259, n375);
not  g1432 (n1592, n224);
buf  g1433 (n1222, n113);
not  g1434 (n813, n409);
buf  g1435 (n1329, n416);
buf  g1436 (n1644, n195);
buf  g1437 (n963, n409);
not  g1438 (n434, n281);
buf  g1439 (n1556, n344);
buf  g1440 (n679, n271);
buf  g1441 (n1250, n122);
not  g1442 (n838, n345);
not  g1443 (n1327, n385);
buf  g1444 (n1639, n399);
not  g1445 (n1251, n273);
buf  g1446 (n1100, n397);
buf  g1447 (n528, n222);
buf  g1448 (n675, n388);
buf  g1449 (n849, n416);
not  g1450 (n1033, n384);
buf  g1451 (n444, n385);
not  g1452 (n972, n355);
buf  g1453 (n1375, n304);
buf  g1454 (n630, n304);
not  g1455 (n677, n392);
not  g1456 (n1195, n402);
not  g1457 (n606, n260);
not  g1458 (n713, n327);
not  g1459 (n985, n223);
not  g1460 (n1039, n115);
buf  g1461 (n1368, n226);
buf  g1462 (n723, n347);
not  g1463 (n530, n117);
buf  g1464 (n1059, n120);
buf  g1465 (n871, n184);
not  g1466 (n1589, n290);
buf  g1467 (n1348, n350);
buf  g1468 (n1065, n298);
not  g1469 (n534, n319);
not  g1470 (n958, n348);
not  g1471 (n1439, n111);
not  g1472 (n1004, n312);
buf  g1473 (n1527, n369);
buf  g1474 (n1324, n214);
buf  g1475 (n1009, n244);
buf  g1476 (n979, n382);
buf  g1477 (n648, n174);
not  g1478 (n546, n220);
buf  g1479 (n1169, n155);
not  g1480 (n1437, n182);
buf  g1481 (n1464, n413);
buf  g1482 (n1005, n163);
buf  g1483 (n1335, n237);
buf  g1484 (n1661, n251);
not  g1485 (n1528, n370);
buf  g1486 (n1476, n271);
not  g1487 (n1228, n264);
not  g1488 (n860, n384);
buf  g1489 (n1603, n139);
buf  g1490 (n1574, n216);
not  g1491 (n881, n141);
buf  g1492 (n622, n192);
not  g1493 (n1583, n191);
buf  g1494 (n600, n150);
not  g1495 (n1466, n306);
not  g1496 (n906, n139);
not  g1497 (n661, n316);
buf  g1498 (n1146, n234);
not  g1499 (n508, n309);
not  g1500 (n904, n144);
buf  g1501 (n1123, n166);
not  g1502 (n1172, n250);
not  g1503 (n1289, n217);
buf  g1504 (n1393, n162);
buf  g1505 (n964, n228);
buf  g1506 (n1094, n204);
not  g1507 (n786, n356);
not  g1508 (n824, n292);
not  g1509 (n1258, n189);
not  g1510 (n1366, n347);
buf  g1511 (n465, n203);
buf  g1512 (n1071, n174);
not  g1513 (n469, n407);
buf  g1514 (n900, n391);
buf  g1515 (n682, n347);
buf  g1516 (n1106, n165);
buf  g1517 (n837, n193);
buf  g1518 (n1113, n126);
buf  g1519 (n1270, n235);
not  g1520 (n625, n129);
not  g1521 (n552, n205);
buf  g1522 (n577, n150);
not  g1523 (n863, n232);
not  g1524 (n829, n349);
buf  g1525 (n1675, n254);
buf  g1526 (n1552, n368);
not  g1527 (n1101, n240);
not  g1528 (n1445, n310);
buf  g1529 (n804, n116);
buf  g1530 (n1276, n343);
buf  g1531 (n1683, n178);
buf  g1532 (n1384, n166);
buf  g1533 (n1413, n233);
buf  g1534 (n803, n178);
buf  g1535 (n1436, n274);
buf  g1536 (n1632, n192);
buf  g1537 (n519, n232);
not  g1538 (n1061, n357);
buf  g1539 (n696, n346);
buf  g1540 (n1490, n404);
not  g1541 (n612, n377);
buf  g1542 (n645, n125);
buf  g1543 (n1538, n225);
not  g1544 (n1607, n399);
not  g1545 (n1216, n334);
not  g1546 (n1468, n381);
buf  g1547 (n1429, n396);
buf  g1548 (n1679, n180);
not  g1549 (n1599, n329);
buf  g1550 (n451, n156);
not  g1551 (n1212, n290);
buf  g1552 (n506, n108);
buf  g1553 (n1048, n112);
buf  g1554 (n1318, n246);
buf  g1555 (n1505, n273);
buf  g1556 (n974, n215);
not  g1557 (n490, n245);
buf  g1558 (n517, n156);
buf  g1559 (n1395, n291);
buf  g1560 (n697, n409);
buf  g1561 (n961, n408);
buf  g1562 (n1363, n312);
buf  g1563 (n1304, n209);
buf  g1564 (n698, n291);
not  g1565 (n745, n276);
not  g1566 (n765, n282);
buf  g1567 (n1397, n199);
not  g1568 (n1072, n417);
buf  g1569 (n1536, n169);
not  g1570 (n781, n251);
buf  g1571 (n555, n349);
not  g1572 (n1183, n419);
buf  g1573 (n913, n291);
buf  g1574 (n1338, n237);
buf  g1575 (n633, n400);
not  g1576 (n758, n141);
not  g1577 (n969, n299);
not  g1578 (n889, n171);
not  g1579 (n1513, n394);
not  g1580 (n1103, n322);
not  g1581 (n1542, n401);
not  g1582 (n1541, n140);
not  g1583 (n1504, n349);
not  g1584 (n759, n354);
buf  g1585 (n536, n134);
buf  g1586 (n1470, n292);
not  g1587 (n1621, n315);
not  g1588 (n463, n219);
not  g1589 (n1668, n410);
buf  g1590 (n1595, n188);
buf  g1591 (n789, n145);
buf  g1592 (n1319, n144);
buf  g1593 (n927, n325);
buf  g1594 (n740, n325);
not  g1595 (n650, n280);
buf  g1596 (n1090, n122);
buf  g1597 (n774, n405);
buf  g1598 (n1035, n147);
buf  g1599 (n1572, n234);
buf  g1600 (n1127, n263);
buf  g1601 (n1104, n172);
not  g1602 (n1678, n191);
buf  g1603 (n966, n393);
not  g1604 (n1451, n124);
buf  g1605 (n1390, n161);
not  g1606 (n1042, n145);
buf  g1607 (n1459, n201);
not  g1608 (n1322, n166);
buf  g1609 (n1373, n129);
buf  g1610 (n1194, n341);
not  g1611 (n480, n177);
not  g1612 (n1239, n200);
buf  g1613 (n1178, n211);
buf  g1614 (n1007, n414);
buf  g1615 (n1252, n374);
buf  g1616 (n1264, n387);
not  g1617 (n560, n257);
not  g1618 (n613, n264);
not  g1619 (n1043, n131);
not  g1620 (n1509, n361);
not  g1621 (n533, n130);
buf  g1622 (n1495, n158);
buf  g1623 (n1562, n418);
buf  g1624 (n1474, n409);
buf  g1625 (n1611, n199);
not  g1626 (n514, n242);
not  g1627 (n557, n197);
not  g1628 (n1243, n263);
buf  g1629 (n912, n404);
not  g1630 (n468, n217);
not  g1631 (n695, n257);
not  g1632 (n1677, n298);
not  g1633 (n1379, n415);
buf  g1634 (n1499, n368);
buf  g1635 (n1314, n275);
buf  g1636 (n908, n282);
not  g1637 (n507, n410);
not  g1638 (n957, n406);
not  g1639 (n1095, n314);
not  g1640 (n1418, n304);
not  g1641 (n1233, n224);
not  g1642 (n1164, n160);
not  g1643 (n1245, n305);
buf  g1644 (n923, n129);
buf  g1645 (n749, n186);
not  g1646 (n433, n206);
buf  g1647 (n1647, n125);
buf  g1648 (n601, n293);
not  g1649 (n1016, n232);
not  g1650 (n1083, n126);
not  g1651 (n484, n343);
buf  g1652 (n989, n188);
buf  g1653 (n1013, n298);
buf  g1654 (n1317, n212);
not  g1655 (n869, n132);
not  g1656 (n641, n283);
not  g1657 (n1432, n230);
buf  g1658 (n551, n403);
nand g1659 (n2067, n1513, n1101, n1555, n1449);
nor  g1660 (n1763, n1336, n1481, n1395, n465);
or   g1661 (n1957, n1551, n1597, n1331, n1093);
or   g1662 (n2052, n633, n1506, n1317, n1478);
xor  g1663 (n1887, n1167, n1548, n1504, n1480);
and  g1664 (n1971, n1065, n1551, n1516, n651);
and  g1665 (n1848, n1457, n1261, n1371, n1495);
or   g1666 (n1973, n1404, n1333, n1601, n457);
xnor g1667 (n1907, n935, n1554, n1530, n1348);
xnor g1668 (n2054, n1016, n1351, n1339, n894);
xnor g1669 (n1923, n1631, n1301, n618, n479);
nand g1670 (n1731, n1284, n1466, n1282, n1294);
xor  g1671 (n1772, n1435, n1352, n1155, n1362);
and  g1672 (n1691, n1438, n1424, n503, n1453);
xor  g1673 (n1719, n1073, n620, n1109, n734);
xnor g1674 (n1819, n1171, n1622, n1491, n1627);
nor  g1675 (n2198, n1268, n1546, n1088, n1349);
nand g1676 (n2011, n667, n548, n1587, n927);
and  g1677 (n1916, n1531, n594, n1020, n792);
nand g1678 (n1889, n1486, n743, n945, n1582);
xnor g1679 (n1783, n552, n1454, n1527, n1453);
nand g1680 (n1687, n433, n1308, n1372, n1574);
or   g1681 (n1744, n839, n900, n431, n622);
xor  g1682 (n1801, n1503, n841, n1176, n1524);
xor  g1683 (n2091, n1389, n1631, n933, n1406);
or   g1684 (n1754, n1576, n1493, n753, n1314);
and  g1685 (n2004, n1542, n1592, n1490, n1163);
and  g1686 (n1846, n721, n1459, n1402, n1017);
xnor g1687 (n2169, n492, n1427, n1080, n1495);
nand g1688 (n2134, n1258, n1351, n1297, n673);
nand g1689 (n1758, n1518, n1461, n899, n1594);
xnor g1690 (n2143, n1346, n1442, n652, n1437);
or   g1691 (n1770, n1005, n1374, n1463, n1056);
or   g1692 (n2020, n1226, n1476, n1002, n1429);
nand g1693 (n2016, n1501, n1014, n1074, n1190);
and  g1694 (n1990, n1561, n1558, n1424, n1347);
xor  g1695 (n2101, n575, n1316, n807, n1436);
nand g1696 (n1905, n1379, n1402, n1623, n1598);
xor  g1697 (n1958, n1477, n504, n1616, n1330);
xnor g1698 (n1824, n901, n1578, n1280, n1177);
nand g1699 (n1688, n1045, n1631, n1515, n885);
nor  g1700 (n1982, n832, n1575, n1572, n1483);
nand g1701 (n1978, n1090, n1390, n1417, n664);
nor  g1702 (n2234, n775, n543, n691, n1453);
and  g1703 (n2042, n719, n1568, n876, n1299);
nor  g1704 (n1767, n1291, n941, n1572, n1289);
and  g1705 (n1829, n970, n1536, n1108, n973);
or   g1706 (n2074, n1293, n1500, n1419, n1591);
or   g1707 (n2235, n610, n1431, n1625, n1352);
or   g1708 (n1720, n1576, n956, n1443, n1084);
nand g1709 (n1791, n992, n1548, n685, n1114);
or   g1710 (n2160, n1315, n1538, n1519, n1464);
nand g1711 (n1712, n1546, n1260, n924, n1218);
nor  g1712 (n2099, n1335, n511, n451, n1486);
or   g1713 (n2034, n1285, n1308, n704, n1530);
nand g1714 (n1797, n506, n1414, n1460, n1173);
xnor g1715 (n2253, n1309, n650, n905, n1574);
and  g1716 (n2210, n1158, n1488, n1192, n1474);
nand g1717 (n1868, n1142, n1449, n1465, n1105);
and  g1718 (n2216, n982, n1341, n1319, n637);
xnor g1719 (n2230, n1611, n1441, n442, n1492);
or   g1720 (n1816, n1361, n1013, n1015, n1029);
nor  g1721 (n2113, n1363, n1254, n1450, n1301);
and  g1722 (n1793, n1343, n1350, n1356, n874);
or   g1723 (n2015, n1426, n1311, n484, n623);
nand g1724 (n2121, n1577, n1552, n1299, n1432);
xnor g1725 (n2238, n564, n1011, n1312, n1574);
or   g1726 (n2153, n1345, n1535, n1369, n1289);
or   g1727 (n1997, n831, n1609, n1237, n801);
nand g1728 (n2199, n1083, n1630, n1277, n1505);
nand g1729 (n1778, n1310, n436, n1387, n1570);
nor  g1730 (n2060, n508, n1403, n1428, n1325);
and  g1731 (n1896, n742, n953, n1514, n1304);
or   g1732 (n1689, n425, n1554, n1532, n1327);
nor  g1733 (n1937, n1587, n1235, n1605, n1371);
or   g1734 (n1922, n1308, n1354, n1434, n1496);
or   g1735 (n2162, n1394, n1420, n1324, n1374);
xnor g1736 (n2186, n1416, n556, n1531, n811);
and  g1737 (n2028, n1502, n1041, n1606, n1497);
xor  g1738 (n1821, n1157, n1449, n489, n1577);
nand g1739 (n1912, n606, n1077, n1436, n1485);
xnor g1740 (n1796, n1357, n1411, n805, n1630);
nor  g1741 (n1962, n1225, n1297, n538, n1612);
xnor g1742 (n2254, n1613, n706, n1197, n1358);
nor  g1743 (n2148, n1599, n1344, n1170, n1443);
nor  g1744 (n1949, n1617, n1547, n1602, n1341);
xor  g1745 (n2263, n1269, n1505, n454, n1509);
nor  g1746 (n2239, n1427, n1260, n1411, n1563);
nor  g1747 (n1950, n1353, n1319, n1075, n946);
nor  g1748 (n1710, n1378, n1597, n870, n1344);
or   g1749 (n2041, n939, n1413, n1442, n1382);
xnor g1750 (n2055, n1266, n1256, n452, n1447);
xor  g1751 (n2040, n1637, n1315, n1607, n605);
nor  g1752 (n1959, n1407, n861, n1322, n755);
nand g1753 (n1968, n473, n1383, n851, n1463);
nand g1754 (n1795, n1595, n940, n824, n1317);
nor  g1755 (n2140, n1524, n1184, n770, n1304);
xor  g1756 (n2025, n1445, n1287, n1295, n1332);
xor  g1757 (n1882, n1541, n979, n1111, n1585);
xnor g1758 (n1749, n642, n972, n786, n1498);
and  g1759 (n2069, n1568, n1362, n1551, n678);
and  g1760 (n2137, n1421, n1470, n1624, n1346);
xor  g1761 (n2217, n1186, n607, n1201, n1362);
nand g1762 (n1727, n1276, n1286, n1498, n1486);
nand g1763 (n1946, n590, n1320, n1460, n1570);
xor  g1764 (n2264, n1459, n1321, n576, n1636);
or   g1765 (n1713, n1472, n1396, n1366, n544);
nand g1766 (n1789, n1543, n1370, n1462, n1456);
xnor g1767 (n1881, n1430, n1433, n1605, n891);
and  g1768 (n2076, n539, n1343, n1553, n806);
xnor g1769 (n1951, n1409, n916, n1168, n1467);
xor  g1770 (n2065, n1281, n788, n1387, n875);
xor  g1771 (n2211, n1004, n1602, n1421, n580);
xor  g1772 (n2100, n1405, n1622, n1507, n1361);
nor  g1773 (n1876, n1489, n1347, n698, n1484);
nand g1774 (n2071, n493, n1390, n681, n1099);
or   g1775 (n2173, n1538, n1307, n1613, n1559);
nand g1776 (n2251, n1141, n1106, n1386, n1283);
xnor g1777 (n1790, n1265, n1569, n1373, n1290);
nor  g1778 (n2119, n553, n1546, n1418, n1007);
nand g1779 (n2127, n1516, n1633, n1266, n1430);
nand g1780 (n1947, n1472, n1275, n991, n925);
or   g1781 (n2064, n684, n1130, n888, n1331);
and  g1782 (n2267, n1292, n1317, n1438, n1406);
nor  g1783 (n2261, n1599, n1332, n1365, n817);
and  g1784 (n2195, n1620, n1350, n877, n596);
xnor g1785 (n2102, n513, n1556, n1282, n1441);
nor  g1786 (n1836, n1326, n777, n581, n579);
xnor g1787 (n1804, n782, n1087, n1537, n1530);
or   g1788 (n1705, n1471, n1224, n1351, n1464);
nor  g1789 (n2247, n1521, n577, n1280, n993);
xor  g1790 (n2266, n957, n1427, n774, n822);
nor  g1791 (n2168, n1081, n1250, n1293, n922);
nand g1792 (n1847, n1040, n1428, n1249, n613);
xnor g1793 (n2026, n522, n1439, n646, n1564);
nand g1794 (n2213, n920, n1274, n1466, n1603);
xor  g1795 (n2024, n1381, n1304, n938, n1571);
xor  g1796 (n1835, n597, n879, n441, n1323);
nor  g1797 (n1747, n1328, n1446, n1600, n1291);
or   g1798 (n1808, n1259, n1589, n733, n1301);
xor  g1799 (n2039, n1464, n1179, n1381, n591);
and  g1800 (n1779, n1501, n668, n1631, n1588);
and  g1801 (n1964, n1232, n448, n981, n1591);
xnor g1802 (n2125, n1372, n1581, n833, n1263);
and  g1803 (n1942, n1627, n1508, n1321, n450);
or   g1804 (n1776, n1612, n1296, n1213, n1270);
and  g1805 (n1817, n1510, n1431, n1586, n679);
or   g1806 (n1883, n1009, n1583, n1104, n1220);
nand g1807 (n2132, n1518, n1419, n1262, n727);
or   g1808 (n1732, n1251, n948, n1506, n1468);
nand g1809 (n2077, n1455, n750, n1162, n1512);
xor  g1810 (n1904, n1563, n1560, n752, n1608);
or   g1811 (n1910, n1590, n793, n532, n1440);
nor  g1812 (n2124, n1398, n1618, n796, n1502);
or   g1813 (n2030, n1520, n1368, n1433, n1635);
nand g1814 (n2059, n1128, n531, n1405, n1608);
and  g1815 (n2237, n1469, n1615, n424, n826);
or   g1816 (n1865, n1629, n1553, n1601, n1443);
and  g1817 (n2104, n1551, n1324, n1449, n896);
xnor g1818 (n1833, n1096, n1154, n1385, n1276);
xor  g1819 (n1726, n558, n1578, n1288, n1301);
nor  g1820 (n1786, n1366, n759, n1513, n440);
xor  g1821 (n2171, n1425, n736, n1438, n1384);
nand g1822 (n1806, n1542, n1422, n803, n1524);
and  g1823 (n2110, n1493, n804, n1337, n621);
or   g1824 (n1760, n675, n1429, n1627, n1576);
nor  g1825 (n1730, n745, n632, n760, n1606);
xnor g1826 (n2009, n1501, n1438, n707, n1475);
xor  g1827 (n1834, n1425, n789, n802, n1305);
xor  g1828 (n1998, n1359, n855, n871, n857);
or   g1829 (n1755, n978, n820, n829, n1418);
nor  g1830 (n2215, n1457, n1169, n1064, n1477);
xnor g1831 (n1828, n1612, n819, n1461, n456);
nand g1832 (n1897, n1510, n1102, n1479, n1351);
xnor g1833 (n1826, n971, n1352, n491, n1329);
xnor g1834 (n2079, n1513, n1148, n1265, n1512);
and  g1835 (n2192, n1478, n1472, n1454, n1327);
nand g1836 (n2201, n1441, n1430, n1119, n1479);
and  g1837 (n1850, n889, n1637, n533, n1496);
or   g1838 (n2120, n1360, n602, n914, n1620);
and  g1839 (n1980, n1203, n1525, n1440, n986);
xnor g1840 (n1707, n1318, n1429, n1393, n1604);
nor  g1841 (n2133, n630, n604, n1537, n1223);
xnor g1842 (n2174, n701, n1611, n1434, n1079);
xor  g1843 (n1831, n917, n475, n911, n969);
or   g1844 (n2207, n1582, n1284, n1406, n497);
or   g1845 (n1722, n1591, n1571, n1446, n1614);
or   g1846 (n1872, n1617, n1603, n955, n1306);
nand g1847 (n1827, n1393, n1413, n1404, n1422);
xor  g1848 (n1753, n1517, n1282, n1637, n1621);
nand g1849 (n1921, n1483, n868, n1069, n1497);
or   g1850 (n1878, n1536, n1399, n1116, n1144);
nand g1851 (n1953, n1423, n1019, n732, n1529);
nor  g1852 (n1736, n674, n1435, n989, n1346);
or   g1853 (n2172, n848, n1255, n1302, n988);
xnor g1854 (n2088, n1509, n1616, n1370, n1279);
and  g1855 (n1724, n1322, n1120, n1450, n1408);
xnor g1856 (n2194, n1535, n1440, n1487, n1341);
and  g1857 (n2033, n1473, n1389, n963, n1299);
xor  g1858 (n2008, n740, n1420, n1295, n444);
or   g1859 (n2051, n1630, n616, n1137, n1523);
xnor g1860 (n2191, n1334, n530, n514, n1611);
nand g1861 (n1810, n1567, n1188, n1342, n1370);
nand g1862 (n1952, n731, n476, n1337, n1262);
xor  g1863 (n1867, n747, n1284, n960, n1208);
and  g1864 (n1870, n1609, n1624, n1596, n1474);
xnor g1865 (n1812, n1364, n852, n483, n1458);
or   g1866 (n1874, n722, n542, n735, n1565);
and  g1867 (n2188, n1348, n937, n1586, n1523);
or   g1868 (n2094, n1594, n1476, n1550, n1303);
or   g1869 (n1841, n561, n1433, n1451, n1487);
nand g1870 (n2184, n1558, n1467, n1380, n1343);
nand g1871 (n2243, n1558, n1270, n1006, n611);
nand g1872 (n2061, n1287, n560, n994, n999);
nand g1873 (n2145, n1042, n1533, n1626, n429);
nor  g1874 (n1869, n1356, n1604, n1412);
and  g1875 (n1879, n959, n509, n1288, n1471);
xor  g1876 (n2129, n641, n1359, n962, n1354);
nor  g1877 (n2111, n723, n1413, n1469, n566);
nor  g1878 (n2106, n1561, n1423, n1509, n821);
xnor g1879 (n1734, n729, n1319, n1180, n1475);
nor  g1880 (n1764, n1396, n1480, n1085, n1635);
nor  g1881 (n1769, n1637, n1357, n1124, n1214);
nor  g1882 (n1794, n1450, n1340, n884, n791);
xor  g1883 (n2157, n1417, n1037, n694, n1428);
and  g1884 (n2103, n1526, n485, n1602, n1187);
nor  g1885 (n2190, n1451, n1018, n1446, n1476);
nor  g1886 (n2013, n1121, n463, n1579, n928);
or   g1887 (n1774, n563, n499, n1492, n699);
and  g1888 (n1773, n1127, n1332, n1291, n1381);
nor  g1889 (n1860, n1543, n1508, n1557, n1525);
nor  g1890 (n1935, n1092, n1385, n1563, n1401);
nor  g1891 (n1920, n1369, n1589, n1067, n1437);
xor  g1892 (n1977, n1425, n520, n1580, n1532);
nor  g1893 (n2175, n682, n764, n1397, n748);
nand g1894 (n1924, n1262, n1526, n1385, n1593);
xnor g1895 (n1994, n1397, n1269, n647, n1634);
and  g1896 (n2115, n1624, n426, n1467, n1437);
or   g1897 (n2268, n1598, n1529, n1383, n1518);
nor  g1898 (n2223, n1276, n464, n1216, n1022);
xnor g1899 (n1766, n1330, n1378, n1635, n1552);
and  g1900 (n2043, n1393, n1497, n779, n1456);
and  g1901 (n2189, n1434, n1517, n1465, n1115);
nand g1902 (n1886, n1509, n1123, n1600, n1134);
nand g1903 (n2149, n1375, n1089, n769, n626);
nand g1904 (n2056, n809, n523, n1181, n1452);
nor  g1905 (n2108, n1524, n1363, n1447, n1361);
nor  g1906 (n2224, n432, n1515, n1580, n625);
and  g1907 (n1866, n1585, n1519, n893, n1200);
and  g1908 (n1700, n1613, n1566, n1583, n818);
and  g1909 (n1820, n1391, n460, n1481, n1444);
xnor g1910 (n1785, n1588, n1610, n1194, n985);
or   g1911 (n1792, n1335, n1071, n430, n1317);
and  g1912 (n1961, n495, n1287, n459, n1462);
xnor g1913 (n1757, n980, n517, n1440, n624);
or   g1914 (n1908, n1569, n1507, n1389, n1150);
and  g1915 (n1803, n1139, n1554, n1532, n1283);
xor  g1916 (n1721, n1426, n1341, n1353, n1527);
nand g1917 (n2090, n741, n1270, n1451, n1054);
xnor g1918 (n2236, n1277, n466, n1326, n1521);
xnor g1919 (n2126, n1100, n1336, n932, n1146);
xnor g1920 (n2166, n1564, n669, n1183, n1435);
and  g1921 (n1832, n1407, n1634, n1138, n1178);
nand g1922 (n1902, n1366, n1136, n1307, n1582);
and  g1923 (n1843, n1455, n800, n1242, n705);
nand g1924 (n1798, n1504, n1293, n1588, n1614);
xor  g1925 (n1740, n1319, n614, n1300, n1521);
nand g1926 (n1733, n1193, n1566, n1601, n1495);
nor  g1927 (n2142, n644, n998, n1356, n1402);
or   g1928 (n2000, n1586, n1375, n481, n1159);
nand g1929 (n1884, n1633, n1373, n655, n435);
xnor g1930 (n1926, n1217, n1408, n1118, n1097);
xnor g1931 (n1861, n968, n1313, n1472, n1269);
xnor g1932 (n1984, n1394, n768, n449, n1350);
xnor g1933 (n2176, n648, n1161, n659, n1499);
nand g1934 (n1837, n1403, n1323, n907, n813);
nand g1935 (n1745, n665, n1247, n1326, n1629);
nand g1936 (n1940, n926, n850, n525, n536);
xnor g1937 (n1913, n1615, n1132, n825, n1542);
nand g1938 (n2063, n1617, n1282, n1285, n1395);
or   g1939 (n1989, n726, n1288, n1284, n1326);
and  g1940 (n1856, n1596, n1231, n1129, n1547);
or   g1941 (n2159, n1391, n1636, n1447, n662);
or   g1942 (n1914, n1061, n562, n1415, n1576);
nor  g1943 (n1782, n1363, n1347, n1585, n1452);
nand g1944 (n1751, n1479, n1619, n1567, n1503);
and  g1945 (n1974, n1406, n1368, n1160, n467);
xnor g1946 (n2170, n1416, n930, n1327, n585);
nor  g1947 (n1859, n814, n1377, n983, n1030);
and  g1948 (n1943, n863, n1542, n1314, n501);
xor  g1949 (n1741, n1210, n1052, n615, n1353);
xnor g1950 (n1852, n1410, n1366, n529, n1202);
xor  g1951 (n2087, n1523, n794, n1522, n1315);
and  g1952 (n1871, n619, n1293, n1596, n1349);
xnor g1953 (n2130, n881, n1415, n1199, n943);
or   g1954 (n2098, n1579, n1376, n695, n919);
or   g1955 (n2155, n835, n1380, n515, n510);
nor  g1956 (n1877, n570, n1625, n1550, n1435);
xor  g1957 (n1988, n1055, n847, n1583, n903);
nand g1958 (n1919, n512, n1567, n1574, n1259);
and  g1959 (n1761, n1318, n1309, n1489, n1605);
xnor g1960 (n2123, n537, n816, n1432, n1310);
or   g1961 (n2109, n1503, n787, n1516, n1315);
or   g1962 (n1706, n844, n1261, n1527, n1575);
nand g1963 (n2032, n1414, n1590, n1264, n1484);
xnor g1964 (n1701, n1593, n628, n1534, n1300);
nand g1965 (n1956, n1335, n798, n1174, n572);
and  g1966 (n1742, n1555, n478, n1416, n1384);
xor  g1967 (n1845, n573, n1444, n661, n1485);
xor  g1968 (n2116, n1469, n1328, n1400, n1236);
and  g1969 (n1807, n1338, n1432, n1043, n1372);
nor  g1970 (n2049, n1035, n1498, n1491, n1175);
nor  g1971 (n2227, n1329, n1454, n567, n773);
and  g1972 (n1685, n952, n1384, n1499, n587);
and  g1973 (n1686, n589, n795, n1047, n1454);
nor  g1974 (n2085, n1364, n490, n1404, n744);
nor  g1975 (n1818, n1433, n1505, n1283, n1545);
nor  g1976 (n2163, n1484, n1588, n1482, n627);
xnor g1977 (n1825, n1233, n1511, n1418, n1318);
xor  g1978 (n2156, n1596, n1382, n540, n1526);
and  g1979 (n1941, n810, n1613, n1620, n1303);
nor  g1980 (n1853, n535, n1632, n1053, n672);
nor  g1981 (n1822, n1547, n1422, n1320, n895);
xnor g1982 (n2018, n1409, n737, n890, n1410);
xor  g1983 (n1800, n1458, n1271, n1492, n1562);
or   g1984 (n2178, n1525, n588, n1500, n471);
and  g1985 (n1917, n645, n1280, n1488, n1389);
nor  g1986 (n1909, n1535, n873, n1310, n1265);
and  g1987 (n1955, n1023, n1471, n1530, n1365);
nand g1988 (n2225, n1581, n1582, n1323, n1298);
nand g1989 (n2057, n1367, n1275, n1632, n1415);
xor  g1990 (n2154, n555, n1427, n1513, n1633);
and  g1991 (n2078, n1267, n1409, n1580, n1360);
and  g1992 (n2053, n446, n494, n853, n658);
and  g1993 (n2081, n1522, n1514, n601, n593);
xor  g1994 (n1934, n1473, n1541, n1448, n1535);
nand g1995 (n1781, n1333, n1512, n710, n987);
xor  g1996 (n2045, n1298, n1552, n1277, n1402);
xor  g1997 (n2257, n686, n516, n977, n996);
nand g1998 (n2035, n1470, n1607, n1529, n1196);
xor  g1999 (n1738, n1205, n1364, n1297, n1305);
nand g2000 (n2062, n1559, n715, n797, n683);
nand g2001 (n1694, n1592, n1290, n1345, n1439);
and  g2002 (n1892, n1424, n763, n1348, n1589);
and  g2003 (n2246, n785, n1603, n842, n1330);
and  g2004 (n2221, n1375, n486, n1367, n1560);
xnor g2005 (n2259, n1477, n912, n690, n1416);
nor  g2006 (n1933, n1528, n1603, n638, n1278);
xnor g2007 (n1901, n1539, n660, n799, n1610);
xnor g2008 (n1996, n1500, n1281, n1570, n1633);
and  g2009 (n2244, n1549, n1091, n1540, n815);
nand g2010 (n2075, n1520, n1384, n838, n1593);
xor  g2011 (n2084, n966, n1621, n1325, n1622);
or   g2012 (n2206, n428, n856, n1597, n1461);
and  g2013 (n1750, n1595, n1273, n1514, n1333);
nor  g2014 (n1809, n902, n1206, n670, n1300);
or   g2015 (n2152, n906, n1605, n872, n1198);
nand g2016 (n2072, n1024, n1487, n830, n546);
nor  g2017 (n1775, n1281, n964, n1609, n666);
nand g2018 (n2019, n1403, n1274, n1289, n689);
nor  g2019 (n2167, n849, n1209, n1555, n1463);
and  g2020 (n2144, n1534, n1295, n739, n559);
nor  g2021 (n2196, n1313, n1352, n1271, n1463);
and  g2022 (n1802, n600, n1562, n1572, n1635);
xnor g2023 (n1975, n1547, n954, n1426, n1165);
and  g2024 (n2248, n1423, n676, n1291, n1034);
nand g2025 (n1788, n629, n472, n1536, n1606);
nand g2026 (n2023, n1117, n1240, n1344, n1541);
or   g2027 (n1880, n1354, n639, n1339, n1468);
nand g2028 (n1752, n1333, n1394, n840, n1131);
or   g2029 (n2031, n653, n1399, n1468, n761);
or   g2030 (n1697, n1219, n1031, n1571, n1010);
xnor g2031 (n2233, n1526, n934, n1307, n1257);
and  g2032 (n1844, n1369, n1457, n1544, n1528);
xor  g2033 (n2105, n692, n1286, n1539, n1428);
xor  g2034 (n1900, n1540, n1248, n1412, n1584);
nand g2035 (n2262, n1149, n1488, n1336, n1044);
and  g2036 (n2001, n843, n1628, n1338, n1365);
xor  g2037 (n1746, n554, n1078, n1587, n1314);
or   g2038 (n2250, n1361, n445, n1436, n1518);
xor  g2039 (n1711, n1556, n1057, n1381, n1355);
or   g2040 (n1911, n1485, n1522, n1275, n1459);
nor  g2041 (n1890, n1368, n1398, n1618, n1479);
xnor g2042 (n2029, n502, n1145, n1520, n772);
nor  g2043 (n1979, n1182, n1422, n1172, n1424);
and  g2044 (n1999, n557, n1471, n1358, n524);
nor  g2045 (n2118, n1512, n1441, n974, n1459);
nor  g2046 (n2245, n812, n1553, n1271, n1490);
nand g2047 (n1759, n1221, n1540, n488, n1469);
xnor g2048 (n1944, n860, n915, n498, n1609);
nor  g2049 (n1885, n1565, n1388, n1519, n1420);
nand g2050 (n2017, n1355, n534, n1628, n1545);
xor  g2051 (n2037, n865, n1417, n643, n1156);
or   g2052 (n1851, n1545, n1355, n1374, n1133);
xor  g2053 (n1970, n1379, n1425, n1305, n1614);
nor  g2054 (n1839, n671, n1296, n1230, n1227);
nor  g2055 (n2220, n1465, n1349, n677, n1439);
xnor g2056 (n2027, n1398, n1063, n738, n1443);
and  g2057 (n2222, n714, n1458, n1126, n551);
or   g2058 (n2046, n1046, n1277, n1272, n1460);
nand g2059 (n2092, n1306, n1376, n1533, n1204);
nand g2060 (n2114, n1632, n862, n1616, n1280);
nor  g2061 (n2012, n1500, n1464, n612, n1536);
xnor g2062 (n2165, n1537, n1152, n474, n1539);
nor  g2063 (n2135, n1508, n1415, n1147, n1008);
or   g2064 (n1893, n1303, n1570, n1094, n1332);
xor  g2065 (n1915, n749, n1565, n1466, n1386);
and  g2066 (n1715, n1294, n1294, n1610, n1245);
xnor g2067 (n2089, n1598, n1039, n1388, n1481);
xnor g2068 (n1842, n918, n1619, n1413, n1252);
and  g2069 (n1993, n1510, n1504, n1311, n1329);
nand g2070 (n1728, n1295, n1553, n711, n595);
xor  g2071 (n1992, n1390, n1564, n1525, n1426);
xor  g2072 (n1954, n976, n1511, n892, n1060);
or   g2073 (n1894, n1343, n1026, n1458, n1358);
or   g2074 (n1976, n1281, n1334, n1001, n1408);
or   g2075 (n1830, n1482, n586, n1501, n1452);
xnor g2076 (n1864, n1495, n1586, n1571, n1215);
nand g2077 (n1698, n1494, n1593, n1594, n1507);
xor  g2078 (n2204, n1490, n1625, n921, n867);
xor  g2079 (n2068, n1337, n1483, n1316, n1532);
or   g2080 (n2200, n1279, n1558, n923, n469);
nand g2081 (n2139, n1353, n1290, n1299, n1191);
xor  g2082 (n1756, n1626, n1623, n1557, n584);
or   g2083 (n2151, n1481, n1493, n582, n1380);
and  g2084 (n1765, n931, n967, n437, n1357);
or   g2085 (n2047, n1508, n756, n1618, n780);
xnor g2086 (n2208, n1400, n1385, n1401, n1334);
or   g2087 (n1771, n1534, n521, n1275, n1268);
and  g2088 (n1777, n1556, n1401, n1618, n720);
xor  g2089 (n1873, n1383, n1480, n1491, n1450);
nand g2090 (n1967, n913, n656, n887, n1340);
or   g2091 (n2205, n1447, n1600, n1496, n1414);
xor  g2092 (n1823, n1480, n1338, n1395, n1021);
xor  g2093 (n1704, n1316, n1595, n640, n1302);
xor  g2094 (n2086, n1456, n1573, n1189, n1304);
or   g2095 (n1716, n1451, n1594, n965, n990);
or   g2096 (n2209, n1414, n878, n1461, n1246);
and  g2097 (n1938, n1517, n1626, n1625, n1342);
and  g2098 (n1995, n1453, n480, n1457, n1239);
xnor g2099 (n1805, n1566, n1330, n598, n1604);
nor  g2100 (n1985, n1347, n1360, n1368, n864);
and  g2101 (n2141, n1311, n693, n1550, n725);
nand g2102 (n1991, n708, n1391, n1578, n1504);
nor  g2103 (n2229, n1392, n1411, n898, n712);
or   g2104 (n2260, n1405, n470, n1068, n1515);
nor  g2105 (n2038, n1541, n1544, n1511, n1288);
xor  g2106 (n2083, n1499, n1379, n1066, n1455);
and  g2107 (n1936, n1322, n1485, n482, n1496);
xor  g2108 (n2240, n1392, n1418, n1497, n1599);
xor  g2109 (n2212, n443, n866, n1626, n1421);
nand g2110 (n1799, n519, n1308, n717, n599);
and  g2111 (n1787, n1318, n950, n1430, n1483);
and  g2112 (n1714, n578, n757, n1578, n1484);
and  g2113 (n1702, n1569, n680, n1321, n1278);
nor  g2114 (n2131, n1397, n1376, n1567, n1493);
nor  g2115 (n1849, n1475, n713, n1337, n1392);
nand g2116 (n1906, n1393, n949, n1573, n631);
nor  g2117 (n1875, n1399, n434, n1462, n1456);
xor  g2118 (n2231, n1211, n1522, n1552, n1486);
or   g2119 (n1903, n568, n1369, n1306, n1412);
nor  g2120 (n1743, n1027, n1448, n1290, n500);
xnor g2121 (n1895, n439, n565, n1624, n702);
nor  g2122 (n2181, n1579, n1263, n1628, n1267);
and  g2123 (n1929, n1587, n1620, n716, n1601);
xor  g2124 (n2095, n1573, n1298, n1356, n1151);
and  g2125 (n1723, n1382, n728, n1434, n1059);
xor  g2126 (n1925, n1533, n854, n1506, n1153);
or   g2127 (n1855, n1348, n1357, n1610, n1494);
nand g2128 (n1862, n1538, n1549, n1629, n1095);
nor  g2129 (n2158, n1309, n1452, n1444, n1549);
or   g2130 (n1784, n574, n1506, n1437, n1238);
or   g2131 (n2117, n1540, n1373, n1207, n1360);
and  g2132 (n2249, n746, n1545, n1565, n1546);
xor  g2133 (n2080, n1365, n1354, n1292, n1442);
nor  g2134 (n1703, n1329, n778, n1359, n1421);
or   g2135 (n1972, n1488, n1498, n1607, n1564);
nor  g2136 (n2242, n1327, n1442, n1373, n1076);
and  g2137 (n2180, n762, n1112, n528, n1420);
xnor g2138 (n2193, n1544, n1264, n1038, n1274);
nand g2139 (n2138, n1579, n1260, n709, n1334);
nor  g2140 (n1931, n751, n837, n1519, n1520);
and  g2141 (n1768, n1561, n1432, n1185, n1627);
xnor g2142 (n1930, n1289, n724, n1345, n1367);
and  g2143 (n2147, n1589, n1279, n1473, n1229);
and  g2144 (n2203, n462, n1363, n1272, n1263);
nor  g2145 (n1960, n1478, n608, n1598, n781);
or   g2146 (n2058, n1276, n1324, n1412, n1303);
xor  g2147 (n1854, n1487, n1387, n703, n1272);
and  g2148 (n1735, n1516, n571, n908, n1331);
or   g2149 (n2070, n487, n1296, n1474, n1320);
nor  g2150 (n2128, n1342, n1062, n1244, n1409);
nor  g2151 (n2002, n1417, n1292, n697, n1448);
nor  g2152 (n2093, n834, n1591, n1468, n1359);
and  g2153 (n1928, n1377, n1378, n541, n1110);
nand g2154 (n1983, n808, n1241, n1419, n583);
xor  g2155 (n2050, n1355, n758, n1475, n783);
xor  g2156 (n1725, n1311, n1113, n995, n1367);
nand g2157 (n1737, n1371, n1575, n1557, n975);
or   g2158 (n2183, n1410, n505, n1273, n1503);
nand g2159 (n1981, n1375, n1572, n942, n1543);
and  g2160 (n2010, n654, n1527, n1590, n882);
xor  g2161 (n2177, n886, n1467, n1568, n636);
xnor g2162 (n1986, n1557, n1554, n1103, n1345);
nor  g2163 (n1780, n1510, n904, n427, n823);
nor  g2164 (n2150, n1278, n1634, n1583, n1122);
nand g2165 (n2036, n827, n1405, n880, n1349);
and  g2166 (n2003, n1548, n1445, n1028, n1600);
xor  g2167 (n2218, n1316, n1386, n1302, n1597);
or   g2168 (n2082, n1344, n1636, n1592, n1608);
or   g2169 (n2185, n1476, n569, n1602, n550);
nand g2170 (n1965, n1195, n1395, n1268, n1340);
nand g2171 (n2097, n1297, n958, n1261, n1058);
xnor g2172 (n2136, n468, n1556, n1292, n1164);
or   g2173 (n1813, n1478, n1374, n1511, n1350);
and  g2174 (n2066, n1364, n1531, n1577, n1489);
or   g2175 (n1888, n910, n1302, n1372, n859);
and  g2176 (n1898, n1234, n1377, n1439, n1555);
xor  g2177 (n2214, n1595, n1294, n1607, n1569);
xor  g2178 (n1927, n730, n1323, n1462, n947);
xor  g2179 (n2258, n518, n1346, n1537, n845);
xnor g2180 (n1932, n1621, n1135, n696, n1446);
xnor g2181 (n1695, n1310, n461, n1531, n1383);
and  g2182 (n2256, n1407, n1266, n1125, n1617);
nand g2183 (n2241, n1392, n1328, n1621, n1382);
and  g2184 (n2187, n1470, n1000, n1314, n1051);
and  g2185 (n2228, n883, n1507, n1502, n1243);
or   g2186 (n2146, n1222, n1410, n1563, n1494);
or   g2187 (n1815, n1036, n1575, n1505, n1490);
nor  g2188 (n2112, n1401, n1376, n1286, n507);
xor  g2189 (n2096, n1253, n1499, n1400, n1273);
and  g2190 (n2006, n1285, n1379, n1400, n1423);
or   g2191 (n1693, n936, n657, n858, n609);
or   g2192 (n2265, n1592, n1404, n1477, n836);
or   g2193 (n1969, n1629, n1049, n1491, n634);
and  g2194 (n1729, n688, n1548, n1397, n1259);
or   g2195 (n2226, n1391, n1470, n1562, n1313);
xor  g2196 (n1838, n1312, n1370, n1358, n1336);
xnor g2197 (n2107, n1212, n1140, n1562, n951);
nor  g2198 (n2022, n1387, n828, n1429, n1003);
and  g2199 (n1692, n1307, n1634, n1533, n592);
or   g2200 (n1863, n1300, n1561, n687, n1577);
xnor g2201 (n1966, n1070, n1448, n766, n649);
nor  g2202 (n2255, n1465, n547, n1632, n1581);
nand g2203 (n2164, n527, n1396, n1338, n1419);
and  g2204 (n2197, n790, n1408, n869, n1528);
and  g2205 (n2122, n1072, n718, n1538, n846);
or   g2206 (n1696, n1298, n1584, n1616, n1544);
xnor g2207 (n1899, n1573, n1313, n771, n1328);
or   g2208 (n1708, n1466, n1445, n1528, n438);
nor  g2209 (n1814, n1517, n1431, n477, n1407);
nand g2210 (n2021, n1619, n1033, n1559, n1630);
xor  g2211 (n1762, n663, n1390, n1585, n1568);
or   g2212 (n2073, n1287, n1482, n1560, n1143);
and  g2213 (n1717, n1581, n944, n1306, n1534);
or   g2214 (n1718, n1321, n1521, n617, n1515);
and  g2215 (n1858, n423, n1309, n767, n1482);
xnor g2216 (n1840, n1331, n700, n455, n1622);
and  g2217 (n2232, n1615, n1394, n1523, n1543);
and  g2218 (n2179, n1098, n447, n1444, n1305);
xnor g2219 (n2005, n1279, n1608, n1283, n1082);
nor  g2220 (n1857, n1550, n784, n1339, n1050);
xor  g2221 (n2161, n1580, n1614, n526, n1396);
or   g2222 (n1939, n1549, n1362, n776, n1431);
xnor g2223 (n1690, n1606, n1398, n1559, n1460);
and  g2224 (n2048, n1411, n1436, n1590, n1342);
nand g2225 (n1891, n1494, n1285, n1086, n1228);
nand g2226 (n1987, n1399, n1584, n1386, n1012);
nand g2227 (n1948, n1403, n1623, n961, n1489);
or   g2228 (n1945, n1636, n909, n1286, n1377);
xnor g2229 (n2182, n1474, n458, n1048, n635);
nand g2230 (n2014, n603, n929, n1502, n1032);
and  g2231 (n2219, n997, n1325, n1539, n1445);
nand g2232 (n1739, n1320, n1492, n1312, n453);
nand g2233 (n1748, n1296, n1267, n1628, n1312);
xnor g2234 (n2007, n1380, n897, n1455, n1566);
nand g2235 (n2252, n1612, n549, n1378, n1278);
and  g2236 (n1811, n1584, n1340, n1325, n1514);
xor  g2237 (n1699, n1025, n496, n754, n984);
nand g2238 (n1709, n1388, n1264, n1166, n545);
or   g2239 (n2202, n1560, n1335, n1619, n1388);
nand g2240 (n2044, n1324, n1599, n1623, n1529);
and  g2241 (n1963, n1611, n1371, n1339, n1473);
nand g2242 (n1918, n1107, n765, n1615, n1322);
not  g2243 (n2275, n1736);
not  g2244 (n2303, n1701);
not  g2245 (n2278, n1695);
buf  g2246 (n2272, n1723);
not  g2247 (n2296, n1801);
buf  g2248 (n2288, n1763);
buf  g2249 (n2313, n1714);
buf  g2250 (n2328, n1782);
buf  g2251 (n2326, n1765);
buf  g2252 (n2289, n1848);
buf  g2253 (n2271, n1740);
not  g2254 (n2323, n1775);
buf  g2255 (n2287, n1831);
not  g2256 (n2314, n1692);
buf  g2257 (n2306, n1803);
not  g2258 (n2305, n1724);
not  g2259 (n2291, n1698);
buf  g2260 (n2317, n1757);
buf  g2261 (n2281, n1824);
not  g2262 (n2297, n1716);
not  g2263 (n2292, n1713);
not  g2264 (n2273, n1835);
buf  g2265 (n2319, n1709);
not  g2266 (n2274, n1784);
and  g2267 (n2283, n1794, n1762, n1727, n1797);
xnor g2268 (n2312, n1753, n1838, n1821, n1845);
nor  g2269 (n2322, n1688, n1705, n1818, n1697);
nand g2270 (n2277, n1707, n1843, n1820, n1702);
nand g2271 (n2325, n1844, n1770, n1777, n1706);
xor  g2272 (n2321, n1836, n1816, n1790, n1788);
and  g2273 (n2316, n1834, n1850, n1754, n1822);
xnor g2274 (n2285, n1833, n1800, n1729, n1718);
xor  g2275 (n2293, n1774, n1773, n1819, n1793);
nand g2276 (n2270, n1852, n1847, n1733, n1725);
or   g2277 (n2311, n1791, n1840, n1826, n1813);
nand g2278 (n2269, n1812, n1696, n1738, n1804);
and  g2279 (n2299, n1712, n1828, n1783, n1719);
xnor g2280 (n2298, n1715, n1717, n1810, n1722);
xnor g2281 (n2309, n1741, n1743, n1778, n1750);
xnor g2282 (n2280, n1798, n1690, n1846, n1785);
nor  g2283 (n2301, n1825, n1815, n1809, n1699);
xor  g2284 (n2294, n1689, n1787, n1829, n1772);
and  g2285 (n2284, n1830, n1720, n1841, n1807);
or   g2286 (n2318, n1764, n1742, n1756, n1710);
nand g2287 (n2295, n1759, n1823, n1711, n1761);
xor  g2288 (n2324, n1817, n1795, n1769, n1731);
nand g2289 (n2286, n1780, n1732, n1748, n1746);
nor  g2290 (n2307, n1728, n1726, n1745, n1693);
nor  g2291 (n2282, n1708, n1694, n1839, n1849);
or   g2292 (n2279, n1703, n1811, n1808, n1766);
nor  g2293 (n2320, n1751, n1827, n1771, n1832);
or   g2294 (n2302, n1851, n1735, n1747, n1734);
xnor g2295 (n2304, n1767, n1686, n1837, n1842);
and  g2296 (n2300, n1755, n1758, n1737, n1744);
xnor g2297 (n2308, n1802, n1814, n1752, n1760);
or   g2298 (n2276, n1749, n1691, n1776, n1768);
nor  g2299 (n2310, n1786, n1685, n1779, n1721);
xnor g2300 (n2315, n1700, n1806, n1792, n1739);
nor  g2301 (n2327, n1781, n1730, n1687, n1796);
nor  g2302 (n2290, n1805, n1704, n1789, n1799);
not  g2303 (n2331, n2278);
not  g2304 (n2335, n2283);
buf  g2305 (n2333, n2285);
not  g2306 (n2329, n2274);
buf  g2307 (n2336, n2282);
buf  g2308 (n2334, n2275);
and  g2309 (n2337, n2272, n2280, n2269, n2273);
nand g2310 (n2332, n2276, n2271, n2279, n2270);
or   g2311 (n2330, n2277, n2286, n2284, n2281);
not  g2312 (n2346, n2329);
not  g2313 (n2347, n2332);
not  g2314 (n2357, n2330);
not  g2315 (n2345, n2333);
buf  g2316 (n2338, n2332);
buf  g2317 (n2355, n2329);
buf  g2318 (n2353, n2330);
buf  g2319 (n2348, n2331);
buf  g2320 (n2352, n2331);
buf  g2321 (n2354, n2331);
buf  g2322 (n2356, n2330);
not  g2323 (n2349, n2332);
buf  g2324 (n2344, n2331);
not  g2325 (n2340, n2333);
not  g2326 (n2341, n2329);
not  g2327 (n2339, n2332);
not  g2328 (n2350, n2329);
not  g2329 (n2351, n2330);
not  g2330 (n2342, n2333);
buf  g2331 (n2343, n2333);
buf  g2332 (n2374, n2287);
not  g2333 (n2359, n2356);
buf  g2334 (n2371, n2347);
not  g2335 (n2372, n2350);
xnor g2336 (n2375, n2336, n422);
or   g2337 (n2363, n2345, n2348, n1638, n2336);
and  g2338 (n2364, n2354, n21, n2335, n2334);
nor  g2339 (n2360, n2340, n22, n2336, n2352);
nand g2340 (n2365, n2355, n1853, n2342, n2341);
xor  g2341 (n2368, n2349, n2337, n1638, n2357);
xnor g2342 (n2366, n2288, n2343, n2338, n2344);
xnor g2343 (n2373, n2335, n21, n2352);
nor  g2344 (n2361, n1639, n2335, n2339, n2351);
nor  g2345 (n2370, n2346, n2334, n2354, n2356);
nand g2346 (n2362, n2355, n1638, n2337, n22);
xor  g2347 (n2358, n2337, n1639, n2334);
or   g2348 (n2367, n22, n2353, n2334);
and  g2349 (n2369, n2357, n2335, n1638, n2336);
buf  g2350 (n2381, n106);
buf  g2351 (n2384, n2373);
buf  g2352 (n2379, n2375);
not  g2353 (n2383, n2368);
buf  g2354 (n2386, n2359);
buf  g2355 (n2388, n2362);
buf  g2356 (n2380, n2372);
buf  g2357 (n2391, n2364);
buf  g2358 (n2377, n2365);
buf  g2359 (n2376, n105);
buf  g2360 (n2378, n2370);
not  g2361 (n2389, n2363);
nand g2362 (n2382, n2369, n2367, n106);
and  g2363 (n2390, n2360, n2361, n105);
xor  g2364 (n2387, n2371, n2374, n2366);
xnor g2365 (n2385, n2358, n105);
or   g2366 (n2392, n2378, n2379, n2376, n2377);
buf  g2367 (n2394, n2392);
or   g2368 (n2393, n2392, n23, n22);
not  g2369 (n2395, n2394);
not  g2370 (n2400, n2394);
buf  g2371 (n2397, n2393);
buf  g2372 (n2398, n2394);
not  g2373 (n2396, n2394);
buf  g2374 (n2399, n2393);
not  g2375 (n2401, n2393);
not  g2376 (n2403, n2398);
buf  g2377 (n2402, n2398);
buf  g2378 (n2407, n2396);
not  g2379 (n2405, n2395);
and  g2380 (n2404, n2395, n2397, n2398);
and  g2381 (n2406, n2397, n2396, n2395);
not  g2382 (n2409, n1641);
xnor g2383 (n2411, n2406, n1640, n2405);
and  g2384 (n2408, n2407, n1639, n1640, n2403);
xnor g2385 (n2410, n1640, n1640, n2404, n2402);
xor  g2386 (n2412, n1855, n1854, n1856, n2408);
and  g2387 (n2413, n2412, n2294, n2289, n2292);
nor  g2388 (n2414, n2290, n2293, n2412, n2291);
not  g2389 (n2418, n2414);
not  g2390 (n2415, n2413);
not  g2391 (n2421, n2414);
buf  g2392 (n2422, n2414);
buf  g2393 (n2417, n2413);
not  g2394 (n2416, n2413);
not  g2395 (n2419, n2413);
buf  g2396 (n2420, n2414);
nor  g2397 (n2433, n2420, n2417);
nor  g2398 (n2434, n1641, n25);
xnor g2399 (n2435, n25, n2422);
xnor g2400 (n2436, n2417, n25);
xor  g2401 (n2439, n23, n2418);
nand g2402 (n2424, n2419, n2381);
or   g2403 (n2431, n2419, n2380);
nor  g2404 (n2423, n2296, n2422);
nor  g2405 (n2425, n2295, n2415);
xor  g2406 (n2430, n2420, n2421);
or   g2407 (n2428, n2297, n23);
nand g2408 (n2429, n24, n2422);
xnor g2409 (n2437, n25, n2421);
xnor g2410 (n2426, n2415, n24);
buf  g2411 (n2440, n2416);
nor  g2412 (n2427, n24, n1641);
nand g2413 (n2438, n2418, n24);
xnor g2414 (n2432, n2421, n23);
not  g2415 (n2456, n2430);
not  g2416 (n2449, n2434);
buf  g2417 (n2452, n2428);
not  g2418 (n2446, n2431);
not  g2419 (n2448, n2438);
not  g2420 (n2450, n2423);
buf  g2421 (n2451, n2425);
not  g2422 (n2442, n2427);
not  g2423 (n2455, n2437);
not  g2424 (n2447, n2432);
not  g2425 (n2453, n2435);
buf  g2426 (n2445, n2426);
buf  g2427 (n2441, n2433);
not  g2428 (n2454, n2429);
buf  g2429 (n2443, n2436);
buf  g2430 (n2444, n2424);
nor  g2431 (n2457, n2456, n2451, n2453);
xor  g2432 (n2465, n2451, n2456, n2454);
xor  g2433 (n2464, n2456, n2451, n2382, n2445);
xor  g2434 (n2460, n2454, n2455, n2450);
and  g2435 (n2466, n2441, n2453, n2442, n2452);
nor  g2436 (n2461, n2387, n2455, n2452, n2449);
or   g2437 (n2459, n2446, n2385, n2444, n2455);
and  g2438 (n2458, n2454, n2383, n2386, n2453);
or   g2439 (n2463, n2452, n2447, n2453, n2448);
nand g2440 (n2462, n2454, n2384, n2452, n2443);
buf  g2441 (n2473, n2460);
not  g2442 (n2474, n2463);
buf  g2443 (n2471, n2461);
not  g2444 (n2468, n2398);
buf  g2445 (n2470, n2459);
xor  g2446 (n2467, n2466, n1641, n1642);
or   g2447 (n2469, n2465, n1642, n2464);
nand g2448 (n2472, n2462, n2399, n1642);
nand g2449 (n2483, n2472, n1870);
xor  g2450 (n2490, n2400, n1858);
xor  g2451 (n2481, n2468, n2472);
buf  g2452 (n2486, n2469);
xor  g2453 (n2491, n1857, n1860);
and  g2454 (n2494, n1866, n1859);
or   g2455 (n2476, n1862, n1864);
nand g2456 (n2493, n1868, n2401);
nand g2457 (n2478, n2473, n2471);
xnor g2458 (n2487, n2471, n2473);
and  g2459 (n2480, n2474, n2468);
buf  g2460 (n2492, n2470);
or   g2461 (n2489, n1865, n1863);
nand g2462 (n2475, n1871, n2399);
or   g2463 (n2479, n2470, n1867);
nand g2464 (n2485, n2400, n2467);
xor  g2465 (n2495, n2400, n2467);
nor  g2466 (n2482, n2399, n2472);
xor  g2467 (n2477, n2467, n1872);
nand g2468 (n2498, n2474, n2400);
and  g2469 (n2484, n2469, n2401);
or   g2470 (n2488, n2473, n2471);
nor  g2471 (n2497, n2474, n2468);
xnor g2472 (n2496, n1869, n1861);
buf  g2473 (n2501, n2475);
not  g2474 (n2507, n2482);
buf  g2475 (n2502, n2479);
not  g2476 (n2504, n2477);
not  g2477 (n2500, n2481);
not  g2478 (n2508, n2483);
buf  g2479 (n2499, n2480);
not  g2480 (n2506, n2484);
not  g2481 (n2505, n2476);
not  g2482 (n2503, n2478);
xnor g2483 (n2521, n2504, n2500, n2501, n2320);
nor  g2484 (n2520, n2507, n2502, n2508, n2309);
nor  g2485 (n2516, n2307, n2305, n2504, n2315);
nand g2486 (n2525, n2501, n2501, n2505, n2324);
xnor g2487 (n2524, n2507, n2500, n2298, n2505);
xnor g2488 (n2515, n2303, n2505, n2302);
xor  g2489 (n2513, n2311, n2300, n2502, n2319);
xnor g2490 (n2517, n2313, n2322, n2308, n2318);
or   g2491 (n2522, n2299, n2503, n2506, n2314);
and  g2492 (n2510, n2316, n2508, n2506, n2503);
and  g2493 (n2518, n2503, n2506, n2502, n2312);
nand g2494 (n2512, n2499, n2500, n2301, n2321);
xnor g2495 (n2519, n2503, n2504, n2323, n2499);
nor  g2496 (n2509, n2500, n2325, n2317, n2502);
xnor g2497 (n2511, n2507, n2506, n2310, n2499);
xor  g2498 (n2514, n2501, n2507, n2304, n2508);
xnor g2499 (n2523, n2306, n2504, n2508, n2499);
buf  g2500 (n2540, n1887);
not  g2501 (n2530, n1886);
and  g2502 (n2532, n2328, n2408);
nand g2503 (n2535, n1882, n2326, n2411, n1881);
nand g2504 (n2539, n2408, n2327, n2509, n2514);
and  g2505 (n2536, n2516, n2409, n2524, n2513);
xor  g2506 (n2537, n1880, n2409, n2411, n2410);
xnor g2507 (n2528, n1877, n2525, n2337, n1874);
xor  g2508 (n2529, n2410, n1879, n2515, n2522);
nand g2509 (n2531, n1885, n1878, n1888, n1873);
xnor g2510 (n2527, n1875, n2410, n1883, n1884);
or   g2511 (n2534, n2411, n2510, n2521, n2511);
nor  g2512 (n2538, n2410, n2408, n1876, n2411);
xnor g2513 (n2526, n2517, n2518, n2409);
xnor g2514 (n2533, n2512, n2520, n2519, n2523);
buf  g2515 (n2547, n1896);
buf  g2516 (n2543, n1901);
buf  g2517 (n2548, n1892);
not  g2518 (n2542, n1890);
buf  g2519 (n2545, n2529);
not  g2520 (n2556, n1893);
not  g2521 (n2551, n2528);
not  g2522 (n2549, n2535);
not  g2523 (n2555, n2536);
nor  g2524 (n2552, n1900, n2532, n2531, n1891);
nand g2525 (n2553, n1898, n2530, n2533, n1906);
nand g2526 (n2554, n2537, n1902, n1905, n2540);
and  g2527 (n2544, n1908, n1907, n1903, n2526);
xor  g2528 (n2546, n1895, n2527, n2538, n2539);
xnor g2529 (n2541, n1904, n2534, n1894, n1889);
nand g2530 (n2550, n2412, n2540, n1897, n1899);
nor  g2531 (n2590, n2545, n1665, n1662, n1660);
nand g2532 (n2587, n1672, n1659, n1683, n1649);
xor  g2533 (n2608, n2546, n1670, n1661);
nor  g2534 (n2572, n1684, n1678, n1653, n1647);
xor  g2535 (n2581, n2547, n1651, n2552, n1678);
xor  g2536 (n2592, n1682, n1648, n1677, n2391);
xnor g2537 (n2582, n1668, n1659, n2556, n2544);
xor  g2538 (n2579, n1664, n1653, n2543, n1643);
xnor g2539 (n2560, n1657, n1660, n1648, n1654);
xnor g2540 (n2607, n1679, n1672, n1677, n1647);
and  g2541 (n2584, n1659, n1909, n2551, n2489);
nor  g2542 (n2567, n1661, n2552, n1649, n1663);
and  g2543 (n2602, n2546, n1667, n2495, n2547);
or   g2544 (n2586, n2550, n1680, n1651, n2556);
xor  g2545 (n2611, n2553, n2496, n1666, n1673);
nor  g2546 (n2615, n1676, n2542, n1649, n1670);
nor  g2547 (n2594, n1684, n2553, n1666, n1650);
xor  g2548 (n2620, n2546, n2485, n1684, n1683);
nand g2549 (n2616, n2541, n1650, n2544, n2555);
nor  g2550 (n2565, n1680, n1674, n2545);
nand g2551 (n2618, n1666, n2543, n2549, n1665);
and  g2552 (n2617, n1681, n1653, n1676, n1663);
xor  g2553 (n2557, n1656, n1679, n1673, n1671);
and  g2554 (n2561, n1643, n2494, n2556, n1652);
or   g2555 (n2609, n2548, n1662, n1681, n2545);
nand g2556 (n2596, n2551, n1652, n2553, n1653);
or   g2557 (n2595, n1667, n1662, n1651, n1645);
or   g2558 (n2599, n2550, n1669, n1675, n1651);
xor  g2559 (n2558, n1649, n1674, n2541, n1645);
or   g2560 (n2601, n2554, n2390, n2541, n1676);
or   g2561 (n2604, n2555, n2548, n2486, n1660);
xor  g2562 (n2568, n1645, n1668, n1676, n1683);
or   g2563 (n2570, n1658, n2550, n1657, n1674);
nand g2564 (n2605, n1663, n1656, n1654, n2495);
and  g2565 (n2563, n2547, n1667, n1657, n2552);
xor  g2566 (n2575, n1669, n1645, n1680, n2542);
or   g2567 (n2610, n1654, n2544, n2554, n1660);
nor  g2568 (n2603, n2542, n2542, n1668, n1679);
xnor g2569 (n2585, n1664, n1644, n1673, n1675);
xnor g2570 (n2564, n1681, n1646, n1652, n1678);
xor  g2571 (n2566, n1655, n2548, n1674, n2554);
nor  g2572 (n2574, n1671, n1654, n1661, n1683);
xor  g2573 (n2571, n1659, n2554, n1677, n1668);
or   g2574 (n2562, n1666, n2552, n1664, n2496);
nor  g2575 (n2589, n1657, n1658, n1655, n2549);
nor  g2576 (n2613, n1673, n2493, n1665, n1669);
nor  g2577 (n2600, n2495, n1647, n2488, n1682);
or   g2578 (n2583, n1665, n2551, n1670, n1644);
xor  g2579 (n2614, n2492, n2548, n2551, n1643);
or   g2580 (n2580, n1675, n1648, n1646, n1681);
xor  g2581 (n2606, n2543, n1663, n1643, n1650);
xor  g2582 (n2578, n2389, n2495, n1672);
xnor g2583 (n2576, n2555, n2493, n2549, n2388);
nand g2584 (n2577, n2541, n1644, n1650);
or   g2585 (n2597, n1647, n1680, n2487, n1646);
or   g2586 (n2588, n1682, n2549, n1655, n1678);
xor  g2587 (n2559, n1664, n1646, n2550, n1661);
nand g2588 (n2573, n2556, n1682, n1675, n2491);
xor  g2589 (n2591, n1671, n1655, n1656, n2555);
xnor g2590 (n2612, n2543, n1671, n2544, n2490);
nand g2591 (n2593, n1652, n2553, n2496, n1677);
nor  g2592 (n2619, n1662, n1658, n1669, n2547);
and  g2593 (n2598, n1684, n2494, n1648, n1679);
and  g2594 (n2569, n1656, n2546, n1667, n1658);
or   g2595 (n2677, n2087, n2085, n1938, n2606);
nand g2596 (n2622, n2594, n2044, n2221, n2176);
xor  g2597 (n2715, n2093, n2192, n2012, n1977);
or   g2598 (n2638, n2143, n2051, n2108, n2572);
nand g2599 (n2680, n2096, n2594, n2159, n1982);
nand g2600 (n2727, n2580, n2605, n2040, n2567);
xor  g2601 (n2707, n2614, n2147, n2042, n2039);
and  g2602 (n2662, n2109, n2114, n2581, n2161);
nand g2603 (n2722, n2239, n2223, n2617, n1966);
or   g2604 (n2667, n2104, n2025, n2247, n2002);
xnor g2605 (n2628, n2575, n2153, n2243, n1912);
nand g2606 (n2669, n2217, n2257, n2615, n2244);
xnor g2607 (n2639, n2105, n2057, n2584, n2035);
nor  g2608 (n2731, n2249, n2578, n2256, n2056);
or   g2609 (n2718, n2082, n1994, n2194, n2053);
nor  g2610 (n2642, n2229, n2614, n2561, n2140);
or   g2611 (n2655, n2066, n2148, n2033, n2260);
or   g2612 (n2735, n2602, n2618, n2565, n2001);
nand g2613 (n2635, n1942, n2185, n2052, n2571);
nor  g2614 (n2630, n2186, n1988, n1932, n2055);
nor  g2615 (n2661, n2589, n1923, n2585, n2224);
nor  g2616 (n2656, n2162, n1975, n2157, n2058);
xnor g2617 (n2621, n2102, n2582, n2592, n2599);
or   g2618 (n2732, n2591, n2619, n1976, n2575);
and  g2619 (n2676, n2022, n2198, n2191, n2007);
or   g2620 (n2721, n2015, n2258, n2596, n2567);
xnor g2621 (n2706, n2240, n2227, n2248, n2602);
or   g2622 (n2645, n2073, n2593, n2216, n2171);
or   g2623 (n2650, n1951, n2173, n2600, n2251);
and  g2624 (n2685, n1998, n2078, n2094, n1979);
xor  g2625 (n2703, n2195, n2564, n2031, n2152);
xor  g2626 (n2651, n2142, n2620, n2235, n2580);
xnor g2627 (n2654, n2577, n2242, n2168, n2589);
xor  g2628 (n2710, n2010, n2156, n2180, n2061);
and  g2629 (n2670, n2196, n2069, n2588, n1983);
and  g2630 (n2708, n2184, n2189, n2107, n2144);
xnor g2631 (n2728, n2263, n1969, n2129, n2212);
nor  g2632 (n2701, n1944, n2214, n2604, n2182);
nand g2633 (n2647, n2219, n2027, n1913, n2136);
or   g2634 (n2664, n2587, n2106, n1958, n2597);
or   g2635 (n2631, n2172, n1987, n2034, n2618);
or   g2636 (n2657, n2588, n2097, n2111, n2193);
nand g2637 (n2733, n2578, n1930, n2586, n2112);
nor  g2638 (n2692, n2146, n2037, n2086, n2074);
nor  g2639 (n2713, n1949, n2201, n1963, n1939);
or   g2640 (n2725, n2593, n2583, n2181, n2236);
and  g2641 (n2689, n2576, n2026, n2117, n2041);
or   g2642 (n2720, n1972, n1943, n2200, n2590);
xor  g2643 (n2644, n2150, n1911, n2072, n1996);
nand g2644 (n2665, n2211, n2003, n2611, n2265);
and  g2645 (n2712, n1964, n2253, n2178, n1971);
and  g2646 (n2729, n2579, n2127, n1992, n2563);
xor  g2647 (n2653, n2131, n1959, n2226, n2209);
xnor g2648 (n2686, n1929, n1921, n2154, n2213);
xor  g2649 (n2693, n2016, n2206, n2163, n1937);
nand g2650 (n2632, n2067, n2014, n2017, n1981);
or   g2651 (n2640, n2569, n1945, n2151, n2603);
nor  g2652 (n2698, n1985, n2177, n1956, n2116);
and  g2653 (n2679, n2255, n2080, n2188, n2092);
and  g2654 (n2737, n2075, n1993, n1980, n2573);
xor  g2655 (n2678, n2208, n2581, n2113, n1925);
nand g2656 (n2682, n2230, n2081, n2128, n2098);
nand g2657 (n2700, n1920, n2601, n2613, n2063);
xor  g2658 (n2683, n1940, n1991, n2101, n2079);
nor  g2659 (n2624, n1933, n2124, n1955, n2577);
and  g2660 (n2646, n2557, n2175, n2570, n2234);
nand g2661 (n2658, n1990, n2076, n2570, n2254);
nor  g2662 (n2696, n1914, n2062, n2615, n2169);
and  g2663 (n2716, n2077, n2245, n1968, n2585);
xnor g2664 (n2740, n2220, n2103, n2586, n2558);
and  g2665 (n2649, n2203, n2006, n2091, n1950);
xnor g2666 (n2709, n2609, n2610, n2572, n2587);
or   g2667 (n2705, n2207, n2048, n2164, n2599);
xor  g2668 (n2637, n2021, n2167, n2238, n2598);
or   g2669 (n2636, n2008, n2204, n2232, n2083);
xor  g2670 (n2687, n2605, n2607, n2590, n2099);
and  g2671 (n2714, n1924, n2562, n2043, n1973);
nor  g2672 (n2734, n2218, n2574, n1965, n2609);
nand g2673 (n2626, n2011, n2046, n2582, n2250);
xnor g2674 (n2668, n2134, n2612, n2210, n2559);
xnor g2675 (n2726, n2122, n2174, n2613, n2120);
nand g2676 (n2730, n1967, n1989, n1926, n1978);
xor  g2677 (n2694, n2579, n2565, n2030, n1986);
and  g2678 (n2739, n2132, n2560, n2597, n1953);
and  g2679 (n2697, n2619, n2133, n1960, n2566);
xor  g2680 (n2699, n2569, n2029, n1974, n2568);
and  g2681 (n2695, n2205, n2050, n2600, n2024);
and  g2682 (n2623, n2141, n2158, n1962, n2065);
and  g2683 (n2627, n2121, n2267, n2118, n2179);
nor  g2684 (n2629, n2606, n2088, n2126, n2009);
xnor g2685 (n2723, n1928, n2584, n1922, n1957);
xnor g2686 (n2675, n2123, n1948, n2222, n2607);
and  g2687 (n2738, n2612, n2036, n2603, n2090);
xor  g2688 (n2674, n2237, n2047, n2119, n2028);
and  g2689 (n2711, n2145, n1918, n2135, n1995);
nand g2690 (n2719, n2049, n2020, n2054, n2608);
and  g2691 (n2625, n1941, n2611, n2266, n2264);
xor  g2692 (n2643, n2576, n2595, n2095, n2023);
and  g2693 (n2688, n2013, n2160, n2598, n2000);
xnor g2694 (n2691, n2608, n2166, n1915, n2170);
nor  g2695 (n2663, n2130, n2583, n1931, n2241);
xnor g2696 (n2736, n2060, n2268, n1936, n2616);
nand g2697 (n2724, n2591, n2610, n2592, n2125);
xnor g2698 (n2704, n1916, n2138, n2573, n2620);
xnor g2699 (n2648, n2604, n2089, n2616, n2262);
nand g2700 (n2652, n2566, n2137, n2233, n1919);
xor  g2701 (n2634, n1954, n2574, n1970, n2019);
nor  g2702 (n2672, n2190, n2202, n2068, n2004);
xor  g2703 (n2671, n1946, n2100, n1984, n2115);
nor  g2704 (n2690, n2187, n2199, n2045, n2070);
nand g2705 (n2684, n2231, n2246, n2571, n1934);
xor  g2706 (n2633, n1997, n2183, n1961, n2197);
xnor g2707 (n2641, n2005, n2064, n2059, n1927);
or   g2708 (n2659, n1999, n2568, n2071, n2617);
nand g2709 (n2717, n2018, n422, n2165, n2252);
nand g2710 (n2681, n2596, n1952, n2215, n2155);
nand g2711 (n2702, n2110, n2038, n2149, n2601);
xor  g2712 (n2660, n2032, n2228, n1910, n2225);
xor  g2713 (n2666, n2139, n2259, n2084, n1917);
nor  g2714 (n2673, n2261, n2595, n1947, n1935);
xnor g2715 (n2744, n2696, n2725, n2649, n2648);
nor  g2716 (n2748, n2665, n2673, n2675, n2632);
nand g2717 (n2742, n2656, n2726, n2623, n2722);
or   g2718 (n2761, n2662, n2497, n2697, n2723);
or   g2719 (n2743, n2627, n2737, n2657, n2706);
xor  g2720 (n2768, n2651, n2637, n2661, n2669);
and  g2721 (n2755, n2715, n2653, n2659, n2680);
or   g2722 (n2766, n2672, n2695, n2644, n2497);
xor  g2723 (n2756, n2704, n2733, n2708, n2724);
and  g2724 (n2759, n2686, n2688, n2711, n2727);
nand g2725 (n2771, n2676, n2641, n2645, n2698);
xor  g2726 (n2746, n2713, n2646, n2626, n2679);
or   g2727 (n2760, n2714, n2716, n2689, n2734);
nand g2728 (n2753, n2692, n2732, n2712, n2710);
nand g2729 (n2770, n2701, n2498, n2643, n2684);
xor  g2730 (n2747, n2683, n2674, n2728, n2634);
or   g2731 (n2752, n2658, n2631, n2736, n2666);
xnor g2732 (n2763, n2670, n2630, n2622, n2735);
xor  g2733 (n2751, n2740, n2642, n2647, n2635);
nor  g2734 (n2749, n2655, n2678, n2729, n2439);
nand g2735 (n2741, n2738, n2731, n2694, n2633);
and  g2736 (n2764, n2401, n2650, n2624, n2700);
xor  g2737 (n2774, n2730, n2639, n2690, n2628);
nor  g2738 (n2773, n2440, n106, n2739, n2691);
and  g2739 (n2767, n2497, n2681, n2677, n2703);
xor  g2740 (n2765, n2717, n2740, n2401, n2663);
xor  g2741 (n2754, n2496, n2707, n2654, n2660);
xor  g2742 (n2757, n2682, n2687, n2671, n2664);
or   g2743 (n2745, n2497, n2699, n2702, n2640);
or   g2744 (n2762, n2719, n2705, n2720, n2721);
xor  g2745 (n2758, n2440, n2668, n2638, n2625);
xnor g2746 (n2769, n2709, n2685, n2636, n2629);
and  g2747 (n2772, n2693, n2667, n2718, n2498);
or   g2748 (n2750, n2652, n2498, n106);
endmodule
