

module Stat_1000_105
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n518,
  n382,
  n542,
  n459,
  n399,
  n425,
  n435,
  n390,
  n407,
  n445,
  n383,
  n362,
  n487,
  n553,
  n426,
  n403,
  n917,
  n915,
  n1022,
  n1019,
  n1023,
  n1030,
  n1024,
  n1028,
  n1032,
  n1025,
  n1020,
  n1031,
  n1021,
  n1027,
  n1026,
  n1029,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n518;
  output n382;
  output n542;
  output n459;
  output n399;
  output n425;
  output n435;
  output n390;
  output n407;
  output n445;
  output n383;
  output n362;
  output n487;
  output n553;
  output n426;
  output n403;
  output n917;
  output n915;
  output n1022;
  output n1019;
  output n1023;
  output n1030;
  output n1024;
  output n1028;
  output n1032;
  output n1025;
  output n1020;
  output n1031;
  output n1021;
  output n1027;
  output n1026;
  output n1029;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n400;
  wire n401;
  wire n402;
  wire n404;
  wire n405;
  wire n406;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n916;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n63,
    n1
  );


  buf
  g1
  (
    n50,
    n11
  );


  buf
  g2
  (
    n43,
    n10
  );


  buf
  g3
  (
    n105,
    n20
  );


  not
  g4
  (
    n70,
    n18
  );


  not
  g5
  (
    KeyWire_0_23,
    n10
  );


  not
  g6
  (
    n44,
    n19
  );


  not
  g7
  (
    n109,
    n7
  );


  not
  g8
  (
    KeyWire_0_40,
    n15
  );


  buf
  g9
  (
    n71,
    n8
  );


  buf
  g10
  (
    n79,
    n13
  );


  buf
  g11
  (
    n60,
    n19
  );


  not
  g12
  (
    n95,
    n13
  );


  buf
  g13
  (
    n83,
    n3
  );


  not
  g14
  (
    n34,
    n5
  );


  not
  g15
  (
    KeyWire_0_24,
    n12
  );


  buf
  g16
  (
    n38,
    n18
  );


  buf
  g17
  (
    n67,
    n14
  );


  not
  g18
  (
    KeyWire_0_2,
    n15
  );


  not
  g19
  (
    n81,
    n15
  );


  not
  g20
  (
    n47,
    n16
  );


  not
  g21
  (
    n96,
    n19
  );


  not
  g22
  (
    n94,
    n6
  );


  not
  g23
  (
    n80,
    n18
  );


  buf
  g24
  (
    n39,
    n4
  );


  not
  g25
  (
    n84,
    n5
  );


  buf
  g26
  (
    n59,
    n5
  );


  not
  g27
  (
    n89,
    n8
  );


  buf
  g28
  (
    n88,
    n5
  );


  buf
  g29
  (
    n75,
    n6
  );


  buf
  g30
  (
    n46,
    n21
  );


  not
  g31
  (
    n49,
    n11
  );


  not
  g32
  (
    KeyWire_0_34,
    n4
  );


  buf
  g33
  (
    n92,
    n6
  );


  not
  g34
  (
    KeyWire_0_37,
    n7
  );


  buf
  g35
  (
    n48,
    n9
  );


  not
  g36
  (
    n85,
    n15
  );


  buf
  g37
  (
    n55,
    n13
  );


  not
  g38
  (
    n104,
    n10
  );


  buf
  g39
  (
    n86,
    n17
  );


  not
  g40
  (
    n52,
    n17
  );


  not
  g41
  (
    n82,
    n14
  );


  not
  g42
  (
    n114,
    n10
  );


  buf
  g43
  (
    n53,
    n14
  );


  buf
  g44
  (
    n97,
    n16
  );


  not
  g45
  (
    n57,
    n8
  );


  not
  g46
  (
    n111,
    n17
  );


  not
  g47
  (
    n91,
    n9
  );


  buf
  g48
  (
    n77,
    n20
  );


  buf
  g49
  (
    n69,
    n11
  );


  buf
  g50
  (
    n68,
    n7
  );


  not
  g51
  (
    n99,
    n9
  );


  buf
  g52
  (
    n90,
    n11
  );


  not
  g53
  (
    n73,
    n21
  );


  not
  g54
  (
    n33,
    n12
  );


  not
  g55
  (
    n36,
    n3
  );


  buf
  g56
  (
    n72,
    n3
  );


  not
  g57
  (
    n101,
    n2
  );


  not
  g58
  (
    n45,
    n14
  );


  buf
  g59
  (
    n40,
    n16
  );


  not
  g60
  (
    n58,
    n19
  );


  not
  g61
  (
    n51,
    n6
  );


  buf
  g62
  (
    n42,
    n12
  );


  buf
  g63
  (
    n108,
    n4
  );


  not
  g64
  (
    n41,
    n1
  );


  not
  g65
  (
    n54,
    n7
  );


  buf
  g66
  (
    n78,
    n2
  );


  not
  g67
  (
    n100,
    n13
  );


  buf
  g68
  (
    n102,
    n9
  );


  not
  g69
  (
    n103,
    n8
  );


  not
  g70
  (
    n66,
    n18
  );


  not
  g71
  (
    n93,
    n17
  );


  buf
  g72
  (
    n76,
    n20
  );


  not
  g73
  (
    n37,
    n2
  );


  not
  g74
  (
    n56,
    n3
  );


  buf
  g75
  (
    n87,
    n16
  );


  buf
  g76
  (
    n61,
    n20
  );


  not
  g77
  (
    n64,
    n1
  );


  not
  g78
  (
    n106,
    n1
  );


  not
  g79
  (
    n74,
    n12
  );


  buf
  g80
  (
    n98,
    n4
  );


  buf
  g81
  (
    n62,
    n2
  );


  not
  g82
  (
    KeyWire_0_39,
    n62
  );


  not
  g83
  (
    n312,
    n90
  );


  not
  g84
  (
    n245,
    n83
  );


  not
  g85
  (
    n220,
    n48
  );


  buf
  g86
  (
    n134,
    n88
  );


  not
  g87
  (
    n284,
    n45
  );


  not
  g88
  (
    n208,
    n40
  );


  not
  g89
  (
    n353,
    n58
  );


  buf
  g90
  (
    n299,
    n72
  );


  not
  g91
  (
    n189,
    n51
  );


  not
  g92
  (
    n146,
    n60
  );


  buf
  g93
  (
    n230,
    n92
  );


  not
  g94
  (
    n244,
    n44
  );


  not
  g95
  (
    n117,
    n37
  );


  not
  g96
  (
    n168,
    n61
  );


  buf
  g97
  (
    n211,
    n50
  );


  not
  g98
  (
    n276,
    n36
  );


  not
  g99
  (
    n138,
    n40
  );


  not
  g100
  (
    n232,
    n37
  );


  not
  g101
  (
    n300,
    n49
  );


  not
  g102
  (
    n221,
    n39
  );


  buf
  g103
  (
    KeyWire_0_28,
    n38
  );


  not
  g104
  (
    n185,
    n75
  );


  buf
  g105
  (
    n354,
    n93
  );


  not
  g106
  (
    n147,
    n66
  );


  buf
  g107
  (
    n273,
    n44
  );


  not
  g108
  (
    n202,
    n53
  );


  buf
  g109
  (
    n278,
    n45
  );


  buf
  g110
  (
    n125,
    n62
  );


  not
  g111
  (
    n324,
    n68
  );


  buf
  g112
  (
    n256,
    n68
  );


  buf
  g113
  (
    n348,
    n76
  );


  not
  g114
  (
    n148,
    n49
  );


  not
  g115
  (
    n281,
    n47
  );


  buf
  g116
  (
    n274,
    n35
  );


  buf
  g117
  (
    n163,
    n82
  );


  buf
  g118
  (
    n293,
    n45
  );


  not
  g119
  (
    n340,
    n83
  );


  not
  g120
  (
    n235,
    n66
  );


  buf
  g121
  (
    KeyWire_0_36,
    n37
  );


  buf
  g122
  (
    n155,
    n56
  );


  buf
  g123
  (
    n135,
    n90
  );


  buf
  g124
  (
    n257,
    n72
  );


  not
  g125
  (
    n305,
    n53
  );


  buf
  g126
  (
    n292,
    n85
  );


  buf
  g127
  (
    n227,
    n49
  );


  not
  g128
  (
    n175,
    n60
  );


  not
  g129
  (
    n171,
    n66
  );


  buf
  g130
  (
    n314,
    n86
  );


  not
  g131
  (
    n250,
    n42
  );


  buf
  g132
  (
    n166,
    n86
  );


  not
  g133
  (
    n344,
    n75
  );


  not
  g134
  (
    n150,
    n55
  );


  not
  g135
  (
    n294,
    n94
  );


  not
  g136
  (
    n204,
    n88
  );


  not
  g137
  (
    n201,
    n65
  );


  not
  g138
  (
    n288,
    n93
  );


  not
  g139
  (
    n167,
    n52
  );


  buf
  g140
  (
    n270,
    n77
  );


  buf
  g141
  (
    n228,
    n67
  );


  not
  g142
  (
    n269,
    n61
  );


  not
  g143
  (
    n341,
    n82
  );


  buf
  g144
  (
    n213,
    n79
  );


  buf
  g145
  (
    n283,
    n63
  );


  buf
  g146
  (
    n309,
    n89
  );


  buf
  g147
  (
    n291,
    n52
  );


  buf
  g148
  (
    n161,
    n69
  );


  not
  g149
  (
    n355,
    n93
  );


  not
  g150
  (
    KeyWire_0_16,
    n41
  );


  buf
  g151
  (
    n303,
    n34
  );


  not
  g152
  (
    n311,
    n68
  );


  not
  g153
  (
    n209,
    n60
  );


  buf
  g154
  (
    n219,
    n59
  );


  not
  g155
  (
    n304,
    n86
  );


  buf
  g156
  (
    n237,
    n88
  );


  not
  g157
  (
    n131,
    n36
  );


  not
  g158
  (
    n316,
    n72
  );


  buf
  g159
  (
    n308,
    n41
  );


  not
  g160
  (
    n216,
    n47
  );


  buf
  g161
  (
    n328,
    n89
  );


  buf
  g162
  (
    n258,
    n84
  );


  not
  g163
  (
    n319,
    n42
  );


  not
  g164
  (
    n289,
    n67
  );


  buf
  g165
  (
    n122,
    n74
  );


  not
  g166
  (
    n149,
    n39
  );


  not
  g167
  (
    n129,
    n63
  );


  buf
  g168
  (
    n287,
    n44
  );


  not
  g169
  (
    n279,
    n74
  );


  not
  g170
  (
    n121,
    n51
  );


  not
  g171
  (
    n246,
    n43
  );


  not
  g172
  (
    n141,
    n54
  );


  not
  g173
  (
    n295,
    n38
  );


  not
  g174
  (
    n140,
    n94
  );


  not
  g175
  (
    n158,
    n74
  );


  buf
  g176
  (
    n322,
    n34
  );


  not
  g177
  (
    n180,
    n56
  );


  buf
  g178
  (
    n210,
    n85
  );


  not
  g179
  (
    n315,
    n63
  );


  not
  g180
  (
    n212,
    n90
  );


  not
  g181
  (
    n162,
    n56
  );


  not
  g182
  (
    n137,
    n48
  );


  not
  g183
  (
    n261,
    n73
  );


  buf
  g184
  (
    n152,
    n78
  );


  not
  g185
  (
    n238,
    n39
  );


  buf
  g186
  (
    KeyWire_0_53,
    n91
  );


  not
  g187
  (
    n133,
    n47
  );


  buf
  g188
  (
    n164,
    n77
  );


  not
  g189
  (
    n192,
    n65
  );


  buf
  g190
  (
    n351,
    n77
  );


  buf
  g191
  (
    n318,
    n70
  );


  buf
  g192
  (
    n115,
    n61
  );


  not
  g193
  (
    n145,
    n79
  );


  buf
  g194
  (
    n203,
    n75
  );


  not
  g195
  (
    n259,
    n81
  );


  not
  g196
  (
    n242,
    n90
  );


  not
  g197
  (
    n290,
    n86
  );


  not
  g198
  (
    n345,
    n70
  );


  not
  g199
  (
    n241,
    n36
  );


  not
  g200
  (
    n251,
    n53
  );


  buf
  g201
  (
    n225,
    n59
  );


  buf
  g202
  (
    n275,
    n54
  );


  buf
  g203
  (
    n332,
    n76
  );


  buf
  g204
  (
    n126,
    n48
  );


  buf
  g205
  (
    n352,
    n58
  );


  buf
  g206
  (
    n123,
    n91
  );


  not
  g207
  (
    n174,
    n50
  );


  not
  g208
  (
    n195,
    n63
  );


  not
  g209
  (
    n179,
    n80
  );


  not
  g210
  (
    n249,
    n69
  );


  not
  g211
  (
    n338,
    n71
  );


  buf
  g212
  (
    n160,
    n42
  );


  not
  g213
  (
    n306,
    n38
  );


  buf
  g214
  (
    n247,
    n60
  );


  buf
  g215
  (
    n262,
    n64
  );


  buf
  g216
  (
    n196,
    n48
  );


  not
  g217
  (
    n254,
    n67
  );


  buf
  g218
  (
    n159,
    n33
  );


  not
  g219
  (
    n265,
    n84
  );


  buf
  g220
  (
    n243,
    n46
  );


  not
  g221
  (
    n165,
    n55
  );


  not
  g222
  (
    n329,
    n91
  );


  buf
  g223
  (
    n142,
    n53
  );


  buf
  g224
  (
    n178,
    n64
  );


  buf
  g225
  (
    n120,
    n62
  );


  buf
  g226
  (
    n337,
    n92
  );


  not
  g227
  (
    KeyWire_0_19,
    n35
  );


  buf
  g228
  (
    n184,
    n73
  );


  not
  g229
  (
    n233,
    n37
  );


  buf
  g230
  (
    n151,
    n85
  );


  not
  g231
  (
    n218,
    n43
  );


  not
  g232
  (
    n214,
    n66
  );


  buf
  g233
  (
    n325,
    n83
  );


  not
  g234
  (
    n177,
    n92
  );


  not
  g235
  (
    n143,
    n87
  );


  not
  g236
  (
    n130,
    n57
  );


  not
  g237
  (
    n224,
    n43
  );


  buf
  g238
  (
    n191,
    n80
  );


  not
  g239
  (
    n154,
    n58
  );


  buf
  g240
  (
    n116,
    n80
  );


  not
  g241
  (
    n286,
    n71
  );


  not
  g242
  (
    KeyWire_0_62,
    n87
  );


  buf
  g243
  (
    n200,
    n35
  );


  buf
  g244
  (
    n326,
    n73
  );


  not
  g245
  (
    n268,
    n57
  );


  buf
  g246
  (
    KeyWire_0_60,
    n41
  );


  buf
  g247
  (
    n124,
    n59
  );


  not
  g248
  (
    n298,
    n42
  );


  buf
  g249
  (
    n334,
    n65
  );


  not
  g250
  (
    n183,
    n88
  );


  not
  g251
  (
    n190,
    n81
  );


  buf
  g252
  (
    n248,
    n71
  );


  buf
  g253
  (
    n206,
    n46
  );


  buf
  g254
  (
    n207,
    n71
  );


  not
  g255
  (
    n347,
    n39
  );


  buf
  g256
  (
    n217,
    n50
  );


  buf
  g257
  (
    n157,
    n33
  );


  not
  g258
  (
    n277,
    n73
  );


  not
  g259
  (
    n313,
    n81
  );


  buf
  g260
  (
    KeyWire_0_32,
    n52
  );


  not
  g261
  (
    KeyWire_0_54,
    n55
  );


  not
  g262
  (
    n139,
    n79
  );


  buf
  g263
  (
    KeyWire_0_50,
    n34
  );


  not
  g264
  (
    n282,
    n94
  );


  not
  g265
  (
    n188,
    n82
  );


  not
  g266
  (
    n172,
    n46
  );


  not
  g267
  (
    n343,
    n78
  );


  buf
  g268
  (
    n310,
    n70
  );


  buf
  g269
  (
    n222,
    n61
  );


  buf
  g270
  (
    n255,
    n82
  );


  not
  g271
  (
    n331,
    n35
  );


  buf
  g272
  (
    n156,
    n94
  );


  not
  g273
  (
    n285,
    n87
  );


  buf
  g274
  (
    n170,
    n89
  );


  buf
  g275
  (
    n327,
    n38
  );


  not
  g276
  (
    n128,
    n75
  );


  buf
  g277
  (
    n223,
    n62
  );


  not
  g278
  (
    n229,
    n77
  );


  not
  g279
  (
    n119,
    n43
  );


  buf
  g280
  (
    n215,
    n50
  );


  buf
  g281
  (
    KeyWire_0_30,
    n49
  );


  buf
  g282
  (
    n187,
    n74
  );


  not
  g283
  (
    n350,
    n34
  );


  not
  g284
  (
    n271,
    n84
  );


  not
  g285
  (
    n240,
    n46
  );


  buf
  g286
  (
    n323,
    n76
  );


  not
  g287
  (
    n253,
    n93
  );


  buf
  g288
  (
    n349,
    n64
  );


  buf
  g289
  (
    n176,
    n36
  );


  not
  g290
  (
    KeyWire_0_25,
    n41
  );


  not
  g291
  (
    n301,
    n68
  );


  not
  g292
  (
    n205,
    n64
  );


  not
  g293
  (
    n267,
    n52
  );


  not
  g294
  (
    n321,
    n33
  );


  not
  g295
  (
    n280,
    n54
  );


  not
  g296
  (
    n297,
    n56
  );


  not
  g297
  (
    n186,
    n69
  );


  buf
  g298
  (
    n336,
    n80
  );


  buf
  g299
  (
    n136,
    n92
  );


  not
  g300
  (
    n335,
    n51
  );


  buf
  g301
  (
    n194,
    n65
  );


  not
  g302
  (
    n197,
    n47
  );


  buf
  g303
  (
    n198,
    n70
  );


  buf
  g304
  (
    n173,
    n76
  );


  not
  g305
  (
    n302,
    n55
  );


  not
  g306
  (
    n193,
    n78
  );


  not
  g307
  (
    n144,
    n58
  );


  not
  g308
  (
    n234,
    n44
  );


  buf
  g309
  (
    n252,
    n40
  );


  buf
  g310
  (
    n317,
    n51
  );


  buf
  g311
  (
    n330,
    n69
  );


  buf
  g312
  (
    n199,
    n91
  );


  not
  g313
  (
    n182,
    n78
  );


  buf
  g314
  (
    n260,
    n40
  );


  buf
  g315
  (
    n356,
    n67
  );


  buf
  g316
  (
    n320,
    n87
  );


  buf
  g317
  (
    n342,
    n84
  );


  buf
  g318
  (
    n153,
    n54
  );


  not
  g319
  (
    n339,
    n72
  );


  not
  g320
  (
    n239,
    n95
  );


  nand
  g321
  (
    n263,
    n81,
    n79
  );


  and
  g322
  (
    n236,
    n57,
    n83,
    n45,
    n85
  );


  xnor
  g323
  (
    n307,
    n33,
    n89,
    n59,
    n57
  );


  or
  g324
  (
    n397,
    n213,
    n137,
    n305,
    n248
  );


  and
  g325
  (
    n360,
    n272,
    n231,
    n227,
    n151
  );


  nor
  g326
  (
    n419,
    n133,
    n165,
    n317,
    n163
  );


  nand
  g327
  (
    n505,
    n147,
    n301,
    n180,
    n313
  );


  or
  g328
  (
    n441,
    n212,
    n163,
    n215,
    n198
  );


  and
  g329
  (
    n506,
    n196,
    n237,
    n174,
    n173
  );


  nor
  g330
  (
    n547,
    n224,
    n232,
    n193,
    n168
  );


  nand
  g331
  (
    KeyWire_0_47,
    n195,
    n219,
    n137,
    n259
  );


  xnor
  g332
  (
    n518,
    n220,
    n264,
    n139,
    n224
  );


  or
  g333
  (
    n434,
    n190,
    n284,
    n289,
    n279
  );


  and
  g334
  (
    n359,
    n194,
    n237,
    n135,
    n244
  );


  xnor
  g335
  (
    KeyWire_0_57,
    n313,
    n202,
    n198,
    n226
  );


  nand
  g336
  (
    n494,
    n138,
    n139,
    n301,
    n160
  );


  and
  g337
  (
    n430,
    n282,
    n164,
    n188,
    n211
  );


  or
  g338
  (
    n414,
    n209,
    n208,
    n293,
    n229
  );


  nand
  g339
  (
    n386,
    n208,
    n300,
    n232,
    n296
  );


  xnor
  g340
  (
    n501,
    n201,
    n268,
    n159,
    n175
  );


  nand
  g341
  (
    n527,
    n217,
    n125,
    n199,
    n184
  );


  xor
  g342
  (
    n504,
    n274,
    n305,
    n284,
    n291
  );


  nand
  g343
  (
    n377,
    n241,
    n292,
    n255,
    n141
  );


  xor
  g344
  (
    n517,
    n287,
    n157,
    n145,
    n308
  );


  and
  g345
  (
    n471,
    n320,
    n264,
    n207,
    n314
  );


  or
  g346
  (
    n451,
    n237,
    n249,
    n159,
    n162
  );


  nand
  g347
  (
    n442,
    n303,
    n199,
    n157,
    n178
  );


  xnor
  g348
  (
    n523,
    n228,
    n214,
    n136,
    n300
  );


  xor
  g349
  (
    n492,
    n183,
    n154,
    n287,
    n115
  );


  nand
  g350
  (
    n387,
    n131,
    n251,
    n268,
    n219
  );


  xnor
  g351
  (
    n555,
    n168,
    n133,
    n259,
    n295
  );


  and
  g352
  (
    KeyWire_0_33,
    n158,
    n191,
    n314,
    n186
  );


  xor
  g353
  (
    n393,
    n179,
    n141,
    n310,
    n166
  );


  or
  g354
  (
    n440,
    n149,
    n215,
    n218,
    n221
  );


  nand
  g355
  (
    n454,
    n191,
    n162,
    n278,
    n159
  );


  xnor
  g356
  (
    n367,
    n195,
    n148,
    n228,
    n185
  );


  xnor
  g357
  (
    n533,
    n265,
    n263,
    n233,
    n246
  );


  nand
  g358
  (
    n467,
    n204,
    n309,
    n130,
    n301
  );


  xnor
  g359
  (
    n540,
    n221,
    n254,
    n175,
    n281
  );


  nand
  g360
  (
    n511,
    n283,
    n171,
    n162,
    n252
  );


  and
  g361
  (
    n398,
    n253,
    n186,
    n286,
    n257
  );


  nor
  g362
  (
    n390,
    n284,
    n188,
    n219,
    n250
  );


  or
  g363
  (
    n401,
    n127,
    n304,
    n143,
    n243
  );


  xor
  g364
  (
    n381,
    n149,
    n160,
    n144,
    n261
  );


  nor
  g365
  (
    n427,
    n194,
    n223,
    n163,
    n191
  );


  or
  g366
  (
    n514,
    n296,
    n258,
    n138,
    n247
  );


  nand
  g367
  (
    n509,
    n272,
    n258,
    n318,
    n224
  );


  nand
  g368
  (
    n510,
    n178,
    n307,
    n214,
    n204
  );


  and
  g369
  (
    n546,
    n156,
    n203,
    n245,
    n239
  );


  xnor
  g370
  (
    n415,
    n274,
    n178,
    n194,
    n279
  );


  xor
  g371
  (
    n469,
    n149,
    n312,
    n217,
    n235
  );


  xor
  g372
  (
    n529,
    n253,
    n316,
    n269,
    n281
  );


  nor
  g373
  (
    n416,
    n221,
    n147,
    n297,
    n293
  );


  or
  g374
  (
    KeyWire_0_29,
    n262,
    n130,
    n267,
    n192
  );


  nand
  g375
  (
    n538,
    n183,
    n260,
    n294,
    n118
  );


  xor
  g376
  (
    n537,
    n267,
    n176,
    n315,
    n233
  );


  xor
  g377
  (
    n425,
    n261,
    n212,
    n216,
    n161
  );


  and
  g378
  (
    KeyWire_0_41,
    n311,
    n249,
    n209,
    n164
  );


  xor
  g379
  (
    n443,
    n292,
    n250,
    n147,
    n311
  );


  and
  g380
  (
    n524,
    n256,
    n140,
    n224,
    n226
  );


  or
  g381
  (
    n502,
    n128,
    n320,
    n206,
    n171
  );


  and
  g382
  (
    KeyWire_0_6,
    n117,
    n275,
    n201,
    n161
  );


  nor
  g383
  (
    n431,
    n315,
    n304,
    n167,
    n264
  );


  xor
  g384
  (
    n358,
    n300,
    n185,
    n126,
    n306
  );


  nand
  g385
  (
    n519,
    n226,
    n289,
    n190,
    n189
  );


  and
  g386
  (
    n531,
    n251,
    n273,
    n218,
    n208
  );


  or
  g387
  (
    n495,
    n173,
    n127,
    n144,
    n235
  );


  nand
  g388
  (
    n521,
    n275,
    n299,
    n242,
    n123
  );


  or
  g389
  (
    n460,
    n261,
    n264,
    n212,
    n294
  );


  xor
  g390
  (
    n410,
    n197,
    n195,
    n296,
    n265
  );


  xor
  g391
  (
    n497,
    n145,
    n305,
    n126,
    n221
  );


  and
  g392
  (
    n468,
    n129,
    n267,
    n225,
    n287
  );


  xor
  g393
  (
    n421,
    n306,
    n182,
    n127,
    n277
  );


  xnor
  g394
  (
    n449,
    n293,
    n161,
    n309,
    n240
  );


  xnor
  g395
  (
    n473,
    n176,
    n172,
    n120,
    n255
  );


  xnor
  g396
  (
    n369,
    n171,
    n183,
    n204,
    n124
  );


  and
  g397
  (
    n459,
    n306,
    n148,
    n193,
    n200
  );


  or
  g398
  (
    n428,
    n177,
    n174,
    n181,
    n286
  );


  nand
  g399
  (
    n450,
    n239,
    n266,
    n136,
    n257
  );


  xnor
  g400
  (
    n404,
    n231,
    n164,
    n292,
    n163
  );


  nand
  g401
  (
    n389,
    n236,
    n230,
    n176,
    n273
  );


  xor
  g402
  (
    n462,
    n123,
    n271,
    n243,
    n155
  );


  xor
  g403
  (
    n516,
    n238,
    n188,
    n260,
    n120
  );


  nand
  g404
  (
    n361,
    n253,
    n148,
    n230,
    n220
  );


  or
  g405
  (
    n500,
    n190,
    n172,
    n151,
    n316
  );


  nand
  g406
  (
    n370,
    n146,
    n238,
    n244,
    n302
  );


  xor
  g407
  (
    n423,
    n251,
    n254,
    n185,
    n261
  );


  nand
  g408
  (
    n508,
    n227,
    n231,
    n137,
    n271
  );


  or
  g409
  (
    n545,
    n247,
    n263,
    n206,
    n205
  );


  nand
  g410
  (
    n422,
    n281,
    n270,
    n218,
    n257
  );


  nor
  g411
  (
    n452,
    n246,
    n270,
    n303,
    n248
  );


  nand
  g412
  (
    n405,
    n288,
    n284,
    n238,
    n234
  );


  xor
  g413
  (
    n528,
    n279,
    n216,
    n241,
    n135
  );


  xnor
  g414
  (
    n493,
    n202,
    n310,
    n134,
    n203
  );


  nand
  g415
  (
    n382,
    n289,
    n267,
    n247,
    n311
  );


  xnor
  g416
  (
    n526,
    n280,
    n256,
    n207,
    n158
  );


  xnor
  g417
  (
    KeyWire_0_44,
    n303,
    n211,
    n229,
    n225
  );


  and
  g418
  (
    n472,
    n242,
    n190,
    n157,
    n238
  );


  and
  g419
  (
    n543,
    n318,
    n150,
    n302,
    n256
  );


  and
  g420
  (
    n515,
    n154,
    n281,
    n260,
    n191
  );


  xor
  g421
  (
    KeyWire_0_20,
    n150,
    n129,
    n298,
    n179
  );


  xnor
  g422
  (
    n384,
    n246,
    n239,
    n198,
    n236
  );


  or
  g423
  (
    n498,
    n148,
    n288,
    n184,
    n205
  );


  and
  g424
  (
    n365,
    n182,
    n226,
    n280,
    n275
  );


  xor
  g425
  (
    n550,
    n188,
    n175,
    n210,
    n259
  );


  nand
  g426
  (
    n433,
    n130,
    n162,
    n248,
    n202
  );


  xor
  g427
  (
    n484,
    n176,
    n174,
    n132,
    n156
  );


  xnor
  g428
  (
    n513,
    n259,
    n244,
    n166,
    n199
  );


  xnor
  g429
  (
    n407,
    n311,
    n151,
    n132,
    n203
  );


  xnor
  g430
  (
    n392,
    n201,
    n192,
    n256,
    n207
  );


  nor
  g431
  (
    n503,
    n193,
    n297,
    n302,
    n116
  );


  xor
  g432
  (
    n388,
    n195,
    n287,
    n266,
    n225
  );


  and
  g433
  (
    n378,
    n179,
    n199,
    n169,
    n309
  );


  nor
  g434
  (
    n463,
    n159,
    n143,
    n152,
    n296
  );


  xor
  g435
  (
    n432,
    n135,
    n160,
    n133,
    n245
  );


  xor
  g436
  (
    n489,
    n167,
    n140,
    n293,
    n228
  );


  nand
  g437
  (
    n487,
    n134,
    n128,
    n197,
    n304
  );


  xor
  g438
  (
    n525,
    n157,
    n155,
    n222,
    n170
  );


  xnor
  g439
  (
    n448,
    n165,
    n169,
    n290,
    n317
  );


  xor
  g440
  (
    n399,
    n234,
    n185,
    n166,
    n319
  );


  nor
  g441
  (
    n379,
    n142,
    n265,
    n282,
    n290
  );


  nand
  g442
  (
    n554,
    n135,
    n285,
    n160,
    n312
  );


  xor
  g443
  (
    n458,
    n131,
    n297,
    n254,
    n242
  );


  xor
  g444
  (
    n411,
    n290,
    n230,
    n181,
    n215
  );


  xnor
  g445
  (
    n391,
    n172,
    n275,
    n165,
    n164
  );


  xnor
  g446
  (
    n486,
    n121,
    n314,
    n235,
    n260
  );


  xor
  g447
  (
    n402,
    n245,
    n262,
    n292,
    n145
  );


  or
  g448
  (
    n542,
    n187,
    n181,
    n299,
    n205
  );


  nor
  g449
  (
    n474,
    n270,
    n258,
    n288,
    n172
  );


  xnor
  g450
  (
    n453,
    n282,
    n298,
    n269,
    n247
  );


  and
  g451
  (
    n373,
    n317,
    n147,
    n268,
    n228
  );


  nor
  g452
  (
    KeyWire_0_35,
    n215,
    n126,
    n273,
    n282
  );


  xor
  g453
  (
    n444,
    n126,
    n149,
    n173,
    n153
  );


  and
  g454
  (
    KeyWire_0_27,
    n143,
    n181,
    n271,
    n312
  );


  xnor
  g455
  (
    n374,
    n183,
    n277,
    n189,
    n216
  );


  xnor
  g456
  (
    n412,
    n309,
    n182,
    n294,
    n202
  );


  nor
  g457
  (
    n400,
    n318,
    n258,
    n180,
    n156
  );


  nor
  g458
  (
    n541,
    n187,
    n280,
    n205,
    n312
  );


  xnor
  g459
  (
    n480,
    n206,
    n142,
    n121,
    n129
  );


  nand
  g460
  (
    n465,
    n294,
    n276,
    n307,
    n150
  );


  nor
  g461
  (
    n408,
    n189,
    n252,
    n239,
    n169
  );


  xor
  g462
  (
    n520,
    n142,
    n140,
    n222,
    n223
  );


  and
  g463
  (
    n475,
    n132,
    n317,
    n129,
    n196
  );


  nand
  g464
  (
    n551,
    n319,
    n158,
    n115,
    n127
  );


  or
  g465
  (
    n534,
    n268,
    n223,
    n308,
    n177
  );


  xnor
  g466
  (
    n488,
    n222,
    n209,
    n186,
    n136
  );


  xnor
  g467
  (
    n438,
    n213,
    n285,
    n130,
    n194
  );


  nor
  g468
  (
    n417,
    n243,
    n316,
    n234,
    n170
  );


  nor
  g469
  (
    n548,
    n290,
    n316,
    n236,
    n279
  );


  or
  g470
  (
    n366,
    n241,
    n236,
    n174,
    n122
  );


  nand
  g471
  (
    n395,
    n263,
    n295,
    n125,
    n198
  );


  or
  g472
  (
    n544,
    n214,
    n201,
    n237,
    n273
  );


  and
  g473
  (
    n485,
    n168,
    n146,
    n301,
    n308
  );


  nand
  g474
  (
    n530,
    n278,
    n276,
    n227,
    n308
  );


  nor
  g475
  (
    n357,
    n182,
    n184,
    n298,
    n150
  );


  or
  g476
  (
    n457,
    n153,
    n289,
    n213,
    n138
  );


  or
  g477
  (
    n536,
    n178,
    n167,
    n291,
    n165
  );


  nor
  g478
  (
    n549,
    n142,
    n229,
    n200,
    n197
  );


  nor
  g479
  (
    n437,
    n118,
    n153,
    n291,
    n251
  );


  or
  g480
  (
    KeyWire_0_5,
    n179,
    n153,
    n154,
    n197
  );


  xnor
  g481
  (
    n418,
    n233,
    n231,
    n319,
    n134
  );


  nand
  g482
  (
    n522,
    n192,
    n288,
    n180,
    n286
  );


  nand
  g483
  (
    n380,
    n119,
    n146,
    n240,
    n277
  );


  nand
  g484
  (
    n385,
    n152,
    n269,
    n141,
    n136
  );


  nor
  g485
  (
    n464,
    n246,
    n196,
    n277,
    n243
  );


  nand
  g486
  (
    n371,
    n204,
    n128,
    n313,
    n170
  );


  xnor
  g487
  (
    n447,
    n116,
    n143,
    n156,
    n171
  );


  xor
  g488
  (
    n507,
    n210,
    n214,
    n310,
    n207
  );


  or
  g489
  (
    n439,
    n274,
    n257,
    n139,
    n161
  );


  nor
  g490
  (
    n496,
    n240,
    n170,
    n193,
    n285
  );


  xnor
  g491
  (
    n461,
    n232,
    n291,
    n285,
    n300
  );


  or
  g492
  (
    n479,
    n152,
    n184,
    n269,
    n212
  );


  xnor
  g493
  (
    n409,
    n280,
    n304,
    n154,
    n177
  );


  nor
  g494
  (
    n406,
    n245,
    n283,
    n265,
    n252
  );


  xor
  g495
  (
    n477,
    n145,
    n196,
    n255,
    n319
  );


  xnor
  g496
  (
    KeyWire_0_10,
    n248,
    n298,
    n235,
    n295
  );


  xnor
  g497
  (
    n535,
    n305,
    n180,
    n225,
    n217
  );


  or
  g498
  (
    n499,
    n169,
    n262,
    n263,
    n166
  );


  xor
  g499
  (
    n426,
    n250,
    n167,
    n271,
    n315
  );


  xor
  g500
  (
    n375,
    n187,
    n152,
    n217,
    n318
  );


  xor
  g501
  (
    n436,
    n302,
    n177,
    n299,
    n283
  );


  xor
  g502
  (
    n372,
    n262,
    n131,
    n144,
    n133
  );


  nor
  g503
  (
    n363,
    n232,
    n266,
    n134,
    n155
  );


  or
  g504
  (
    n456,
    n227,
    n229,
    n295,
    n315
  );


  and
  g505
  (
    n455,
    n233,
    n140,
    n203,
    n230
  );


  nor
  g506
  (
    n413,
    n208,
    n216,
    n146,
    n234
  );


  nor
  g507
  (
    n394,
    n187,
    n220,
    n117,
    n306
  );


  or
  g508
  (
    n478,
    n283,
    n137,
    n173,
    n254
  );


  or
  g509
  (
    n403,
    n250,
    n192,
    n278,
    n122
  );


  and
  g510
  (
    n466,
    n297,
    n314,
    n244,
    n249
  );


  xor
  g511
  (
    n446,
    n223,
    n252,
    n274,
    n151
  );


  xor
  g512
  (
    n481,
    n313,
    n286,
    n303,
    n200
  );


  and
  g513
  (
    n445,
    n128,
    n200,
    n242,
    n276
  );


  nand
  g514
  (
    n476,
    n131,
    n144,
    n218,
    n138
  );


  xor
  g515
  (
    n424,
    n158,
    n272,
    n307,
    n141
  );


  and
  g516
  (
    n429,
    n220,
    n175,
    n206,
    n189
  );


  and
  g517
  (
    n368,
    n278,
    n210,
    n186,
    n240
  );


  xnor
  g518
  (
    n553,
    n209,
    n213,
    n310,
    n249
  );


  xnor
  g519
  (
    n383,
    n119,
    n241,
    n139,
    n211
  );


  nand
  g520
  (
    n491,
    n255,
    n270,
    n210,
    n299
  );


  xor
  g521
  (
    n532,
    n124,
    n132,
    n222,
    n272
  );


  and
  g522
  (
    n482,
    n168,
    n211,
    n219,
    n155
  );


  nand
  g523
  (
    n556,
    n307,
    n276,
    n266,
    n253
  );


  or
  g524
  (
    n620,
    n457,
    n547,
    n371,
    n29
  );


  nand
  g525
  (
    n648,
    n520,
    n540,
    n449,
    n337
  );


  xnor
  g526
  (
    n756,
    n443,
    n348,
    n415,
    n416
  );


  xor
  g527
  (
    n608,
    n326,
    n438,
    n423,
    n502
  );


  xor
  g528
  (
    n565,
    n497,
    n488,
    n462,
    n518
  );


  nor
  g529
  (
    n715,
    n334,
    n468,
    n439,
    n329
  );


  xnor
  g530
  (
    n662,
    n367,
    n517,
    n321,
    n432
  );


  and
  g531
  (
    n577,
    n329,
    n498,
    n371,
    n433
  );


  and
  g532
  (
    n622,
    n400,
    n364,
    n22,
    n424
  );


  or
  g533
  (
    n694,
    n387,
    n449,
    n473,
    n339
  );


  and
  g534
  (
    n769,
    n543,
    n434,
    n437,
    n499
  );


  and
  g535
  (
    n579,
    n472,
    n369,
    n389,
    n476
  );


  or
  g536
  (
    n619,
    n26,
    n385,
    n544,
    n333
  );


  nand
  g537
  (
    n617,
    n553,
    n471,
    n425,
    n331
  );


  xnor
  g538
  (
    n661,
    n328,
    n467,
    n505
  );


  xnor
  g539
  (
    n765,
    n459,
    n456,
    n523,
    n439
  );


  nor
  g540
  (
    n712,
    n546,
    n548,
    n516,
    n531
  );


  nand
  g541
  (
    KeyWire_0_9,
    n531,
    n334,
    n365,
    n28
  );


  or
  g542
  (
    n768,
    n450,
    n468,
    n401,
    n540
  );


  nor
  g543
  (
    n777,
    n343,
    n403,
    n395,
    n459
  );


  and
  g544
  (
    n735,
    n482,
    n403,
    n343,
    n523
  );


  and
  g545
  (
    n586,
    n542,
    n427,
    n446,
    n526
  );


  or
  g546
  (
    n611,
    n101,
    n473,
    n407,
    n511
  );


  nor
  g547
  (
    n754,
    n410,
    n479,
    n495,
    n430
  );


  xor
  g548
  (
    n666,
    n447,
    n552,
    n99,
    n453
  );


  and
  g549
  (
    n567,
    n346,
    n472,
    n426,
    n386
  );


  nand
  g550
  (
    n750,
    n437,
    n491,
    n492,
    n400
  );


  nand
  g551
  (
    n651,
    n471,
    n530,
    n439
  );


  xnor
  g552
  (
    n612,
    n370,
    n544,
    n502,
    n500
  );


  and
  g553
  (
    n560,
    n407,
    n330,
    n446,
    n99
  );


  nor
  g554
  (
    n582,
    n536,
    n419,
    n511,
    n490
  );


  and
  g555
  (
    n701,
    n541,
    n521,
    n24,
    n554
  );


  xor
  g556
  (
    n587,
    n497,
    n493,
    n400,
    n31
  );


  and
  g557
  (
    n600,
    n518,
    n407,
    n503,
    n533
  );


  nand
  g558
  (
    n594,
    n411,
    n490,
    n369,
    n541
  );


  xor
  g559
  (
    n685,
    n469,
    n320,
    n100,
    n444
  );


  xor
  g560
  (
    n734,
    n445,
    n397,
    n327,
    n496
  );


  xnor
  g561
  (
    n656,
    n358,
    n367,
    n525,
    n451
  );


  xnor
  g562
  (
    n650,
    n553,
    n510,
    n343,
    n397
  );


  and
  g563
  (
    n705,
    n419,
    n378,
    n362,
    n390
  );


  or
  g564
  (
    n764,
    n97,
    n535,
    n100,
    n329
  );


  or
  g565
  (
    n590,
    n330,
    n329,
    n442,
    n545
  );


  nand
  g566
  (
    n606,
    n515,
    n489,
    n498,
    n516
  );


  xor
  g567
  (
    KeyWire_0_59,
    n453,
    n403,
    n537,
    n493
  );


  nor
  g568
  (
    n779,
    n411,
    n528,
    n448,
    n434
  );


  and
  g569
  (
    n647,
    n494,
    n396,
    n394,
    n552
  );


  xor
  g570
  (
    n737,
    n440,
    n537,
    n346,
    n349
  );


  xor
  g571
  (
    KeyWire_0_3,
    n489,
    n405,
    n402,
    n521
  );


  xor
  g572
  (
    n566,
    n323,
    n30,
    n455,
    n373
  );


  or
  g573
  (
    n706,
    n31,
    n401,
    n548,
    n449
  );


  and
  g574
  (
    KeyWire_0_46,
    n372,
    n400,
    n551,
    n408
  );


  xnor
  g575
  (
    n760,
    n410,
    n450,
    n527
  );


  and
  g576
  (
    n634,
    n420,
    n461,
    n440,
    n30
  );


  nand
  g577
  (
    n595,
    n96,
    n430,
    n435,
    n462
  );


  nand
  g578
  (
    n716,
    n342,
    n494,
    n395,
    n382
  );


  nand
  g579
  (
    n564,
    n414,
    n24,
    n337,
    n442
  );


  nor
  g580
  (
    KeyWire_0_43,
    n491,
    n523,
    n381,
    n412
  );


  nand
  g581
  (
    n676,
    n339,
    n388,
    n359,
    n428
  );


  nor
  g582
  (
    n641,
    n413,
    n463,
    n535,
    n29
  );


  or
  g583
  (
    n758,
    n27,
    n478,
    n96,
    n336
  );


  and
  g584
  (
    n708,
    n527,
    n465,
    n22,
    n393
  );


  or
  g585
  (
    n767,
    n494,
    n528,
    n423,
    n475
  );


  nor
  g586
  (
    n751,
    n339,
    n417,
    n404,
    n493
  );


  nor
  g587
  (
    n629,
    n433,
    n429,
    n21,
    n381
  );


  nor
  g588
  (
    n729,
    n546,
    n406,
    n460
  );


  xor
  g589
  (
    n783,
    n375,
    n399,
    n471,
    n514
  );


  and
  g590
  (
    n605,
    n408,
    n447,
    n415,
    n409
  );


  xnor
  g591
  (
    n589,
    n404,
    n483,
    n418,
    n332
  );


  and
  g592
  (
    n730,
    n459,
    n549,
    n357,
    n534
  );


  nor
  g593
  (
    n621,
    n422,
    n506,
    n366,
    n398
  );


  nor
  g594
  (
    KeyWire_0_0,
    n446,
    n425,
    n344,
    n380
  );


  and
  g595
  (
    n693,
    n463,
    n501,
    n505,
    n525
  );


  nand
  g596
  (
    n578,
    n328,
    n451,
    n396,
    n462
  );


  or
  g597
  (
    n686,
    n374,
    n435,
    n527,
    n455
  );


  or
  g598
  (
    n563,
    n516,
    n473,
    n320,
    n423
  );


  xnor
  g599
  (
    n644,
    n331,
    n538,
    n532,
    n443
  );


  xor
  g600
  (
    n725,
    n488,
    n514,
    n444,
    n501
  );


  or
  g601
  (
    n678,
    n348,
    n495,
    n508,
    n532
  );


  xnor
  g602
  (
    n721,
    n403,
    n518,
    n321,
    n501
  );


  xnor
  g603
  (
    n742,
    n422,
    n513,
    n424,
    n551
  );


  or
  g604
  (
    n616,
    n443,
    n483,
    n467,
    n493
  );


  nand
  g605
  (
    n575,
    n409,
    n456,
    n455,
    n542
  );


  xor
  g606
  (
    KeyWire_0_45,
    n321,
    n521,
    n445,
    n330
  );


  xnor
  g607
  (
    n630,
    n486,
    n518,
    n443,
    n497
  );


  nor
  g608
  (
    n749,
    n504,
    n411,
    n341,
    n398
  );


  xnor
  g609
  (
    n649,
    n431,
    n479,
    n532,
    n23
  );


  nand
  g610
  (
    n741,
    n337,
    n498,
    n531,
    n417
  );


  and
  g611
  (
    n573,
    n470,
    n340,
    n458,
    n539
  );


  or
  g612
  (
    n763,
    n368,
    n31,
    n524,
    n464
  );


  or
  g613
  (
    KeyWire_0_61,
    n499,
    n473,
    n505,
    n446
  );


  nand
  g614
  (
    KeyWire_0_22,
    n445,
    n543,
    n453,
    n402
  );


  or
  g615
  (
    n574,
    n484,
    n455,
    n447,
    n338
  );


  and
  g616
  (
    KeyWire_0_26,
    n531,
    n543,
    n469,
    n472
  );


  xnor
  g617
  (
    n632,
    n441,
    n448,
    n454,
    n341
  );


  or
  g618
  (
    n633,
    n537,
    n99,
    n440,
    n429
  );


  or
  g619
  (
    n562,
    n492,
    n466,
    n512,
    n442
  );


  xnor
  g620
  (
    n727,
    n418,
    n533,
    n492,
    n396
  );


  or
  g621
  (
    n696,
    n429,
    n401,
    n344,
    n477
  );


  and
  g622
  (
    n736,
    n536,
    n525,
    n30,
    n503
  );


  nand
  g623
  (
    n603,
    n441,
    n523,
    n549,
    n345
  );


  nand
  g624
  (
    KeyWire_0_4,
    n333,
    n515,
    n343,
    n451
  );


  xor
  g625
  (
    n709,
    n342,
    n519,
    n347,
    n529
  );


  nand
  g626
  (
    n739,
    n325,
    n421,
    n513
  );


  nor
  g627
  (
    n609,
    n376,
    n477,
    n480,
    n461
  );


  xor
  g628
  (
    n628,
    n437,
    n422,
    n485,
    n508
  );


  xor
  g629
  (
    n703,
    n97,
    n338,
    n495,
    n472
  );


  xnor
  g630
  (
    n627,
    n522,
    n420,
    n524,
    n431
  );


  nand
  g631
  (
    KeyWire_0_38,
    n508,
    n468,
    n529,
    n341
  );


  nand
  g632
  (
    n688,
    n417,
    n96,
    n509,
    n422
  );


  xnor
  g633
  (
    n680,
    n342,
    n509,
    n437,
    n541
  );


  or
  g634
  (
    n770,
    n504,
    n530,
    n525
  );


  xor
  g635
  (
    n669,
    n25,
    n402,
    n483
  );


  nor
  g636
  (
    n720,
    n474,
    n504,
    n360,
    n480
  );


  nand
  g637
  (
    n635,
    n499,
    n486,
    n325,
    n517
  );


  nand
  g638
  (
    n642,
    n477,
    n427,
    n332,
    n374
  );


  xnor
  g639
  (
    n675,
    n331,
    n390,
    n496,
    n398
  );


  and
  g640
  (
    n668,
    n373,
    n512,
    n460,
    n524
  );


  and
  g641
  (
    n569,
    n344,
    n101,
    n413,
    n428
  );


  xor
  g642
  (
    n583,
    n545,
    n550,
    n542,
    n485
  );


  xnor
  g643
  (
    n673,
    n25,
    n475,
    n532,
    n330
  );


  or
  g644
  (
    n724,
    n509,
    n378,
    n438,
    n368
  );


  xor
  g645
  (
    n719,
    n24,
    n551,
    n510,
    n102
  );


  xnor
  g646
  (
    n618,
    n456,
    n95,
    n444,
    n397
  );


  nor
  g647
  (
    n599,
    n384,
    n482,
    n545,
    n503
  );


  or
  g648
  (
    KeyWire_0_1,
    n470,
    n511,
    n29,
    n456
  );


  or
  g649
  (
    n753,
    n361,
    n526,
    n500,
    n372
  );


  xor
  g650
  (
    n652,
    n364,
    n539,
    n322,
    n418
  );


  and
  g651
  (
    n643,
    n384,
    n419,
    n334,
    n548
  );


  nor
  g652
  (
    n707,
    n462,
    n370,
    n460,
    n435
  );


  nor
  g653
  (
    n657,
    n98,
    n332,
    n336,
    n491
  );


  nand
  g654
  (
    n782,
    n481,
    n380,
    n467,
    n375
  );


  xor
  g655
  (
    n744,
    n348,
    n552,
    n410,
    n506
  );


  or
  g656
  (
    n593,
    n510,
    n449,
    n102,
    n508
  );


  or
  g657
  (
    n740,
    n331,
    n22,
    n539,
    n24
  );


  and
  g658
  (
    n674,
    n538,
    n528,
    n444,
    n428
  );


  xor
  g659
  (
    n568,
    n513,
    n522,
    n427,
    n486
  );


  or
  g660
  (
    n762,
    n545,
    n358,
    n416,
    n487
  );


  nor
  g661
  (
    n723,
    n346,
    n481,
    n338,
    n552
  );


  or
  g662
  (
    n759,
    n347,
    n460,
    n327,
    n506
  );


  or
  g663
  (
    n717,
    n379,
    n438,
    n491,
    n359
  );


  nor
  g664
  (
    n683,
    n471,
    n475,
    n534,
    n28
  );


  xnor
  g665
  (
    n679,
    n101,
    n98,
    n326,
    n379
  );


  xnor
  g666
  (
    n646,
    n447,
    n549,
    n543,
    n345
  );


  xor
  g667
  (
    n580,
    n515,
    n463,
    n334,
    n404
  );


  and
  g668
  (
    KeyWire_0_18,
    n414,
    n429,
    n326,
    n457
  );


  nand
  g669
  (
    n581,
    n31,
    n32,
    n464,
    n554
  );


  xor
  g670
  (
    n601,
    n490,
    n335,
    n533,
    n463
  );


  and
  g671
  (
    KeyWire_0_56,
    n480,
    n405,
    n487,
    n396
  );


  xor
  g672
  (
    n614,
    n324,
    n499,
    n551,
    n410
  );


  and
  g673
  (
    n772,
    n27,
    n496,
    n520,
    n454
  );


  nor
  g674
  (
    n626,
    n436,
    n328,
    n489,
    n496
  );


  and
  g675
  (
    n692,
    n480,
    n100,
    n433,
    n534
  );


  and
  g676
  (
    n761,
    n482,
    n442,
    n340,
    n452
  );


  or
  g677
  (
    n636,
    n519,
    n327,
    n476,
    n424
  );


  xor
  g678
  (
    n638,
    n478,
    n507,
    n502,
    n30
  );


  xnor
  g679
  (
    n691,
    n479,
    n448,
    n324,
    n452
  );


  xor
  g680
  (
    n597,
    n519,
    n399,
    n393,
    n395
  );


  nand
  g681
  (
    n766,
    n417,
    n528,
    n486,
    n101
  );


  nand
  g682
  (
    n745,
    n324,
    n539,
    n546,
    n412
  );


  or
  g683
  (
    n698,
    n494,
    n340,
    n500,
    n428
  );


  nand
  g684
  (
    n584,
    n519,
    n535,
    n498,
    n28
  );


  xnor
  g685
  (
    n610,
    n363,
    n484,
    n406,
    n21
  );


  xor
  g686
  (
    n728,
    n506,
    n507,
    n500,
    n404
  );


  nand
  g687
  (
    n558,
    n341,
    n464,
    n323,
    n465
  );


  xor
  g688
  (
    n660,
    n322,
    n509,
    n420,
    n522
  );


  nor
  g689
  (
    n684,
    n524,
    n415,
    n438,
    n454
  );


  xor
  g690
  (
    n592,
    n432,
    n481,
    n469,
    n391
  );


  nor
  g691
  (
    n714,
    n398,
    n515,
    n477,
    n490
  );


  and
  g692
  (
    n718,
    n399,
    n448,
    n345,
    n349
  );


  nor
  g693
  (
    n780,
    n492,
    n392,
    n323,
    n324
  );


  xor
  g694
  (
    n771,
    n347,
    n344,
    n389,
    n466
  );


  xor
  g695
  (
    n604,
    n526,
    n336,
    n432,
    n408
  );


  xnor
  g696
  (
    n591,
    n414,
    n95,
    n452,
    n100
  );


  or
  g697
  (
    n623,
    n453,
    n411,
    n335,
    n365
  );


  nand
  g698
  (
    n561,
    n474,
    n25,
    n517,
    n497
  );


  nand
  g699
  (
    n654,
    n26,
    n395,
    n550,
    n388
  );


  xnor
  g700
  (
    KeyWire_0_21,
    n335,
    n409,
    n439,
    n445
  );


  xnor
  g701
  (
    n624,
    n452,
    n360,
    n327,
    n383
  );


  and
  g702
  (
    n570,
    n461,
    n458,
    n541,
    n337
  );


  or
  g703
  (
    n640,
    n99,
    n435,
    n514,
    n454
  );


  or
  g704
  (
    n748,
    n501,
    n421,
    n431,
    n28
  );


  nor
  g705
  (
    n755,
    n464,
    n465,
    n336,
    n357
  );


  or
  g706
  (
    n690,
    n507,
    n489,
    n502,
    n366
  );


  nand
  g707
  (
    n598,
    n413,
    n458,
    n436,
    n511
  );


  nor
  g708
  (
    n559,
    n32,
    n419,
    n26,
    n425
  );


  nand
  g709
  (
    n697,
    n512,
    n325,
    n468,
    n363
  );


  nor
  g710
  (
    n775,
    n459,
    n426,
    n96,
    n485
  );


  nand
  g711
  (
    n738,
    n25,
    n97,
    n430,
    n326
  );


  xor
  g712
  (
    n639,
    n516,
    n478,
    n26,
    n482
  );


  and
  g713
  (
    n615,
    n550,
    n430,
    n547,
    n554
  );


  nand
  g714
  (
    n713,
    n32,
    n322,
    n547,
    n361
  );


  nand
  g715
  (
    n663,
    n377,
    n391,
    n457,
    n538
  );


  nand
  g716
  (
    n743,
    n348,
    n394,
    n333,
    n23
  );


  and
  g717
  (
    n572,
    n451,
    n323,
    n409,
    n520
  );


  or
  g718
  (
    n710,
    n434,
    n421,
    n414,
    n426
  );


  xor
  g719
  (
    n747,
    n423,
    n416,
    n550,
    n476
  );


  xnor
  g720
  (
    n576,
    n475,
    n529,
    n335,
    n440
  );


  nor
  g721
  (
    n670,
    n549,
    n32,
    n362,
    n397
  );


  nor
  g722
  (
    n571,
    n547,
    n97,
    n377,
    n420
  );


  nor
  g723
  (
    n700,
    n481,
    n479,
    n544,
    n469
  );


  xor
  g724
  (
    n699,
    n465,
    n553,
    n421,
    n349
  );


  xor
  g725
  (
    n681,
    n533,
    n376,
    n347,
    n536
  );


  nand
  g726
  (
    n757,
    n441,
    n425,
    n540,
    n488
  );


  nand
  g727
  (
    n613,
    n383,
    n333,
    n548,
    n520
  );


  xnor
  g728
  (
    n645,
    n441,
    n487,
    n98,
    n434
  );


  nor
  g729
  (
    n731,
    n495,
    n424,
    n466,
    n488
  );


  nand
  g730
  (
    n596,
    n457,
    n485,
    n514,
    n385
  );


  and
  g731
  (
    n711,
    n427,
    n436,
    n484,
    n503
  );


  or
  g732
  (
    n722,
    n433,
    n392,
    n415,
    n535
  );


  nand
  g733
  (
    n625,
    n458,
    n412,
    n401,
    n483
  );


  xnor
  g734
  (
    KeyWire_0_7,
    n470,
    n461,
    n538,
    n431
  );


  and
  g735
  (
    n655,
    n405,
    n27,
    n321,
    n349
  );


  and
  g736
  (
    n672,
    n487,
    n529,
    n544,
    n416
  );


  and
  g737
  (
    n774,
    n325,
    n406,
    n328,
    n474
  );


  nor
  g738
  (
    n689,
    n436,
    n399,
    n27,
    n405
  );


  or
  g739
  (
    n665,
    n432,
    n426,
    n484,
    n534
  );


  nand
  g740
  (
    n682,
    n470,
    n474,
    n408,
    n540
  );


  nand
  g741
  (
    n671,
    n412,
    n342,
    n478,
    n23
  );


  nand
  g742
  (
    n557,
    n450,
    n23,
    n322,
    n339
  );


  nor
  g743
  (
    n658,
    n387,
    n467,
    n29,
    n382
  );


  and
  g744
  (
    n588,
    n95,
    n526,
    n476,
    n332
  );


  nand
  g745
  (
    n773,
    n527,
    n407,
    n536,
    n542
  );


  nor
  g746
  (
    n704,
    n386,
    n546,
    n504,
    n340
  );


  xor
  g747
  (
    n607,
    n98,
    n512,
    n510,
    n466
  );


  xor
  g748
  (
    n781,
    n346,
    n522,
    n413,
    n418
  );


  nor
  g749
  (
    n677,
    n345,
    n507,
    n553,
    n537
  );


  and
  g750
  (
    n733,
    n338,
    n22,
    n517,
    n521
  );


  or
  g751
  (
    n793,
    n686,
    n629,
    n617,
    n626
  );


  and
  g752
  (
    n822,
    n668,
    n580,
    n619,
    n620
  );


  or
  g753
  (
    n808,
    n670,
    n678,
    n567,
    n689
  );


  xnor
  g754
  (
    n827,
    n651,
    n594,
    n624,
    n593
  );


  or
  g755
  (
    n812,
    n608,
    n105,
    n690,
    n637
  );


  and
  g756
  (
    n825,
    n667,
    n577,
    n589,
    n106
  );


  or
  g757
  (
    n785,
    n672,
    n102,
    n639,
    n566
  );


  xor
  g758
  (
    n818,
    n681,
    n633,
    n606,
    n604
  );


  nand
  g759
  (
    n819,
    n602,
    n103,
    n582,
    n568
  );


  xor
  g760
  (
    KeyWire_0_52,
    n659,
    n572,
    n614,
    n350
  );


  or
  g761
  (
    n817,
    n352,
    n682,
    n103,
    n585
  );


  and
  g762
  (
    n811,
    n104,
    n597,
    n351,
    n592
  );


  xnor
  g763
  (
    n829,
    n687,
    n674,
    n352,
    n575
  );


  xor
  g764
  (
    n788,
    n685,
    n646,
    n605,
    n350
  );


  or
  g765
  (
    n790,
    n611,
    n105,
    n662,
    n688
  );


  xnor
  g766
  (
    n797,
    n654,
    n105,
    n621,
    n600
  );


  xor
  g767
  (
    n820,
    n644,
    n652,
    n667,
    n627
  );


  and
  g768
  (
    n798,
    n607,
    n658,
    n691,
    n622
  );


  and
  g769
  (
    n828,
    n107,
    n676,
    n673
  );


  xor
  g770
  (
    n815,
    n636,
    n351,
    n686,
    n649
  );


  xnor
  g771
  (
    n802,
    n102,
    n685,
    n578,
    n642
  );


  nand
  g772
  (
    n804,
    n671,
    n591,
    n681,
    n647
  );


  nor
  g773
  (
    n807,
    n668,
    n106,
    n351,
    n666
  );


  nor
  g774
  (
    n794,
    n571,
    n352,
    n623,
    n596
  );


  xor
  g775
  (
    n830,
    n573,
    n692,
    n590,
    n584
  );


  nor
  g776
  (
    n787,
    n616,
    n350,
    n680,
    n625
  );


  xnor
  g777
  (
    KeyWire_0_8,
    n628,
    n613,
    n678,
    n107
  );


  nor
  g778
  (
    n809,
    n640,
    n565,
    n105,
    n103
  );


  and
  g779
  (
    n800,
    n660,
    n672,
    n609,
    n691
  );


  nor
  g780
  (
    n805,
    n650,
    n618,
    n684,
    n631
  );


  or
  g781
  (
    n816,
    n630,
    n574,
    n106,
    n599
  );


  nor
  g782
  (
    n796,
    n103,
    n583,
    n641,
    n653
  );


  nand
  g783
  (
    n823,
    n648,
    n104,
    n576,
    n684
  );


  nor
  g784
  (
    n814,
    n569,
    n595,
    n673,
    n682
  );


  xor
  g785
  (
    n813,
    n689,
    n645,
    n670,
    n665
  );


  or
  g786
  (
    KeyWire_0_55,
    n104,
    n677,
    n692,
    n581
  );


  xor
  g787
  (
    n824,
    n107,
    n352,
    n615,
    n688
  );


  and
  g788
  (
    KeyWire_0_63,
    n351,
    n675,
    n669,
    n601
  );


  or
  g789
  (
    n826,
    n598,
    n683,
    n579,
    n632
  );


  nor
  g790
  (
    n789,
    n104,
    n107,
    n664,
    n612
  );


  xnor
  g791
  (
    n786,
    n661,
    n106,
    n663,
    n677
  );


  nor
  g792
  (
    n803,
    n669,
    n655,
    n603,
    n680
  );


  xor
  g793
  (
    KeyWire_0_49,
    n657,
    n638,
    n635,
    n679
  );


  nor
  g794
  (
    n810,
    n690,
    n634,
    n610,
    n675
  );


  nand
  g795
  (
    KeyWire_0_11,
    n656,
    n588,
    n587,
    n683
  );


  xnor
  g796
  (
    n791,
    n687,
    n674,
    n586,
    n643
  );


  xnor
  g797
  (
    n801,
    n570,
    n350,
    n671,
    n679
  );


  buf
  g798
  (
    n875,
    n798
  );


  not
  g799
  (
    n864,
    n794
  );


  buf
  g800
  (
    n840,
    n109
  );


  buf
  g801
  (
    n847,
    n805
  );


  buf
  g802
  (
    n859,
    n804
  );


  buf
  g803
  (
    n862,
    n793
  );


  buf
  g804
  (
    n865,
    n114
  );


  buf
  g805
  (
    n869,
    n112
  );


  not
  g806
  (
    n844,
    n113
  );


  buf
  g807
  (
    n831,
    n787
  );


  not
  g808
  (
    n832,
    n108
  );


  not
  g809
  (
    n866,
    n113
  );


  buf
  g810
  (
    KeyWire_0_14,
    n111
  );


  buf
  g811
  (
    n860,
    n113
  );


  buf
  g812
  (
    n876,
    n806
  );


  buf
  g813
  (
    n849,
    n787
  );


  buf
  g814
  (
    n845,
    n795
  );


  buf
  g815
  (
    n872,
    n791
  );


  not
  g816
  (
    n871,
    n801
  );


  buf
  g817
  (
    n868,
    n803
  );


  not
  g818
  (
    n834,
    n790
  );


  buf
  g819
  (
    n878,
    n808
  );


  not
  g820
  (
    n873,
    n785
  );


  not
  g821
  (
    n877,
    n795
  );


  not
  g822
  (
    n880,
    n802
  );


  buf
  g823
  (
    n870,
    n109
  );


  buf
  g824
  (
    n838,
    n112
  );


  not
  g825
  (
    n848,
    n803
  );


  buf
  g826
  (
    KeyWire_0_15,
    n801
  );


  not
  g827
  (
    n835,
    n788
  );


  buf
  g828
  (
    n857,
    n797
  );


  not
  g829
  (
    n861,
    n793
  );


  buf
  g830
  (
    n867,
    n788
  );


  not
  g831
  (
    n841,
    n112
  );


  not
  g832
  (
    n837,
    n108
  );


  not
  g833
  (
    n858,
    n110
  );


  not
  g834
  (
    n853,
    n792
  );


  not
  g835
  (
    KeyWire_0_12,
    n792
  );


  buf
  g836
  (
    n850,
    n807
  );


  buf
  g837
  (
    n843,
    n791
  );


  xnor
  g838
  (
    n839,
    n796,
    n789
  );


  nor
  g839
  (
    n856,
    n112,
    n808,
    n790,
    n108
  );


  nand
  g840
  (
    n852,
    n802,
    n809,
    n786,
    n789
  );


  nand
  g841
  (
    n851,
    n109,
    n806,
    n108,
    n796
  );


  and
  g842
  (
    n863,
    n109,
    n799,
    n804,
    n785
  );


  nor
  g843
  (
    n879,
    n797,
    n114,
    n786,
    n111
  );


  nor
  g844
  (
    n842,
    n807,
    n110,
    n111
  );


  xor
  g845
  (
    n855,
    n784,
    n110,
    n805,
    n798
  );


  nand
  g846
  (
    n854,
    n113,
    n800,
    n794
  );


  xnor
  g847
  (
    n833,
    n799,
    n111,
    n114
  );


  nor
  g848
  (
    n915,
    n856,
    n864,
    n847,
    n870
  );


  xnor
  g849
  (
    n884,
    n849,
    n854,
    n846,
    n862
  );


  xnor
  g850
  (
    n886,
    n851,
    n853,
    n849,
    n836
  );


  and
  g851
  (
    n885,
    n872,
    n859,
    n869,
    n842
  );


  nor
  g852
  (
    n900,
    n849,
    n861,
    n854,
    n871
  );


  nor
  g853
  (
    n911,
    n832,
    n831,
    n833,
    n843
  );


  nand
  g854
  (
    n904,
    n850,
    n856,
    n852,
    n869
  );


  or
  g855
  (
    KeyWire_0_17,
    n835,
    n852,
    n844,
    n865
  );


  xnor
  g856
  (
    n896,
    n864,
    n833,
    n834
  );


  nand
  g857
  (
    n914,
    n864,
    n834,
    n866,
    n863
  );


  xnor
  g858
  (
    n891,
    n845,
    n861,
    n841,
    n865
  );


  nor
  g859
  (
    n916,
    n848,
    n859,
    n845,
    n870
  );


  xnor
  g860
  (
    n890,
    n860,
    n849,
    n832,
    n855
  );


  xor
  g861
  (
    n881,
    n862,
    n855,
    n837,
    n840
  );


  or
  g862
  (
    n919,
    n863,
    n848,
    n861,
    n868
  );


  nor
  g863
  (
    n920,
    n854,
    n845,
    n855,
    n862
  );


  xor
  g864
  (
    n905,
    n838,
    n852,
    n864,
    n843
  );


  nand
  g865
  (
    n902,
    n857,
    n843,
    n842,
    n868
  );


  nand
  g866
  (
    n899,
    n867,
    n865,
    n844,
    n850
  );


  nand
  g867
  (
    n922,
    n850,
    n869,
    n834,
    n836
  );


  xor
  g868
  (
    n913,
    n867,
    n871,
    n851,
    n866
  );


  or
  g869
  (
    n907,
    n839,
    n861,
    n853,
    n847
  );


  or
  g870
  (
    n906,
    n841,
    n857,
    n858
  );


  and
  g871
  (
    n888,
    n863,
    n859,
    n832,
    n836
  );


  or
  g872
  (
    n912,
    n870,
    n860,
    n835,
    n837
  );


  xor
  g873
  (
    n882,
    n848,
    n846,
    n868,
    n872
  );


  nor
  g874
  (
    n889,
    n866,
    n837,
    n853,
    n839
  );


  nand
  g875
  (
    n883,
    n840,
    n835,
    n859,
    n872
  );


  or
  g876
  (
    n887,
    n843,
    n841,
    n872,
    n858
  );


  xnor
  g877
  (
    n894,
    n871,
    n839,
    n850,
    n848
  );


  xor
  g878
  (
    n909,
    n835,
    n836,
    n860,
    n866
  );


  xnor
  g879
  (
    n895,
    n871,
    n851,
    n831,
    n870
  );


  xnor
  g880
  (
    n892,
    n833,
    n838,
    n869,
    n840
  );


  nand
  g881
  (
    n898,
    n842,
    n854,
    n834,
    n857
  );


  nand
  g882
  (
    n921,
    n867,
    n852,
    n858,
    n841
  );


  and
  g883
  (
    n901,
    n846,
    n855,
    n844
  );


  or
  g884
  (
    n893,
    n867,
    n858,
    n860,
    n863
  );


  nand
  g885
  (
    n917,
    n847,
    n862,
    n840,
    n873
  );


  or
  g886
  (
    n897,
    n865,
    n851,
    n837,
    n838
  );


  xor
  g887
  (
    n918,
    n868,
    n845,
    n839,
    n856
  );


  or
  g888
  (
    n908,
    n853,
    n832,
    n873,
    n842
  );


  xnor
  g889
  (
    n910,
    n847,
    n846,
    n838,
    n856
  );


  xnor
  g890
  (
    n936,
    n885,
    n353,
    n878,
    n715
  );


  nand
  g891
  (
    n925,
    n877,
    n874,
    n719,
    n704
  );


  xnor
  g892
  (
    n931,
    n880,
    n915,
    n917,
    n721
  );


  xnor
  g893
  (
    n932,
    n725,
    n353,
    n900,
    n724
  );


  xor
  g894
  (
    n955,
    n896,
    n724,
    n708,
    n701
  );


  nand
  g895
  (
    n949,
    n877,
    n722,
    n721,
    n711
  );


  nand
  g896
  (
    n937,
    n909,
    n875,
    n700,
    n879
  );


  or
  g897
  (
    n959,
    n695,
    n356,
    n702,
    n694
  );


  and
  g898
  (
    n961,
    n874,
    n918,
    n702,
    n876
  );


  nand
  g899
  (
    n951,
    n879,
    n895,
    n723,
    n556
  );


  or
  g900
  (
    n926,
    n355,
    n875,
    n697,
    n889
  );


  nor
  g901
  (
    KeyWire_0_13,
    n884,
    n904,
    n696,
    n717
  );


  xor
  g902
  (
    n956,
    n877,
    n353,
    n693,
    n901
  );


  xor
  g903
  (
    n940,
    n880,
    n712,
    n911
  );


  or
  g904
  (
    n927,
    n880,
    n707,
    n716,
    n710
  );


  xor
  g905
  (
    n948,
    n354,
    n709,
    n718,
    n903
  );


  nand
  g906
  (
    n953,
    n908,
    n899,
    n878,
    n913
  );


  and
  g907
  (
    n933,
    n879,
    n716,
    n887,
    n556
  );


  xor
  g908
  (
    n943,
    n696,
    n705,
    n888,
    n706
  );


  nor
  g909
  (
    n928,
    n704,
    n922,
    n700,
    n698
  );


  or
  g910
  (
    n935,
    n897,
    n722,
    n919,
    n723
  );


  nand
  g911
  (
    n962,
    n891,
    n906,
    n709,
    n698
  );


  nor
  g912
  (
    n934,
    n910,
    n555,
    n705,
    n898
  );


  xnor
  g913
  (
    n923,
    n878,
    n878,
    n355,
    n894
  );


  nand
  g914
  (
    n947,
    n720,
    n354,
    n876
  );


  nor
  g915
  (
    n960,
    n905,
    n556,
    n880,
    n356
  );


  nand
  g916
  (
    n954,
    n875,
    n916,
    n694,
    n902
  );


  xnor
  g917
  (
    n924,
    n714,
    n355,
    n877,
    n875
  );


  or
  g918
  (
    n939,
    n717,
    n713,
    n555
  );


  nand
  g919
  (
    n929,
    n719,
    n879,
    n695,
    n715
  );


  xnor
  g920
  (
    n942,
    n714,
    n876,
    n873,
    n893
  );


  nor
  g921
  (
    KeyWire_0_51,
    n554,
    n883,
    n706,
    n707
  );


  xnor
  g922
  (
    n944,
    n720,
    n701,
    n555,
    n699
  );


  xor
  g923
  (
    n938,
    n699,
    n873,
    n555,
    n556
  );


  xor
  g924
  (
    n958,
    n708,
    n718,
    n892,
    n356
  );


  nand
  g925
  (
    n952,
    n874,
    n693,
    n354,
    n912
  );


  and
  g926
  (
    n930,
    n354,
    n921,
    n703,
    n356
  );


  or
  g927
  (
    n957,
    n886,
    n874,
    n355,
    n907
  );


  nand
  g928
  (
    n946,
    n914,
    n890,
    n920,
    n697
  );


  and
  g929
  (
    n945,
    n710,
    n711,
    n353,
    n703
  );


  nor
  g930
  (
    n1010,
    n941,
    n930,
    n827,
    n748
  );


  and
  g931
  (
    n987,
    n732,
    n764,
    n932,
    n774
  );


  nor
  g932
  (
    KeyWire_0_48,
    n933,
    n761,
    n951,
    n952
  );


  nand
  g933
  (
    n1016,
    n955,
    n753,
    n778,
    n777
  );


  xnor
  g934
  (
    n977,
    n742,
    n823,
    n819,
    n945
  );


  or
  g935
  (
    n998,
    n953,
    n735,
    n947,
    n959
  );


  xnor
  g936
  (
    n969,
    n775,
    n812,
    n954,
    n952
  );


  or
  g937
  (
    n979,
    n811,
    n778,
    n751,
    n735
  );


  xor
  g938
  (
    n972,
    n934,
    n779,
    n936,
    n738
  );


  xor
  g939
  (
    n964,
    n926,
    n768,
    n781,
    n772
  );


  or
  g940
  (
    n986,
    n809,
    n738,
    n938,
    n759
  );


  xor
  g941
  (
    n1001,
    n825,
    n943,
    n762,
    n814
  );


  or
  g942
  (
    n993,
    n755,
    n754,
    n816,
    n744
  );


  xor
  g943
  (
    n1003,
    n780,
    n743,
    n820,
    n948
  );


  nor
  g944
  (
    n980,
    n741,
    n771,
    n824,
    n773
  );


  xor
  g945
  (
    n971,
    n731,
    n820,
    n828,
    n783
  );


  xor
  g946
  (
    n1015,
    n960,
    n810,
    n734,
    n782
  );


  and
  g947
  (
    n997,
    n955,
    n775,
    n821,
    n928
  );


  and
  g948
  (
    n1012,
    n727,
    n773,
    n761,
    n956
  );


  nor
  g949
  (
    n978,
    n756,
    n827,
    n829,
    n822
  );


  xnor
  g950
  (
    n983,
    n729,
    n925,
    n733,
    n817
  );


  nor
  g951
  (
    n1000,
    n733,
    n757,
    n931,
    n772
  );


  xnor
  g952
  (
    n1018,
    n740,
    n754,
    n760,
    n826
  );


  xnor
  g953
  (
    n985,
    n755,
    n927,
    n781,
    n828
  );


  xor
  g954
  (
    n996,
    n748,
    n825,
    n935,
    n951
  );


  xnor
  g955
  (
    n1009,
    n745,
    n741,
    n771,
    n830
  );


  xnor
  g956
  (
    n992,
    n962,
    n818,
    n817,
    n739
  );


  and
  g957
  (
    n1013,
    n929,
    n760,
    n937,
    n737
  );


  and
  g958
  (
    n994,
    n746,
    n756,
    n774,
    n757
  );


  or
  g959
  (
    n1006,
    n822,
    n734,
    n946,
    n777
  );


  or
  g960
  (
    n968,
    n942,
    n766,
    n725,
    n826
  );


  or
  g961
  (
    n963,
    n766,
    n769,
    n758,
    n816
  );


  xnor
  g962
  (
    n1007,
    n954,
    n780,
    n749,
    n763
  );


  xnor
  g963
  (
    n990,
    n949,
    n783,
    n744,
    n823
  );


  and
  g964
  (
    n975,
    n812,
    n811,
    n818,
    n739
  );


  nor
  g965
  (
    n1008,
    n813,
    n737,
    n939,
    n751
  );


  xor
  g966
  (
    n974,
    n728,
    n747,
    n829,
    n957
  );


  and
  g967
  (
    n988,
    n815,
    n829,
    n923,
    n727
  );


  and
  g968
  (
    n1017,
    n736,
    n828,
    n731,
    n776
  );


  nor
  g969
  (
    KeyWire_0_31,
    n747,
    n813,
    n764,
    n752
  );


  xor
  g970
  (
    n984,
    n762,
    n940,
    n948,
    n827
  );


  nor
  g971
  (
    n1005,
    n749,
    n829,
    n726
  );


  and
  g972
  (
    KeyWire_0_42,
    n830,
    n770,
    n736,
    n776
  );


  xnor
  g973
  (
    n965,
    n759,
    n830,
    n959,
    n769
  );


  xor
  g974
  (
    n966,
    n824,
    n746,
    n830,
    n752
  );


  xor
  g975
  (
    n989,
    n949,
    n740,
    n770,
    n958
  );


  nand
  g976
  (
    n1004,
    n767,
    n810,
    n730,
    n815
  );


  xnor
  g977
  (
    n982,
    n729,
    n758,
    n742,
    n950
  );


  nor
  g978
  (
    n970,
    n768,
    n950,
    n765,
    n728
  );


  xnor
  g979
  (
    n999,
    n814,
    n767,
    n753,
    n782
  );


  nor
  g980
  (
    n1011,
    n956,
    n962,
    n961
  );


  xor
  g981
  (
    n1014,
    n750,
    n953,
    n819,
    n924
  );


  and
  g982
  (
    n973,
    n827,
    n730,
    n957,
    n743
  );


  and
  g983
  (
    n1002,
    n944,
    n763,
    n821,
    n960
  );


  and
  g984
  (
    n991,
    n958,
    n750,
    n745,
    n765
  );


  nand
  g985
  (
    n967,
    n828,
    n947,
    n779,
    n732
  );


  or
  g986
  (
    KeyWire_0_58,
    n967,
    n1008,
    n977,
    n1006
  );


  nand
  g987
  (
    n1027,
    n985,
    n1011,
    n997,
    n1004
  );


  nor
  g988
  (
    n1031,
    n995,
    n1002,
    n1000,
    n966
  );


  xor
  g989
  (
    n1029,
    n980,
    n989,
    n1003,
    n964
  );


  xor
  g990
  (
    n1024,
    n994,
    n1005,
    n1007,
    n1012
  );


  and
  g991
  (
    n1032,
    n976,
    n1013,
    n983,
    n998
  );


  xor
  g992
  (
    n1022,
    n992,
    n990,
    n969,
    n968
  );


  and
  g993
  (
    n1030,
    n1018,
    n986,
    n970,
    n1015
  );


  and
  g994
  (
    n1025,
    n1014,
    n988,
    n1001,
    n978
  );


  and
  g995
  (
    n1020,
    n972,
    n982,
    n971,
    n987
  );


  xor
  g996
  (
    n1023,
    n984,
    n981,
    n991,
    n999
  );


  xnor
  g997
  (
    n1019,
    n1010,
    n1017,
    n974,
    n965
  );


  xor
  g998
  (
    n1021,
    n979,
    n1009,
    n973,
    n1016
  );


  xnor
  g999
  (
    n1028,
    n963,
    n996,
    n993,
    n975
  );


  xnor
  KeyGate_0_0
  (
    n637,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n631,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n107,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n585,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n726,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n396,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n435,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n776,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n806,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n602,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n512,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n795,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n874,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n950,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n836,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n846,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n264,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n903,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n667,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n226,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n470,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n687,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n664,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n110,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n65,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n181,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n653,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n483,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n132,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n364,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n333,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n981,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n169,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n376,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n35,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n362,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n266,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n113,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n746,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n296,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n112,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n490,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n995,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n778,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n420,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n752,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n702,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n539,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n976,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n792,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n346,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n941,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n799,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n127,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n272,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n784,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n695,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n552,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n1026,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n732,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n118,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n659,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n231,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n821,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

