// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1375_21_1 written by SynthGen on 2021/06/15 15:04:53
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1375_21_1 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21,
 n899, n912, n919, n930, n909, n936, n907, n924,
 n937, n904, n927, n902, n934, n931, n985, n1020,
 n1045, n1037, n1042, n1040, n1019, n1041, n1039, n1031,
 n1022, n1032, n1035, n1046, n1038, n1348, n1382, n1386,
 n1383, n1384, n1379, n1388, n1380, n1387, n1389, n1381,
 n1378, n1396, n1394, n1395, n1393);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21;

output n899, n912, n919, n930, n909, n936, n907, n924,
 n937, n904, n927, n902, n934, n931, n985, n1020,
 n1045, n1037, n1042, n1040, n1019, n1041, n1039, n1031,
 n1022, n1032, n1035, n1046, n1038, n1348, n1382, n1386,
 n1383, n1384, n1379, n1388, n1380, n1387, n1389, n1381,
 n1378, n1396, n1394, n1395, n1393;

wire n22, n23, n24, n25, n26, n27, n28, n29,
 n30, n31, n32, n33, n34, n35, n36, n37,
 n38, n39, n40, n41, n42, n43, n44, n45,
 n46, n47, n48, n49, n50, n51, n52, n53,
 n54, n55, n56, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n67, n68, n69,
 n70, n71, n72, n73, n74, n75, n76, n77,
 n78, n79, n80, n81, n82, n83, n84, n85,
 n86, n87, n88, n89, n90, n91, n92, n93,
 n94, n95, n96, n97, n98, n99, n100, n101,
 n102, n103, n104, n105, n106, n107, n108, n109,
 n110, n111, n112, n113, n114, n115, n116, n117,
 n118, n119, n120, n121, n122, n123, n124, n125,
 n126, n127, n128, n129, n130, n131, n132, n133,
 n134, n135, n136, n137, n138, n139, n140, n141,
 n142, n143, n144, n145, n146, n147, n148, n149,
 n150, n151, n152, n153, n154, n155, n156, n157,
 n158, n159, n160, n161, n162, n163, n164, n165,
 n166, n167, n168, n169, n170, n171, n172, n173,
 n174, n175, n176, n177, n178, n179, n180, n181,
 n182, n183, n184, n185, n186, n187, n188, n189,
 n190, n191, n192, n193, n194, n195, n196, n197,
 n198, n199, n200, n201, n202, n203, n204, n205,
 n206, n207, n208, n209, n210, n211, n212, n213,
 n214, n215, n216, n217, n218, n219, n220, n221,
 n222, n223, n224, n225, n226, n227, n228, n229,
 n230, n231, n232, n233, n234, n235, n236, n237,
 n238, n239, n240, n241, n242, n243, n244, n245,
 n246, n247, n248, n249, n250, n251, n252, n253,
 n254, n255, n256, n257, n258, n259, n260, n261,
 n262, n263, n264, n265, n266, n267, n268, n269,
 n270, n271, n272, n273, n274, n275, n276, n277,
 n278, n279, n280, n281, n282, n283, n284, n285,
 n286, n287, n288, n289, n290, n291, n292, n293,
 n294, n295, n296, n297, n298, n299, n300, n301,
 n302, n303, n304, n305, n306, n307, n308, n309,
 n310, n311, n312, n313, n314, n315, n316, n317,
 n318, n319, n320, n321, n322, n323, n324, n325,
 n326, n327, n328, n329, n330, n331, n332, n333,
 n334, n335, n336, n337, n338, n339, n340, n341,
 n342, n343, n344, n345, n346, n347, n348, n349,
 n350, n351, n352, n353, n354, n355, n356, n357,
 n358, n359, n360, n361, n362, n363, n364, n365,
 n366, n367, n368, n369, n370, n371, n372, n373,
 n374, n375, n376, n377, n378, n379, n380, n381,
 n382, n383, n384, n385, n386, n387, n388, n389,
 n390, n391, n392, n393, n394, n395, n396, n397,
 n398, n399, n400, n401, n402, n403, n404, n405,
 n406, n407, n408, n409, n410, n411, n412, n413,
 n414, n415, n416, n417, n418, n419, n420, n421,
 n422, n423, n424, n425, n426, n427, n428, n429,
 n430, n431, n432, n433, n434, n435, n436, n437,
 n438, n439, n440, n441, n442, n443, n444, n445,
 n446, n447, n448, n449, n450, n451, n452, n453,
 n454, n455, n456, n457, n458, n459, n460, n461,
 n462, n463, n464, n465, n466, n467, n468, n469,
 n470, n471, n472, n473, n474, n475, n476, n477,
 n478, n479, n480, n481, n482, n483, n484, n485,
 n486, n487, n488, n489, n490, n491, n492, n493,
 n494, n495, n496, n497, n498, n499, n500, n501,
 n502, n503, n504, n505, n506, n507, n508, n509,
 n510, n511, n512, n513, n514, n515, n516, n517,
 n518, n519, n520, n521, n522, n523, n524, n525,
 n526, n527, n528, n529, n530, n531, n532, n533,
 n534, n535, n536, n537, n538, n539, n540, n541,
 n542, n543, n544, n545, n546, n547, n548, n549,
 n550, n551, n552, n553, n554, n555, n556, n557,
 n558, n559, n560, n561, n562, n563, n564, n565,
 n566, n567, n568, n569, n570, n571, n572, n573,
 n574, n575, n576, n577, n578, n579, n580, n581,
 n582, n583, n584, n585, n586, n587, n588, n589,
 n590, n591, n592, n593, n594, n595, n596, n597,
 n598, n599, n600, n601, n602, n603, n604, n605,
 n606, n607, n608, n609, n610, n611, n612, n613,
 n614, n615, n616, n617, n618, n619, n620, n621,
 n622, n623, n624, n625, n626, n627, n628, n629,
 n630, n631, n632, n633, n634, n635, n636, n637,
 n638, n639, n640, n641, n642, n643, n644, n645,
 n646, n647, n648, n649, n650, n651, n652, n653,
 n654, n655, n656, n657, n658, n659, n660, n661,
 n662, n663, n664, n665, n666, n667, n668, n669,
 n670, n671, n672, n673, n674, n675, n676, n677,
 n678, n679, n680, n681, n682, n683, n684, n685,
 n686, n687, n688, n689, n690, n691, n692, n693,
 n694, n695, n696, n697, n698, n699, n700, n701,
 n702, n703, n704, n705, n706, n707, n708, n709,
 n710, n711, n712, n713, n714, n715, n716, n717,
 n718, n719, n720, n721, n722, n723, n724, n725,
 n726, n727, n728, n729, n730, n731, n732, n733,
 n734, n735, n736, n737, n738, n739, n740, n741,
 n742, n743, n744, n745, n746, n747, n748, n749,
 n750, n751, n752, n753, n754, n755, n756, n757,
 n758, n759, n760, n761, n762, n763, n764, n765,
 n766, n767, n768, n769, n770, n771, n772, n773,
 n774, n775, n776, n777, n778, n779, n780, n781,
 n782, n783, n784, n785, n786, n787, n788, n789,
 n790, n791, n792, n793, n794, n795, n796, n797,
 n798, n799, n800, n801, n802, n803, n804, n805,
 n806, n807, n808, n809, n810, n811, n812, n813,
 n814, n815, n816, n817, n818, n819, n820, n821,
 n822, n823, n824, n825, n826, n827, n828, n829,
 n830, n831, n832, n833, n834, n835, n836, n837,
 n838, n839, n840, n841, n842, n843, n844, n845,
 n846, n847, n848, n849, n850, n851, n852, n853,
 n854, n855, n856, n857, n858, n859, n860, n861,
 n862, n863, n864, n865, n866, n867, n868, n869,
 n870, n871, n872, n873, n874, n875, n876, n877,
 n878, n879, n880, n881, n882, n883, n884, n885,
 n886, n887, n888, n889, n890, n891, n892, n893,
 n894, n895, n896, n897, n898, n900, n901, n903,
 n905, n906, n908, n910, n911, n913, n914, n915,
 n916, n917, n918, n920, n921, n922, n923, n925,
 n926, n928, n929, n932, n933, n935, n938, n939,
 n940, n941, n942, n943, n944, n945, n946, n947,
 n948, n949, n950, n951, n952, n953, n954, n955,
 n956, n957, n958, n959, n960, n961, n962, n963,
 n964, n965, n966, n967, n968, n969, n970, n971,
 n972, n973, n974, n975, n976, n977, n978, n979,
 n980, n981, n982, n983, n984, n986, n987, n988,
 n989, n990, n991, n992, n993, n994, n995, n996,
 n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
 n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
 n1013, n1014, n1015, n1016, n1017, n1018, n1021, n1023,
 n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1033,
 n1034, n1036, n1043, n1044, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
 n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
 n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
 n1372, n1373, n1374, n1375, n1376, n1377, n1385, n1390,
 n1391, n1392;

not  g0 (n53, n1);
buf  g1 (n54, n17);
buf  g2 (n71, n15);
buf  g3 (n79, n2);
buf  g4 (n57, n14);
not  g5 (n69, n6);
not  g6 (n99, n14);
not  g7 (n50, n12);
buf  g8 (n64, n3);
buf  g9 (n45, n10);
buf  g10 (n31, n21);
buf  g11 (n70, n17);
buf  g12 (n66, n7);
not  g13 (n27, n1);
not  g14 (n101, n20);
not  g15 (n36, n4);
not  g16 (n95, n13);
buf  g17 (n37, n4);
not  g18 (n23, n4);
not  g19 (n38, n11);
buf  g20 (n26, n19);
buf  g21 (n74, n17);
buf  g22 (n56, n13);
buf  g23 (n41, n18);
buf  g24 (n80, n18);
not  g25 (n102, n11);
buf  g26 (n67, n3);
buf  g27 (n75, n16);
not  g28 (n100, n9);
buf  g29 (n68, n6);
not  g30 (n65, n20);
not  g31 (n103, n7);
buf  g32 (n32, n5);
buf  g33 (n78, n12);
not  g34 (n58, n11);
not  g35 (n92, n3);
buf  g36 (n89, n21);
not  g37 (n87, n5);
buf  g38 (n24, n12);
not  g39 (n22, n10);
not  g40 (n90, n20);
buf  g41 (n25, n10);
not  g42 (n73, n13);
not  g43 (n60, n19);
buf  g44 (n84, n2);
not  g45 (n93, n8);
not  g46 (n88, n1);
buf  g47 (n63, n21);
not  g48 (n97, n19);
buf  g49 (n33, n14);
buf  g50 (n76, n8);
not  g51 (n82, n8);
not  g52 (n98, n10);
not  g53 (n77, n14);
buf  g54 (n46, n13);
buf  g55 (n44, n2);
not  g56 (n30, n16);
not  g57 (n62, n8);
buf  g58 (n86, n7);
not  g59 (n47, n18);
not  g60 (n40, n17);
not  g61 (n91, n5);
buf  g62 (n83, n15);
not  g63 (n59, n15);
buf  g64 (n39, n3);
buf  g65 (n72, n12);
buf  g66 (n85, n16);
buf  g67 (n61, n21);
buf  g68 (n104, n1);
not  g69 (n105, n18);
buf  g70 (n55, n16);
not  g71 (n29, n11);
not  g72 (n52, n9);
buf  g73 (n48, n6);
buf  g74 (n34, n6);
not  g75 (n51, n7);
not  g76 (n96, n2);
not  g77 (n28, n19);
buf  g78 (n43, n9);
buf  g79 (n49, n4);
not  g80 (n42, n15);
not  g81 (n35, n20);
not  g82 (n81, n5);
not  g83 (n94, n9);
buf  g84 (n188, n83);
buf  g85 (n224, n56);
buf  g86 (n225, n82);
buf  g87 (n242, n32);
buf  g88 (n382, n66);
not  g89 (n386, n44);
buf  g90 (n288, n39);
buf  g91 (n227, n60);
not  g92 (n365, n86);
not  g93 (n243, n84);
buf  g94 (n377, n89);
buf  g95 (n159, n35);
not  g96 (n289, n60);
not  g97 (n371, n54);
not  g98 (n317, n78);
not  g99 (n276, n45);
not  g100 (n133, n66);
not  g101 (n108, n67);
buf  g102 (n249, n26);
not  g103 (n362, n89);
not  g104 (n143, n57);
buf  g105 (n292, n28);
not  g106 (n393, n90);
not  g107 (n303, n70);
not  g108 (n168, n68);
not  g109 (n346, n77);
buf  g110 (n154, n82);
not  g111 (n172, n98);
not  g112 (n384, n81);
not  g113 (n403, n48);
buf  g114 (n182, n45);
buf  g115 (n389, n38);
buf  g116 (n241, n87);
not  g117 (n201, n73);
not  g118 (n174, n41);
buf  g119 (n200, n57);
buf  g120 (n264, n100);
not  g121 (n397, n75);
buf  g122 (n301, n100);
buf  g123 (n162, n79);
buf  g124 (n266, n44);
not  g125 (n245, n62);
not  g126 (n323, n62);
buf  g127 (n205, n32);
buf  g128 (n165, n99);
not  g129 (n274, n51);
not  g130 (n146, n92);
not  g131 (n291, n58);
buf  g132 (n373, n80);
not  g133 (n329, n81);
buf  g134 (n420, n44);
buf  g135 (n171, n92);
buf  g136 (n216, n72);
buf  g137 (n214, n94);
not  g138 (n107, n43);
buf  g139 (n111, n52);
buf  g140 (n271, n26);
buf  g141 (n331, n43);
not  g142 (n151, n39);
not  g143 (n232, n30);
not  g144 (n211, n43);
buf  g145 (n226, n34);
not  g146 (n370, n84);
not  g147 (n192, n57);
buf  g148 (n358, n53);
buf  g149 (n110, n24);
not  g150 (n234, n85);
buf  g151 (n353, n38);
buf  g152 (n186, n34);
not  g153 (n410, n49);
not  g154 (n209, n93);
not  g155 (n124, n33);
not  g156 (n144, n31);
not  g157 (n220, n85);
not  g158 (n170, n97);
not  g159 (n388, n53);
buf  g160 (n212, n49);
buf  g161 (n324, n72);
buf  g162 (n175, n25);
not  g163 (n375, n63);
buf  g164 (n251, n50);
not  g165 (n176, n83);
not  g166 (n374, n64);
buf  g167 (n217, n29);
not  g168 (n153, n57);
buf  g169 (n126, n93);
buf  g170 (n137, n33);
buf  g171 (n263, n29);
not  g172 (n296, n79);
not  g173 (n202, n76);
buf  g174 (n412, n58);
buf  g175 (n204, n60);
not  g176 (n235, n61);
not  g177 (n414, n40);
buf  g178 (n284, n25);
not  g179 (n173, n44);
buf  g180 (n307, n35);
not  g181 (n299, n24);
buf  g182 (n339, n53);
not  g183 (n319, n41);
not  g184 (n312, n74);
buf  g185 (n309, n89);
not  g186 (n277, n56);
buf  g187 (n113, n26);
not  g188 (n394, n55);
not  g189 (n421, n83);
not  g190 (n240, n49);
not  g191 (n161, n97);
not  g192 (n341, n47);
not  g193 (n247, n94);
not  g194 (n318, n27);
buf  g195 (n194, n73);
buf  g196 (n123, n40);
buf  g197 (n304, n85);
not  g198 (n295, n82);
buf  g199 (n298, n23);
not  g200 (n351, n88);
not  g201 (n334, n45);
buf  g202 (n239, n29);
not  g203 (n340, n91);
buf  g204 (n206, n58);
not  g205 (n290, n85);
not  g206 (n286, n82);
buf  g207 (n333, n51);
not  g208 (n155, n36);
buf  g209 (n366, n91);
buf  g210 (n409, n77);
not  g211 (n136, n61);
not  g212 (n253, n23);
not  g213 (n342, n71);
buf  g214 (n268, n59);
buf  g215 (n367, n51);
not  g216 (n387, n80);
not  g217 (n140, n37);
buf  g218 (n158, n35);
not  g219 (n407, n33);
buf  g220 (n352, n50);
buf  g221 (n197, n64);
buf  g222 (n281, n95);
not  g223 (n326, n50);
buf  g224 (n308, n68);
not  g225 (n280, n86);
buf  g226 (n125, n76);
buf  g227 (n395, n22);
buf  g228 (n230, n36);
not  g229 (n398, n64);
not  g230 (n213, n68);
not  g231 (n190, n31);
buf  g232 (n355, n92);
buf  g233 (n385, n37);
buf  g234 (n369, n34);
buf  g235 (n218, n88);
not  g236 (n343, n47);
buf  g237 (n167, n99);
not  g238 (n166, n43);
buf  g239 (n347, n27);
not  g240 (n294, n97);
buf  g241 (n272, n52);
buf  g242 (n325, n23);
not  g243 (n160, n100);
buf  g244 (n273, n25);
buf  g245 (n164, n99);
buf  g246 (n223, n58);
not  g247 (n238, n99);
buf  g248 (n219, n74);
not  g249 (n418, n24);
buf  g250 (n256, n69);
buf  g251 (n415, n67);
not  g252 (n364, n38);
not  g253 (n114, n92);
not  g254 (n129, n45);
not  g255 (n178, n70);
buf  g256 (n344, n42);
not  g257 (n121, n54);
buf  g258 (n348, n90);
not  g259 (n116, n41);
buf  g260 (n328, n67);
buf  g261 (n285, n49);
buf  g262 (n270, n28);
buf  g263 (n399, n51);
buf  g264 (n180, n90);
buf  g265 (n181, n74);
buf  g266 (n314, n83);
buf  g267 (n198, n48);
not  g268 (n336, n22);
not  g269 (n354, n63);
not  g270 (n231, n96);
not  g271 (n305, n31);
buf  g272 (n332, n86);
not  g273 (n260, n27);
not  g274 (n112, n52);
buf  g275 (n302, n61);
buf  g276 (n119, n59);
not  g277 (n222, n42);
not  g278 (n132, n48);
buf  g279 (n177, n53);
not  g280 (n402, n98);
buf  g281 (n128, n22);
not  g282 (n233, n59);
buf  g283 (n117, n87);
not  g284 (n138, n22);
buf  g285 (n248, n80);
buf  g286 (n149, n24);
not  g287 (n156, n77);
buf  g288 (n141, n71);
buf  g289 (n163, n35);
buf  g290 (n316, n32);
buf  g291 (n311, n69);
not  g292 (n131, n94);
buf  g293 (n215, n100);
buf  g294 (n378, n95);
not  g295 (n338, n25);
not  g296 (n255, n65);
buf  g297 (n221, n34);
not  g298 (n269, n46);
not  g299 (n356, n46);
buf  g300 (n145, n69);
buf  g301 (n115, n79);
not  g302 (n310, n96);
not  g303 (n405, n23);
not  g304 (n246, n73);
not  g305 (n416, n36);
not  g306 (n287, n60);
not  g307 (n127, n91);
buf  g308 (n392, n36);
buf  g309 (n148, n70);
not  g310 (n120, n76);
not  g311 (n404, n56);
buf  g312 (n380, n69);
buf  g313 (n349, n39);
not  g314 (n390, n95);
not  g315 (n361, n81);
buf  g316 (n419, n94);
buf  g317 (n147, n73);
buf  g318 (n122, n95);
not  g319 (n261, n52);
buf  g320 (n282, n66);
buf  g321 (n279, n98);
not  g322 (n293, n87);
buf  g323 (n363, n90);
buf  g324 (n259, n47);
not  g325 (n391, n89);
not  g326 (n228, n78);
buf  g327 (n134, n61);
buf  g328 (n229, n74);
not  g329 (n401, n62);
buf  g330 (n152, n46);
not  g331 (n306, n68);
not  g332 (n262, n59);
buf  g333 (n327, n75);
buf  g334 (n345, n30);
not  g335 (n360, n88);
buf  g336 (n372, n77);
buf  g337 (n169, n55);
not  g338 (n139, n91);
not  g339 (n195, n63);
buf  g340 (n383, n72);
not  g341 (n297, n31);
buf  g342 (n265, n40);
not  g343 (n109, n84);
not  g344 (n237, n65);
buf  g345 (n320, n40);
buf  g346 (n275, n96);
not  g347 (n376, n41);
not  g348 (n254, n65);
not  g349 (n207, n30);
not  g350 (n357, n78);
buf  g351 (n196, n37);
not  g352 (n184, n80);
buf  g353 (n335, n71);
not  g354 (n118, n32);
not  g355 (n157, n75);
not  g356 (n413, n93);
not  g357 (n278, n62);
not  g358 (n408, n28);
buf  g359 (n359, n55);
not  g360 (n300, n54);
not  g361 (n396, n29);
buf  g362 (n208, n26);
buf  g363 (n185, n39);
buf  g364 (n142, n47);
not  g365 (n236, n79);
buf  g366 (n406, n28);
buf  g367 (n210, n98);
not  g368 (n106, n27);
buf  g369 (n135, n42);
not  g370 (n252, n65);
not  g371 (n130, n76);
not  g372 (n379, n72);
not  g373 (n187, n64);
buf  g374 (n267, n71);
not  g375 (n191, n63);
not  g376 (n330, n50);
buf  g377 (n313, n97);
buf  g378 (n150, n96);
not  g379 (n258, n42);
buf  g380 (n337, n54);
not  g381 (n189, n46);
buf  g382 (n381, n87);
not  g383 (n368, n30);
not  g384 (n411, n67);
not  g385 (n179, n55);
buf  g386 (n283, n93);
not  g387 (n315, n38);
buf  g388 (n250, n37);
buf  g389 (n203, n33);
not  g390 (n400, n81);
not  g391 (n199, n66);
buf  g392 (n322, n48);
not  g393 (n417, n78);
not  g394 (n244, n75);
not  g395 (n193, n84);
buf  g396 (n257, n70);
not  g397 (n183, n88);
buf  g398 (n350, n56);
buf  g399 (n321, n86);
buf  g400 (n682, n114);
not  g401 (n646, n112);
buf  g402 (n439, n362);
buf  g403 (n514, n334);
not  g404 (n571, n366);
not  g405 (n434, n354);
buf  g406 (n516, n167);
buf  g407 (n618, n388);
buf  g408 (n607, n341);
buf  g409 (n426, n138);
not  g410 (n648, n179);
buf  g411 (n495, n133);
not  g412 (n501, n202);
not  g413 (n531, n360);
not  g414 (n603, n140);
not  g415 (n544, n315);
not  g416 (n552, n261);
not  g417 (n471, n332);
buf  g418 (n521, n364);
not  g419 (n524, n207);
not  g420 (n649, n312);
buf  g421 (n468, n132);
buf  g422 (n507, n407);
not  g423 (n575, n178);
not  g424 (n678, n142);
not  g425 (n556, n397);
not  g426 (n609, n378);
not  g427 (n467, n347);
not  g428 (n481, n117);
not  g429 (n592, n295);
buf  g430 (n526, n335);
not  g431 (n657, n352);
not  g432 (n593, n344);
not  g433 (n611, n335);
not  g434 (n605, n181);
not  g435 (n587, n404);
not  g436 (n557, n369);
not  g437 (n632, n118);
not  g438 (n479, n240);
buf  g439 (n631, n330);
not  g440 (n606, n325);
buf  g441 (n596, n338);
buf  g442 (n643, n393);
buf  g443 (n687, n239);
buf  g444 (n652, n407);
buf  g445 (n469, n334);
not  g446 (n608, n283);
buf  g447 (n505, n213);
not  g448 (n542, n317);
not  g449 (n681, n353);
buf  g450 (n441, n122);
buf  g451 (n513, n245);
buf  g452 (n431, n287);
buf  g453 (n494, n298);
not  g454 (n500, n119);
buf  g455 (n625, n212);
not  g456 (n437, n136);
not  g457 (n663, n227);
buf  g458 (n601, n311);
not  g459 (n496, n199);
buf  g460 (n658, n339);
buf  g461 (n466, n147);
not  g462 (n474, n221);
not  g463 (n641, n351);
not  g464 (n644, n344);
not  g465 (n622, n350);
buf  g466 (n543, n129);
buf  g467 (n547, n375);
not  g468 (n538, n222);
not  g469 (n623, n346);
buf  g470 (n489, n231);
buf  g471 (n440, n347);
not  g472 (n511, n300);
buf  g473 (n655, n405);
not  g474 (n667, n110);
not  g475 (n512, n367);
buf  g476 (n450, n219);
buf  g477 (n560, n113);
buf  g478 (n662, n206);
not  g479 (n515, n277);
buf  g480 (n568, n236);
not  g481 (n503, n137);
buf  g482 (n435, n395);
not  g483 (n443, n337);
buf  g484 (n537, n196);
buf  g485 (n457, n190);
buf  g486 (n425, n338);
not  g487 (n533, n372);
not  g488 (n452, n187);
buf  g489 (n429, n220);
not  g490 (n616, n305);
not  g491 (n642, n125);
buf  g492 (n619, n402);
not  g493 (n665, n408);
not  g494 (n588, n280);
buf  g495 (n666, n378);
buf  g496 (n480, n210);
buf  g497 (n454, n390);
not  g498 (n430, n211);
buf  g499 (n630, n345);
buf  g500 (n580, n370);
buf  g501 (n549, n173);
buf  g502 (n576, n318);
buf  g503 (n462, n238);
not  g504 (n573, n352);
buf  g505 (n520, n184);
buf  g506 (n484, n276);
buf  g507 (n554, n158);
not  g508 (n647, n278);
not  g509 (n422, n313);
not  g510 (n566, n385);
buf  g511 (n614, n365);
not  g512 (n685, n349);
buf  g513 (n536, n169);
buf  g514 (n672, n356);
buf  g515 (n629, n229);
not  g516 (n659, n248);
not  g517 (n436, n265);
buf  g518 (n493, n328);
not  g519 (n651, n371);
not  g520 (n562, n194);
not  g521 (n669, n208);
buf  g522 (n519, n145);
buf  g523 (n530, n180);
not  g524 (n504, n403);
buf  g525 (n491, n291);
not  g526 (n639, n381);
buf  g527 (n578, n348);
not  g528 (n645, n148);
not  g529 (n428, n398);
not  g530 (n442, n364);
buf  g531 (n626, n242);
not  g532 (n445, n215);
not  g533 (n423, n201);
not  g534 (n463, n128);
not  g535 (n564, n124);
not  g536 (n595, n290);
not  g537 (n477, n127);
buf  g538 (n532, n406);
buf  g539 (n490, n392);
not  g540 (n502, n224);
not  g541 (n535, n324);
buf  g542 (n527, n348);
buf  g543 (n448, n108);
buf  g544 (n499, n374);
not  g545 (n460, n175);
buf  g546 (n584, n350);
not  g547 (n604, n320);
not  g548 (n598, n397);
not  g549 (n546, n268);
buf  g550 (n483, n170);
not  g551 (n541, n408);
not  g552 (n615, n337);
buf  g553 (n555, n304);
not  g554 (n599, n382);
not  g555 (n432, n342);
not  g556 (n508, n116);
buf  g557 (n633, n303);
not  g558 (n487, n259);
buf  g559 (n656, n256);
buf  g560 (n581, n131);
not  g561 (n600, n404);
buf  g562 (n677, n271);
not  g563 (n574, n356);
not  g564 (n563, n310);
buf  g565 (n680, n339);
not  g566 (n640, n216);
buf  g567 (n451, n361);
buf  g568 (n482, n177);
buf  g569 (n637, n323);
not  g570 (n497, n243);
buf  g571 (n558, n361);
buf  g572 (n638, n151);
not  g573 (n522, n359);
not  g574 (n438, n262);
not  g575 (n617, n385);
not  g576 (n540, n355);
not  g577 (n433, n260);
not  g578 (n528, n363);
not  g579 (n453, n376);
not  g580 (n449, n164);
buf  g581 (n594, n407);
buf  g582 (n679, n368);
not  g583 (n498, n139);
buf  g584 (n523, n284);
not  g585 (n661, n264);
buf  g586 (n675, n153);
buf  g587 (n613, n299);
not  g588 (n553, n327);
buf  g589 (n660, n154);
not  g590 (n488, n393);
buf  g591 (n534, n267);
buf  g592 (n591, n270);
not  g593 (n475, n343);
not  g594 (n473, n340);
buf  g595 (n458, n357);
buf  g596 (n634, n282);
buf  g597 (n561, n149);
buf  g598 (n650, n106);
buf  g599 (n654, n121);
buf  g600 (n465, n193);
buf  g601 (n670, n228);
buf  g602 (n628, n292);
buf  g603 (n559, n134);
not  g604 (n570, n297);
not  g605 (n674, n362);
not  g606 (n586, n165);
buf  g607 (n583, n186);
not  g608 (n673, n218);
not  g609 (n517, n203);
not  g610 (n492, n126);
not  g611 (n525, n109);
buf  g612 (n636, n322);
buf  g613 (n461, n189);
not  g614 (n518, n301);
buf  g615 (n621, n257);
buf  g616 (n459, n263);
buf  g617 (n565, n353);
buf  g618 (n550, n285);
buf  g619 (n486, n384);
not  g620 (n446, n369);
buf  g621 (n635, n402);
or   g622 (n620, n396, n253, n377, n269);
xor  g623 (n476, n326, n333, n401, n185);
or   g624 (n456, n281, n168, n143, n255);
and  g625 (n567, n400, n123, n373, n357);
xnor g626 (n470, n226, n409, n198, n365);
and  g627 (n551, n404, n174, n381, n246);
nand g628 (n447, n249, n374, n405, n368);
xnor g629 (n529, n192, n237, n341, n252);
nor  g630 (n506, n191, n359, n386, n406);
and  g631 (n539, n209, n273, n346, n157);
nand g632 (n624, n316, n195, n396, n391);
nand g633 (n590, n241, n244, n286, n409);
nand g634 (n653, n107, n384, n306, n399);
and  g635 (n577, n379, n161, n247, n403);
nor  g636 (n478, n115, n345, n389, n183);
or   g637 (n612, n225, n250, n205, n373);
nand g638 (n464, n266, n376, n160, n351);
xnor g639 (n548, n159, n336, n367, n370);
xnor g640 (n572, n355, n294, n156, n296);
nor  g641 (n676, n288, n400, n401, n223);
xnor g642 (n569, n146, n130, n171, n387);
xnor g643 (n427, n197, n204, n394, n354);
and  g644 (n668, n360, n407, n389, n398);
or   g645 (n683, n234, n233, n406, n387);
xnor g646 (n627, n319, n163, n141, n214);
xnor g647 (n545, n406, n403, n371, n358);
or   g648 (n585, n382, n399, n230, n342);
and  g649 (n424, n232, n386, n358, n380);
and  g650 (n510, n274, n377, n343, n172);
and  g651 (n472, n408, n314, n135, n394);
nand g652 (n610, n289, n402, n200, n308);
nor  g653 (n485, n144, n363, n176, n395);
xor  g654 (n455, n408, n120, n409, n279);
and  g655 (n579, n235, n182, n372, n392);
nand g656 (n444, n410, n272, n383, n150);
nor  g657 (n664, n340, n309, n275, n307);
nor  g658 (n686, n254, n403, n111, n258);
nor  g659 (n684, n333, n390, n366, n379);
and  g660 (n671, n321, n405, n383, n375);
xor  g661 (n582, n331, n388, n336, n293);
xor  g662 (n597, n405, n329, n409, n402);
xnor g663 (n509, n166, n188, n155, n380);
xnor g664 (n602, n162, n152, n302, n404);
nand g665 (n589, n217, n251, n391, n349);
not  g666 (n739, n437);
buf  g667 (n894, n563);
not  g668 (n831, n653);
not  g669 (n825, n453);
not  g670 (n784, n585);
not  g671 (n764, n657);
buf  g672 (n893, n481);
not  g673 (n719, n627);
buf  g674 (n800, n520);
not  g675 (n758, n608);
not  g676 (n720, n645);
not  g677 (n803, n440);
not  g678 (n850, n677);
not  g679 (n691, n681);
buf  g680 (n810, n517);
buf  g681 (n717, n503);
not  g682 (n716, n479);
buf  g683 (n703, n499);
buf  g684 (n834, n564);
not  g685 (n860, n508);
buf  g686 (n756, n589);
buf  g687 (n793, n626);
not  g688 (n752, n556);
not  g689 (n757, n471);
buf  g690 (n726, n594);
buf  g691 (n852, n560);
not  g692 (n744, n588);
not  g693 (n829, n436);
not  g694 (n796, n603);
not  g695 (n725, n493);
buf  g696 (n806, n612);
buf  g697 (n778, n635);
not  g698 (n724, n613);
buf  g699 (n817, n557);
not  g700 (n705, n485);
not  g701 (n730, n551);
buf  g702 (n813, n428);
buf  g703 (n842, n678);
not  g704 (n839, n680);
buf  g705 (n847, n624);
not  g706 (n741, n592);
buf  g707 (n708, n455);
buf  g708 (n878, n611);
buf  g709 (n690, n480);
not  g710 (n771, n649);
not  g711 (n801, n558);
buf  g712 (n820, n658);
buf  g713 (n743, n625);
not  g714 (n699, n682);
buf  g715 (n856, n675);
not  g716 (n869, n464);
buf  g717 (n854, n661);
not  g718 (n875, n559);
not  g719 (n688, n568);
not  g720 (n692, n526);
not  g721 (n713, n514);
not  g722 (n892, n476);
not  g723 (n866, n482);
not  g724 (n740, n561);
not  g725 (n823, n498);
buf  g726 (n824, n474);
not  g727 (n779, n430);
not  g728 (n762, n622);
buf  g729 (n853, n570);
buf  g730 (n870, n527);
not  g731 (n751, n667);
not  g732 (n765, n542);
not  g733 (n873, n660);
buf  g734 (n728, n549);
not  g735 (n867, n484);
not  g736 (n868, n576);
not  g737 (n738, n650);
buf  g738 (n855, n633);
buf  g739 (n807, n490);
buf  g740 (n750, n664);
buf  g741 (n763, n466);
buf  g742 (n710, n615);
buf  g743 (n812, n423);
buf  g744 (n837, n541);
buf  g745 (n818, n656);
not  g746 (n721, n492);
buf  g747 (n732, n593);
buf  g748 (n695, n602);
not  g749 (n693, n616);
not  g750 (n883, n426);
buf  g751 (n889, n652);
buf  g752 (n887, n583);
not  g753 (n698, n427);
not  g754 (n707, n506);
not  g755 (n845, n463);
buf  g756 (n706, n424);
buf  g757 (n736, n601);
buf  g758 (n787, n548);
not  g759 (n772, n491);
not  g760 (n742, n575);
not  g761 (n888, n504);
not  g762 (n773, n523);
buf  g763 (n872, n515);
not  g764 (n895, n665);
not  g765 (n841, n619);
not  g766 (n882, n647);
buf  g767 (n804, n473);
not  g768 (n737, n641);
not  g769 (n799, n441);
not  g770 (n766, n530);
not  g771 (n702, n555);
buf  g772 (n808, n571);
buf  g773 (n879, n552);
not  g774 (n770, n574);
not  g775 (n788, n553);
buf  g776 (n822, n509);
not  g777 (n722, n655);
buf  g778 (n826, n648);
not  g779 (n749, n569);
not  g780 (n715, n431);
not  g781 (n851, n606);
not  g782 (n733, n467);
buf  g783 (n783, n525);
not  g784 (n798, n511);
not  g785 (n760, n469);
not  g786 (n767, n489);
buf  g787 (n754, n435);
buf  g788 (n886, n600);
buf  g789 (n857, n605);
buf  g790 (n811, n590);
buf  g791 (n775, n434);
buf  g792 (n774, n634);
not  g793 (n761, n668);
not  g794 (n858, n477);
not  g795 (n880, n538);
buf  g796 (n846, n618);
not  g797 (n863, n629);
not  g798 (n838, n519);
not  g799 (n791, n572);
buf  g800 (n833, n614);
buf  g801 (n689, n544);
buf  g802 (n727, n443);
buf  g803 (n821, n659);
not  g804 (n797, n591);
buf  g805 (n802, n573);
not  g806 (n814, n598);
not  g807 (n753, n550);
buf  g808 (n694, n540);
not  g809 (n884, n518);
buf  g810 (n729, n512);
buf  g811 (n781, n654);
not  g812 (n792, n579);
buf  g813 (n769, n496);
not  g814 (n697, n566);
buf  g815 (n874, n513);
buf  g816 (n734, n584);
buf  g817 (n864, n596);
buf  g818 (n731, n529);
buf  g819 (n777, n522);
not  g820 (n861, n500);
buf  g821 (n890, n539);
buf  g822 (n789, n444);
buf  g823 (n723, n458);
not  g824 (n844, n617);
not  g825 (n832, n488);
not  g826 (n755, n537);
not  g827 (n881, n578);
buf  g828 (n805, n439);
not  g829 (n876, n432);
buf  g830 (n816, n676);
buf  g831 (n891, n679);
not  g832 (n840, n565);
buf  g833 (n711, n532);
not  g834 (n859, n586);
buf  g835 (n786, n638);
not  g836 (n848, n630);
not  g837 (n745, n483);
not  g838 (n849, n607);
not  g839 (n794, n448);
buf  g840 (n704, n599);
not  g841 (n843, n581);
not  g842 (n862, n609);
not  g843 (n835, n459);
not  g844 (n748, n632);
not  g845 (n700, n666);
not  g846 (n795, n545);
not  g847 (n759, n494);
not  g848 (n877, n644);
not  g849 (n776, n478);
buf  g850 (n701, n487);
not  g851 (n718, n639);
buf  g852 (n827, n495);
not  g853 (n782, n502);
not  g854 (n865, n623);
not  g855 (n696, n451);
nand g856 (n790, n580, n533, n673);
nand g857 (n746, n462, n636, n449, n468);
and  g858 (n809, n457, n642, n446, n567);
nand g859 (n735, n628, n456, n450, n442);
and  g860 (n815, n497, n597, n507, n587);
nand g861 (n836, n670, n640, n546, n547);
nand g862 (n768, n669, n674, n470, n554);
xor  g863 (n819, n643, n460, n528, n510);
and  g864 (n747, n663, n620, n662, n505);
xnor g865 (n780, n672, n433, n671, n425);
and  g866 (n714, n543, n534, n536, n637);
nor  g867 (n830, n465, n595, n631, n454);
nor  g868 (n709, n461, n472, n531, n429);
xor  g869 (n871, n452, n610, n438, n447);
xnor g870 (n885, n577, n524, n486, n475);
xnor g871 (n785, n535, n604, n445, n521);
nor  g872 (n712, n646, n516, n422, n501);
nand g873 (n828, n651, n621, n582, n562);
nor  g874 (n935, n800, n736, n755, n784);
and  g875 (n909, n803, n748, n706, n771);
and  g876 (n904, n761, n689, n747, n843);
nor  g877 (n903, n854, n715, n798, n769);
or   g878 (n921, n860, n815, n764, n704);
nor  g879 (n896, n775, n808, n794, n716);
and  g880 (n924, n714, n858, n745, n718);
xor  g881 (n912, n735, n719, n795, n778);
or   g882 (n906, n834, n836, n844, n780);
or   g883 (n913, n767, n851, n691, n862);
nand g884 (n930, n744, n773, n785, n741);
nand g885 (n937, n807, n845, n841, n731);
xor  g886 (n922, n738, n837, n753, n855);
and  g887 (n914, n824, n701, n853, n816);
nor  g888 (n899, n835, n768, n765, n840);
xnor g889 (n939, n712, n802, n713, n734);
and  g890 (n932, n789, n705, n825, n696);
nand g891 (n927, n781, n821, n856, n700);
or   g892 (n928, n758, n702, n693, n742);
nor  g893 (n925, n770, n833, n721, n805);
xnor g894 (n910, n838, n814, n711, n848);
nor  g895 (n915, n688, n810, n818, n850);
and  g896 (n918, n828, n766, n754, n760);
nor  g897 (n929, n697, n792, n827, n710);
or   g898 (n938, n722, n787, n732, n817);
or   g899 (n936, n774, n762, n757, n791);
xnor g900 (n908, n726, n857, n799, n729);
or   g901 (n900, n783, n699, n698, n786);
or   g902 (n917, n743, n777, n820, n782);
and  g903 (n919, n846, n752, n790, n852);
xnor g904 (n933, n695, n728, n859, n723);
nor  g905 (n916, n779, n806, n724, n819);
xnor g906 (n926, n831, n772, n708, n730);
nand g907 (n923, n826, n822, n717, n751);
xor  g908 (n920, n740, n739, n830, n813);
and  g909 (n902, n863, n788, n749, n793);
nand g910 (n905, n756, n750, n811, n759);
xor  g911 (n897, n709, n829, n804, n727);
xnor g912 (n931, n707, n849, n861, n832);
or   g913 (n898, n823, n703, n763, n733);
and  g914 (n901, n809, n776, n720, n801);
xor  g915 (n934, n737, n842, n847, n797);
or   g916 (n907, n694, n746, n812, n690);
xor  g917 (n911, n839, n796, n725, n692);
buf  g918 (n961, n930);
buf  g919 (n947, n936);
buf  g920 (n943, n931);
not  g921 (n951, n920);
not  g922 (n965, n925);
buf  g923 (n960, n913);
not  g924 (n950, n915);
buf  g925 (n955, n928);
buf  g926 (n958, n934);
buf  g927 (n956, n911);
buf  g928 (n967, n919);
not  g929 (n962, n912);
buf  g930 (n953, n922);
not  g931 (n964, n926);
not  g932 (n940, n937);
not  g933 (n945, n918);
buf  g934 (n948, n933);
not  g935 (n941, n932);
not  g936 (n963, n935);
buf  g937 (n944, n924);
buf  g938 (n952, n917);
buf  g939 (n942, n921);
buf  g940 (n966, n927);
not  g941 (n969, n929);
buf  g942 (n946, n938);
buf  g943 (n949, n914);
buf  g944 (n957, n923);
buf  g945 (n968, n939);
not  g946 (n959, n910);
not  g947 (n954, n916);
nand g948 (n973, n957, n940, n962);
and  g949 (n988, n957, n942, n959);
nand g950 (n985, n958, n966, n963, n954);
xnor g951 (n983, n954, n949, n941, n961);
or   g952 (n976, n949, n946, n944, n945);
xnor g953 (n981, n956, n941, n962, n964);
nand g954 (n977, n945, n952, n959);
or   g955 (n979, n945, n961, n949, n947);
or   g956 (n971, n964, n962, n963, n946);
xor  g957 (n978, n942, n948, n940);
nor  g958 (n974, n943, n955, n946);
nor  g959 (n996, n960, n956, n965, n944);
xor  g960 (n970, n963, n960, n948, n956);
and  g961 (n980, n954, n950, n960, n966);
or   g962 (n990, n951, n943, n940, n949);
nor  g963 (n989, n966, n958, n944, n947);
xor  g964 (n984, n946, n955, n943, n957);
xnor g965 (n992, n952, n950, n957, n948);
nor  g966 (n994, n953, n942, n951, n965);
or   g967 (n995, n960, n964, n963, n940);
nor  g968 (n986, n958, n953, n964, n961);
xor  g969 (n975, n944, n952, n953, n959);
nor  g970 (n982, n965, n941, n956, n951);
xnor g971 (n987, n953, n947, n955);
nand g972 (n993, n945, n943, n961, n941);
nand g973 (n991, n950, n962, n954, n958);
and  g974 (n972, n950, n951, n959, n965);
buf  g975 (n1008, n985);
buf  g976 (n1011, n980);
not  g977 (n999, n982);
buf  g978 (n998, n978);
not  g979 (n1002, n989);
not  g980 (n1009, n984);
not  g981 (n1000, n988);
not  g982 (n1015, n983);
not  g983 (n1003, n979);
buf  g984 (n997, n972);
buf  g985 (n1013, n976);
buf  g986 (n1005, n973);
not  g987 (n1006, n981);
buf  g988 (n1001, n986);
buf  g989 (n1014, n990);
not  g990 (n1007, n971);
buf  g991 (n1010, n977);
not  g992 (n1004, n975);
not  g993 (n1012, n987);
buf  g994 (n1016, n974);
buf  g995 (n1024, n866);
buf  g996 (n1040, n410);
buf  g997 (n1023, n1000);
not  g998 (n1022, n870);
or   g999 (n1030, n1000, n1004);
nor  g1000 (n1028, n1015, n1010, n969, n999);
or   g1001 (n1043, n1008, n1012, n1014);
nand g1002 (n1044, n999, n967, n968, n1002);
xor  g1003 (n1046, n998, n1005, n997, n1009);
nand g1004 (n1034, n1011, n1007, n867, n1010);
xor  g1005 (n1035, n968, n1008, n1000, n1005);
nand g1006 (n1021, n966, n1009, n1003, n871);
xor  g1007 (n1018, n1015, n967, n1001, n1012);
xnor g1008 (n1025, n969, n1003, n997, n998);
xor  g1009 (n1033, n410, n1005, n1015, n968);
or   g1010 (n1029, n872, n1004, n1003, n1001);
nor  g1011 (n1027, n1013, n1006, n998, n1004);
xor  g1012 (n1026, n1012, n969, n1007);
and  g1013 (n1041, n1012, n1013, n868, n869);
and  g1014 (n1031, n1014, n1003, n1002, n1016);
nand g1015 (n1038, n967, n873, n1002, n1001);
xor  g1016 (n1019, n864, n1011, n1016, n1010);
xor  g1017 (n1032, n969, n1006, n1016, n1015);
nand g1018 (n1045, n410, n1013, n1009, n1011);
nor  g1019 (n1036, n999, n1014, n1013, n1008);
xnor g1020 (n1039, n1000, n1005, n1009, n967);
or   g1021 (n1020, n997, n999, n1010, n1011);
and  g1022 (n1037, n1002, n1016, n1004, n1008);
xnor g1023 (n1042, n997, n998, n1006, n968);
and  g1024 (n1017, n865, n1006, n1007, n1001);
not  g1025 (n1050, n1034);
not  g1026 (n1047, n1031);
not  g1027 (n1048, n1033);
buf  g1028 (n1049, n1032);
nor  g1029 (n1056, n104, n1041);
nand g1030 (n1051, n1047, n883);
xnor g1031 (n1057, n1049, n1047, n1050, n1036);
or   g1032 (n1064, n1040, n101, n1048, n686);
nor  g1033 (n1058, n1049, n102, n1050, n685);
xor  g1034 (n1055, n875, n887, n411, n1049);
nor  g1035 (n1052, n102, n411, n1047, n877);
nor  g1036 (n1060, n411, n879, n885, n683);
nand g1037 (n1054, n103, n684, n411, n1049);
or   g1038 (n1063, n101, n1048, n1039, n1050);
and  g1039 (n1053, n876, n882, n101, n103);
nor  g1040 (n1066, n1035, n102, n888, n880);
or   g1041 (n1065, n881, n884, n874, n878);
and  g1042 (n1059, n103, n412, n1050, n886);
and  g1043 (n1061, n1038, n1037, n102, n101);
xnor g1044 (n1062, n1048, n1048, n103, n1047);
not  g1045 (n1081, n1054);
buf  g1046 (n1072, n1056);
not  g1047 (n1068, n1057);
not  g1048 (n1080, n1060);
not  g1049 (n1071, n1061);
buf  g1050 (n1074, n1053);
buf  g1051 (n1085, n1058);
not  g1052 (n1067, n1063);
not  g1053 (n1078, n1058);
buf  g1054 (n1083, n1061);
not  g1055 (n1070, n1057);
not  g1056 (n1069, n1060);
not  g1057 (n1075, n1062);
not  g1058 (n1084, n1059);
not  g1059 (n1077, n1052);
buf  g1060 (n1082, n1062);
buf  g1061 (n1073, n1055);
buf  g1062 (n1076, n1051);
not  g1063 (n1079, n1059);
buf  g1064 (n1086, n1056);
not  g1065 (n1141, n1074);
not  g1066 (n1126, n1083);
buf  g1067 (n1107, n1068);
not  g1068 (n1145, n1075);
not  g1069 (n1101, n1072);
buf  g1070 (n1096, n1082);
not  g1071 (n1124, n1086);
buf  g1072 (n1116, n1071);
not  g1073 (n1132, n1077);
buf  g1074 (n1114, n415);
buf  g1075 (n1148, n1074);
buf  g1076 (n1098, n415);
buf  g1077 (n1106, n1076);
not  g1078 (n1146, n412);
not  g1079 (n1117, n1086);
not  g1080 (n1122, n1069);
buf  g1081 (n1092, n1076);
not  g1082 (n1120, n1073);
buf  g1083 (n1139, n1067);
not  g1084 (n1108, n1071);
not  g1085 (n1129, n1080);
not  g1086 (n1094, n1069);
buf  g1087 (n1089, n1085);
not  g1088 (n1112, n416);
not  g1089 (n1093, n1083);
buf  g1090 (n1128, n413);
buf  g1091 (n1118, n1071);
not  g1092 (n1109, n412);
not  g1093 (n1138, n1068);
buf  g1094 (n1097, n1073);
buf  g1095 (n1123, n414);
not  g1096 (n1100, n1072);
not  g1097 (n1090, n412);
not  g1098 (n1111, n417);
buf  g1099 (n1125, n1075);
buf  g1100 (n1091, n1084);
buf  g1101 (n1147, n1068);
not  g1102 (n1102, n1067);
not  g1103 (n1143, n1078);
buf  g1104 (n1113, n1079);
not  g1105 (n1144, n1085);
buf  g1106 (n1119, n1082);
buf  g1107 (n1133, n415);
not  g1108 (n1136, n413);
not  g1109 (n1121, n418);
buf  g1110 (n1115, n1067);
buf  g1111 (n1137, n418);
xnor g1112 (n1095, n1069, n1072);
nor  g1113 (n1131, n1082, n1069, n1075);
nand g1114 (n1142, n1068, n1079, n1083, n1080);
or   g1115 (n1105, n1079, n413, n1081, n1073);
xor  g1116 (n1140, n1070, n1070, n1076, n414);
xnor g1117 (n1088, n1085, n417, n1074);
and  g1118 (n1087, n1083, n1085, n1073, n1077);
or   g1119 (n1134, n1067, n416, n1072, n1078);
xnor g1120 (n1103, n414, n1084, n1077, n415);
and  g1121 (n1099, n1071, n1078, n1082);
nand g1122 (n1127, n1086, n1074, n1081, n1080);
or   g1123 (n1104, n416, n416, n417, n1086);
and  g1124 (n1110, n1080, n1070, n1076, n1084);
xor  g1125 (n1130, n413, n1077, n1079, n1070);
nor  g1126 (n1135, n1084, n414, n1081);
buf  g1127 (n1169, n1138);
not  g1128 (n1192, n1112);
buf  g1129 (n1150, n1145);
not  g1130 (n1202, n1105);
not  g1131 (n1196, n1132);
buf  g1132 (n1171, n1100);
buf  g1133 (n1176, n1107);
buf  g1134 (n1182, n1130);
not  g1135 (n1164, n1134);
buf  g1136 (n1149, n1123);
buf  g1137 (n1205, n1110);
not  g1138 (n1201, n1122);
not  g1139 (n1179, n1115);
not  g1140 (n1186, n1101);
buf  g1141 (n1191, n1140);
buf  g1142 (n1190, n1090);
buf  g1143 (n1188, n1094);
buf  g1144 (n1154, n1088);
buf  g1145 (n1168, n1095);
not  g1146 (n1194, n1091);
buf  g1147 (n1181, n1103);
not  g1148 (n1199, n1127);
not  g1149 (n1174, n1124);
buf  g1150 (n1200, n1135);
not  g1151 (n1156, n1116);
buf  g1152 (n1189, n1125);
not  g1153 (n1184, n1108);
buf  g1154 (n1153, n1133);
not  g1155 (n1152, n1137);
not  g1156 (n1162, n1121);
not  g1157 (n1204, n1129);
not  g1158 (n1187, n1114);
buf  g1159 (n1163, n1099);
buf  g1160 (n1173, n1144);
not  g1161 (n1151, n1126);
not  g1162 (n1177, n1141);
not  g1163 (n1207, n1111);
buf  g1164 (n1157, n1136);
buf  g1165 (n1208, n1089);
not  g1166 (n1158, n1120);
buf  g1167 (n1165, n1131);
not  g1168 (n1180, n1128);
not  g1169 (n1195, n1102);
not  g1170 (n1193, n1097);
buf  g1171 (n1159, n1139);
not  g1172 (n1197, n1109);
buf  g1173 (n1161, n1098);
buf  g1174 (n1203, n1087);
buf  g1175 (n1185, n1146);
buf  g1176 (n1170, n1093);
buf  g1177 (n1166, n1142);
not  g1178 (n1183, n1092);
buf  g1179 (n1167, n1118);
buf  g1180 (n1206, n1119);
buf  g1181 (n1178, n1096);
buf  g1182 (n1155, n1143);
buf  g1183 (n1172, n1106);
buf  g1184 (n1160, n1113);
buf  g1185 (n1198, n1104);
buf  g1186 (n1175, n1117);
not  g1187 (n1317, n1164);
buf  g1188 (n1255, n1184);
buf  g1189 (n1220, n1156);
buf  g1190 (n1313, n1185);
buf  g1191 (n1318, n1160);
buf  g1192 (n1242, n1203);
buf  g1193 (n1229, n1180);
not  g1194 (n1214, n1201);
not  g1195 (n1291, n1198);
not  g1196 (n1305, n1189);
buf  g1197 (n1278, n1176);
not  g1198 (n1212, n1159);
not  g1199 (n1267, n1168);
not  g1200 (n1233, n1167);
buf  g1201 (n1259, n1178);
not  g1202 (n1222, n1183);
buf  g1203 (n1323, n1154);
not  g1204 (n1262, n1191);
buf  g1205 (n1271, n1181);
not  g1206 (n1249, n1174);
not  g1207 (n1269, n1163);
not  g1208 (n1321, n1206);
buf  g1209 (n1211, n1169);
buf  g1210 (n1247, n1174);
not  g1211 (n1314, n1188);
not  g1212 (n1244, n1165);
not  g1213 (n1284, n1173);
not  g1214 (n1260, n1157);
not  g1215 (n1251, n1184);
not  g1216 (n1275, n1179);
not  g1217 (n1258, n1197);
buf  g1218 (n1307, n1169);
not  g1219 (n1236, n1149);
buf  g1220 (n1300, n1197);
not  g1221 (n1218, n1200);
buf  g1222 (n1293, n1173);
not  g1223 (n1315, n1154);
not  g1224 (n1235, n1168);
buf  g1225 (n1266, n1195);
buf  g1226 (n1243, n1205);
buf  g1227 (n1324, n1165);
buf  g1228 (n1209, n1155);
not  g1229 (n1253, n1201);
buf  g1230 (n1219, n1173);
not  g1231 (n1295, n1152);
not  g1232 (n1273, n1200);
not  g1233 (n1282, n1200);
buf  g1234 (n1292, n1180);
not  g1235 (n1246, n1178);
not  g1236 (n1263, n1199);
buf  g1237 (n1250, n1205);
not  g1238 (n1264, n1181);
buf  g1239 (n1304, n1162);
buf  g1240 (n1277, n1188);
buf  g1241 (n1234, n1180);
buf  g1242 (n1289, n1156);
not  g1243 (n1215, n1208);
not  g1244 (n1257, n1203);
buf  g1245 (n1268, n1151);
not  g1246 (n1241, n1171);
not  g1247 (n1316, n1149);
not  g1248 (n1281, n418);
not  g1249 (n1224, n1187);
buf  g1250 (n1302, n1179);
not  g1251 (n1221, n1162);
buf  g1252 (n1311, n1167);
not  g1253 (n1279, n1190);
not  g1254 (n1276, n1191);
not  g1255 (n1294, n1204);
buf  g1256 (n1238, n1176);
buf  g1257 (n1310, n1192);
not  g1258 (n1240, n1158);
buf  g1259 (n1227, n1161);
nor  g1260 (n1237, n1194, n1199, n1190);
xnor g1261 (n1290, n1206, n1159, n1150);
xnor g1262 (n1239, n1194, n1185, n1206, n1178);
and  g1263 (n1245, n1158, n1203, n1166, n1202);
xor  g1264 (n1231, n1157, n1170, n1180, n1169);
xor  g1265 (n1256, n1205, n1155);
xor  g1266 (n1312, n1201, n1175, n1157, n1163);
nand g1267 (n1223, n1196, n1177, n1161, n1159);
xnor g1268 (n1248, n1195, n1187, n1189, n1163);
nand g1269 (n1297, n1169, n1176, n1196, n1170);
nand g1270 (n1225, n1153, n1164, n1171, n1162);
or   g1271 (n1287, n1160, n1193, n1207, n1189);
nor  g1272 (n1283, n1158, n1182, n1175, n1152);
or   g1273 (n1274, n1186, n1183, n1198, n1154);
xor  g1274 (n1301, n1176, n1198, n1193, n1202);
or   g1275 (n1226, n1192, n1188, n1195, n1205);
nand g1276 (n1217, n1191, n1183, n1192, n1200);
xnor g1277 (n1272, n1182, n1192, n1202, n1152);
nor  g1278 (n1296, n1163, n1197, n1153, n1151);
xnor g1279 (n1320, n1153, n1177, n1170, n1171);
or   g1280 (n1252, n1161, n1181, n1167, n1195);
or   g1281 (n1308, n1168, n1158, n1204, n1165);
and  g1282 (n1213, n1194, n1043, n1156, n1166);
nor  g1283 (n1298, n1193, n1149, n1164, n1194);
nand g1284 (n1280, n1154, n1208, n1150, n1185);
nand g1285 (n1288, n1172, n1202, n1177, n1042);
or   g1286 (n1306, n1190, n1207, n1181, n1178);
xnor g1287 (n1210, n1208, n1166, n1150, n1186);
xor  g1288 (n1309, n1183, n1201, n1177, n1149);
xnor g1289 (n1228, n1164, n1167, n1208, n1184);
or   g1290 (n1286, n1151, n1193, n1196, n1153);
xnor g1291 (n1216, n1157, n1199, n1151, n1159);
xor  g1292 (n1261, n1171, n1182, n1203, n1168);
nand g1293 (n1322, n1161, n1173, n1197, n1172);
xnor g1294 (n1285, n1206, n1152, n1190, n1175);
or   g1295 (n1254, n1198, n1182, n1187, n1207);
nor  g1296 (n1232, n1185, n1170, n1188, n1160);
nor  g1297 (n1265, n1150, n1184, n1175, n1199);
nand g1298 (n1270, n1172, n1174, n1187, n1186);
nor  g1299 (n1230, n1186, n1207, n1166, n1156);
or   g1300 (n1319, n1165, n1189, n1204, n1172);
nand g1301 (n1303, n1179, n1174, n1191, n1204);
or   g1302 (n1299, n1179, n1160, n1196, n1162);
xor  g1303 (n1340, n1299, n1296, n1267, n1227);
xor  g1304 (n1345, n1271, n1266, n1255, n1246);
xor  g1305 (n1343, n1286, n1279, n1215, n1234);
xor  g1306 (n1346, n1218, n1213, n1256, n1211);
and  g1307 (n1325, n1217, n1250, n1239, n1241);
nand g1308 (n1337, n1275, n1298, n1238, n1225);
and  g1309 (n1328, n1210, n1281, n1285, n1291);
xor  g1310 (n1332, n1287, n1315, n1223, n1252);
xnor g1311 (n1347, n1236, n1214, n1249, n1282);
or   g1312 (n1351, n1297, n1314, n1309, n1243);
nand g1313 (n1327, n1306, n1212, n1226, n1219);
xnor g1314 (n1334, n1284, n1277, n1251, n1295);
xnor g1315 (n1336, n1235, n1294, n1244, n1240);
nor  g1316 (n1342, n1216, n1272, n1248, n1224);
or   g1317 (n1341, n1289, n1293, n1230, n1312);
nor  g1318 (n1335, n1245, n1260, n1262, n1247);
or   g1319 (n1349, n1242, n1237, n1263, n1276);
nor  g1320 (n1348, n1253, n1283, n1232, n1310);
and  g1321 (n1338, n1261, n1264, n1292, n1270);
and  g1322 (n1326, n1313, n1302, n1233, n1273);
and  g1323 (n1330, n1274, n1278, n1268, n1316);
and  g1324 (n1329, n1259, n1280, n1308, n1228);
xor  g1325 (n1339, n1305, n1258, n1222, n1231);
xnor g1326 (n1350, n1269, n1311, n1301, n1304);
xnor g1327 (n1331, n1257, n1221, n1209, n1220);
xor  g1328 (n1344, n1303, n1265, n1290, n1307);
nand g1329 (n1333, n1254, n1300, n1288, n1229);
not  g1330 (n1353, n1319);
buf  g1331 (n1367, n1336);
buf  g1332 (n1371, n1330);
buf  g1333 (n1355, n1064);
not  g1334 (n1362, n1326);
not  g1335 (n1373, n1147);
buf  g1336 (n1365, n1351);
not  g1337 (n1352, n1344);
not  g1338 (n1359, n1338);
not  g1339 (n1358, n1340);
buf  g1340 (n1366, n1318);
not  g1341 (n1368, n1335);
not  g1342 (n1372, n894);
not  g1343 (n1363, n1348);
nand g1344 (n1377, n1064, n1349);
xnor g1345 (n1354, n1347, n1317, n895, n418);
xor  g1346 (n1357, n1339, n1334, n1350, n1065);
and  g1347 (n1356, n1321, n1343, n891, n1341);
xor  g1348 (n1376, n1324, n1327, n893, n1066);
xnor g1349 (n1370, n1331, n1346, n1322, n996);
xnor g1350 (n1364, n1045, n687, n889, n1342);
and  g1351 (n1369, n890, n1044, n1320, n1066);
xnor g1352 (n1361, n992, n993, n995, n1332);
xnor g1353 (n1374, n1329, n1333, n1328, n892);
xnor g1354 (n1375, n1046, n1323, n1337, n1065);
nor  g1355 (n1360, n991, n1063, n994, n1345);
nand g1356 (n1379, n1358, n1373, n1377, n1356);
nand g1357 (n1383, n1355, n1360, n1371, n1369);
and  g1358 (n1380, n1366, n1365, n1359, n1357);
or   g1359 (n1387, n1368, n1376, n1358);
xor  g1360 (n1381, n1359, n1364, n1369, n1372);
xor  g1361 (n1386, n1360, n1354, n1352, n1363);
nand g1362 (n1388, n1362, n1373, n1364, n1365);
or   g1363 (n1382, n1368, n1377, n1363, n1361);
nor  g1364 (n1389, n1367, n1370, n1371, n1374);
nor  g1365 (n1384, n1372, n1366, n1367, n1357);
and  g1366 (n1378, n1362, n1374, n1370, n1361);
nor  g1367 (n1385, n1353, n1375, n419);
xor  g1368 (n1390, n1148, n1389);
nand g1369 (n1392, n105, n105, n104, n1390);
and  g1370 (n1391, n1390, n104, n105);
xor  g1371 (n1394, n420, n1392, n421);
xnor g1372 (n1393, n419, n105, n421, n420);
or   g1373 (n1396, n420, n1391);
nor  g1374 (n1395, n419, n419, n1392, n421);
endmodule
