

module Stat_1664_71_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n1356,
  n1348,
  n1346,
  n1350,
  n1353,
  n1354,
  n1345,
  n1349,
  n1667,
  n1670,
  n1662,
  n1663,
  n1664,
  n1668,
  n1671,
  n1665,
  n1672,
  n1669,
  n1684,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1356;output n1348;output n1346;output n1350;output n1353;output n1354;output n1345;output n1349;output n1667;output n1670;output n1662;output n1663;output n1664;output n1668;output n1671;output n1665;output n1672;output n1669;output n1684;
  wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1347;wire n1351;wire n1352;wire n1355;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1666;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  buf
  g0
  (
    n34,
    n6
  );


  buf
  g1
  (
    n25,
    n7
  );


  buf
  g2
  (
    n30,
    n1
  );


  not
  g3
  (
    n40,
    n5
  );


  buf
  g4
  (
    n27,
    n7
  );


  not
  g5
  (
    n28,
    n3
  );


  buf
  g6
  (
    n31,
    n8
  );


  not
  g7
  (
    n42,
    n9
  );


  not
  g8
  (
    n29,
    n7
  );


  not
  g9
  (
    n43,
    n3
  );


  buf
  g10
  (
    n22,
    n1
  );


  buf
  g11
  (
    n23,
    n6
  );


  not
  g12
  (
    n32,
    n5
  );


  buf
  g13
  (
    n35,
    n1
  );


  buf
  g14
  (
    n36,
    n7
  );


  nand
  g15
  (
    n37,
    n1,
    n4
  );


  and
  g16
  (
    n39,
    n6,
    n8
  );


  and
  g17
  (
    n24,
    n5,
    n8
  );


  xor
  g18
  (
    n44,
    n3,
    n4
  );


  buf
  g19
  (
    n38,
    n2
  );


  and
  g20
  (
    n21,
    n4,
    n2
  );


  xor
  g21
  (
    n26,
    n4,
    n6
  );


  and
  g22
  (
    n33,
    n8,
    n3
  );


  nand
  g23
  (
    n41,
    n2,
    n5
  );


  buf
  g24
  (
    n50,
    n22
  );


  not
  g25
  (
    n54,
    n21
  );


  not
  g26
  (
    n53,
    n22
  );


  not
  g27
  (
    n49,
    n22
  );


  not
  g28
  (
    n46,
    n21
  );


  buf
  g29
  (
    n45,
    n22
  );


  buf
  g30
  (
    n48,
    n23
  );


  buf
  g31
  (
    n51,
    n21
  );


  not
  g32
  (
    KeyWire_0_15,
    n23
  );


  buf
  g33
  (
    n47,
    n21
  );


  not
  g34
  (
    n57,
    n45
  );


  not
  g35
  (
    n61,
    n45
  );


  not
  g36
  (
    n58,
    n46
  );


  buf
  g37
  (
    n64,
    n46
  );


  not
  g38
  (
    n65,
    n46
  );


  buf
  g39
  (
    n59,
    n47
  );


  not
  g40
  (
    n55,
    n45
  );


  buf
  g41
  (
    n56,
    n45
  );


  buf
  g42
  (
    n63,
    n47
  );


  buf
  g43
  (
    n60,
    n47
  );


  buf
  g44
  (
    n66,
    n46
  );


  buf
  g45
  (
    n62,
    n47
  );


  buf
  g46
  (
    n102,
    n26
  );


  buf
  g47
  (
    n93,
    n26
  );


  not
  g48
  (
    n67,
    n65
  );


  not
  g49
  (
    KeyWire_0_28,
    n27
  );


  not
  g50
  (
    n86,
    n35
  );


  not
  g51
  (
    n76,
    n24
  );


  not
  g52
  (
    n74,
    n24
  );


  not
  g53
  (
    n105,
    n28
  );


  not
  g54
  (
    n72,
    n62
  );


  not
  g55
  (
    n99,
    n23
  );


  buf
  g56
  (
    n87,
    n64
  );


  not
  g57
  (
    n84,
    n60
  );


  not
  g58
  (
    n96,
    n60
  );


  buf
  g59
  (
    n94,
    n27
  );


  not
  g60
  (
    n68,
    n40
  );


  buf
  g61
  (
    KeyWire_0_10,
    n34
  );


  buf
  g62
  (
    n104,
    n62
  );


  buf
  g63
  (
    n100,
    n58
  );


  not
  g64
  (
    n75,
    n31
  );


  not
  g65
  (
    n82,
    n40
  );


  not
  g66
  (
    n73,
    n30
  );


  buf
  g67
  (
    n107,
    n59
  );


  xnor
  g68
  (
    n83,
    n30,
    n32
  );


  xor
  g69
  (
    n108,
    n25,
    n65,
    n60,
    n33
  );


  or
  g70
  (
    n113,
    n35,
    n61,
    n60,
    n37
  );


  or
  g71
  (
    n110,
    n31,
    n34,
    n32,
    n37
  );


  nand
  g72
  (
    n89,
    n57,
    n39,
    n66,
    n29
  );


  nor
  g73
  (
    n98,
    n30,
    n38,
    n57,
    n35
  );


  and
  g74
  (
    n103,
    n35,
    n31,
    n28,
    n24
  );


  nand
  g75
  (
    n79,
    n25,
    n39,
    n27,
    n34
  );


  nor
  g76
  (
    n95,
    n26,
    n58,
    n36,
    n40
  );


  nor
  g77
  (
    n85,
    n63,
    n64,
    n32
  );


  nand
  g78
  (
    n101,
    n34,
    n62,
    n55
  );


  nor
  g79
  (
    n88,
    n40,
    n55,
    n36
  );


  nand
  g80
  (
    n91,
    n59,
    n29,
    n56,
    n30
  );


  nand
  g81
  (
    n109,
    n39,
    n61,
    n27,
    n38
  );


  or
  g82
  (
    n106,
    n65,
    n23,
    n33,
    n38
  );


  and
  g83
  (
    n71,
    n63,
    n66,
    n55,
    n29
  );


  and
  g84
  (
    n70,
    n41,
    n41,
    n32,
    n59
  );


  xnor
  g85
  (
    n81,
    n29,
    n28,
    n64,
    n56
  );


  nand
  g86
  (
    n97,
    n24,
    n26,
    n61
  );


  and
  g87
  (
    n92,
    n28,
    n59,
    n63,
    n37
  );


  nand
  g88
  (
    n69,
    n36,
    n56,
    n31,
    n33
  );


  nand
  g89
  (
    n112,
    n36,
    n39,
    n33,
    n25
  );


  and
  g90
  (
    n111,
    n56,
    n63,
    n66,
    n37
  );


  or
  g91
  (
    n80,
    n25,
    n57,
    n58
  );


  and
  g92
  (
    n90,
    n65,
    n58,
    n38,
    n66
  );


  not
  g93
  (
    n119,
    n81
  );


  buf
  g94
  (
    n162,
    n75
  );


  buf
  g95
  (
    n143,
    n77
  );


  buf
  g96
  (
    n134,
    n82
  );


  not
  g97
  (
    n177,
    n83
  );


  not
  g98
  (
    n188,
    n74
  );


  buf
  g99
  (
    n147,
    n68
  );


  not
  g100
  (
    n153,
    n86
  );


  not
  g101
  (
    n172,
    n85
  );


  buf
  g102
  (
    n199,
    n87
  );


  not
  g103
  (
    n137,
    n81
  );


  buf
  g104
  (
    n174,
    n71
  );


  not
  g105
  (
    n123,
    n71
  );


  not
  g106
  (
    n168,
    n76
  );


  not
  g107
  (
    n132,
    n70
  );


  buf
  g108
  (
    n175,
    n79
  );


  not
  g109
  (
    n193,
    n72
  );


  buf
  g110
  (
    n133,
    n84
  );


  buf
  g111
  (
    n186,
    n76
  );


  buf
  g112
  (
    n176,
    n72
  );


  buf
  g113
  (
    n166,
    n80
  );


  not
  g114
  (
    n131,
    n74
  );


  buf
  g115
  (
    n192,
    n73
  );


  buf
  g116
  (
    n144,
    n79
  );


  not
  g117
  (
    n122,
    n87
  );


  not
  g118
  (
    n126,
    n84
  );


  not
  g119
  (
    n115,
    n81
  );


  buf
  g120
  (
    n169,
    n81
  );


  not
  g121
  (
    n142,
    n67
  );


  not
  g122
  (
    n165,
    n83
  );


  buf
  g123
  (
    n150,
    n69
  );


  buf
  g124
  (
    n130,
    n70
  );


  not
  g125
  (
    n163,
    n69
  );


  buf
  g126
  (
    n159,
    n77
  );


  not
  g127
  (
    n141,
    n80
  );


  buf
  g128
  (
    n161,
    n73
  );


  not
  g129
  (
    n197,
    n80
  );


  buf
  g130
  (
    n185,
    n71
  );


  buf
  g131
  (
    n183,
    n77
  );


  not
  g132
  (
    n195,
    n87
  );


  not
  g133
  (
    KeyWire_0_3,
    n67
  );


  buf
  g134
  (
    n151,
    n86
  );


  buf
  g135
  (
    n149,
    n80
  );


  not
  g136
  (
    n120,
    n68
  );


  not
  g137
  (
    n191,
    n70
  );


  buf
  g138
  (
    n158,
    n75
  );


  not
  g139
  (
    n124,
    n70
  );


  not
  g140
  (
    n154,
    n84
  );


  buf
  g141
  (
    n114,
    n78
  );


  buf
  g142
  (
    n116,
    n79
  );


  not
  g143
  (
    n184,
    n82
  );


  not
  g144
  (
    n152,
    n82
  );


  buf
  g145
  (
    n139,
    n85
  );


  not
  g146
  (
    n187,
    n86
  );


  buf
  g147
  (
    n117,
    n78
  );


  buf
  g148
  (
    n125,
    n79
  );


  buf
  g149
  (
    n189,
    n86
  );


  not
  g150
  (
    n138,
    n85
  );


  not
  g151
  (
    n118,
    n69
  );


  not
  g152
  (
    n160,
    n69
  );


  not
  g153
  (
    n171,
    n68
  );


  not
  g154
  (
    n140,
    n82
  );


  buf
  g155
  (
    n190,
    n74
  );


  buf
  g156
  (
    n194,
    n73
  );


  buf
  g157
  (
    n129,
    n88
  );


  buf
  g158
  (
    n128,
    n83
  );


  buf
  g159
  (
    n145,
    n84
  );


  not
  g160
  (
    n198,
    n87
  );


  buf
  g161
  (
    n167,
    n88
  );


  buf
  g162
  (
    n121,
    n76
  );


  buf
  g163
  (
    n157,
    n77
  );


  not
  g164
  (
    n155,
    n78
  );


  not
  g165
  (
    n170,
    n83
  );


  buf
  g166
  (
    n182,
    n67
  );


  buf
  g167
  (
    n146,
    n78
  );


  not
  g168
  (
    n178,
    n74
  );


  buf
  g169
  (
    n196,
    n67
  );


  buf
  g170
  (
    n148,
    n76
  );


  buf
  g171
  (
    n127,
    n75
  );


  buf
  g172
  (
    n173,
    n73
  );


  buf
  g173
  (
    n164,
    n85
  );


  not
  g174
  (
    n179,
    n72
  );


  buf
  g175
  (
    n180,
    n75
  );


  not
  g176
  (
    n156,
    n72
  );


  buf
  g177
  (
    n181,
    n68
  );


  not
  g178
  (
    n136,
    n71
  );


  buf
  g179
  (
    n224,
    n115
  );


  not
  g180
  (
    n241,
    n118
  );


  buf
  g181
  (
    n229,
    n123
  );


  not
  g182
  (
    n244,
    n120
  );


  buf
  g183
  (
    n230,
    n118
  );


  not
  g184
  (
    n213,
    n121
  );


  buf
  g185
  (
    n211,
    n116
  );


  buf
  g186
  (
    n219,
    n125
  );


  not
  g187
  (
    n248,
    n125
  );


  not
  g188
  (
    n220,
    n117
  );


  not
  g189
  (
    n239,
    n126
  );


  buf
  g190
  (
    n215,
    n115
  );


  not
  g191
  (
    n223,
    n116
  );


  buf
  g192
  (
    n249,
    n122
  );


  buf
  g193
  (
    n206,
    n119
  );


  not
  g194
  (
    n242,
    n122
  );


  not
  g195
  (
    n210,
    n127
  );


  buf
  g196
  (
    n237,
    n127
  );


  not
  g197
  (
    n225,
    n123
  );


  buf
  g198
  (
    n204,
    n114
  );


  buf
  g199
  (
    n201,
    n122
  );


  buf
  g200
  (
    n233,
    n126
  );


  not
  g201
  (
    n222,
    n117
  );


  buf
  g202
  (
    n207,
    n114
  );


  not
  g203
  (
    n203,
    n127
  );


  buf
  g204
  (
    n231,
    n124
  );


  buf
  g205
  (
    n235,
    n120
  );


  buf
  g206
  (
    n226,
    n114
  );


  buf
  g207
  (
    n232,
    n124
  );


  not
  g208
  (
    n236,
    n121
  );


  buf
  g209
  (
    n247,
    n122
  );


  buf
  g210
  (
    n227,
    n124
  );


  not
  g211
  (
    n208,
    n124
  );


  not
  g212
  (
    n214,
    n123
  );


  not
  g213
  (
    n209,
    n123
  );


  buf
  g214
  (
    n205,
    n120
  );


  not
  g215
  (
    n245,
    n127
  );


  buf
  g216
  (
    n221,
    n114
  );


  buf
  g217
  (
    n228,
    n115
  );


  not
  g218
  (
    n202,
    n119
  );


  buf
  g219
  (
    n238,
    n116
  );


  buf
  g220
  (
    n216,
    n120
  );


  not
  g221
  (
    n240,
    n126
  );


  not
  g222
  (
    n217,
    n117
  );


  not
  g223
  (
    n243,
    n116
  );


  not
  g224
  (
    n212,
    n119
  );


  buf
  g225
  (
    n246,
    n115
  );


  buf
  g226
  (
    n234,
    n119
  );


  nor
  g227
  (
    n218,
    n125,
    n126,
    n117,
    n118
  );


  or
  g228
  (
    n200,
    n118,
    n121,
    n125
  );


  not
  g229
  (
    n251,
    n226
  );


  not
  g230
  (
    n304,
    n245
  );


  buf
  g231
  (
    n278,
    n232
  );


  not
  g232
  (
    n281,
    n215
  );


  buf
  g233
  (
    n264,
    n229
  );


  buf
  g234
  (
    n311,
    n222
  );


  buf
  g235
  (
    n254,
    n241
  );


  buf
  g236
  (
    n293,
    n247
  );


  not
  g237
  (
    n328,
    n202
  );


  buf
  g238
  (
    n290,
    n229
  );


  buf
  g239
  (
    n283,
    n240
  );


  buf
  g240
  (
    n268,
    n219
  );


  buf
  g241
  (
    n310,
    n204
  );


  buf
  g242
  (
    KeyWire_0_0,
    n204
  );


  not
  g243
  (
    n299,
    n235
  );


  buf
  g244
  (
    n312,
    n203
  );


  not
  g245
  (
    n329,
    n200
  );


  not
  g246
  (
    n272,
    n205
  );


  buf
  g247
  (
    n289,
    n202
  );


  buf
  g248
  (
    n314,
    n228
  );


  not
  g249
  (
    n282,
    n212
  );


  buf
  g250
  (
    n285,
    n226
  );


  not
  g251
  (
    n259,
    n230
  );


  buf
  g252
  (
    n321,
    n205
  );


  buf
  g253
  (
    n295,
    n211
  );


  buf
  g254
  (
    n260,
    n53
  );


  buf
  g255
  (
    n327,
    n211
  );


  not
  g256
  (
    n257,
    n248
  );


  buf
  g257
  (
    n325,
    n227
  );


  nor
  g258
  (
    n305,
    n10,
    n240,
    n207
  );


  nor
  g259
  (
    n258,
    n232,
    n209,
    n213,
    n234
  );


  and
  g260
  (
    n308,
    n204,
    n218,
    n241,
    n208
  );


  xnor
  g261
  (
    n300,
    n207,
    n215,
    n204,
    n231
  );


  or
  g262
  (
    n330,
    n205,
    n221,
    n48,
    n11
  );


  and
  g263
  (
    n261,
    n218,
    n239,
    n233,
    n228
  );


  nand
  g264
  (
    n274,
    n243,
    n219,
    n210,
    n213
  );


  xnor
  g265
  (
    n324,
    n233,
    n48,
    n200,
    n50
  );


  and
  g266
  (
    n270,
    n218,
    n214,
    n210,
    n249
  );


  nor
  g267
  (
    n317,
    n217,
    n52,
    n246,
    n10
  );


  xnor
  g268
  (
    n307,
    n239,
    n222,
    n244,
    n216
  );


  xor
  g269
  (
    n280,
    n233,
    n244,
    n237,
    n209
  );


  xnor
  g270
  (
    n318,
    n231,
    n224,
    n212,
    n213
  );


  xor
  g271
  (
    n269,
    n53,
    n10,
    n240,
    n245
  );


  nor
  g272
  (
    n301,
    n212,
    n202,
    n213,
    n205
  );


  nor
  g273
  (
    n276,
    n237,
    n50,
    n9,
    n249
  );


  or
  g274
  (
    n253,
    n52,
    n49,
    n203,
    n10
  );


  nand
  g275
  (
    n288,
    n247,
    n244,
    n245,
    n52
  );


  xor
  g276
  (
    n302,
    n54,
    n223,
    n228,
    n207
  );


  xnor
  g277
  (
    n322,
    n210,
    n246,
    n242,
    n227
  );


  or
  g278
  (
    n255,
    n227,
    n214,
    n202,
    n220
  );


  nand
  g279
  (
    n266,
    n206,
    n49,
    n52,
    n231
  );


  xor
  g280
  (
    n252,
    n223,
    n237,
    n238,
    n54
  );


  nand
  g281
  (
    n284,
    n201,
    n221,
    n243,
    n49
  );


  xnor
  g282
  (
    n271,
    n206,
    n9,
    n234,
    n222
  );


  nor
  g283
  (
    n309,
    n224,
    n220,
    n48
  );


  or
  g284
  (
    n275,
    n200,
    n245,
    n50,
    n235
  );


  and
  g285
  (
    n292,
    n236,
    n221,
    n215,
    n219
  );


  or
  g286
  (
    n256,
    n208,
    n210,
    n235,
    n234
  );


  xor
  g287
  (
    n297,
    n249,
    n200,
    n53,
    n225
  );


  or
  g288
  (
    n306,
    n216,
    n238,
    n50,
    n249
  );


  nand
  g289
  (
    n296,
    n11,
    n229,
    n241,
    n203
  );


  nand
  g290
  (
    n326,
    n217,
    n234,
    n232,
    n218
  );


  and
  g291
  (
    n323,
    n247,
    n9,
    n224,
    n239
  );


  xor
  g292
  (
    n265,
    n208,
    n233,
    n236,
    n49
  );


  nand
  g293
  (
    n298,
    n247,
    n206,
    n237,
    n238
  );


  nor
  g294
  (
    n262,
    n222,
    n225,
    n208,
    n51
  );


  nand
  g295
  (
    n263,
    n239,
    n209,
    n248,
    n240
  );


  xor
  g296
  (
    n277,
    n217,
    n223,
    n244,
    n238
  );


  nor
  g297
  (
    n279,
    n230,
    n219,
    n225,
    n242
  );


  and
  g298
  (
    n267,
    n203,
    n220,
    n221,
    n242
  );


  nor
  g299
  (
    n319,
    n248,
    n212,
    n225,
    n227
  );


  xor
  g300
  (
    n294,
    n211,
    n214,
    n230,
    n217
  );


  xor
  g301
  (
    n250,
    n216,
    n51,
    n248,
    n246
  );


  xor
  g302
  (
    n315,
    n243,
    n229,
    n230,
    n88
  );


  or
  g303
  (
    n316,
    n201,
    n236,
    n226,
    n207
  );


  nor
  g304
  (
    n273,
    n246,
    n231,
    n226,
    n48
  );


  and
  g305
  (
    n287,
    n201,
    n236,
    n243,
    n215
  );


  xnor
  g306
  (
    n320,
    n242,
    n223,
    n224,
    n241
  );


  xnor
  g307
  (
    n313,
    n206,
    n201,
    n232,
    n209
  );


  xnor
  g308
  (
    n303,
    n228,
    n235,
    n53,
    n51
  );


  nand
  g309
  (
    n286,
    n211,
    n214,
    n216,
    n51
  );


  xnor
  g310
  (
    n362,
    n325,
    n141,
    n133,
    n268
  );


  nor
  g311
  (
    n360,
    n275,
    n309,
    n144,
    n328
  );


  nand
  g312
  (
    n369,
    n154,
    n253,
    n315,
    n308
  );


  nor
  g313
  (
    n381,
    n279,
    n267,
    n134,
    n325
  );


  and
  g314
  (
    n402,
    n159,
    n141,
    n146,
    n327
  );


  xor
  g315
  (
    n351,
    n326,
    n142,
    n261,
    n255
  );


  nand
  g316
  (
    n427,
    n286,
    n148,
    n128,
    n152
  );


  xnor
  g317
  (
    n388,
    n288,
    n160,
    n302,
    n307
  );


  nor
  g318
  (
    n345,
    n274,
    n296,
    n259,
    n263
  );


  nor
  g319
  (
    n363,
    n286,
    n322,
    n328,
    n136
  );


  nand
  g320
  (
    n431,
    n271,
    n263,
    n276,
    n142
  );


  nor
  g321
  (
    n336,
    n300,
    n300,
    n287,
    n313
  );


  xnor
  g322
  (
    n403,
    n278,
    n136,
    n150
  );


  and
  g323
  (
    n334,
    n151,
    n254,
    n318,
    n326
  );


  xnor
  g324
  (
    n348,
    n138,
    n322,
    n327,
    n281
  );


  xor
  g325
  (
    n342,
    n155,
    n156,
    n281,
    n309
  );


  xor
  g326
  (
    n359,
    n330,
    n276,
    n287,
    n262
  );


  nor
  g327
  (
    n424,
    n133,
    n128,
    n329,
    n264
  );


  xnor
  g328
  (
    n335,
    n273,
    n156,
    n297,
    n280
  );


  or
  g329
  (
    n434,
    n313,
    n256,
    n140,
    n136
  );


  nor
  g330
  (
    n408,
    n144,
    n272,
    n320,
    n258
  );


  nor
  g331
  (
    n442,
    n286,
    n282,
    n295,
    n275
  );


  or
  g332
  (
    n357,
    n149,
    n293,
    n260,
    n278
  );


  nand
  g333
  (
    n382,
    n150,
    n324,
    n327,
    n266
  );


  or
  g334
  (
    n346,
    n328,
    n251,
    n260,
    n303
  );


  and
  g335
  (
    n340,
    n151,
    n270,
    n153,
    n264
  );


  nand
  g336
  (
    n374,
    n280,
    n159,
    n138,
    n283
  );


  or
  g337
  (
    n349,
    n139,
    n308,
    n147,
    n155
  );


  or
  g338
  (
    n371,
    n137,
    n258,
    n297,
    n292
  );


  xor
  g339
  (
    n358,
    n146,
    n280,
    n131,
    n314
  );


  and
  g340
  (
    n430,
    n254,
    n321,
    n316,
    n264
  );


  xnor
  g341
  (
    n422,
    n250,
    n259,
    n304,
    n134
  );


  or
  g342
  (
    n433,
    n132,
    n314,
    n160
  );


  xor
  g343
  (
    n419,
    n300,
    n254,
    n317,
    n255
  );


  xnor
  g344
  (
    n428,
    n311,
    n150,
    n281,
    n282
  );


  nor
  g345
  (
    n387,
    n304,
    n293,
    n276,
    n157
  );


  nand
  g346
  (
    n333,
    n258,
    n140,
    n308,
    n301
  );


  or
  g347
  (
    n331,
    n295,
    n143,
    n255,
    n257
  );


  xnor
  g348
  (
    n404,
    n294,
    n154,
    n143,
    n275
  );


  or
  g349
  (
    n410,
    n137,
    n319,
    n129,
    n261
  );


  xnor
  g350
  (
    n375,
    n272,
    n283,
    n298,
    n285
  );


  nand
  g351
  (
    n414,
    n290,
    n130,
    n302,
    n329
  );


  nor
  g352
  (
    n361,
    n301,
    n279,
    n254,
    n297
  );


  xnor
  g353
  (
    n385,
    n289,
    n290,
    n129,
    n309
  );


  nor
  g354
  (
    n379,
    n152,
    n312,
    n292,
    n158
  );


  xnor
  g355
  (
    n441,
    n298,
    n317,
    n284,
    n133
  );


  nor
  g356
  (
    n343,
    n304,
    n266,
    n269,
    n152
  );


  xor
  g357
  (
    n332,
    n288,
    n271,
    n299,
    n287
  );


  nor
  g358
  (
    n391,
    n268,
    n145,
    n153,
    n315
  );


  nand
  g359
  (
    n377,
    n289,
    n146,
    n328,
    n132
  );


  and
  g360
  (
    n365,
    n295,
    n321,
    n283,
    n128
  );


  xnor
  g361
  (
    n390,
    n325,
    n305,
    n263,
    n274
  );


  and
  g362
  (
    n405,
    n316,
    n312,
    n318,
    n324
  );


  and
  g363
  (
    n370,
    n252,
    n159,
    n325,
    n156
  );


  nor
  g364
  (
    n354,
    n320,
    n273,
    n250,
    n257
  );


  or
  g365
  (
    n435,
    n252,
    n147,
    n267,
    n274
  );


  xnor
  g366
  (
    n440,
    n282,
    n154,
    n268,
    n263
  );


  nor
  g367
  (
    n356,
    n330,
    n157,
    n291,
    n266
  );


  or
  g368
  (
    n398,
    n276,
    n131,
    n319,
    n320
  );


  nand
  g369
  (
    n439,
    n145,
    n131,
    n141,
    n267
  );


  and
  g370
  (
    n384,
    n326,
    n251,
    n306,
    n319
  );


  or
  g371
  (
    n426,
    n291,
    n329,
    n140,
    n256
  );


  and
  g372
  (
    n355,
    n312,
    n273,
    n136,
    n261
  );


  nor
  g373
  (
    n401,
    n327,
    n156,
    n272,
    n330
  );


  or
  g374
  (
    n400,
    n289,
    n284,
    n145,
    n296
  );


  xor
  g375
  (
    n397,
    n129,
    n316,
    n252,
    n155
  );


  or
  g376
  (
    n406,
    n307,
    n267,
    n260,
    n143
  );


  xnor
  g377
  (
    n411,
    n269,
    n310,
    n317,
    n291
  );


  xnor
  g378
  (
    n353,
    n310,
    n320,
    n145,
    n277
  );


  or
  g379
  (
    n380,
    n142,
    n314,
    n253,
    n153
  );


  nor
  g380
  (
    n407,
    n251,
    n149,
    n296,
    n140
  );


  and
  g381
  (
    n373,
    n290,
    n287,
    n285
  );


  nand
  g382
  (
    n395,
    n298,
    n310,
    n264,
    n283
  );


  nand
  g383
  (
    n350,
    n255,
    n147,
    n292,
    n301
  );


  or
  g384
  (
    n372,
    n142,
    n149,
    n312,
    n257
  );


  or
  g385
  (
    n367,
    n305,
    n258,
    n318,
    n157
  );


  or
  g386
  (
    n386,
    n323,
    n130,
    n139,
    n296
  );


  nand
  g387
  (
    n432,
    n271,
    n285,
    n262,
    n269
  );


  xor
  g388
  (
    n368,
    n323,
    n139,
    n270,
    n277
  );


  nand
  g389
  (
    n399,
    n290,
    n279,
    n256,
    n271
  );


  xnor
  g390
  (
    n337,
    n307,
    n281,
    n305,
    n137
  );


  xor
  g391
  (
    n366,
    n155,
    n293,
    n270,
    n132
  );


  and
  g392
  (
    n352,
    n288,
    n299,
    n130,
    n324
  );


  and
  g393
  (
    n421,
    n307,
    n315,
    n330,
    n304
  );


  and
  g394
  (
    n347,
    n294,
    n137,
    n297,
    n149
  );


  nor
  g395
  (
    n393,
    n286,
    n324,
    n152,
    n323
  );


  nor
  g396
  (
    n413,
    n157,
    n153,
    n299,
    n306
  );


  nor
  g397
  (
    n443,
    n311,
    n250,
    n143,
    n141
  );


  xnor
  g398
  (
    n444,
    n273,
    n160,
    n158,
    n139
  );


  and
  g399
  (
    n338,
    n278,
    n144,
    n313,
    n131
  );


  nor
  g400
  (
    n416,
    n148,
    n311,
    n251,
    n259
  );


  xnor
  g401
  (
    n389,
    n294,
    n309,
    n158
  );


  xor
  g402
  (
    n417,
    n277,
    n311,
    n310,
    n322
  );


  and
  g403
  (
    n344,
    n129,
    n146,
    n314,
    n289
  );


  and
  g404
  (
    n425,
    n130,
    n148,
    n302,
    n132
  );


  and
  g405
  (
    n437,
    n265,
    n323,
    n135,
    n259
  );


  xor
  g406
  (
    n339,
    n265,
    n303,
    n266,
    n279
  );


  nand
  g407
  (
    n378,
    n275,
    n300,
    n316,
    n301
  );


  nor
  g408
  (
    n383,
    n256,
    n135,
    n270,
    n292
  );


  xor
  g409
  (
    n409,
    n278,
    n326,
    n272,
    n154
  );


  xor
  g410
  (
    n429,
    n134,
    n151,
    n269,
    n265
  );


  xor
  g411
  (
    n376,
    n321,
    n298,
    n306,
    n262
  );


  nor
  g412
  (
    n396,
    n128,
    n303,
    n299,
    n144
  );


  nor
  g413
  (
    n418,
    n329,
    n288,
    n317,
    n293
  );


  xor
  g414
  (
    n412,
    n318,
    n250,
    n313,
    n253
  );


  xor
  g415
  (
    n423,
    n253,
    n159,
    n261,
    n284
  );


  nand
  g416
  (
    n394,
    n302,
    n308,
    n252,
    n135
  );


  nand
  g417
  (
    n364,
    n280,
    n282,
    n277,
    n294
  );


  or
  g418
  (
    n341,
    n315,
    n265,
    n322,
    n260
  );


  xor
  g419
  (
    n438,
    n133,
    n284,
    n306,
    n138
  );


  nor
  g420
  (
    n420,
    n303,
    n134,
    n135,
    n151
  );


  nand
  g421
  (
    n392,
    n147,
    n274,
    n148,
    n321
  );


  xnor
  g422
  (
    n415,
    n138,
    n268,
    n319,
    n291
  );


  xnor
  g423
  (
    n436,
    n262,
    n257,
    n305,
    n295
  );


  buf
  g424
  (
    n449,
    n336
  );


  buf
  g425
  (
    n451,
    n336
  );


  nand
  g426
  (
    n450,
    n341,
    n331,
    n338
  );


  xor
  g427
  (
    n448,
    n339,
    n332,
    n331
  );


  nand
  g428
  (
    n447,
    n335,
    n338,
    n340,
    n333
  );


  xnor
  g429
  (
    n458,
    n341,
    n334,
    n342,
    n331
  );


  nand
  g430
  (
    n456,
    n336,
    n335
  );


  or
  g431
  (
    KeyWire_0_17,
    n339,
    n339,
    n333,
    n342
  );


  and
  g432
  (
    n453,
    n338,
    n335,
    n331,
    n334
  );


  nor
  g433
  (
    n445,
    n332,
    n340,
    n341,
    n337
  );


  nand
  g434
  (
    n446,
    n341,
    n337,
    n333
  );


  and
  g435
  (
    n457,
    n337,
    n332,
    n343,
    n340
  );


  xor
  g436
  (
    n455,
    n338,
    n342,
    n334
  );


  nand
  g437
  (
    n454,
    n339,
    n340,
    n342,
    n337
  );


  not
  g438
  (
    n461,
    n448
  );


  not
  g439
  (
    n465,
    n447
  );


  not
  g440
  (
    n467,
    n445
  );


  buf
  g441
  (
    n459,
    n446
  );


  buf
  g442
  (
    n464,
    n445
  );


  not
  g443
  (
    n460,
    n449
  );


  not
  g444
  (
    n466,
    n446
  );


  buf
  g445
  (
    n462,
    n448
  );


  not
  g446
  (
    n463,
    n447
  );


  not
  g447
  (
    n479,
    n459
  );


  not
  g448
  (
    n476,
    n461
  );


  not
  g449
  (
    n469,
    n462
  );


  buf
  g450
  (
    n481,
    n461
  );


  not
  g451
  (
    n484,
    n462
  );


  not
  g452
  (
    n474,
    n465
  );


  buf
  g453
  (
    n471,
    n463
  );


  not
  g454
  (
    n490,
    n461
  );


  not
  g455
  (
    n488,
    n459
  );


  buf
  g456
  (
    n482,
    n462
  );


  buf
  g457
  (
    n487,
    n464
  );


  not
  g458
  (
    n477,
    n463
  );


  not
  g459
  (
    n486,
    n460
  );


  not
  g460
  (
    n470,
    n464
  );


  not
  g461
  (
    n485,
    n459
  );


  buf
  g462
  (
    n475,
    n460
  );


  buf
  g463
  (
    n493,
    n465
  );


  not
  g464
  (
    n468,
    n463
  );


  buf
  g465
  (
    n492,
    n464
  );


  not
  g466
  (
    n472,
    n462
  );


  buf
  g467
  (
    n473,
    n464
  );


  buf
  g468
  (
    n483,
    n463
  );


  buf
  g469
  (
    n491,
    n460
  );


  not
  g470
  (
    n478,
    n461
  );


  buf
  g471
  (
    n480,
    n465
  );


  buf
  g472
  (
    n489,
    n465
  );


  buf
  g473
  (
    n500,
    n471
  );


  not
  g474
  (
    n499,
    n470
  );


  not
  g475
  (
    n494,
    n468
  );


  not
  g476
  (
    n497,
    n471
  );


  buf
  g477
  (
    n505,
    n471
  );


  buf
  g478
  (
    n495,
    n470
  );


  buf
  g479
  (
    n504,
    n469
  );


  buf
  g480
  (
    n501,
    n468
  );


  buf
  g481
  (
    n502,
    n468
  );


  buf
  g482
  (
    n496,
    n471
  );


  not
  g483
  (
    n503,
    n468
  );


  not
  g484
  (
    n498,
    n469
  );


  and
  g485
  (
    n506,
    n469,
    n470
  );


  buf
  g486
  (
    n527,
    n497
  );


  buf
  g487
  (
    n507,
    n498
  );


  buf
  g488
  (
    n512,
    n495
  );


  not
  g489
  (
    n514,
    n494
  );


  buf
  g490
  (
    n520,
    n497
  );


  buf
  g491
  (
    n521,
    n496
  );


  buf
  g492
  (
    n510,
    n497
  );


  not
  g493
  (
    n517,
    n496
  );


  not
  g494
  (
    n528,
    n496
  );


  buf
  g495
  (
    n513,
    n494
  );


  not
  g496
  (
    n524,
    n498
  );


  not
  g497
  (
    n525,
    n498
  );


  not
  g498
  (
    n516,
    n499
  );


  not
  g499
  (
    n509,
    n495
  );


  buf
  g500
  (
    n523,
    n497
  );


  buf
  g501
  (
    n511,
    n499
  );


  not
  g502
  (
    n508,
    n494
  );


  not
  g503
  (
    n522,
    n496
  );


  not
  g504
  (
    n526,
    n498
  );


  not
  g505
  (
    n519,
    n495
  );


  buf
  g506
  (
    n518,
    n495
  );


  not
  g507
  (
    n515,
    n494
  );


  not
  g508
  (
    n529,
    n511
  );


  not
  g509
  (
    n535,
    n511
  );


  not
  g510
  (
    n536,
    n510
  );


  not
  g511
  (
    n534,
    n510
  );


  not
  g512
  (
    n530,
    n507
  );


  not
  g513
  (
    n533,
    n507
  );


  not
  g514
  (
    n537,
    n507
  );


  not
  g515
  (
    n539,
    n509
  );


  not
  g516
  (
    n538,
    n508
  );


  and
  g517
  (
    n531,
    n507,
    n511,
    n509
  );


  xor
  g518
  (
    n532,
    n511,
    n510,
    n509
  );


  nand
  g519
  (
    n575,
    n113,
    n100,
    n97,
    n107
  );


  or
  g520
  (
    n546,
    n499,
    n112,
    n102,
    n529
  );


  or
  g521
  (
    n557,
    n90,
    n90,
    n539,
    n89
  );


  xor
  g522
  (
    n542,
    n91,
    n109,
    n103
  );


  xnor
  g523
  (
    n552,
    n91,
    n500,
    n92,
    n106
  );


  nor
  g524
  (
    n556,
    n343,
    n90,
    n112,
    n92
  );


  xor
  g525
  (
    n569,
    n104,
    n41,
    n501,
    n101
  );


  nand
  g526
  (
    n554,
    n530,
    n110,
    n537
  );


  or
  g527
  (
    n579,
    n103,
    n43,
    n536,
    n94
  );


  nor
  g528
  (
    n571,
    n106,
    n533,
    n531
  );


  and
  g529
  (
    n563,
    n500,
    n42,
    n105,
    n102
  );


  nand
  g530
  (
    n545,
    n42,
    n106,
    n108,
    n112
  );


  xor
  g531
  (
    n555,
    n538,
    n536,
    n105,
    n345
  );


  nor
  g532
  (
    KeyWire_0_18,
    n539,
    n107,
    n98,
    n112
  );


  or
  g533
  (
    n566,
    n89,
    n103,
    n538,
    n96
  );


  or
  g534
  (
    n564,
    n101,
    n110,
    n41,
    n113
  );


  and
  g535
  (
    n560,
    n500,
    n44,
    n100
  );


  xor
  g536
  (
    n549,
    n100,
    n501,
    n43,
    n97
  );


  nand
  g537
  (
    n576,
    n538,
    n107,
    n99,
    n97
  );


  nor
  g538
  (
    n582,
    n95,
    n343,
    n345,
    n106
  );


  and
  g539
  (
    n559,
    n539,
    n532,
    n531,
    n529
  );


  or
  g540
  (
    n553,
    n531,
    n111,
    n93,
    n533
  );


  nor
  g541
  (
    n562,
    n42,
    n100,
    n108,
    n107
  );


  nor
  g542
  (
    n561,
    n536,
    n111,
    n89,
    n108
  );


  nor
  g543
  (
    n543,
    n101,
    n95,
    n537,
    n113
  );


  xor
  g544
  (
    n577,
    n91,
    n92,
    n95,
    n96
  );


  nor
  g545
  (
    n581,
    n104,
    n103,
    n529,
    n111
  );


  xnor
  g546
  (
    n547,
    n99,
    n501,
    n93,
    n109
  );


  or
  g547
  (
    n540,
    n537,
    n102,
    n98,
    n43
  );


  nand
  g548
  (
    n580,
    n499,
    n535,
    n102,
    n530
  );


  or
  g549
  (
    n583,
    n98,
    n531,
    n44,
    n539
  );


  nor
  g550
  (
    n541,
    n99,
    n44,
    n96,
    n111
  );


  nor
  g551
  (
    n544,
    n344,
    n93,
    n95,
    n538
  );


  or
  g552
  (
    n551,
    n530,
    n344,
    n343,
    n534
  );


  and
  g553
  (
    n558,
    n92,
    n88,
    n536,
    n105
  );


  nor
  g554
  (
    n578,
    n98,
    n91,
    n534,
    n530
  );


  xor
  g555
  (
    n572,
    n104,
    n97,
    n535,
    n534
  );


  nor
  g556
  (
    n565,
    n344,
    n99,
    n533,
    n529
  );


  and
  g557
  (
    KeyWire_0_24,
    n535,
    n532,
    n101,
    n537
  );


  or
  g558
  (
    n570,
    n42,
    n94,
    n532,
    n89
  );


  and
  g559
  (
    n574,
    n344,
    n110,
    n532,
    n93
  );


  nand
  g560
  (
    n550,
    n105,
    n90,
    n534,
    n108
  );


  xor
  g561
  (
    n573,
    n94,
    n535,
    n96,
    n104
  );


  xor
  g562
  (
    n568,
    n94,
    n109,
    n500,
    n43
  );


  nand
  g563
  (
    n599,
    n170,
    n167,
    n174,
    n547
  );


  or
  g564
  (
    n598,
    n544,
    n548,
    n173,
    n177
  );


  xor
  g565
  (
    n597,
    n174,
    n557,
    n546,
    n170
  );


  nand
  g566
  (
    n593,
    n166,
    n175,
    n165,
    n549
  );


  nand
  g567
  (
    n588,
    n177,
    n172,
    n164,
    n165
  );


  nor
  g568
  (
    n584,
    n550,
    n556,
    n162,
    n563
  );


  or
  g569
  (
    n585,
    n168,
    n173,
    n176,
    n162
  );


  and
  g570
  (
    n604,
    n164,
    n551,
    n554,
    n177
  );


  or
  g571
  (
    n603,
    n166,
    n163,
    n174,
    n164
  );


  xor
  g572
  (
    n605,
    n171,
    n170,
    n555,
    n161
  );


  xnor
  g573
  (
    n589,
    n161,
    n543,
    n165,
    n163
  );


  nor
  g574
  (
    n591,
    n175,
    n545,
    n176,
    n169
  );


  xnor
  g575
  (
    n601,
    n172,
    n178,
    n167,
    n170
  );


  nand
  g576
  (
    n594,
    n166,
    n542,
    n163,
    n171
  );


  or
  g577
  (
    n596,
    n162,
    n552,
    n176,
    n173
  );


  nor
  g578
  (
    n592,
    n178,
    n162,
    n174,
    n171
  );


  or
  g579
  (
    n595,
    n176,
    n165,
    n166,
    n177
  );


  and
  g580
  (
    n587,
    n168,
    n168,
    n178,
    n562
  );


  xor
  g581
  (
    n586,
    n173,
    n171,
    n167,
    n559
  );


  or
  g582
  (
    n590,
    n558,
    n172,
    n161,
    n164
  );


  xor
  g583
  (
    n607,
    n168,
    n169,
    n564,
    n561
  );


  and
  g584
  (
    n602,
    n161,
    n169,
    n175,
    n167
  );


  or
  g585
  (
    KeyWire_0_1,
    n169,
    n172,
    n560,
    n175
  );


  nor
  g586
  (
    n606,
    n540,
    n553,
    n163,
    n541
  );


  buf
  g587
  (
    n647,
    n598
  );


  buf
  g588
  (
    n643,
    n589
  );


  not
  g589
  (
    n645,
    n346
  );


  buf
  g590
  (
    n618,
    n346
  );


  not
  g591
  (
    n639,
    n601
  );


  buf
  g592
  (
    n629,
    n585
  );


  not
  g593
  (
    n626,
    n594
  );


  not
  g594
  (
    n633,
    n593
  );


  not
  g595
  (
    n648,
    n592
  );


  buf
  g596
  (
    n640,
    n590
  );


  not
  g597
  (
    n649,
    n587
  );


  buf
  g598
  (
    n628,
    n593
  );


  not
  g599
  (
    n637,
    n596
  );


  not
  g600
  (
    n612,
    n596
  );


  not
  g601
  (
    n641,
    n607
  );


  not
  g602
  (
    n613,
    n606
  );


  not
  g603
  (
    n621,
    n594
  );


  buf
  g604
  (
    n615,
    n602
  );


  not
  g605
  (
    n609,
    n601
  );


  not
  g606
  (
    n619,
    n607
  );


  buf
  g607
  (
    n617,
    n600
  );


  not
  g608
  (
    n642,
    n595
  );


  not
  g609
  (
    n620,
    n591
  );


  buf
  g610
  (
    n627,
    n591
  );


  buf
  g611
  (
    n632,
    n604
  );


  buf
  g612
  (
    n616,
    n345
  );


  buf
  g613
  (
    n630,
    n604
  );


  not
  g614
  (
    n631,
    n599
  );


  not
  g615
  (
    n608,
    n600
  );


  buf
  g616
  (
    n644,
    n589
  );


  buf
  g617
  (
    n638,
    n606
  );


  buf
  g618
  (
    n634,
    n590
  );


  buf
  g619
  (
    KeyWire_0_14,
    n605
  );


  buf
  g620
  (
    n624,
    n597
  );


  not
  g621
  (
    n636,
    n599
  );


  buf
  g622
  (
    n635,
    n592
  );


  not
  g623
  (
    n614,
    n588
  );


  not
  g624
  (
    n650,
    n584
  );


  not
  g625
  (
    n646,
    n603
  );


  buf
  g626
  (
    n623,
    n603
  );


  buf
  g627
  (
    n610,
    n602
  );


  buf
  g628
  (
    n611,
    n595
  );


  nor
  g629
  (
    n651,
    n598,
    n605
  );


  or
  g630
  (
    n622,
    n345,
    n607,
    n597,
    n586
  );


  or
  g631
  (
    n664,
    n620,
    n623,
    n631,
    n632
  );


  xnor
  g632
  (
    n655,
    n615,
    n617,
    n633,
    n611
  );


  or
  g633
  (
    n665,
    n608,
    n622,
    n628,
    n613
  );


  xor
  g634
  (
    KeyWire_0_27,
    n629,
    n611,
    n631,
    n622
  );


  xor
  g635
  (
    n661,
    n631,
    n634,
    n621,
    n613
  );


  nor
  g636
  (
    n668,
    n617,
    n619,
    n614,
    n616
  );


  nand
  g637
  (
    n662,
    n627,
    n610,
    n611,
    n614
  );


  or
  g638
  (
    KeyWire_0_29,
    n608,
    n630,
    n614,
    n622
  );


  nor
  g639
  (
    n663,
    n608,
    n610,
    n612,
    n624
  );


  nor
  g640
  (
    n675,
    n628,
    n626,
    n632,
    n621
  );


  nor
  g641
  (
    n659,
    n612,
    n625,
    n624,
    n634
  );


  xor
  g642
  (
    n671,
    n627,
    n632,
    n628
  );


  xor
  g643
  (
    n669,
    n615,
    n618,
    n623,
    n617
  );


  xor
  g644
  (
    n667,
    n617,
    n628,
    n609,
    n614
  );


  xnor
  g645
  (
    n677,
    n627,
    n624,
    n622,
    n630
  );


  and
  g646
  (
    n678,
    n612,
    n610,
    n621,
    n618
  );


  xor
  g647
  (
    n670,
    n610,
    n623,
    n620,
    n625
  );


  xor
  g648
  (
    n674,
    n612,
    n618,
    n616,
    n621
  );


  xor
  g649
  (
    n673,
    n633,
    n613,
    n634,
    n629
  );


  nand
  g650
  (
    n654,
    n609,
    n620,
    n623,
    n616
  );


  xor
  g651
  (
    n652,
    n630,
    n626,
    n615,
    n609
  );


  and
  g652
  (
    n660,
    n626,
    n611,
    n624,
    n615
  );


  nor
  g653
  (
    n666,
    n620,
    n625,
    n631,
    n634
  );


  nor
  g654
  (
    n676,
    n618,
    n630,
    n633,
    n626
  );


  or
  g655
  (
    n656,
    n616,
    n619,
    n633
  );


  or
  g656
  (
    n658,
    n629,
    n627,
    n609,
    n619
  );


  xnor
  g657
  (
    n653,
    n625,
    n608,
    n613,
    n629
  );


  nand
  g658
  (
    n679,
    n655,
    n658,
    n657,
    n652
  );


  nor
  g659
  (
    n680,
    n653,
    n654,
    n659,
    n656
  );


  buf
  g660
  (
    n683,
    n679
  );


  not
  g661
  (
    n681,
    n679
  );


  buf
  g662
  (
    n682,
    n679
  );


  nand
  g663
  (
    n686,
    n682,
    n683
  );


  and
  g664
  (
    n685,
    n683,
    n683,
    n682,
    n681
  );


  nor
  g665
  (
    n684,
    n682,
    n681
  );


  buf
  g666
  (
    n688,
    n684
  );


  not
  g667
  (
    n689,
    n346
  );


  xor
  g668
  (
    n691,
    n348,
    n349,
    n684,
    n686
  );


  or
  g669
  (
    n690,
    n347,
    n346,
    n348,
    n349
  );


  and
  g670
  (
    n687,
    n348,
    n685,
    n686,
    n347
  );


  xor
  g671
  (
    n692,
    n685,
    n348,
    n347
  );


  not
  g672
  (
    n693,
    n687
  );


  buf
  g673
  (
    n694,
    n688
  );


  not
  g674
  (
    n697,
    n691
  );


  not
  g675
  (
    n695,
    n690
  );


  xnor
  g676
  (
    n696,
    n691,
    n689,
    n692
  );


  and
  g677
  (
    n698,
    n358,
    n353,
    n360,
    n696
  );


  nor
  g678
  (
    n707,
    n355,
    n351,
    n694,
    n354
  );


  and
  g679
  (
    n708,
    n356,
    n352,
    n357,
    n353
  );


  xor
  g680
  (
    n709,
    n354,
    n352,
    n359,
    n361
  );


  nand
  g681
  (
    n702,
    n694,
    n358,
    n362,
    n695
  );


  xor
  g682
  (
    n703,
    n693,
    n697,
    n357
  );


  xnor
  g683
  (
    n699,
    n359,
    n355,
    n352,
    n353
  );


  or
  g684
  (
    n706,
    n693,
    n354,
    n360,
    n696
  );


  or
  g685
  (
    n704,
    n356,
    n695,
    n355,
    n360
  );


  xnor
  g686
  (
    n715,
    n693,
    n350,
    n362
  );


  xor
  g687
  (
    n714,
    n349,
    n349,
    n695,
    n362
  );


  nor
  g688
  (
    n700,
    n352,
    n358,
    n353,
    n360
  );


  xor
  g689
  (
    n711,
    n350,
    n354,
    n357,
    n351
  );


  xnor
  g690
  (
    n710,
    n356,
    n357,
    n695,
    n696
  );


  nand
  g691
  (
    n712,
    n693,
    n355,
    n358,
    n359
  );


  nand
  g692
  (
    n701,
    n696,
    n694,
    n351,
    n361
  );


  or
  g693
  (
    n713,
    n694,
    n356,
    n361,
    n351
  );


  xnor
  g694
  (
    n705,
    n361,
    n359,
    n697,
    n350
  );


  buf
  g695
  (
    n719,
    n699
  );


  not
  g696
  (
    n717,
    n698
  );


  not
  g697
  (
    n716,
    n698
  );


  not
  g698
  (
    n721,
    n698
  );


  buf
  g699
  (
    n720,
    n698
  );


  buf
  g700
  (
    n718,
    n699
  );


  or
  g701
  (
    n732,
    n505,
    n506,
    n721,
    n13
  );


  xnor
  g702
  (
    n739,
    n13,
    n506,
    n580
  );


  or
  g703
  (
    n730,
    n719,
    n13,
    n14,
    n721
  );


  or
  g704
  (
    n722,
    n566,
    n16,
    n717,
    n502
  );


  nand
  g705
  (
    n735,
    n15,
    n567,
    n719,
    n717
  );


  and
  g706
  (
    n734,
    n720,
    n503,
    n718,
    n501
  );


  nand
  g707
  (
    n731,
    n505,
    n15,
    n716,
    n721
  );


  xor
  g708
  (
    n736,
    n12,
    n720,
    n502,
    n571
  );


  nand
  g709
  (
    n744,
    n583,
    n506,
    n504,
    n720
  );


  nand
  g710
  (
    n740,
    n721,
    n503,
    n574,
    n502
  );


  xnor
  g711
  (
    n728,
    n16,
    n716,
    n505,
    n17
  );


  xnor
  g712
  (
    n727,
    n579,
    n575,
    n16,
    n565
  );


  or
  g713
  (
    n725,
    n14,
    n11,
    n13,
    n503
  );


  nor
  g714
  (
    n743,
    n15,
    n576,
    n568,
    n573
  );


  xor
  g715
  (
    n737,
    n717,
    n17,
    n686,
    n716
  );


  or
  g716
  (
    n726,
    n582,
    n569,
    n505,
    n717
  );


  xor
  g717
  (
    n729,
    n12,
    n716,
    n719,
    n577
  );


  xor
  g718
  (
    n733,
    n581,
    n578,
    n718
  );


  and
  g719
  (
    n741,
    n17,
    n719,
    n503,
    n504
  );


  xnor
  g720
  (
    n724,
    n718,
    n502,
    n12,
    n16
  );


  xor
  g721
  (
    n723,
    n572,
    n12,
    n14
  );


  nor
  g722
  (
    n742,
    n11,
    n504,
    n720,
    n697
  );


  nand
  g723
  (
    n738,
    n570,
    n504,
    n15,
    n686
  );


  buf
  g724
  (
    n747,
    n722
  );


  not
  g725
  (
    n774,
    n731
  );


  not
  g726
  (
    n767,
    n734
  );


  buf
  g727
  (
    n778,
    n723
  );


  not
  g728
  (
    n762,
    n733
  );


  buf
  g729
  (
    n757,
    n730
  );


  buf
  g730
  (
    n754,
    n726
  );


  buf
  g731
  (
    n764,
    n724
  );


  buf
  g732
  (
    n761,
    n732
  );


  buf
  g733
  (
    n786,
    n723
  );


  not
  g734
  (
    n782,
    n731
  );


  not
  g735
  (
    n775,
    n723
  );


  not
  g736
  (
    n784,
    n729
  );


  not
  g737
  (
    n776,
    n729
  );


  buf
  g738
  (
    n779,
    n732
  );


  buf
  g739
  (
    n777,
    n728
  );


  buf
  g740
  (
    n789,
    n734
  );


  not
  g741
  (
    n770,
    n724
  );


  buf
  g742
  (
    n787,
    n724
  );


  not
  g743
  (
    n781,
    n726
  );


  not
  g744
  (
    n755,
    n730
  );


  not
  g745
  (
    n766,
    n722
  );


  buf
  g746
  (
    n745,
    n727
  );


  not
  g747
  (
    n753,
    n726
  );


  buf
  g748
  (
    n763,
    n732
  );


  buf
  g749
  (
    n760,
    n733
  );


  buf
  g750
  (
    n772,
    n725
  );


  not
  g751
  (
    n769,
    n734
  );


  buf
  g752
  (
    n758,
    n725
  );


  not
  g753
  (
    n785,
    n727
  );


  not
  g754
  (
    n751,
    n733
  );


  not
  g755
  (
    n788,
    n728
  );


  buf
  g756
  (
    n783,
    n730
  );


  not
  g757
  (
    n750,
    n724
  );


  buf
  g758
  (
    n765,
    n730
  );


  not
  g759
  (
    n780,
    n734
  );


  buf
  g760
  (
    n759,
    n727
  );


  not
  g761
  (
    n771,
    n725
  );


  not
  g762
  (
    n768,
    n732
  );


  buf
  g763
  (
    n752,
    n733
  );


  buf
  g764
  (
    n746,
    n731
  );


  not
  g765
  (
    n773,
    n725
  );


  and
  g766
  (
    n756,
    n726,
    n731
  );


  and
  g767
  (
    n748,
    n728,
    n722,
    n729,
    n727
  );


  nand
  g768
  (
    n749,
    n728,
    n729,
    n723,
    n722
  );


  or
  g769
  (
    n806,
    n761,
    n758,
    n760,
    n762
  );


  and
  g770
  (
    n795,
    n757,
    n762,
    n749
  );


  or
  g771
  (
    n809,
    n752,
    n762,
    n747,
    n764
  );


  xor
  g772
  (
    n796,
    n748,
    n757,
    n755,
    n759
  );


  nor
  g773
  (
    n797,
    n745,
    n748,
    n763
  );


  nand
  g774
  (
    n804,
    n747,
    n745,
    n755,
    n762
  );


  or
  g775
  (
    n808,
    n750,
    n749,
    n754
  );


  xor
  g776
  (
    n801,
    n759,
    n752,
    n745,
    n758
  );


  xor
  g777
  (
    n798,
    n750,
    n753,
    n763,
    n747
  );


  xor
  g778
  (
    n803,
    n760,
    n748,
    n753,
    n746
  );


  xor
  g779
  (
    n800,
    n751,
    n751,
    n757,
    n756
  );


  xnor
  g780
  (
    n805,
    n756,
    n761,
    n764
  );


  and
  g781
  (
    n792,
    n748,
    n749,
    n758,
    n754
  );


  xor
  g782
  (
    n793,
    n764,
    n756,
    n750,
    n753
  );


  xnor
  g783
  (
    n802,
    n759,
    n746,
    n751,
    n745
  );


  or
  g784
  (
    n790,
    n758,
    n750,
    n761,
    n755
  );


  nor
  g785
  (
    n791,
    n760,
    n752,
    n751,
    n754
  );


  nor
  g786
  (
    n794,
    n746,
    n761,
    n755,
    n747
  );


  and
  g787
  (
    n799,
    n763,
    n756,
    n746,
    n752
  );


  and
  g788
  (
    n807,
    n760,
    n757,
    n753,
    n759
  );


  and
  g789
  (
    n810,
    n800,
    n795,
    n792,
    n801
  );


  or
  g790
  (
    n815,
    n702,
    n800,
    n701
  );


  or
  g791
  (
    KeyWire_0_19,
    n710,
    n799,
    n707,
    n795
  );


  nand
  g792
  (
    n814,
    n797,
    n700,
    n707,
    n793
  );


  or
  g793
  (
    n812,
    n797,
    n791,
    n794,
    n793
  );


  nor
  g794
  (
    n823,
    n798,
    n796,
    n790,
    n709
  );


  or
  g795
  (
    n817,
    n708,
    n706,
    n701
  );


  or
  g796
  (
    n816,
    n704,
    n702,
    n705
  );


  nand
  g797
  (
    n825,
    n701,
    n702,
    n708
  );


  or
  g798
  (
    KeyWire_0_11,
    n703,
    n796,
    n798,
    n705
  );


  xor
  g799
  (
    n822,
    n710,
    n700,
    n699,
    n709
  );


  nand
  g800
  (
    n811,
    n704,
    n703,
    n794,
    n702
  );


  and
  g801
  (
    n819,
    n699,
    n700,
    n703,
    n799
  );


  xor
  g802
  (
    n813,
    n709,
    n708,
    n704
  );


  and
  g803
  (
    n818,
    n700,
    n705,
    n707
  );


  nor
  g804
  (
    n820,
    n709,
    n706,
    n703
  );


  and
  g805
  (
    n834,
    n770,
    n812,
    n813,
    n765
  );


  and
  g806
  (
    n835,
    n812,
    n770,
    n767
  );


  nand
  g807
  (
    n832,
    n773,
    n769,
    n814,
    n816
  );


  nand
  g808
  (
    n827,
    n816,
    n765,
    n767
  );


  nand
  g809
  (
    n826,
    n768,
    n815,
    n772,
    n765
  );


  nor
  g810
  (
    n831,
    n773,
    n765,
    n770,
    n771
  );


  nand
  g811
  (
    n830,
    n769,
    n813,
    n771,
    n768
  );


  nand
  g812
  (
    n837,
    n810,
    n772
  );


  nor
  g813
  (
    n829,
    n771,
    n766,
    n772,
    n768
  );


  and
  g814
  (
    n828,
    n767,
    n769,
    n771
  );


  xnor
  g815
  (
    n836,
    n815,
    n766,
    n811
  );


  nand
  g816
  (
    n833,
    n811,
    n768,
    n814,
    n766
  );


  and
  g817
  (
    n847,
    n449,
    n179,
    n455,
    n178
  );


  nor
  g818
  (
    n843,
    n827,
    n179,
    n829
  );


  nand
  g819
  (
    n845,
    n836,
    n830,
    n837
  );


  xnor
  g820
  (
    n850,
    n831,
    n180,
    n454
  );


  or
  g821
  (
    n854,
    n180,
    n831,
    n182,
    n833
  );


  nor
  g822
  (
    n851,
    n363,
    n450,
    n362,
    n834
  );


  nand
  g823
  (
    n855,
    n831,
    n835,
    n363,
    n179
  );


  nand
  g824
  (
    n853,
    n837,
    n834,
    n827,
    n451
  );


  or
  g825
  (
    n841,
    n452,
    n454,
    n181,
    n364
  );


  or
  g826
  (
    n844,
    n836,
    n181,
    n832,
    n363
  );


  and
  g827
  (
    n852,
    n830,
    n834,
    n829,
    n832
  );


  nor
  g828
  (
    n840,
    n453,
    n452,
    n181
  );


  nor
  g829
  (
    n846,
    n836,
    n826,
    n829,
    n832
  );


  nand
  g830
  (
    n842,
    n179,
    n826,
    n453,
    n455
  );


  nand
  g831
  (
    n849,
    n453,
    n450,
    n837,
    n180
  );


  or
  g832
  (
    n856,
    n836,
    n830,
    n454,
    n835
  );


  or
  g833
  (
    n839,
    n182,
    n364,
    n833,
    n828
  );


  xnor
  g834
  (
    n848,
    n828,
    n833,
    n364
  );


  nor
  g835
  (
    n857,
    n834,
    n363,
    n832,
    n835
  );


  or
  g836
  (
    n838,
    n835,
    n831,
    n451,
    n54
  );


  or
  g837
  (
    n860,
    n844,
    n847,
    n365,
    n375
  );


  nor
  g838
  (
    n863,
    n850,
    n841,
    n374,
    n369
  );


  nand
  g839
  (
    n878,
    n851,
    n370,
    n369
  );


  xor
  g840
  (
    n872,
    n368,
    n839,
    n366,
    n513
  );


  nand
  g841
  (
    n874,
    n367,
    n843,
    n512,
    n374
  );


  nor
  g842
  (
    n862,
    n372,
    n371,
    n366
  );


  nand
  g843
  (
    n868,
    n365,
    n846,
    n368,
    n467
  );


  or
  g844
  (
    n864,
    n512,
    n845,
    n514,
    n849
  );


  xor
  g845
  (
    n877,
    n367,
    n844,
    n514,
    n660
  );


  xnor
  g846
  (
    n871,
    n513,
    n842,
    n371,
    n845
  );


  nand
  g847
  (
    n875,
    n369,
    n366,
    n846,
    n374
  );


  or
  g848
  (
    n870,
    n513,
    n466,
    n371
  );


  xnor
  g849
  (
    n876,
    n840,
    n849,
    n512,
    n374
  );


  xor
  g850
  (
    n873,
    n373,
    n848,
    n367,
    n365
  );


  nand
  g851
  (
    n861,
    n513,
    n367,
    n368,
    n467
  );


  nand
  g852
  (
    n867,
    n512,
    n848,
    n370,
    n467
  );


  and
  g853
  (
    n859,
    n838,
    n366,
    n850,
    n372
  );


  or
  g854
  (
    n865,
    n466,
    n373,
    n375,
    n467
  );


  or
  g855
  (
    n866,
    n373,
    n847,
    n364,
    n368
  );


  nor
  g856
  (
    n858,
    n370,
    n373,
    n372
  );


  nor
  g857
  (
    n869,
    n466,
    n365,
    n369,
    n851
  );


  xnor
  g858
  (
    n915,
    n641,
    n646,
    n636,
    n476
  );


  or
  g859
  (
    n887,
    n859,
    n871,
    n192,
    n873
  );


  and
  g860
  (
    n916,
    n472,
    n869,
    n191,
    n859
  );


  xor
  g861
  (
    n926,
    n489,
    n187,
    n198,
    n481
  );


  and
  g862
  (
    n908,
    n476,
    n481,
    n647,
    n648
  );


  and
  g863
  (
    n914,
    n862,
    n645,
    n863
  );


  xor
  g864
  (
    n950,
    n650,
    n875,
    n489,
    n864
  );


  xor
  g865
  (
    n881,
    n873,
    n641,
    n475,
    n638
  );


  and
  g866
  (
    n895,
    n456,
    n185,
    n869,
    n871
  );


  nor
  g867
  (
    n936,
    n484,
    n190,
    n192,
    n870
  );


  xor
  g868
  (
    n957,
    n199,
    n484,
    n863,
    n680
  );


  nand
  g869
  (
    n937,
    n859,
    n489,
    n864,
    n478
  );


  nor
  g870
  (
    n897,
    n489,
    n484,
    n646,
    n186
  );


  xor
  g871
  (
    n913,
    n376,
    n188,
    n480,
    n195
  );


  xor
  g872
  (
    KeyWire_0_23,
    n871,
    n874,
    n475,
    n642
  );


  xor
  g873
  (
    n933,
    n635,
    n476,
    n473,
    n859
  );


  nor
  g874
  (
    n939,
    n472,
    n475,
    n735,
    n647
  );


  xor
  g875
  (
    n917,
    n869,
    n375,
    n642,
    n190
  );


  nand
  g876
  (
    n894,
    n483,
    n490,
    n198
  );


  nor
  g877
  (
    n954,
    n651,
    n647,
    n635,
    n198
  );


  xnor
  g878
  (
    n921,
    n485,
    n472,
    n189,
    n860
  );


  or
  g879
  (
    n946,
    n642,
    n191,
    n183,
    n486
  );


  xor
  g880
  (
    n922,
    n189,
    n858,
    n479,
    n184
  );


  and
  g881
  (
    n923,
    n877,
    n801,
    n479,
    n194
  );


  nand
  g882
  (
    n888,
    n865,
    n868,
    n644,
    n861
  );


  or
  g883
  (
    n890,
    n644,
    n482,
    n877
  );


  xor
  g884
  (
    n929,
    n649,
    n485,
    n375,
    n806
  );


  or
  g885
  (
    n951,
    n874,
    n804,
    n191,
    n198
  );


  xnor
  g886
  (
    n883,
    n863,
    n199,
    n639,
    n803
  );


  xor
  g887
  (
    n882,
    n483,
    n863,
    n647,
    n491
  );


  xnor
  g888
  (
    n910,
    n194,
    n455,
    n635,
    n860
  );


  nor
  g889
  (
    n909,
    n861,
    n861,
    n475,
    n185
  );


  xor
  g890
  (
    n919,
    n195,
    n872,
    n637,
    n194
  );


  xor
  g891
  (
    n912,
    n188,
    n876,
    n477,
    n191
  );


  nand
  g892
  (
    n947,
    n486,
    n479,
    n869,
    n867
  );


  xnor
  g893
  (
    n911,
    n643,
    n195,
    n637,
    n680
  );


  and
  g894
  (
    n944,
    n484,
    n641,
    n873,
    n192
  );


  or
  g895
  (
    n884,
    n183,
    n488,
    n184,
    n480
  );


  xnor
  g896
  (
    n958,
    n483,
    n182,
    n642,
    n488
  );


  and
  g897
  (
    n948,
    n866,
    n490,
    n864,
    n862
  );


  xnor
  g898
  (
    n885,
    n481,
    n477,
    n867,
    n478
  );


  and
  g899
  (
    n907,
    n803,
    n870,
    n872,
    n639
  );


  and
  g900
  (
    n942,
    n474,
    n376,
    n805,
    n650
  );


  or
  g901
  (
    n903,
    n870,
    n199,
    n474,
    n643
  );


  xor
  g902
  (
    n952,
    n197,
    n193,
    n650,
    n640
  );


  nand
  g903
  (
    n900,
    n189,
    n651,
    n184,
    n188
  );


  xor
  g904
  (
    n920,
    n874,
    n640,
    n638,
    n865
  );


  nor
  g905
  (
    n934,
    n455,
    n866,
    n804,
    n189
  );


  nor
  g906
  (
    n945,
    n194,
    n638,
    n861
  );


  xor
  g907
  (
    n898,
    n187,
    n185,
    n876,
    n636
  );


  xnor
  g908
  (
    n905,
    n474,
    n482,
    n192,
    n183
  );


  nand
  g909
  (
    n949,
    n860,
    n488,
    n199,
    n636
  );


  xor
  g910
  (
    n925,
    n490,
    n644,
    n868
  );


  nor
  g911
  (
    n902,
    n473,
    n866,
    n187,
    n482
  );


  and
  g912
  (
    n904,
    n646,
    n643,
    n183,
    n186
  );


  or
  g913
  (
    n892,
    n806,
    n473,
    n872,
    n196
  );


  nor
  g914
  (
    n940,
    n197,
    n862,
    n481,
    n193
  );


  xnor
  g915
  (
    n938,
    n865,
    n648,
    n649,
    n805
  );


  and
  g916
  (
    n927,
    n486,
    n645,
    n186,
    n196
  );


  nand
  g917
  (
    n932,
    n650,
    n649,
    n184,
    n474
  );


  and
  g918
  (
    n953,
    n649,
    n487,
    n477,
    n486
  );


  nor
  g919
  (
    n896,
    n866,
    n646,
    n858,
    n864
  );


  and
  g920
  (
    n891,
    n477,
    n478,
    n802,
    n858
  );


  xor
  g921
  (
    n943,
    n485,
    n487,
    n867,
    n479
  );


  xor
  g922
  (
    n930,
    n195,
    n651,
    n860,
    n640
  );


  or
  g923
  (
    n955,
    n875,
    n867,
    n480,
    n476
  );


  xnor
  g924
  (
    n935,
    n875,
    n196,
    n802,
    n640
  );


  and
  g925
  (
    n886,
    n480,
    n472,
    n868,
    n877
  );


  and
  g926
  (
    n924,
    n187,
    n186,
    n644,
    n185
  );


  nand
  g927
  (
    n889,
    n491,
    n875,
    n487
  );


  xnor
  g928
  (
    n906,
    n862,
    n636,
    n456,
    n639
  );


  nor
  g929
  (
    n880,
    n188,
    n870,
    n478,
    n639
  );


  nand
  g930
  (
    n901,
    n488,
    n483,
    n641,
    n197
  );


  and
  g931
  (
    n899,
    n871,
    n190,
    n873,
    n648
  );


  and
  g932
  (
    n956,
    n197,
    n473,
    n865,
    n651
  );


  nand
  g933
  (
    n879,
    n872,
    n643,
    n858,
    n485
  );


  and
  g934
  (
    n918,
    n193,
    n196,
    n874,
    n635
  );


  xor
  g935
  (
    n931,
    n193,
    n876,
    n637
  );


  xor
  g936
  (
    n928,
    n456,
    n491,
    n645,
    n190
  );


  nor
  g937
  (
    n941,
    n637,
    n182,
    n648,
    n877
  );


  xnor
  g938
  (
    n971,
    n902,
    n879,
    n897,
    n885
  );


  nand
  g939
  (
    n961,
    n889,
    n907,
    n882,
    n903
  );


  and
  g940
  (
    n964,
    n890,
    n883,
    n891,
    n887
  );


  xnor
  g941
  (
    n959,
    n892,
    n885,
    n896,
    n900
  );


  nand
  g942
  (
    n970,
    n907,
    n883,
    n897,
    n904
  );


  xnor
  g943
  (
    n968,
    n896,
    n894,
    n888
  );


  nor
  g944
  (
    n966,
    n903,
    n886,
    n895,
    n900
  );


  nor
  g945
  (
    n969,
    n899,
    n890,
    n906,
    n895
  );


  xnor
  g946
  (
    n972,
    n881,
    n908,
    n898,
    n888
  );


  xor
  g947
  (
    n962,
    n889,
    n906,
    n901,
    n880
  );


  nand
  g948
  (
    n960,
    n891,
    n884,
    n893,
    n880
  );


  or
  g949
  (
    n973,
    n881,
    n892,
    n893,
    n886
  );


  xor
  g950
  (
    n965,
    n884,
    n887,
    n905,
    n879
  );


  nand
  g951
  (
    n963,
    n902,
    n901,
    n908,
    n898
  );


  and
  g952
  (
    KeyWire_0_22,
    n899,
    n904,
    n905,
    n882
  );


  xor
  g953
  (
    n988,
    n972,
    n515,
    n519,
    n837
  );


  nor
  g954
  (
    n986,
    n519,
    n967,
    n518,
    n516
  );


  nand
  g955
  (
    n983,
    n520,
    n969,
    n712,
    n714
  );


  or
  g956
  (
    n989,
    n963,
    n712,
    n968,
    n710
  );


  or
  g957
  (
    n975,
    n710,
    n960,
    n376,
    n970
  );


  and
  g958
  (
    n977,
    n514,
    n961,
    n973
  );


  and
  g959
  (
    KeyWire_0_5,
    n517,
    n972,
    n456,
    n959
  );


  nor
  g960
  (
    n974,
    n516,
    n518,
    n517
  );


  or
  g961
  (
    n978,
    n714,
    n711,
    n713
  );


  nand
  g962
  (
    n982,
    n518,
    n713,
    n519,
    n516
  );


  nand
  g963
  (
    n984,
    n515,
    n515,
    n971,
    n712
  );


  and
  g964
  (
    n981,
    n711,
    n711,
    n514,
    n517
  );


  or
  g965
  (
    n979,
    n968,
    n713,
    n970,
    n965
  );


  and
  g966
  (
    n985,
    n519,
    n713,
    n969,
    n966
  );


  or
  g967
  (
    n976,
    n515,
    n517,
    n712,
    n516
  );


  nor
  g968
  (
    n980,
    n964,
    n962,
    n376,
    n971
  );


  buf
  g969
  (
    n993,
    n978
  );


  not
  g970
  (
    n1012,
    n975
  );


  buf
  g971
  (
    n1021,
    n974
  );


  not
  g972
  (
    n1001,
    n980
  );


  not
  g973
  (
    n1004,
    n978
  );


  buf
  g974
  (
    n1003,
    n976
  );


  not
  g975
  (
    n1009,
    n980
  );


  buf
  g976
  (
    n1020,
    n977
  );


  buf
  g977
  (
    n997,
    n983
  );


  buf
  g978
  (
    n1019,
    n979
  );


  not
  g979
  (
    n1002,
    n984
  );


  not
  g980
  (
    n1015,
    n982
  );


  not
  g981
  (
    n1010,
    n975
  );


  not
  g982
  (
    n1007,
    n982
  );


  buf
  g983
  (
    n1011,
    n974
  );


  not
  g984
  (
    n1018,
    n981
  );


  not
  g985
  (
    n1013,
    n984
  );


  not
  g986
  (
    n1000,
    n982
  );


  buf
  g987
  (
    n1016,
    n975
  );


  buf
  g988
  (
    n1014,
    n981
  );


  buf
  g989
  (
    n996,
    n980
  );


  buf
  g990
  (
    n991,
    n983
  );


  not
  g991
  (
    n994,
    n981
  );


  buf
  g992
  (
    n1008,
    n979
  );


  not
  g993
  (
    n999,
    n909
  );


  or
  g994
  (
    n992,
    n983,
    n984,
    n981
  );


  or
  g995
  (
    n1005,
    n978,
    n979
  );


  and
  g996
  (
    n995,
    n975,
    n982,
    n980
  );


  or
  g997
  (
    n1017,
    n985,
    n976
  );


  xnor
  g998
  (
    n998,
    n974,
    n976,
    n983
  );


  xor
  g999
  (
    n1006,
    n974,
    n977,
    n984
  );


  xnor
  g1000
  (
    n990,
    n978,
    n977
  );


  buf
  g1001
  (
    n1022,
    n990
  );


  not
  g1002
  (
    n1026,
    n912
  );


  nand
  g1003
  (
    n1024,
    n910,
    n1022
  );


  xor
  g1004
  (
    n1025,
    n1022,
    n911
  );


  or
  g1005
  (
    n1023,
    n1022,
    n909,
    n910
  );


  or
  g1006
  (
    n1031,
    n1026,
    n521,
    n527
  );


  xor
  g1007
  (
    n1039,
    n913,
    n913,
    n1026,
    n1023
  );


  nor
  g1008
  (
    n1033,
    n520,
    n807,
    n522,
    n1026
  );


  nor
  g1009
  (
    n1042,
    n524,
    n809,
    n1025
  );


  xor
  g1010
  (
    n1034,
    n524,
    n457,
    n458,
    n1024
  );


  xor
  g1011
  (
    n1037,
    n526,
    n526,
    n523,
    n521
  );


  nor
  g1012
  (
    n1030,
    n458,
    n523,
    n524,
    n525
  );


  nor
  g1013
  (
    n1041,
    n522,
    n525,
    n458,
    n520
  );


  xnor
  g1014
  (
    n1029,
    n457,
    n1024,
    n527
  );


  or
  g1015
  (
    n1038,
    n522,
    n1024,
    n809,
    n525
  );


  and
  g1016
  (
    n1036,
    n457,
    n1026,
    n527,
    n520
  );


  nor
  g1017
  (
    n1035,
    n457,
    n526,
    n808,
    n807
  );


  or
  g1018
  (
    n1032,
    n521,
    n1023,
    n914,
    n523
  );


  or
  g1019
  (
    n1028,
    n458,
    n1025,
    n1024,
    n808
  );


  xor
  g1020
  (
    n1027,
    n523,
    n526,
    n522,
    n524
  );


  xor
  g1021
  (
    n1040,
    n1025,
    n1023,
    n525
  );


  and
  g1022
  (
    n1075,
    n671,
    n492,
    n385,
    n379
  );


  xnor
  g1023
  (
    n1062,
    n392,
    n380,
    n663,
    n1032
  );


  nand
  g1024
  (
    n1094,
    n383,
    n1028,
    n395,
    n743
  );


  nor
  g1025
  (
    n1065,
    n389,
    n821,
    n387
  );


  and
  g1026
  (
    n1071,
    n1029,
    n820,
    n1031,
    n667
  );


  and
  g1027
  (
    n1060,
    n379,
    n1036,
    n383,
    n1041
  );


  nand
  g1028
  (
    n1087,
    n1038,
    n492,
    n735,
    n394
  );


  nor
  g1029
  (
    n1074,
    n987,
    n381,
    n384,
    n380
  );


  xnor
  g1030
  (
    n1058,
    n820,
    n739,
    n386,
    n1039
  );


  nand
  g1031
  (
    n1067,
    n665,
    n674,
    n818,
    n384
  );


  and
  g1032
  (
    n1080,
    n735,
    n1030,
    n379
  );


  nor
  g1033
  (
    n1093,
    n744,
    n386,
    n743,
    n673
  );


  nor
  g1034
  (
    n1106,
    n822,
    n382,
    n676,
    n390
  );


  or
  g1035
  (
    n1066,
    n389,
    n664,
    n393,
    n381
  );


  nand
  g1036
  (
    n1078,
    n824,
    n822,
    n384,
    n743
  );


  xnor
  g1037
  (
    n1047,
    n1031,
    n396,
    n740
  );


  and
  g1038
  (
    n1083,
    n819,
    n1032,
    n383,
    n738
  );


  nand
  g1039
  (
    n1053,
    n383,
    n822,
    n395,
    n678
  );


  and
  g1040
  (
    n1045,
    n675,
    n823,
    n377,
    n740
  );


  xnor
  g1041
  (
    n1063,
    n1027,
    n741,
    n739,
    n744
  );


  nand
  g1042
  (
    n1085,
    n985,
    n394,
    n1033,
    n382
  );


  nor
  g1043
  (
    n1100,
    n1028,
    n823,
    n737,
    n1034
  );


  nand
  g1044
  (
    n1044,
    n1028,
    n818,
    n738,
    n1035
  );


  xor
  g1045
  (
    n1052,
    n987,
    n673,
    n818,
    n1028
  );


  and
  g1046
  (
    n1104,
    n820,
    n1032,
    n1037,
    n1041
  );


  and
  g1047
  (
    n1061,
    n385,
    n670,
    n391,
    n1040
  );


  nor
  g1048
  (
    n1055,
    n988,
    n393,
    n1042,
    n661
  );


  and
  g1049
  (
    n1101,
    n380,
    n393,
    n395
  );


  or
  g1050
  (
    n1082,
    n391,
    n388,
    n744,
    n1038
  );


  and
  g1051
  (
    n1103,
    n674,
    n396,
    n1032
  );


  and
  g1052
  (
    n1089,
    n1029,
    n1037,
    n735,
    n388
  );


  xnor
  g1053
  (
    n1096,
    n743,
    n736,
    n378,
    n1029
  );


  and
  g1054
  (
    n1092,
    n1034,
    n377,
    n672,
    n741
  );


  nor
  g1055
  (
    n1097,
    n738,
    n1030,
    n988,
    n672
  );


  xor
  g1056
  (
    n1068,
    n989,
    n821,
    n1027,
    n1040
  );


  xnor
  g1057
  (
    n1054,
    n1042,
    n742,
    n380,
    n819
  );


  xnor
  g1058
  (
    n1059,
    n1033,
    n389,
    n1034,
    n385
  );


  xnor
  g1059
  (
    n1105,
    n1029,
    n1038,
    n738,
    n985
  );


  nand
  g1060
  (
    n1057,
    n1031,
    n392,
    n988,
    n396
  );


  and
  g1061
  (
    n1079,
    n675,
    n387,
    n1042,
    n1041
  );


  or
  g1062
  (
    n1084,
    n384,
    n736,
    n378,
    n1035
  );


  nand
  g1063
  (
    n1049,
    n985,
    n388,
    n666
  );


  xnor
  g1064
  (
    n1069,
    n1035,
    n741,
    n822,
    n386
  );


  xnor
  g1065
  (
    n1102,
    n819,
    n381,
    n739,
    n392
  );


  nor
  g1066
  (
    n1086,
    n987,
    n381,
    n741,
    n1031
  );


  nor
  g1067
  (
    n1076,
    n385,
    n1033,
    n1036
  );


  and
  g1068
  (
    n1043,
    n740,
    n394,
    n1038,
    n737
  );


  xor
  g1069
  (
    n1051,
    n736,
    n817,
    n986,
    n491
  );


  or
  g1070
  (
    n1050,
    n668,
    n737,
    n1035,
    n1027
  );


  or
  g1071
  (
    n1088,
    n824,
    n736,
    n382,
    n823
  );


  xor
  g1072
  (
    n1091,
    n823,
    n378,
    n390
  );


  xor
  g1073
  (
    n1056,
    n819,
    n742,
    n397,
    n391
  );


  xor
  g1074
  (
    n1072,
    n382,
    n676,
    n739,
    n821
  );


  xnor
  g1075
  (
    n1099,
    n986,
    n1039,
    n1040,
    n987
  );


  and
  g1076
  (
    n1064,
    n677,
    n1027,
    n986,
    n1040
  );


  or
  g1077
  (
    n1098,
    n1030,
    n387,
    n737,
    n391
  );


  xor
  g1078
  (
    n1048,
    n392,
    n1042,
    n1036,
    n1030
  );


  nand
  g1079
  (
    n1077,
    n817,
    n662,
    n821,
    n1039
  );


  and
  g1080
  (
    n1090,
    n824,
    n1037,
    n393,
    n677
  );


  xor
  g1081
  (
    n1073,
    n378,
    n386,
    n394,
    n742
  );


  xor
  g1082
  (
    n1095,
    n986,
    n1039,
    n1033,
    n377
  );


  and
  g1083
  (
    n1046,
    n1037,
    n988,
    n818,
    n1041
  );


  xnor
  g1084
  (
    n1081,
    n744,
    n1034,
    n820,
    n390
  );


  xor
  g1085
  (
    n1070,
    n389,
    n742,
    n669,
    n377
  );


  nor
  g1086
  (
    n1151,
    n990,
    n1073,
    n1081,
    n1105
  );


  or
  g1087
  (
    n1183,
    n1080,
    n1103,
    n1003,
    n1052
  );


  xor
  g1088
  (
    n1149,
    n1002,
    n1098,
    n1011,
    n1094
  );


  xor
  g1089
  (
    n1144,
    n1076,
    n1020,
    n1090,
    n999
  );


  and
  g1090
  (
    n1160,
    n1010,
    n1102,
    n1003,
    n1099
  );


  xor
  g1091
  (
    n1171,
    n1060,
    n773,
    n1045,
    n1020
  );


  xor
  g1092
  (
    n1128,
    n996,
    n1081,
    n999,
    n1009
  );


  xnor
  g1093
  (
    n1165,
    n1104,
    n1043,
    n1049,
    n995
  );


  and
  g1094
  (
    n1203,
    n997,
    n1096,
    n1066,
    n1000
  );


  or
  g1095
  (
    n1113,
    n1098,
    n998,
    n1090,
    n1008
  );


  nand
  g1096
  (
    n1170,
    n1087,
    n991,
    n1095,
    n1062
  );


  xnor
  g1097
  (
    n1194,
    n1069,
    n1009,
    n1049,
    n1106
  );


  or
  g1098
  (
    n1167,
    n1106,
    n1014,
    n1082,
    n776
  );


  xnor
  g1099
  (
    n1131,
    n1064,
    n1097,
    n995,
    n994
  );


  and
  g1100
  (
    n1158,
    n1013,
    n1011,
    n1021,
    n1018
  );


  and
  g1101
  (
    n1173,
    n1006,
    n1101,
    n1096,
    n1012
  );


  nor
  g1102
  (
    n1200,
    n1062,
    n1092,
    n1043,
    n1067
  );


  or
  g1103
  (
    n1154,
    n1059,
    n1093,
    n1057,
    n995
  );


  xor
  g1104
  (
    n1119,
    n1056,
    n1095,
    n1058,
    n1097
  );


  or
  g1105
  (
    n1198,
    n1083,
    n1012,
    n1018,
    n1106
  );


  nand
  g1106
  (
    n1190,
    n1020,
    n1006,
    n1056,
    n1068
  );


  xor
  g1107
  (
    n1197,
    n1100,
    n1069,
    n1004,
    n1068
  );


  xor
  g1108
  (
    n1111,
    n1007,
    n1008,
    n1012,
    n1105
  );


  nor
  g1109
  (
    n1136,
    n1000,
    n1102,
    n1094,
    n1088
  );


  nor
  g1110
  (
    n1157,
    n1043,
    n1088,
    n1070,
    n1087
  );


  xor
  g1111
  (
    n1118,
    n991,
    n1046,
    n1086,
    n774
  );


  nor
  g1112
  (
    n1115,
    n1047,
    n1089,
    n998,
    n1100
  );


  nor
  g1113
  (
    KeyWire_0_25,
    n1085,
    n775,
    n1046,
    n1053
  );


  nor
  g1114
  (
    n1182,
    n777,
    n1076,
    n1089,
    n1097
  );


  xor
  g1115
  (
    n1179,
    n1079,
    n1087,
    n1006,
    n1053
  );


  or
  g1116
  (
    n1153,
    n1089,
    n1054,
    n1053,
    n992
  );


  nand
  g1117
  (
    n1121,
    n1091,
    n1065,
    n1099,
    n1049
  );


  xnor
  g1118
  (
    n1134,
    n1092,
    n993,
    n1073,
    n1061
  );


  nor
  g1119
  (
    n1143,
    n994,
    n1091,
    n1054,
    n1058
  );


  and
  g1120
  (
    n1116,
    n1014,
    n991,
    n1048,
    n1095
  );


  xor
  g1121
  (
    n1132,
    n1059,
    n774,
    n1075,
    n1094
  );


  xor
  g1122
  (
    n1206,
    n997,
    n997,
    n1019,
    n1083
  );


  xnor
  g1123
  (
    n1188,
    n1084,
    n1061,
    n996,
    n1060
  );


  xnor
  g1124
  (
    n1164,
    n1071,
    n1051,
    n1105,
    n1075
  );


  nor
  g1125
  (
    n1202,
    n1067,
    n1074,
    n1005,
    n1047
  );


  xor
  g1126
  (
    n1141,
    n1017,
    n775,
    n1055,
    n1014
  );


  or
  g1127
  (
    n1125,
    n1006,
    n1063,
    n1051,
    n1016
  );


  xnor
  g1128
  (
    n1129,
    n1044,
    n1017,
    n1064,
    n1050
  );


  xnor
  g1129
  (
    n1193,
    n1057,
    n1077,
    n1072,
    n1010
  );


  nand
  g1130
  (
    n1138,
    n1047,
    n1001,
    n1008,
    n1057
  );


  xnor
  g1131
  (
    n1120,
    n1076,
    n1082,
    n1059,
    n1088
  );


  xor
  g1132
  (
    n1139,
    n1071,
    n1069,
    n1005,
    n992
  );


  xor
  g1133
  (
    n1159,
    n996,
    n1072,
    n1099,
    n774
  );


  nand
  g1134
  (
    n1172,
    n997,
    n1100,
    n1045
  );


  xor
  g1135
  (
    n1123,
    n1000,
    n1084,
    n1081,
    n1009
  );


  xnor
  g1136
  (
    n1133,
    n1062,
    n1002,
    n1049,
    n999
  );


  nand
  g1137
  (
    n1152,
    n1096,
    n1098,
    n1061,
    n1074
  );


  nor
  g1138
  (
    n1201,
    n1007,
    n1080,
    n1021,
    n1093
  );


  nand
  g1139
  (
    n1191,
    n1020,
    n1099,
    n1018,
    n1055
  );


  xor
  g1140
  (
    n1147,
    n1052,
    n1068,
    n1054,
    n1072
  );


  or
  g1141
  (
    n1142,
    n1077,
    n1072,
    n775,
    n1071
  );


  xor
  g1142
  (
    n1166,
    n1104,
    n1078,
    n991,
    n1079
  );


  and
  g1143
  (
    n1137,
    n1060,
    n1044,
    n1010,
    n1063
  );


  xnor
  g1144
  (
    n1156,
    n1092,
    n1004,
    n1066,
    n1044
  );


  and
  g1145
  (
    n1163,
    n1005,
    n1080,
    n1103,
    n1009
  );


  nand
  g1146
  (
    n1122,
    n1053,
    n1064,
    n1062,
    n992
  );


  and
  g1147
  (
    n1114,
    n1102,
    n1011,
    n1066,
    n1073
  );


  xnor
  g1148
  (
    n1162,
    n1017,
    n1070,
    n1086,
    n1085
  );


  nor
  g1149
  (
    n1177,
    n1064,
    n1004,
    n1098,
    n1055
  );


  xnor
  g1150
  (
    n1126,
    n1079,
    n1094,
    n1045,
    n1092
  );


  or
  g1151
  (
    n1148,
    n1069,
    n1083,
    n1061,
    n1001
  );


  xnor
  g1152
  (
    n1112,
    n1074,
    n1082,
    n1060,
    n1052
  );


  nor
  g1153
  (
    n1175,
    n1078,
    n1065,
    n992,
    n1013
  );


  or
  g1154
  (
    n1145,
    n1077,
    n1015,
    n1047,
    n1052
  );


  nand
  g1155
  (
    n1196,
    n996,
    n1004,
    n1104,
    n1050
  );


  and
  g1156
  (
    n1184,
    n1077,
    n1082,
    n1076,
    n1048
  );


  or
  g1157
  (
    n1189,
    n993,
    n773,
    n1008,
    n1075
  );


  xor
  g1158
  (
    n1174,
    n994,
    n1103,
    n1083,
    n1003
  );


  and
  g1159
  (
    n1108,
    n999,
    n1079,
    n1007,
    n1043
  );


  and
  g1160
  (
    n1109,
    n1070,
    n774,
    n1065,
    n1054
  );


  nor
  g1161
  (
    n1150,
    n1103,
    n1019,
    n1016,
    n1050
  );


  and
  g1162
  (
    n1135,
    n776,
    n1101,
    n1087,
    n990
  );


  nand
  g1163
  (
    n1178,
    n1015,
    n1080,
    n1088,
    n1016
  );


  nand
  g1164
  (
    n1195,
    n1058,
    n1078,
    n993,
    n1089
  );


  nand
  g1165
  (
    n1204,
    n1063,
    n1048,
    n777,
    n1055
  );


  xor
  g1166
  (
    n1181,
    n1046,
    n1012,
    n1075,
    n1051
  );


  xnor
  g1167
  (
    n1186,
    n1019,
    n1050,
    n998,
    n1095
  );


  xnor
  g1168
  (
    n1185,
    n1105,
    n1066,
    n1101,
    n1102
  );


  xnor
  g1169
  (
    n1130,
    n1073,
    n1021,
    n1086,
    n1016
  );


  xnor
  g1170
  (
    n1168,
    n1056,
    n998,
    n1091,
    n1104
  );


  or
  g1171
  (
    n1199,
    n1014,
    n1090,
    n1056,
    n1081
  );


  and
  g1172
  (
    n1155,
    n1068,
    n1048,
    n993,
    n1086
  );


  xnor
  g1173
  (
    n1169,
    n777,
    n1018,
    n1090,
    n1051
  );


  xnor
  g1174
  (
    n1140,
    n1100,
    n1010,
    n1085,
    n1101
  );


  xor
  g1175
  (
    n1124,
    n1007,
    n1063,
    n1093,
    n990
  );


  nand
  g1176
  (
    n1107,
    n1071,
    n776,
    n1002,
    n1021
  );


  xnor
  g1177
  (
    n1192,
    n1013,
    n1013,
    n1106,
    n1046
  );


  nor
  g1178
  (
    n1161,
    n776,
    n1019,
    n1078,
    n1059
  );


  and
  g1179
  (
    n1110,
    n1074,
    n1000,
    n1005,
    n995
  );


  xor
  g1180
  (
    n1127,
    n1067,
    n1001,
    n1084
  );


  nor
  g1181
  (
    n1146,
    n1070,
    n1017,
    n1044,
    n775
  );


  and
  g1182
  (
    n1187,
    n1011,
    n1015,
    n994,
    n1067
  );


  and
  g1183
  (
    n1117,
    n1091,
    n1085,
    n1001,
    n1097
  );


  or
  g1184
  (
    n1180,
    n1093,
    n1057,
    n1015,
    n1096
  );


  nor
  g1185
  (
    n1176,
    n1003,
    n1002,
    n1058,
    n1065
  );


  nor
  g1186
  (
    n1211,
    n1126,
    n1133,
    n1136,
    n1110
  );


  nand
  g1187
  (
    n1222,
    n1134,
    n1132,
    n1135,
    n1119
  );


  and
  g1188
  (
    n1219,
    n1110,
    n1127,
    n1138,
    n1122
  );


  xnor
  g1189
  (
    n1215,
    n1125,
    n1138,
    n1115
  );


  xor
  g1190
  (
    n1220,
    n1139,
    n1108,
    n1121,
    n1138
  );


  and
  g1191
  (
    n1208,
    n1120,
    n1112,
    n1108,
    n1140
  );


  and
  g1192
  (
    n1214,
    n1140,
    n1138,
    n1136,
    n1129
  );


  and
  g1193
  (
    n1216,
    n1109,
    n1111,
    n1122,
    n1137
  );


  or
  g1194
  (
    KeyWire_0_20,
    n1116,
    n1133,
    n1128,
    n1130
  );


  nand
  g1195
  (
    n1218,
    n1118,
    n1134,
    n1130,
    n1121
  );


  and
  g1196
  (
    n1227,
    n1111,
    n1123,
    n1124,
    n1139
  );


  and
  g1197
  (
    n1221,
    n1109,
    n1128,
    n1116,
    n1139
  );


  nor
  g1198
  (
    n1209,
    n1140,
    n1131,
    n1137,
    n1107
  );


  nand
  g1199
  (
    n1213,
    n1112,
    n1125,
    n1133,
    n1113
  );


  xnor
  g1200
  (
    n1223,
    n1139,
    n1131,
    n1114
  );


  nor
  g1201
  (
    n1225,
    n1135,
    n1123,
    n1134,
    n1117
  );


  and
  g1202
  (
    n1210,
    n1129,
    n1140,
    n1137,
    n1120
  );


  or
  g1203
  (
    n1224,
    n1137,
    n1126,
    n1119,
    n1107
  );


  xor
  g1204
  (
    n1212,
    n1124,
    n1134,
    n1127,
    n1117
  );


  and
  g1205
  (
    n1207,
    n1135,
    n1136,
    n1118,
    n1113
  );


  and
  g1206
  (
    n1217,
    n1132,
    n1133,
    n1135,
    n1136
  );


  xnor
  g1207
  (
    n1242,
    n786,
    n784,
    n528,
    n777
  );


  nand
  g1208
  (
    n1238,
    n715,
    n1221,
    n878,
    n778
  );


  xnor
  g1209
  (
    n1246,
    n1220,
    n1211,
    n781,
    n825
  );


  xor
  g1210
  (
    n1228,
    n779,
    n1214,
    n528,
    n878
  );


  nand
  g1211
  (
    n1245,
    n785,
    n786,
    n1225,
    n778
  );


  nand
  g1212
  (
    n1231,
    n1216,
    n781,
    n780,
    n1219
  );


  nand
  g1213
  (
    n1248,
    n715,
    n784,
    n1210,
    n782
  );


  or
  g1214
  (
    n1237,
    n528,
    n783,
    n779,
    n789
  );


  nand
  g1215
  (
    n1236,
    n1213,
    n778,
    n786,
    n780
  );


  and
  g1216
  (
    n1247,
    n1223,
    n785,
    n1224,
    n788
  );


  and
  g1217
  (
    n1235,
    n788,
    n714,
    n787,
    n784
  );


  and
  g1218
  (
    n1234,
    n714,
    n784,
    n780,
    n787
  );


  xnor
  g1219
  (
    n1232,
    n789,
    n787,
    n1215,
    n715
  );


  xor
  g1220
  (
    n1229,
    n528,
    n1222,
    n1218,
    n778
  );


  nand
  g1221
  (
    n1240,
    n779,
    n825,
    n1227,
    n783
  );


  nor
  g1222
  (
    n1241,
    n1208,
    n780,
    n783,
    n779
  );


  nand
  g1223
  (
    n1249,
    n782,
    n785,
    n878,
    n1207
  );


  or
  g1224
  (
    n1244,
    n787,
    n1212,
    n1226,
    n824
  );


  and
  g1225
  (
    n1233,
    n782,
    n825,
    n1209,
    n781
  );


  xnor
  g1226
  (
    n1230,
    n715,
    n786,
    n783,
    n1227
  );


  xor
  g1227
  (
    n1243,
    n782,
    n789,
    n785,
    n825
  );


  nand
  g1228
  (
    n1239,
    n1217,
    n788,
    n781
  );


  xnor
  g1229
  (
    n1251,
    n1142,
    n1147,
    n1178,
    n1174
  );


  nor
  g1230
  (
    n1289,
    n1158,
    n1148,
    n1168,
    n1237
  );


  or
  g1231
  (
    n1297,
    n1232,
    n1235,
    n1175,
    n1228
  );


  and
  g1232
  (
    n1265,
    n1150,
    n1154,
    n1237,
    n1168
  );


  xor
  g1233
  (
    n1271,
    n1178,
    n1181,
    n1159,
    n1143
  );


  or
  g1234
  (
    n1279,
    n1241,
    n1152,
    n1156,
    n1166
  );


  nor
  g1235
  (
    n1275,
    n1163,
    n1148,
    n1246,
    n1244
  );


  or
  g1236
  (
    n1270,
    n1234,
    n1163,
    n1240,
    n1146
  );


  nor
  g1237
  (
    n1295,
    n1245,
    n1155,
    n1172,
    n1236
  );


  xnor
  g1238
  (
    n1285,
    n1242,
    n1228,
    n1148,
    n1247
  );


  or
  g1239
  (
    n1312,
    n1242,
    n1160,
    n1153,
    n1149
  );


  or
  g1240
  (
    n1304,
    n1153,
    n1181,
    n1167,
    n1247
  );


  nor
  g1241
  (
    n1264,
    n1180,
    n1143,
    n1159,
    n1173
  );


  or
  g1242
  (
    n1296,
    n1149,
    n1150,
    n1152,
    n1229
  );


  and
  g1243
  (
    n1260,
    n1160,
    n1154,
    n1155,
    n1238
  );


  nand
  g1244
  (
    n1259,
    n1241,
    n1158,
    n1172,
    n1231
  );


  and
  g1245
  (
    n1253,
    n1153,
    n1233,
    n1177,
    n1151
  );


  xor
  g1246
  (
    KeyWire_0_26,
    n1172,
    n1235,
    n1236,
    n1179
  );


  nor
  g1247
  (
    n1288,
    n1161,
    n914,
    n1231,
    n1141
  );


  and
  g1248
  (
    n1282,
    n1164,
    n1245,
    n1249,
    n1244
  );


  nor
  g1249
  (
    n1268,
    n1162,
    n1151,
    n1180,
    n1181
  );


  xor
  g1250
  (
    n1292,
    n1182,
    n1236,
    n1179,
    n1158
  );


  nor
  g1251
  (
    n1281,
    n1146,
    n1175,
    n1242,
    n1173
  );


  xor
  g1252
  (
    n1310,
    n1175,
    n1147,
    n1156,
    n1154
  );


  and
  g1253
  (
    n1298,
    n1161,
    n1157,
    n1160,
    n1234
  );


  xnor
  g1254
  (
    n1284,
    n1237,
    n1247,
    n1238,
    n1240
  );


  and
  g1255
  (
    KeyWire_0_30,
    n1141,
    n1239,
    n1178,
    n1167
  );


  or
  g1256
  (
    n1300,
    n1246,
    n1229,
    n1147
  );


  xor
  g1257
  (
    n1269,
    n1159,
    n1162,
    n1171,
    n1144
  );


  or
  g1258
  (
    n1276,
    n1171,
    n1248,
    n1176,
    n1244
  );


  and
  g1259
  (
    n1262,
    n1230,
    n1181,
    n1233,
    n1174
  );


  nor
  g1260
  (
    n1273,
    n1144,
    n1230,
    n1165,
    n1142
  );


  nand
  g1261
  (
    n1274,
    n1249,
    n1170,
    n1171,
    n1233
  );


  or
  g1262
  (
    n1278,
    n1164,
    n1162,
    n1233,
    n1239
  );


  and
  g1263
  (
    n1305,
    n1175,
    n1238,
    n1176,
    n1146
  );


  nor
  g1264
  (
    n1287,
    n1229,
    n1155,
    n1162,
    n1170
  );


  nand
  g1265
  (
    n1309,
    n1237,
    n1229,
    n1248,
    n1177
  );


  xnor
  g1266
  (
    n1302,
    n1176,
    n1231,
    n1182,
    n1157
  );


  and
  g1267
  (
    n1286,
    n1235,
    n1169,
    n1230,
    n1234
  );


  or
  g1268
  (
    KeyWire_0_6,
    n1179,
    n1243,
    n1150,
    n1144
  );


  xor
  g1269
  (
    n1250,
    n1164,
    n1150,
    n1173,
    n1239
  );


  or
  g1270
  (
    n1293,
    n1144,
    n1230,
    n1149,
    n1156
  );


  xor
  g1271
  (
    n1277,
    n1141,
    n1169,
    n1248,
    n1177
  );


  nor
  g1272
  (
    n1252,
    n1243,
    n1182,
    n1241,
    n1145
  );


  nand
  g1273
  (
    n1313,
    n1178,
    n1247,
    n1246,
    n1161
  );


  nor
  g1274
  (
    n1267,
    n1146,
    n1163,
    n1241,
    n1231
  );


  xnor
  g1275
  (
    n1283,
    n1143,
    n1228,
    n1166,
    n1157
  );


  nor
  g1276
  (
    n1261,
    n1232,
    n1235,
    n1170,
    n1157
  );


  nand
  g1277
  (
    n1307,
    n1168,
    n1180,
    n1148,
    n1166
  );


  xnor
  g1278
  (
    n1266,
    n1174,
    n1159,
    n1176,
    n1249
  );


  and
  g1279
  (
    n1257,
    n1153,
    n1166,
    n1177,
    n1156
  );


  xnor
  g1280
  (
    n1255,
    n1243,
    n1248,
    n1163,
    n1232
  );


  xor
  g1281
  (
    n1301,
    n1173,
    n1167,
    n1170,
    n1234
  );


  nand
  g1282
  (
    n1280,
    n1152,
    n1142,
    n1171,
    n1167
  );


  nand
  g1283
  (
    n1299,
    n1142,
    n1232,
    n1242,
    n1168
  );


  or
  g1284
  (
    n1256,
    n1145,
    n1169,
    n1165,
    n1240
  );


  xnor
  g1285
  (
    n1291,
    n1249,
    n1240,
    n1228,
    n1238
  );


  or
  g1286
  (
    n1306,
    n1155,
    n1164,
    n1245,
    n1243
  );


  nand
  g1287
  (
    n1254,
    n1172,
    n1165,
    n1151
  );


  or
  g1288
  (
    n1308,
    n1239,
    n1245,
    n1161,
    n1160
  );


  xor
  g1289
  (
    n1263,
    n1180,
    n1145,
    n1244,
    n1143
  );


  nand
  g1290
  (
    n1311,
    n1149,
    n1152,
    n1174,
    n1158
  );


  xnor
  g1291
  (
    n1290,
    n1179,
    n1141,
    n1236,
    n1145
  );


  or
  g1292
  (
    n1294,
    n1151,
    n1154,
    n1246,
    n1169
  );


  not
  g1293
  (
    n1326,
    n1301
  );


  buf
  g1294
  (
    n1317,
    n1301
  );


  not
  g1295
  (
    n1315,
    n1274
  );


  not
  g1296
  (
    n1319,
    n1281
  );


  not
  g1297
  (
    n1330,
    n1286
  );


  buf
  g1298
  (
    n1336,
    n1295
  );


  not
  g1299
  (
    n1339,
    n1293
  );


  buf
  g1300
  (
    n1320,
    n1259
  );


  not
  g1301
  (
    n1321,
    n1267
  );


  not
  g1302
  (
    n1314,
    n1250
  );


  buf
  g1303
  (
    n1337,
    n1299
  );


  not
  g1304
  (
    n1340,
    n1255
  );


  buf
  g1305
  (
    n1325,
    n1303
  );


  buf
  g1306
  (
    n1335,
    n1291
  );


  not
  g1307
  (
    n1331,
    n1251
  );


  nand
  g1308
  (
    n1338,
    n1273,
    n1285
  );


  nor
  g1309
  (
    n1344,
    n1272,
    n1292,
    n1270
  );


  xnor
  g1310
  (
    n1322,
    n1275,
    n1253,
    n1268
  );


  xnor
  g1311
  (
    n1324,
    n1304,
    n1264,
    n1276
  );


  nand
  g1312
  (
    n1334,
    n1269,
    n1289,
    n1283
  );


  or
  g1313
  (
    n1342,
    n1304,
    n1284,
    n1278
  );


  nand
  g1314
  (
    n1343,
    n1266,
    n1261,
    n1300
  );


  nand
  g1315
  (
    n1341,
    n1265,
    n1279,
    n1298
  );


  nand
  g1316
  (
    KeyWire_0_21,
    n1252,
    n1299,
    n1256
  );


  or
  g1317
  (
    n1323,
    n1290,
    n1263,
    n1302
  );


  nor
  g1318
  (
    n1332,
    n1300,
    n1271,
    n1302
  );


  nand
  g1319
  (
    n1333,
    n1277,
    n1260,
    n1258
  );


  and
  g1320
  (
    n1316,
    n1296,
    n1298,
    n1282
  );


  nor
  g1321
  (
    n1329,
    n1297,
    n1303,
    n1262
  );


  nor
  g1322
  (
    n1327,
    n1254,
    n1280,
    n1287
  );


  xnor
  g1323
  (
    n1318,
    n1288,
    n1294,
    n1257
  );


  nand
  g1324
  (
    n1353,
    n1328,
    n1315,
    n1314,
    n1316
  );


  nand
  g1325
  (
    n1348,
    n1323,
    n1321,
    n1315,
    n1325
  );


  nand
  g1326
  (
    n1345,
    n1323,
    n1324,
    n1329,
    n1319
  );


  xor
  g1327
  (
    n1350,
    n1327,
    n1317,
    n1324,
    n1320
  );


  and
  g1328
  (
    n1355,
    n1329,
    n1327,
    n1320,
    n1318
  );


  nand
  g1329
  (
    n1356,
    n1322,
    n1325,
    n1324,
    n1321
  );


  and
  g1330
  (
    n1352,
    n1316,
    n1319,
    n1320,
    n1315
  );


  and
  g1331
  (
    n1347,
    n1325,
    n1317,
    n1326,
    n1314
  );


  xor
  g1332
  (
    n1354,
    n1326,
    n1317,
    n1318,
    n1329
  );


  nand
  g1333
  (
    n1349,
    n1328,
    n1328,
    n1323,
    n1321
  );


  xnor
  g1334
  (
    n1351,
    n1326,
    n1316,
    n1322,
    n1314
  );


  nor
  g1335
  (
    n1346,
    n1322,
    n1319,
    n1327,
    n1318
  );


  or
  g1336
  (
    n1359,
    n915,
    n915,
    n1354,
    n1353
  );


  nor
  g1337
  (
    n1357,
    n919,
    n919,
    n917,
    n1356
  );


  xor
  g1338
  (
    n1358,
    n1355,
    n918,
    n920
  );


  and
  g1339
  (
    n1360,
    n917,
    n916,
    n918
  );


  and
  g1340
  (
    n1362,
    n1329,
    n1358,
    n1360,
    n1334
  );


  nor
  g1341
  (
    n1367,
    n1333,
    n1360,
    n1335,
    n1357
  );


  nor
  g1342
  (
    n1371,
    n1331,
    n1331,
    n678,
    n1358
  );


  or
  g1343
  (
    n1363,
    n1360,
    n1357,
    n1332,
    n1331
  );


  xnor
  g1344
  (
    n1373,
    n1330,
    n1358,
    n1359,
    n1335
  );


  xnor
  g1345
  (
    n1372,
    n493,
    n1359
  );


  xor
  g1346
  (
    n1364,
    n1358,
    n1336,
    n1332,
    n1330
  );


  xnor
  g1347
  (
    n1365,
    n492,
    n493,
    n1330,
    n1334
  );


  xor
  g1348
  (
    n1366,
    n1357,
    n1360,
    n680,
    n1336
  );


  nor
  g1349
  (
    n1368,
    n1330,
    n1333,
    n1335,
    n493
  );


  and
  g1350
  (
    n1369,
    n1332,
    n1333,
    n1335,
    n492
  );


  and
  g1351
  (
    n1370,
    n1331,
    n1357,
    n1334,
    n1359
  );


  and
  g1352
  (
    n1361,
    n1336,
    n1332,
    n1333,
    n1334
  );


  xnor
  g1353
  (
    n1395,
    n1366,
    n931,
    n927
  );


  xnor
  g1354
  (
    n1388,
    n931,
    n921,
    n924,
    n941
  );


  xor
  g1355
  (
    n1387,
    n940,
    n920,
    n1362,
    n928
  );


  nor
  g1356
  (
    n1379,
    n924,
    n936,
    n1373,
    n938
  );


  xor
  g1357
  (
    n1402,
    n1362,
    n1363,
    n922,
    n938
  );


  xor
  g1358
  (
    n1392,
    n935,
    n924,
    n927
  );


  xnor
  g1359
  (
    n1377,
    n937,
    n926,
    n1372
  );


  nand
  g1360
  (
    n1404,
    n935,
    n934,
    n932,
    n942
  );


  nand
  g1361
  (
    n1397,
    n1363,
    n943,
    n940,
    n942
  );


  xor
  g1362
  (
    n1389,
    n939,
    n927,
    n928
  );


  xnor
  g1363
  (
    n1403,
    n923,
    n940,
    n938,
    n929
  );


  or
  g1364
  (
    n1375,
    n938,
    n941,
    n932,
    n939
  );


  xor
  g1365
  (
    n1383,
    n1364,
    n1373,
    n932,
    n942
  );


  nor
  g1366
  (
    n1399,
    n935,
    n1365,
    n923,
    n942
  );


  xor
  g1367
  (
    n1384,
    n941,
    n936,
    n929,
    n922
  );


  xnor
  g1368
  (
    n1385,
    n929,
    n1371,
    n926,
    n940
  );


  xor
  g1369
  (
    n1400,
    n926,
    n930,
    n1373,
    n1361
  );


  and
  g1370
  (
    n1382,
    n930,
    n1369,
    n927,
    n939
  );


  nor
  g1371
  (
    n1381,
    n1370,
    n929,
    n936,
    n921
  );


  nor
  g1372
  (
    n1393,
    n934,
    n933,
    n922,
    n1367
  );


  xor
  g1373
  (
    n1378,
    n935,
    n923,
    n921,
    n941
  );


  nand
  g1374
  (
    n1398,
    n921,
    n926,
    n934,
    n1370
  );


  xor
  g1375
  (
    n1386,
    n1371,
    n1368,
    n936,
    n937
  );


  xnor
  g1376
  (
    n1396,
    n937,
    n925,
    n1368
  );


  and
  g1377
  (
    n1391,
    n1371,
    n1373,
    n930,
    n931
  );


  xor
  g1378
  (
    n1380,
    n923,
    n1365,
    n1369,
    n933
  );


  xnor
  g1379
  (
    n1394,
    n937,
    n925,
    n933,
    n934
  );


  nand
  g1380
  (
    n1401,
    n932,
    n1372,
    n1370,
    n933
  );


  xor
  g1381
  (
    n1374,
    n928,
    n925,
    n930,
    n1366
  );


  and
  g1382
  (
    n1390,
    n1367,
    n1369,
    n1368,
    n922
  );


  nand
  g1383
  (
    n1376,
    n1364,
    n920,
    n1361,
    n939
  );


  buf
  g1384
  (
    n1407,
    n1374
  );


  buf
  g1385
  (
    n1405,
    n1376
  );


  nand
  g1386
  (
    n1406,
    n1377,
    n1375
  );


  nor
  g1387
  (
    n1409,
    n1394,
    n1390,
    n1406
  );


  or
  g1388
  (
    n1419,
    n1407,
    n1393
  );


  or
  g1389
  (
    n1408,
    n1407,
    n1389,
    n1398,
    n1380
  );


  xor
  g1390
  (
    n1417,
    n1405,
    n1406,
    n989
  );


  nand
  g1391
  (
    n1410,
    n1391,
    n1394,
    n1395,
    n989
  );


  xnor
  g1392
  (
    n1411,
    n1405,
    n1391,
    n1381,
    n1399
  );


  xnor
  g1393
  (
    n1414,
    n1392,
    n1388,
    n1383,
    n1397
  );


  nor
  g1394
  (
    n1415,
    n878,
    n1405,
    n1387,
    n1392
  );


  or
  g1395
  (
    n1413,
    n1386,
    n1382,
    n1399,
    n1379
  );


  xor
  g1396
  (
    n1418,
    n1396,
    n1385,
    n1384,
    n1407
  );


  xor
  g1397
  (
    n1416,
    n1405,
    n1396,
    n943,
    n989
  );


  nand
  g1398
  (
    n1412,
    n1397,
    n1378,
    n1395,
    n1398
  );


  nand
  g1399
  (
    n1435,
    n1417,
    n1193,
    n1408,
    n1401
  );


  xnor
  g1400
  (
    n1434,
    n1188,
    n1186,
    n1192,
    n1191
  );


  xnor
  g1401
  (
    n1433,
    n1419,
    n1192,
    n1188
  );


  nor
  g1402
  (
    n1422,
    n1414,
    n1189,
    n1187,
    n1193
  );


  nor
  g1403
  (
    n1420,
    n1186,
    n1190,
    n1418
  );


  and
  g1404
  (
    n1427,
    n1187,
    n1188,
    n1400,
    n1193
  );


  nand
  g1405
  (
    n1425,
    n1187,
    n1183,
    n1189,
    n1190
  );


  and
  g1406
  (
    n1426,
    n1183,
    n1186,
    n1417
  );


  xor
  g1407
  (
    n1424,
    n1185,
    n1183,
    n1189,
    n1184
  );


  or
  g1408
  (
    n1430,
    n1419,
    n1189,
    n1184,
    n1413
  );


  xnor
  g1409
  (
    n1432,
    n1190,
    n1400,
    n1416
  );


  xnor
  g1410
  (
    n1428,
    n1191,
    n1409,
    n1192,
    n1184
  );


  xor
  g1411
  (
    n1431,
    n1401,
    n1184,
    n1183,
    n1418
  );


  xor
  g1412
  (
    n1421,
    n1412,
    n1191,
    n1415,
    n1185
  );


  nand
  g1413
  (
    n1423,
    n1182,
    n1187,
    n1192,
    n1410
  );


  xor
  g1414
  (
    n1429,
    n1411,
    n1185,
    n1191
  );


  not
  g1415
  (
    n1443,
    n1309
  );


  buf
  g1416
  (
    n1461,
    n1424
  );


  buf
  g1417
  (
    n1451,
    n1426
  );


  buf
  g1418
  (
    n1436,
    n1427
  );


  not
  g1419
  (
    n1457,
    n1428
  );


  buf
  g1420
  (
    n1438,
    n1425
  );


  not
  g1421
  (
    n1459,
    n1428
  );


  buf
  g1422
  (
    n1440,
    n1306
  );


  not
  g1423
  (
    n1449,
    n1424
  );


  not
  g1424
  (
    n1437,
    n1428
  );


  not
  g1425
  (
    n1456,
    n1420
  );


  buf
  g1426
  (
    n1446,
    n1306
  );


  not
  g1427
  (
    n1441,
    n1421
  );


  buf
  g1428
  (
    n1450,
    n1428
  );


  not
  g1429
  (
    n1439,
    n1422
  );


  buf
  g1430
  (
    n1462,
    n1424
  );


  buf
  g1431
  (
    n1445,
    n1421
  );


  buf
  g1432
  (
    n1458,
    n1426
  );


  nand
  g1433
  (
    n1455,
    n1424,
    n1429,
    n1308,
    n1427
  );


  nor
  g1434
  (
    n1453,
    n1310,
    n1423,
    n1422,
    n1305
  );


  nor
  g1435
  (
    n1442,
    n1429,
    n1309,
    n1420,
    n1425
  );


  nor
  g1436
  (
    n1460,
    n1426,
    n1427,
    n1402,
    n1429
  );


  and
  g1437
  (
    n1447,
    n1420,
    n1421,
    n1423,
    n1426
  );


  and
  g1438
  (
    n1452,
    n1420,
    n1308,
    n1307,
    n1427
  );


  xnor
  g1439
  (
    n1448,
    n1403,
    n1422,
    n1429,
    n1423
  );


  xnor
  g1440
  (
    n1454,
    n1422,
    n1421,
    n1402,
    n1305
  );


  xnor
  g1441
  (
    n1444,
    n1423,
    n1425,
    n1307
  );


  nand
  g1442
  (
    n1468,
    n1446,
    n1436,
    n1452,
    n1444
  );


  xnor
  g1443
  (
    n1467,
    n1451,
    n1448,
    n1450,
    n1446
  );


  xor
  g1444
  (
    n1464,
    n1448,
    n1445,
    n1440,
    n1438
  );


  nand
  g1445
  (
    n1465,
    n1439,
    n1441,
    n1447,
    n1450
  );


  and
  g1446
  (
    n1463,
    n1437,
    n1442,
    n1447,
    n1443
  );


  nand
  g1447
  (
    n1466,
    n1452,
    n1449,
    n1451
  );


  xor
  g1448
  (
    n1488,
    n1312,
    n1463,
    n948,
    n957
  );


  and
  g1449
  (
    n1487,
    n958,
    n945,
    n1311,
    n951
  );


  xnor
  g1450
  (
    n1483,
    n956,
    n1464,
    n951,
    n954
  );


  xor
  g1451
  (
    n1480,
    n956,
    n1466,
    n945,
    n1463
  );


  xnor
  g1452
  (
    n1475,
    n946,
    n956,
    n1467,
    n947
  );


  nand
  g1453
  (
    n1469,
    n1468,
    n949,
    n1465,
    n1311
  );


  or
  g1454
  (
    n1474,
    n954,
    n951,
    n952,
    n949
  );


  nor
  g1455
  (
    n1477,
    n1463,
    n958,
    n955,
    n948
  );


  nor
  g1456
  (
    n1482,
    n1465,
    n944,
    n1466,
    n950
  );


  xnor
  g1457
  (
    n1476,
    n946,
    n1466,
    n1313,
    n950
  );


  or
  g1458
  (
    n1491,
    n1468,
    n954,
    n958,
    n952
  );


  nand
  g1459
  (
    n1484,
    n956,
    n952,
    n953,
    n957
  );


  or
  g1460
  (
    n1492,
    n944,
    n957,
    n1312,
    n1313
  );


  xnor
  g1461
  (
    n1485,
    n1465,
    n951,
    n949,
    n947
  );


  nor
  g1462
  (
    n1486,
    n1465,
    n953,
    n1313,
    n955
  );


  or
  g1463
  (
    n1479,
    n1312,
    n1311,
    n1467,
    n944
  );


  and
  g1464
  (
    n1470,
    n1468,
    n952,
    n945,
    n957
  );


  and
  g1465
  (
    n1472,
    n955,
    n955,
    n1466,
    n948
  );


  or
  g1466
  (
    n1471,
    n949,
    n946,
    n1467,
    n1464
  );


  or
  g1467
  (
    n1473,
    n954,
    n944,
    n958,
    n1468
  );


  xnor
  g1468
  (
    n1490,
    n1464,
    n953,
    n947
  );


  nor
  g1469
  (
    n1481,
    n943,
    n1310,
    n950,
    n946
  );


  and
  g1470
  (
    n1489,
    n950,
    n1463,
    n945,
    n1467
  );


  or
  g1471
  (
    n1478,
    n948,
    n947,
    n1464,
    n943
  );


  xor
  g1472
  (
    n1510,
    n1472,
    n1491,
    n1470
  );


  xor
  g1473
  (
    n1519,
    n1489,
    n1474,
    n1336,
    n1483
  );


  xnor
  g1474
  (
    n1517,
    n1490,
    n1483,
    n1492,
    n1339
  );


  xor
  g1475
  (
    KeyWire_0_7,
    n1483,
    n1337,
    n1486,
    n1480
  );


  nor
  g1476
  (
    n1511,
    n1471,
    n1489,
    n1338,
    n1480
  );


  and
  g1477
  (
    n1508,
    n1476,
    n1478,
    n1454,
    n1339
  );


  nand
  g1478
  (
    n1504,
    n1338,
    n1491,
    n1479,
    n1469
  );


  and
  g1479
  (
    n1512,
    n1341,
    n1456,
    n1475,
    n1472
  );


  xnor
  g1480
  (
    n1520,
    n1474,
    n1478,
    n1479,
    n1486
  );


  nor
  g1481
  (
    n1497,
    n1469,
    n1487,
    n1481,
    n1341
  );


  nor
  g1482
  (
    n1507,
    n1491,
    n1477,
    n1492,
    n1481
  );


  and
  g1483
  (
    n1514,
    n1343,
    n1472,
    n1453,
    n1476
  );


  xnor
  g1484
  (
    n1509,
    n1339,
    n1479,
    n1481,
    n1480
  );


  and
  g1485
  (
    n1495,
    n1340,
    n1344,
    n1489,
    n1455
  );


  nor
  g1486
  (
    n1498,
    n1492,
    n1344,
    n1473,
    n1470
  );


  xor
  g1487
  (
    n1525,
    n1342,
    n1488,
    n1473,
    n1337
  );


  or
  g1488
  (
    n1521,
    n1342,
    n1475,
    n1454,
    n1487
  );


  nor
  g1489
  (
    n1494,
    n1344,
    n1485,
    n1484,
    n1482
  );


  and
  g1490
  (
    n1496,
    n1340,
    n1473,
    n1482,
    n1488
  );


  nor
  g1491
  (
    n1523,
    n1484,
    n1487,
    n1472,
    n1488
  );


  and
  g1492
  (
    n1526,
    n1475,
    n1338,
    n1477,
    n1474
  );


  or
  g1493
  (
    n1522,
    n1486,
    n1476,
    n1478
  );


  or
  g1494
  (
    n1524,
    n1490,
    n1474,
    n1482,
    n1491
  );


  and
  g1495
  (
    n1501,
    n1484,
    n1471,
    n1475,
    n1479
  );


  nand
  g1496
  (
    n1500,
    n1482,
    n1342,
    n1343
  );


  xor
  g1497
  (
    n1506,
    n1340,
    n1485,
    n1488,
    n1341
  );


  or
  g1498
  (
    n1505,
    n1341,
    n1338,
    n1340,
    n1483
  );


  xor
  g1499
  (
    n1503,
    n1478,
    n1469,
    n1481,
    n1487
  );


  and
  g1500
  (
    n1499,
    n1455,
    n1473,
    n1337,
    n1484
  );


  or
  g1501
  (
    n1515,
    n1339,
    n1480,
    n1453,
    n1486
  );


  xor
  g1502
  (
    n1502,
    n1490,
    n1489,
    n1485,
    n1471
  );


  nand
  g1503
  (
    n1518,
    n1471,
    n1344,
    n1342,
    n1343
  );


  xor
  g1504
  (
    n1493,
    n1337,
    n1490,
    n1469,
    n1477
  );


  xnor
  g1505
  (
    n1516,
    n1485,
    n1492,
    n1477,
    n1470
  );


  xor
  g1506
  (
    n1527,
    n406,
    n1524,
    n1513,
    n408
  );


  nor
  g1507
  (
    KeyWire_0_16,
    n1494,
    n1435,
    n435
  );


  and
  g1508
  (
    n1594,
    n400,
    n1495,
    n418,
    n431
  );


  nand
  g1509
  (
    n1529,
    n401,
    n1496,
    n432,
    n1511
  );


  and
  g1510
  (
    KeyWire_0_4,
    n434,
    n424,
    n1523,
    n401
  );


  or
  g1511
  (
    n1544,
    n414,
    n1515,
    n1430,
    n1501
  );


  xnor
  g1512
  (
    n1540,
    n397,
    n442,
    n1508,
    n407
  );


  xnor
  g1513
  (
    n1600,
    n428,
    n416,
    n403,
    n1511
  );


  nor
  g1514
  (
    n1564,
    n441,
    n1514,
    n405,
    n434
  );


  nor
  g1515
  (
    n1560,
    n399,
    n439,
    n1494,
    n1522
  );


  nand
  g1516
  (
    KeyWire_0_31,
    n1518,
    n421,
    n1519,
    n427
  );


  xnor
  g1517
  (
    n1593,
    n1493,
    n1500,
    n1519,
    n409
  );


  nor
  g1518
  (
    n1542,
    n405,
    n1501,
    n1513,
    n411
  );


  xnor
  g1519
  (
    n1531,
    n406,
    n1515,
    n1526,
    n408
  );


  xnor
  g1520
  (
    n1605,
    n1515,
    n1526,
    n410,
    n430
  );


  xor
  g1521
  (
    n1603,
    n1435,
    n1511,
    n426,
    n1518
  );


  xor
  g1522
  (
    n1578,
    n407,
    n422,
    n430,
    n402
  );


  xor
  g1523
  (
    n1576,
    n426,
    n441,
    n1524,
    n1432
  );


  xor
  g1524
  (
    n1547,
    n1495,
    n417,
    n1517,
    n1509
  );


  and
  g1525
  (
    n1565,
    n1434,
    n1516,
    n398,
    n415
  );


  or
  g1526
  (
    KeyWire_0_9,
    n436,
    n400,
    n408,
    n1523
  );


  nor
  g1527
  (
    n1571,
    n1522,
    n432,
    n1508,
    n429
  );


  xnor
  g1528
  (
    n1536,
    n1521,
    n1513,
    n424,
    n425
  );


  xor
  g1529
  (
    n1546,
    n1514,
    n405,
    n425,
    n1507
  );


  xnor
  g1530
  (
    n1587,
    n412,
    n415,
    n1517,
    n1519
  );


  xnor
  g1531
  (
    n1572,
    n436,
    n428,
    n1522,
    n1434
  );


  xor
  g1532
  (
    n1598,
    n1431,
    n414,
    n1521,
    n1510
  );


  and
  g1533
  (
    n1555,
    n1513,
    n1433,
    n427,
    n439
  );


  and
  g1534
  (
    n1588,
    n404,
    n441,
    n424,
    n418
  );


  and
  g1535
  (
    n1539,
    n429,
    n438,
    n416,
    n421
  );


  xnor
  g1536
  (
    n1533,
    n412,
    n1431,
    n19,
    n402
  );


  nand
  g1537
  (
    n1592,
    n1521,
    n430,
    n1434,
    n421
  );


  nor
  g1538
  (
    n1573,
    n423,
    n439,
    n1498,
    n422
  );


  xor
  g1539
  (
    n1590,
    n406,
    n1516,
    n403,
    n18
  );


  or
  g1540
  (
    n1554,
    n422,
    n414,
    n438,
    n1500
  );


  and
  g1541
  (
    n1566,
    n17,
    n407,
    n1510,
    n435
  );


  xor
  g1542
  (
    n1581,
    n437,
    n1430,
    n403,
    n1520
  );


  or
  g1543
  (
    n1538,
    n1431,
    n1525,
    n412
  );


  and
  g1544
  (
    n1589,
    n417,
    n415,
    n1499,
    n1496
  );


  and
  g1545
  (
    n1553,
    n1525,
    n440,
    n411,
    n437
  );


  or
  g1546
  (
    n1559,
    n1431,
    n405,
    n419,
    n1432
  );


  or
  g1547
  (
    n1602,
    n413,
    n400,
    n1510,
    n1512
  );


  nand
  g1548
  (
    n1545,
    n1504,
    n1506,
    n1505,
    n1430
  );


  nor
  g1549
  (
    n1556,
    n1507,
    n1516,
    n411,
    n420
  );


  nor
  g1550
  (
    n1530,
    n1504,
    n431,
    n789,
    n1435
  );


  nor
  g1551
  (
    n1586,
    n1521,
    n1523,
    n1526,
    n432
  );


  or
  g1552
  (
    KeyWire_0_8,
    n1516,
    n431,
    n433,
    n1524
  );


  or
  g1553
  (
    n1541,
    n407,
    n19,
    n421,
    n1493
  );


  xnor
  g1554
  (
    n1563,
    n1497,
    n1512,
    n1517,
    n1498
  );


  xnor
  g1555
  (
    n1567,
    n434,
    n419,
    n409,
    n415
  );


  or
  g1556
  (
    n1597,
    n420,
    n1499,
    n435,
    n399
  );


  nand
  g1557
  (
    n1601,
    n18,
    n1434,
    n432,
    n423
  );


  nor
  g1558
  (
    n1582,
    n436,
    n398,
    n399,
    n401
  );


  nand
  g1559
  (
    n1596,
    n1505,
    n417,
    n397,
    n438
  );


  xnor
  g1560
  (
    KeyWire_0_12,
    n410,
    n1515,
    n1432,
    n440
  );


  nor
  g1561
  (
    n1537,
    n439,
    n403,
    n1517,
    n422
  );


  nand
  g1562
  (
    n1569,
    n1526,
    n428,
    n436,
    n19
  );


  nor
  g1563
  (
    n1591,
    n426,
    n1520,
    n423,
    n1433
  );


  xnor
  g1564
  (
    n1599,
    n425,
    n1430,
    n401,
    n1433
  );


  nand
  g1565
  (
    n1585,
    n406,
    n433,
    n402,
    n1503
  );


  nand
  g1566
  (
    n1562,
    n433,
    n1514,
    n398,
    n429
  );


  and
  g1567
  (
    n1558,
    n18,
    n1502,
    n424,
    n425
  );


  nor
  g1568
  (
    n1551,
    n427,
    n438,
    n400,
    n437
  );


  nor
  g1569
  (
    n1534,
    n413,
    n1509,
    n418,
    n1511
  );


  xnor
  g1570
  (
    n1580,
    n437,
    n1520,
    n413,
    n1512
  );


  nor
  g1571
  (
    n1548,
    n417,
    n1518,
    n413,
    n1522
  );


  and
  g1572
  (
    n1595,
    n440,
    n442,
    n434,
    n1519
  );


  nand
  g1573
  (
    n1561,
    n410,
    n18,
    n404,
    n427
  );


  xnor
  g1574
  (
    n1574,
    n430,
    n412,
    n416,
    n411
  );


  and
  g1575
  (
    n1604,
    n404,
    n1524,
    n429,
    n1518
  );


  nand
  g1576
  (
    n1549,
    n1433,
    n431,
    n442,
    n1502
  );


  xor
  g1577
  (
    n1568,
    n1512,
    n428,
    n1525,
    n414
  );


  nand
  g1578
  (
    n1528,
    n402,
    n1506,
    n441,
    n433
  );


  and
  g1579
  (
    n1557,
    n1497,
    n1514,
    n419,
    n408
  );


  or
  g1580
  (
    n1577,
    n410,
    n420,
    n416,
    n1503
  );


  or
  g1581
  (
    n1552,
    n426,
    n418,
    n399,
    n409
  );


  xor
  g1582
  (
    n1535,
    n1520,
    n404,
    n419,
    n1432
  );


  xor
  g1583
  (
    n1584,
    n420,
    n397,
    n423,
    n435
  );


  or
  g1584
  (
    n1579,
    n440,
    n1523,
    n398,
    n409
  );


  xor
  g1585
  (
    n1606,
    n1530,
    n1528,
    n1529,
    n1527
  );


  or
  g1586
  (
    n1609,
    n853,
    n854,
    n1606,
    n857
  );


  nand
  g1587
  (
    n1607,
    n852,
    n852,
    n1606,
    n857
  );


  nor
  g1588
  (
    n1608,
    n855,
    n1606
  );


  nand
  g1589
  (
    n1610,
    n853,
    n854,
    n856
  );


  xnor
  g1590
  (
    n1612,
    n1533,
    n1608,
    n1609,
    n1404
  );


  xnor
  g1591
  (
    n1614,
    n1607,
    n1534,
    n1608,
    n1532
  );


  nand
  g1592
  (
    n1611,
    n1403,
    n1609,
    n1535,
    n1607
  );


  nand
  g1593
  (
    n1613,
    n1608,
    n1531,
    n1609
  );


  xor
  g1594
  (
    n1618,
    n1539,
    n1538,
    n1614,
    n1541
  );


  and
  g1595
  (
    n1617,
    n1613,
    n20
  );


  xor
  g1596
  (
    n1616,
    n1540,
    n1611,
    n1542,
    n1537
  );


  xor
  g1597
  (
    n1615,
    n20,
    n1536,
    n19,
    n1612
  );


  xor
  g1598
  (
    n1632,
    n1615,
    n1553,
    n1618,
    n1581
  );


  xor
  g1599
  (
    n1624,
    n1616,
    n1575,
    n1586,
    n1552
  );


  and
  g1600
  (
    n1629,
    n1567,
    n1617,
    n1571,
    n1568
  );


  or
  g1601
  (
    n1633,
    n1617,
    n1564,
    n1583,
    n1582
  );


  xor
  g1602
  (
    n1628,
    n1574,
    n1546,
    n1566,
    n1544
  );


  and
  g1603
  (
    n1622,
    n1590,
    n1617,
    n1569,
    n1558
  );


  xnor
  g1604
  (
    n1621,
    n1562,
    n1565,
    n1618,
    n1580
  );


  xor
  g1605
  (
    n1634,
    n1548,
    n1554,
    n1618,
    n1587
  );


  xnor
  g1606
  (
    n1631,
    n1616,
    n1579,
    n1585,
    n1577
  );


  nor
  g1607
  (
    n1630,
    n1556,
    n1616,
    n1588,
    n1543
  );


  xnor
  g1608
  (
    n1620,
    n1560,
    n1549,
    n1576,
    n1557
  );


  xnor
  g1609
  (
    n1626,
    n1615,
    n1573,
    n1584,
    n1555
  );


  xnor
  g1610
  (
    n1627,
    n1563,
    n1570,
    n1561,
    n1589
  );


  or
  g1611
  (
    n1625,
    n1578,
    n1572,
    n1550,
    n1617
  );


  xnor
  g1612
  (
    KeyWire_0_2,
    n1615,
    n1618,
    n1551,
    n1559
  );


  and
  g1613
  (
    n1619,
    n1615,
    n1616,
    n1545,
    n1547
  );


  xor
  g1614
  (
    n1644,
    n1195,
    n1202,
    n1629,
    n1199
  );


  and
  g1615
  (
    n1658,
    n1204,
    n1630,
    n1623,
    n1196
  );


  or
  g1616
  (
    n1641,
    n1202,
    n1621,
    n1201,
    n1631
  );


  nor
  g1617
  (
    n1657,
    n1195,
    n1632,
    n1200,
    n1629
  );


  nand
  g1618
  (
    n1635,
    n1205,
    n1198,
    n1622,
    n1204
  );


  or
  g1619
  (
    n1648,
    n1633,
    n1206,
    n1622
  );


  xnor
  g1620
  (
    n1646,
    n1199,
    n1197,
    n1203,
    n1205
  );


  xor
  g1621
  (
    n1638,
    n1628,
    n1626,
    n1619,
    n1194
  );


  xor
  g1622
  (
    n1645,
    n1200,
    n1195,
    n1194,
    n1620
  );


  or
  g1623
  (
    n1651,
    n1206,
    n1204,
    n1624,
    n1625
  );


  and
  g1624
  (
    n1643,
    n1627,
    n1201,
    n1196,
    n1193
  );


  nand
  g1625
  (
    n1640,
    n1201,
    n1205,
    n1621,
    n1199
  );


  or
  g1626
  (
    n1636,
    n1619,
    n1626,
    n1204,
    n1628
  );


  nand
  g1627
  (
    n1654,
    n1627,
    n1203,
    n1631,
    n1625
  );


  nand
  g1628
  (
    n1649,
    n54,
    n1630,
    n1621,
    n1203
  );


  or
  g1629
  (
    n1653,
    n1205,
    n1622,
    n1202,
    n1620
  );


  nor
  g1630
  (
    n1642,
    n1198,
    n1202,
    n1197,
    n1629
  );


  and
  g1631
  (
    n1647,
    n1623,
    n1623,
    n1201,
    n1624
  );


  nor
  g1632
  (
    n1650,
    n1632,
    n1196,
    n1197,
    n1625
  );


  nand
  g1633
  (
    n1639,
    n1200,
    n1628,
    n1197,
    n1198
  );


  and
  g1634
  (
    n1652,
    n1200,
    n1196,
    n1632,
    n1620
  );


  xnor
  g1635
  (
    n1637,
    n1194,
    n1206,
    n1203,
    n1626
  );


  or
  g1636
  (
    n1656,
    n1630,
    n1194,
    n1627,
    n1624
  );


  nor
  g1637
  (
    KeyWire_0_13,
    n1199,
    n1195,
    n1198,
    n1631
  );


  xnor
  g1638
  (
    n1670,
    n1639,
    n1650,
    n1602,
    n1653
  );


  nand
  g1639
  (
    n1666,
    n1593,
    n1652,
    n1636,
    n1657
  );


  nand
  g1640
  (
    n1665,
    n1460,
    n1647,
    n1458,
    n1656
  );


  nor
  g1641
  (
    n1662,
    n1610,
    n1648,
    n1594,
    n1654
  );


  xnor
  g1642
  (
    n1664,
    n1595,
    n1643,
    n1458,
    n1459
  );


  nand
  g1643
  (
    n1667,
    n1654,
    n1457,
    n1596,
    n1603
  );


  nor
  g1644
  (
    n1660,
    n1597,
    n1655,
    n1641,
    n1635
  );


  nor
  g1645
  (
    n1672,
    n1658,
    n1459,
    n1656,
    n1591
  );


  or
  g1646
  (
    n1661,
    n1460,
    n1640,
    n1644,
    n1653
  );


  nor
  g1647
  (
    n1671,
    n1637,
    n1599,
    n1645,
    n1649
  );


  xor
  g1648
  (
    n1668,
    n1610,
    n1638,
    n1456,
    n1651
  );


  and
  g1649
  (
    n1663,
    n1610,
    n1457,
    n1592,
    n1642
  );


  xor
  g1650
  (
    n1669,
    n1651,
    n1600,
    n1601,
    n1655
  );


  or
  g1651
  (
    n1659,
    n1652,
    n1657,
    n1646,
    n1598
  );


  and
  g1652
  (
    n1674,
    n1669,
    n1634,
    n1670,
    n1633
  );


  xnor
  g1653
  (
    n1673,
    n1404,
    n1671,
    n1672,
    n1633
  );


  xor
  g1654
  (
    n1675,
    n1604,
    n1674,
    n1673,
    n113
  );


  not
  g1655
  (
    n1676,
    n1675
  );


  xnor
  g1656
  (
    n1677,
    n1658,
    n1634
  );


  not
  g1657
  (
    n1678,
    n1676
  );


  nor
  g1658
  (
    n1679,
    n443,
    n1678,
    n442
  );


  nand
  g1659
  (
    n1680,
    n1461,
    n1462
  );


  or
  g1660
  (
    n1682,
    n443,
    n444,
    n1679
  );


  xor
  g1661
  (
    n1683,
    n444,
    n1680,
    n443,
    n1610
  );


  xor
  g1662
  (
    n1681,
    n1677,
    n1680,
    n444,
    n443
  );


  and
  g1663
  (
    n1684,
    n1683,
    n1681,
    n1605,
    n1682
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n291,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n600,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1623,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n135,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1570,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n987,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1303,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1513,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1575,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1543,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n77,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n824,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1550,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1655,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n625,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n52,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1532,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n452,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n567,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n821,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1226,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1328,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n967,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n893,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n548,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n1205,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1272,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n672,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n78,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n657,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1258,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n1583,
    KeyNOTWire_0_31
  );


endmodule

