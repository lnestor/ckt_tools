

module Stat_791_1127
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n810,
  n803,
  n805,
  n797,
  n801,
  n799,
  n795,
  n802,
  n796,
  n806,
  n807,
  n798,
  n809,
  n808,
  n804,
  n794,
  n800,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n810;
  output n803;
  output n805;
  output n797;
  output n801;
  output n799;
  output n795;
  output n802;
  output n796;
  output n806;
  output n807;
  output n798;
  output n809;
  output n808;
  output n804;
  output n794;
  output n800;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n83,
    n4
  );


  not
  g1
  (
    n32,
    n12
  );


  buf
  g2
  (
    n25,
    n3
  );


  buf
  g3
  (
    n29,
    n17
  );


  not
  g4
  (
    n95,
    n19
  );


  buf
  g5
  (
    n93,
    n11
  );


  buf
  g6
  (
    n33,
    n6
  );


  not
  g7
  (
    KeyWire_0_19,
    n16
  );


  buf
  g8
  (
    n62,
    n2
  );


  not
  g9
  (
    n79,
    n9
  );


  not
  g10
  (
    n67,
    n1
  );


  buf
  g11
  (
    n63,
    n9
  );


  not
  g12
  (
    n86,
    n12
  );


  buf
  g13
  (
    n94,
    n2
  );


  not
  g14
  (
    n41,
    n7
  );


  not
  g15
  (
    n91,
    n13
  );


  buf
  g16
  (
    n64,
    n7
  );


  buf
  g17
  (
    n22,
    n8
  );


  buf
  g18
  (
    n56,
    n18
  );


  buf
  g19
  (
    n51,
    n11
  );


  buf
  g20
  (
    n60,
    n4
  );


  not
  g21
  (
    n69,
    n4
  );


  not
  g22
  (
    n45,
    n1
  );


  buf
  g23
  (
    n77,
    n10
  );


  not
  g24
  (
    KeyWire_0_52,
    n18
  );


  buf
  g25
  (
    n52,
    n16
  );


  not
  g26
  (
    KeyWire_0_1,
    n15
  );


  buf
  g27
  (
    n85,
    n1
  );


  buf
  g28
  (
    n40,
    n15
  );


  not
  g29
  (
    n71,
    n4
  );


  buf
  g30
  (
    n68,
    n16
  );


  not
  g31
  (
    KeyWire_0_7,
    n17
  );


  buf
  g32
  (
    n84,
    n2
  );


  buf
  g33
  (
    n80,
    n14
  );


  buf
  g34
  (
    n26,
    n8
  );


  not
  g35
  (
    n72,
    n14
  );


  not
  g36
  (
    KeyWire_0_0,
    n17
  );


  buf
  g37
  (
    n21,
    n18
  );


  not
  g38
  (
    n37,
    n14
  );


  buf
  g39
  (
    n81,
    n12
  );


  not
  g40
  (
    n82,
    n18
  );


  not
  g41
  (
    n28,
    n19
  );


  buf
  g42
  (
    n48,
    n7
  );


  not
  g43
  (
    n42,
    n5
  );


  not
  g44
  (
    n70,
    n3
  );


  not
  g45
  (
    n78,
    n11
  );


  buf
  g46
  (
    n57,
    n17
  );


  not
  g47
  (
    n59,
    n19
  );


  not
  g48
  (
    n76,
    n5
  );


  not
  g49
  (
    n23,
    n13
  );


  not
  g50
  (
    n74,
    n5
  );


  buf
  g51
  (
    n38,
    n7
  );


  not
  g52
  (
    n92,
    n3
  );


  buf
  g53
  (
    n90,
    n13
  );


  not
  g54
  (
    n61,
    n12
  );


  not
  g55
  (
    n27,
    n8
  );


  not
  g56
  (
    n65,
    n9
  );


  not
  g57
  (
    n43,
    n5
  );


  buf
  g58
  (
    n73,
    n14
  );


  not
  g59
  (
    n34,
    n2
  );


  buf
  g60
  (
    n47,
    n6
  );


  buf
  g61
  (
    n50,
    n19
  );


  not
  g62
  (
    n39,
    n11
  );


  buf
  g63
  (
    KeyWire_0_22,
    n13
  );


  buf
  g64
  (
    n88,
    n3
  );


  buf
  g65
  (
    n54,
    n16
  );


  not
  g66
  (
    n35,
    n6
  );


  not
  g67
  (
    n66,
    n15
  );


  not
  g68
  (
    n89,
    n8
  );


  buf
  g69
  (
    n87,
    n10
  );


  buf
  g70
  (
    n44,
    n15
  );


  buf
  g71
  (
    n53,
    n10
  );


  not
  g72
  (
    n49,
    n6
  );


  not
  g73
  (
    n30,
    n9
  );


  not
  g74
  (
    n46,
    n1
  );


  buf
  g75
  (
    n20,
    n10
  );


  not
  g76
  (
    n238,
    n51
  );


  not
  g77
  (
    n159,
    n35
  );


  not
  g78
  (
    n142,
    n39
  );


  buf
  g79
  (
    n361,
    n64
  );


  not
  g80
  (
    n353,
    n75
  );


  buf
  g81
  (
    n310,
    n30
  );


  buf
  g82
  (
    n302,
    n45
  );


  not
  g83
  (
    n119,
    n66
  );


  buf
  g84
  (
    n278,
    n59
  );


  buf
  g85
  (
    n147,
    n41
  );


  not
  g86
  (
    n233,
    n28
  );


  not
  g87
  (
    KeyWire_0_8,
    n32
  );


  not
  g88
  (
    n166,
    n27
  );


  buf
  g89
  (
    n279,
    n81
  );


  buf
  g90
  (
    n306,
    n42
  );


  not
  g91
  (
    n236,
    n41
  );


  buf
  g92
  (
    n124,
    n30
  );


  buf
  g93
  (
    KeyWire_0_6,
    n52
  );


  buf
  g94
  (
    n202,
    n93
  );


  buf
  g95
  (
    n227,
    n25
  );


  not
  g96
  (
    n208,
    n55
  );


  not
  g97
  (
    n311,
    n46
  );


  buf
  g98
  (
    n342,
    n50
  );


  not
  g99
  (
    n234,
    n87
  );


  not
  g100
  (
    n106,
    n78
  );


  not
  g101
  (
    n221,
    n82
  );


  not
  g102
  (
    n171,
    n30
  );


  buf
  g103
  (
    n217,
    n88
  );


  not
  g104
  (
    n99,
    n84
  );


  not
  g105
  (
    n308,
    n29
  );


  buf
  g106
  (
    n101,
    n77
  );


  not
  g107
  (
    n160,
    n47
  );


  buf
  g108
  (
    KeyWire_0_58,
    n43
  );


  not
  g109
  (
    n117,
    n26
  );


  buf
  g110
  (
    n277,
    n69
  );


  not
  g111
  (
    KeyWire_0_13,
    n69
  );


  buf
  g112
  (
    n176,
    n76
  );


  buf
  g113
  (
    n377,
    n27
  );


  buf
  g114
  (
    n275,
    n25
  );


  buf
  g115
  (
    n121,
    n71
  );


  buf
  g116
  (
    n192,
    n76
  );


  not
  g117
  (
    n211,
    n94
  );


  not
  g118
  (
    n112,
    n92
  );


  not
  g119
  (
    n241,
    n61
  );


  buf
  g120
  (
    n287,
    n83
  );


  buf
  g121
  (
    KeyWire_0_5,
    n21
  );


  not
  g122
  (
    n355,
    n70
  );


  not
  g123
  (
    n96,
    n47
  );


  not
  g124
  (
    n304,
    n75
  );


  not
  g125
  (
    n200,
    n82
  );


  not
  g126
  (
    n134,
    n89
  );


  not
  g127
  (
    n137,
    n22
  );


  buf
  g128
  (
    n317,
    n51
  );


  buf
  g129
  (
    n225,
    n70
  );


  not
  g130
  (
    n327,
    n43
  );


  not
  g131
  (
    n296,
    n53
  );


  buf
  g132
  (
    n194,
    n68
  );


  not
  g133
  (
    n395,
    n72
  );


  not
  g134
  (
    n265,
    n95
  );


  buf
  g135
  (
    n324,
    n50
  );


  not
  g136
  (
    KeyWire_0_23,
    n55
  );


  not
  g137
  (
    n183,
    n85
  );


  buf
  g138
  (
    n316,
    n67
  );


  buf
  g139
  (
    n280,
    n71
  );


  not
  g140
  (
    n397,
    n74
  );


  buf
  g141
  (
    KeyWire_0_54,
    n45
  );


  buf
  g142
  (
    n351,
    n88
  );


  buf
  g143
  (
    n152,
    n75
  );


  not
  g144
  (
    n357,
    n21
  );


  not
  g145
  (
    n345,
    n21
  );


  not
  g146
  (
    n141,
    n25
  );


  buf
  g147
  (
    n220,
    n84
  );


  not
  g148
  (
    n281,
    n40
  );


  not
  g149
  (
    n113,
    n29
  );


  not
  g150
  (
    n365,
    n65
  );


  not
  g151
  (
    KeyWire_0_25,
    n65
  );


  buf
  g152
  (
    n340,
    n79
  );


  buf
  g153
  (
    n379,
    n42
  );


  buf
  g154
  (
    n341,
    n64
  );


  buf
  g155
  (
    n254,
    n76
  );


  buf
  g156
  (
    n393,
    n44
  );


  buf
  g157
  (
    n396,
    n80
  );


  buf
  g158
  (
    n100,
    n30
  );


  buf
  g159
  (
    n288,
    n87
  );


  not
  g160
  (
    n179,
    n93
  );


  buf
  g161
  (
    n146,
    n86
  );


  not
  g162
  (
    n102,
    n20
  );


  not
  g163
  (
    n344,
    n93
  );


  buf
  g164
  (
    n381,
    n38
  );


  not
  g165
  (
    n149,
    n32
  );


  not
  g166
  (
    n328,
    n78
  );


  buf
  g167
  (
    n260,
    n79
  );


  not
  g168
  (
    n226,
    n29
  );


  buf
  g169
  (
    n163,
    n37
  );


  buf
  g170
  (
    n116,
    n90
  );


  not
  g171
  (
    n153,
    n56
  );


  not
  g172
  (
    n292,
    n89
  );


  not
  g173
  (
    n283,
    n26
  );


  buf
  g174
  (
    n133,
    n31
  );


  not
  g175
  (
    n253,
    n94
  );


  not
  g176
  (
    n123,
    n63
  );


  not
  g177
  (
    n154,
    n26
  );


  not
  g178
  (
    n122,
    n54
  );


  buf
  g179
  (
    n120,
    n91
  );


  buf
  g180
  (
    n105,
    n81
  );


  buf
  g181
  (
    n191,
    n48
  );


  buf
  g182
  (
    n314,
    n42
  );


  not
  g183
  (
    n323,
    n44
  );


  not
  g184
  (
    KeyWire_0_35,
    n58
  );


  not
  g185
  (
    n293,
    n57
  );


  buf
  g186
  (
    n128,
    n53
  );


  not
  g187
  (
    n243,
    n73
  );


  not
  g188
  (
    n129,
    n37
  );


  buf
  g189
  (
    n130,
    n55
  );


  not
  g190
  (
    n250,
    n43
  );


  buf
  g191
  (
    n228,
    n93
  );


  buf
  g192
  (
    n307,
    n54
  );


  buf
  g193
  (
    n282,
    n91
  );


  buf
  g194
  (
    n334,
    n68
  );


  not
  g195
  (
    n97,
    n50
  );


  buf
  g196
  (
    n242,
    n28
  );


  not
  g197
  (
    n127,
    n85
  );


  not
  g198
  (
    n374,
    n90
  );


  buf
  g199
  (
    n389,
    n49
  );


  buf
  g200
  (
    n337,
    n80
  );


  not
  g201
  (
    n188,
    n94
  );


  buf
  g202
  (
    n162,
    n64
  );


  buf
  g203
  (
    n270,
    n36
  );


  buf
  g204
  (
    n150,
    n86
  );


  buf
  g205
  (
    n204,
    n73
  );


  not
  g206
  (
    n274,
    n24
  );


  not
  g207
  (
    n185,
    n33
  );


  buf
  g208
  (
    n151,
    n21
  );


  buf
  g209
  (
    n165,
    n35
  );


  buf
  g210
  (
    n103,
    n79
  );


  not
  g211
  (
    KeyWire_0_46,
    n20
  );


  not
  g212
  (
    n318,
    n78
  );


  buf
  g213
  (
    n148,
    n37
  );


  not
  g214
  (
    KeyWire_0_44,
    n85
  );


  buf
  g215
  (
    n257,
    n77
  );


  not
  g216
  (
    n376,
    n95
  );


  buf
  g217
  (
    n143,
    n89
  );


  not
  g218
  (
    n138,
    n58
  );


  not
  g219
  (
    n369,
    n47
  );


  not
  g220
  (
    KeyWire_0_28,
    n90
  );


  not
  g221
  (
    n319,
    n51
  );


  buf
  g222
  (
    n230,
    n78
  );


  not
  g223
  (
    n371,
    n37
  );


  buf
  g224
  (
    n300,
    n92
  );


  not
  g225
  (
    n145,
    n56
  );


  not
  g226
  (
    n222,
    n24
  );


  buf
  g227
  (
    n161,
    n83
  );


  not
  g228
  (
    n290,
    n62
  );


  not
  g229
  (
    n356,
    n23
  );


  buf
  g230
  (
    n189,
    n66
  );


  buf
  g231
  (
    n259,
    n22
  );


  not
  g232
  (
    KeyWire_0_27,
    n67
  );


  buf
  g233
  (
    n390,
    n74
  );


  not
  g234
  (
    n244,
    n84
  );


  not
  g235
  (
    n115,
    n61
  );


  not
  g236
  (
    n312,
    n73
  );


  buf
  g237
  (
    n391,
    n46
  );


  not
  g238
  (
    n347,
    n95
  );


  buf
  g239
  (
    n346,
    n75
  );


  buf
  g240
  (
    n173,
    n35
  );


  buf
  g241
  (
    n237,
    n34
  );


  buf
  g242
  (
    n268,
    n92
  );


  not
  g243
  (
    n174,
    n39
  );


  not
  g244
  (
    n180,
    n72
  );


  not
  g245
  (
    n375,
    n87
  );


  not
  g246
  (
    n291,
    n60
  );


  not
  g247
  (
    n240,
    n65
  );


  buf
  g248
  (
    n289,
    n84
  );


  not
  g249
  (
    n322,
    n34
  );


  not
  g250
  (
    n199,
    n53
  );


  not
  g251
  (
    n144,
    n26
  );


  not
  g252
  (
    n219,
    n34
  );


  buf
  g253
  (
    n297,
    n25
  );


  not
  g254
  (
    n198,
    n35
  );


  not
  g255
  (
    n286,
    n34
  );


  buf
  g256
  (
    n256,
    n38
  );


  buf
  g257
  (
    n325,
    n53
  );


  buf
  g258
  (
    n261,
    n45
  );


  buf
  g259
  (
    n246,
    n91
  );


  not
  g260
  (
    n224,
    n57
  );


  buf
  g261
  (
    n104,
    n92
  );


  not
  g262
  (
    n336,
    n71
  );


  not
  g263
  (
    n249,
    n72
  );


  buf
  g264
  (
    n350,
    n33
  );


  not
  g265
  (
    n321,
    n94
  );


  buf
  g266
  (
    n172,
    n49
  );


  buf
  g267
  (
    n186,
    n59
  );


  not
  g268
  (
    n263,
    n73
  );


  buf
  g269
  (
    n181,
    n87
  );


  not
  g270
  (
    n205,
    n58
  );


  buf
  g271
  (
    KeyWire_0_34,
    n52
  );


  buf
  g272
  (
    n339,
    n40
  );


  not
  g273
  (
    n335,
    n68
  );


  buf
  g274
  (
    n284,
    n27
  );


  not
  g275
  (
    n267,
    n74
  );


  buf
  g276
  (
    n332,
    n83
  );


  buf
  g277
  (
    n269,
    n41
  );


  buf
  g278
  (
    KeyWire_0_59,
    n31
  );


  not
  g279
  (
    n329,
    n28
  );


  buf
  g280
  (
    n197,
    n45
  );


  not
  g281
  (
    n372,
    n52
  );


  buf
  g282
  (
    n309,
    n56
  );


  buf
  g283
  (
    n266,
    n23
  );


  not
  g284
  (
    n262,
    n38
  );


  buf
  g285
  (
    n373,
    n70
  );


  not
  g286
  (
    n299,
    n95
  );


  buf
  g287
  (
    n384,
    n22
  );


  buf
  g288
  (
    n175,
    n48
  );


  buf
  g289
  (
    n360,
    n32
  );


  not
  g290
  (
    n212,
    n62
  );


  not
  g291
  (
    n155,
    n48
  );


  not
  g292
  (
    n218,
    n62
  );


  buf
  g293
  (
    n232,
    n67
  );


  not
  g294
  (
    n177,
    n33
  );


  buf
  g295
  (
    n295,
    n69
  );


  not
  g296
  (
    n140,
    n40
  );


  buf
  g297
  (
    n305,
    n47
  );


  buf
  g298
  (
    KeyWire_0_53,
    n62
  );


  not
  g299
  (
    n343,
    n44
  );


  buf
  g300
  (
    n135,
    n82
  );


  buf
  g301
  (
    n348,
    n36
  );


  not
  g302
  (
    n158,
    n90
  );


  buf
  g303
  (
    n215,
    n56
  );


  not
  g304
  (
    n125,
    n55
  );


  not
  g305
  (
    n168,
    n20
  );


  buf
  g306
  (
    n136,
    n50
  );


  not
  g307
  (
    n251,
    n72
  );


  buf
  g308
  (
    n383,
    n64
  );


  not
  g309
  (
    n108,
    n61
  );


  not
  g310
  (
    n207,
    n70
  );


  buf
  g311
  (
    n131,
    n40
  );


  not
  g312
  (
    n213,
    n49
  );


  buf
  g313
  (
    KeyWire_0_14,
    n51
  );


  not
  g314
  (
    n190,
    n61
  );


  buf
  g315
  (
    n354,
    n74
  );


  buf
  g316
  (
    KeyWire_0_12,
    n66
  );


  buf
  g317
  (
    n326,
    n86
  );


  buf
  g318
  (
    n398,
    n23
  );


  buf
  g319
  (
    n206,
    n46
  );


  buf
  g320
  (
    n362,
    n88
  );


  buf
  g321
  (
    n272,
    n58
  );


  not
  g322
  (
    n294,
    n23
  );


  buf
  g323
  (
    n196,
    n76
  );


  buf
  g324
  (
    n182,
    n36
  );


  not
  g325
  (
    n98,
    n83
  );


  not
  g326
  (
    n229,
    n57
  );


  not
  g327
  (
    n255,
    n71
  );


  buf
  g328
  (
    n315,
    n80
  );


  buf
  g329
  (
    n248,
    n43
  );


  not
  g330
  (
    n239,
    n86
  );


  not
  g331
  (
    n118,
    n41
  );


  buf
  g332
  (
    n368,
    n77
  );


  not
  g333
  (
    n338,
    n80
  );


  buf
  g334
  (
    n298,
    n33
  );


  buf
  g335
  (
    n210,
    n59
  );


  buf
  g336
  (
    n252,
    n60
  );


  buf
  g337
  (
    n157,
    n88
  );


  buf
  g338
  (
    n388,
    n31
  );


  not
  g339
  (
    n169,
    n44
  );


  buf
  g340
  (
    n187,
    n77
  );


  buf
  g341
  (
    n386,
    n49
  );


  buf
  g342
  (
    n214,
    n59
  );


  buf
  g343
  (
    n363,
    n22
  );


  buf
  g344
  (
    n264,
    n20
  );


  not
  g345
  (
    n247,
    n31
  );


  buf
  g346
  (
    n330,
    n32
  );


  buf
  g347
  (
    n271,
    n79
  );


  not
  g348
  (
    n195,
    n65
  );


  not
  g349
  (
    n132,
    n68
  );


  buf
  g350
  (
    n366,
    n39
  );


  not
  g351
  (
    n245,
    n48
  );


  buf
  g352
  (
    n273,
    n81
  );


  not
  g353
  (
    KeyWire_0_9,
    n82
  );


  not
  g354
  (
    n216,
    n29
  );


  buf
  g355
  (
    n378,
    n24
  );


  buf
  g356
  (
    n156,
    n63
  );


  not
  g357
  (
    n209,
    n27
  );


  not
  g358
  (
    n167,
    n57
  );


  not
  g359
  (
    n203,
    n63
  );


  not
  g360
  (
    n193,
    n66
  );


  not
  g361
  (
    n184,
    n67
  );


  not
  g362
  (
    n370,
    n42
  );


  not
  g363
  (
    n107,
    n60
  );


  buf
  g364
  (
    KeyWire_0_45,
    n46
  );


  not
  g365
  (
    n359,
    n85
  );


  not
  g366
  (
    n139,
    n60
  );


  not
  g367
  (
    n111,
    n89
  );


  buf
  g368
  (
    n303,
    n54
  );


  not
  g369
  (
    KeyWire_0_47,
    n36
  );


  buf
  g370
  (
    n367,
    n63
  );


  buf
  g371
  (
    n349,
    n24
  );


  not
  g372
  (
    n352,
    n54
  );


  not
  g373
  (
    n235,
    n69
  );


  not
  g374
  (
    n385,
    n52
  );


  buf
  g375
  (
    n333,
    n38
  );


  buf
  g376
  (
    n276,
    n39
  );


  not
  g377
  (
    n164,
    n91
  );


  buf
  g378
  (
    n285,
    n28
  );


  buf
  g379
  (
    n126,
    n81
  );


  not
  g380
  (
    n413,
    n110
  );


  not
  g381
  (
    n402,
    n99
  );


  buf
  g382
  (
    n421,
    n105
  );


  not
  g383
  (
    n412,
    n112
  );


  not
  g384
  (
    n410,
    n119
  );


  not
  g385
  (
    n414,
    n118
  );


  not
  g386
  (
    n401,
    n111
  );


  not
  g387
  (
    n422,
    n97
  );


  buf
  g388
  (
    n423,
    n113
  );


  buf
  g389
  (
    n419,
    n106
  );


  buf
  g390
  (
    n416,
    n114
  );


  buf
  g391
  (
    n405,
    n104
  );


  buf
  g392
  (
    n408,
    n120
  );


  not
  g393
  (
    n403,
    n103
  );


  buf
  g394
  (
    n418,
    n109
  );


  buf
  g395
  (
    n425,
    n121
  );


  not
  g396
  (
    n407,
    n115
  );


  not
  g397
  (
    n404,
    n107
  );


  buf
  g398
  (
    n415,
    n101
  );


  buf
  g399
  (
    n406,
    n108
  );


  not
  g400
  (
    n400,
    n96
  );


  buf
  g401
  (
    n424,
    n116
  );


  buf
  g402
  (
    n420,
    n98
  );


  not
  g403
  (
    n409,
    n117
  );


  buf
  g404
  (
    n411,
    n100
  );


  buf
  g405
  (
    n417,
    n102
  );


  nand
  g406
  (
    n439,
    n404,
    n136,
    n412,
    n400
  );


  or
  g407
  (
    n478,
    n298,
    n402,
    n413,
    n283
  );


  or
  g408
  (
    n472,
    n284,
    n184,
    n421,
    n133
  );


  xnor
  g409
  (
    n429,
    n216,
    n271,
    n182,
    n310
  );


  and
  g410
  (
    n447,
    n400,
    n268,
    n280,
    n402
  );


  or
  g411
  (
    n483,
    n263,
    n173,
    n308,
    n285
  );


  nor
  g412
  (
    KeyWire_0_43,
    n168,
    n277,
    n254,
    n401
  );


  and
  g413
  (
    n498,
    n279,
    n262,
    n410,
    n278
  );


  nor
  g414
  (
    n488,
    n160,
    n304,
    n409,
    n218
  );


  xor
  g415
  (
    n492,
    n420,
    n185,
    n273,
    n187
  );


  and
  g416
  (
    n497,
    n280,
    n276,
    n151,
    n424
  );


  nor
  g417
  (
    KeyWire_0_55,
    n413,
    n417,
    n407,
    n270
  );


  and
  g418
  (
    n450,
    n236,
    n279,
    n241,
    n163
  );


  xnor
  g419
  (
    n487,
    n412,
    n123,
    n164,
    n282
  );


  and
  g420
  (
    n509,
    n417,
    n298,
    n405,
    n191
  );


  nor
  g421
  (
    n519,
    n200,
    n271,
    n423,
    n282
  );


  or
  g422
  (
    n505,
    n289,
    n205,
    n285,
    n291
  );


  xor
  g423
  (
    n463,
    n401,
    n422,
    n282,
    n255
  );


  or
  g424
  (
    n431,
    n304,
    n303,
    n403,
    n188
  );


  nand
  g425
  (
    n434,
    n294,
    n294,
    n175,
    n153
  );


  nor
  g426
  (
    KeyWire_0_41,
    n406,
    n162,
    n194,
    n418
  );


  xor
  g427
  (
    n513,
    n273,
    n222,
    n181,
    n404
  );


  nand
  g428
  (
    n442,
    n285,
    n183,
    n300,
    n281
  );


  nor
  g429
  (
    n476,
    n303,
    n211,
    n210,
    n272
  );


  nand
  g430
  (
    KeyWire_0_16,
    n248,
    n308,
    n295,
    n135
  );


  nor
  g431
  (
    n469,
    n406,
    n253,
    n290,
    n284
  );


  xor
  g432
  (
    n448,
    n301,
    n289,
    n166,
    n228
  );


  and
  g433
  (
    n512,
    n302,
    n128,
    n243,
    n411
  );


  nor
  g434
  (
    n459,
    n408,
    n172,
    n276,
    n233
  );


  xnor
  g435
  (
    n508,
    n169,
    n299,
    n209,
    n401
  );


  and
  g436
  (
    KeyWire_0_38,
    n171,
    n293,
    n154,
    n275
  );


  nand
  g437
  (
    n528,
    n299,
    n280,
    n272,
    n408
  );


  nand
  g438
  (
    n427,
    n401,
    n409,
    n422,
    n299
  );


  nor
  g439
  (
    n467,
    n308,
    n287,
    n425,
    n311
  );


  nor
  g440
  (
    n484,
    n286,
    n275,
    n144,
    n259
  );


  nor
  g441
  (
    n428,
    n293,
    n258,
    n409,
    n279
  );


  or
  g442
  (
    n500,
    n290,
    n275,
    n282,
    n141
  );


  and
  g443
  (
    n433,
    n303,
    n286,
    n414,
    n240
  );


  or
  g444
  (
    n454,
    n158,
    n201,
    n292,
    n249
  );


  xnor
  g445
  (
    n495,
    n420,
    n300,
    n186,
    n285
  );


  nand
  g446
  (
    n494,
    n408,
    n410,
    n306,
    n256
  );


  nor
  g447
  (
    n518,
    n409,
    n221,
    n297,
    n410
  );


  and
  g448
  (
    n435,
    n244,
    n142,
    n230,
    n421
  );


  and
  g449
  (
    KeyWire_0_26,
    n301,
    n261,
    n278,
    n193
  );


  xor
  g450
  (
    KeyWire_0_21,
    n157,
    n203,
    n140,
    n303
  );


  nand
  g451
  (
    n522,
    n264,
    n302,
    n161,
    n130
  );


  nand
  g452
  (
    n457,
    n202,
    n125,
    n235,
    n307
  );


  xor
  g453
  (
    n465,
    n307,
    n299,
    n425,
    n199
  );


  nand
  g454
  (
    n523,
    n405,
    n139,
    n227,
    n421
  );


  nand
  g455
  (
    n515,
    n404,
    n411,
    n155,
    n287
  );


  or
  g456
  (
    n455,
    n407,
    n310,
    n129,
    n296
  );


  nand
  g457
  (
    n480,
    n305,
    n422,
    n419,
    n134
  );


  xnor
  g458
  (
    n426,
    n223,
    n192,
    n416,
    n413
  );


  and
  g459
  (
    n482,
    n265,
    n252,
    n413,
    n246
  );


  nand
  g460
  (
    n443,
    n411,
    n407,
    n293,
    n132
  );


  xor
  g461
  (
    n437,
    n288,
    n311,
    n208,
    n305
  );


  nor
  g462
  (
    n438,
    n250,
    n269,
    n405,
    n415
  );


  nand
  g463
  (
    n502,
    n122,
    n416,
    n420,
    n404
  );


  xor
  g464
  (
    n474,
    n308,
    n311,
    n289,
    n412
  );


  and
  g465
  (
    n514,
    n272,
    n291,
    n302,
    n229
  );


  and
  g466
  (
    n506,
    n287,
    n275,
    n292,
    n137
  );


  or
  g467
  (
    n491,
    n423,
    n204,
    n281,
    n296
  );


  xnor
  g468
  (
    n490,
    n403,
    n274,
    n217,
    n424
  );


  or
  g469
  (
    n511,
    n405,
    n309,
    n415,
    n287
  );


  nand
  g470
  (
    n516,
    n292,
    n283,
    n309,
    n271
  );


  and
  g471
  (
    n496,
    n298,
    n296,
    n274,
    n407
  );


  nand
  g472
  (
    n475,
    n305,
    n257,
    n278,
    n400
  );


  nor
  g473
  (
    n479,
    n239,
    n286,
    n206,
    n138
  );


  nor
  g474
  (
    n481,
    n271,
    n305,
    n302,
    n131
  );


  xnor
  g475
  (
    n458,
    n215,
    n273,
    n306,
    n406
  );


  xor
  g476
  (
    n430,
    n174,
    n415,
    n197,
    n127
  );


  nand
  g477
  (
    n517,
    n304,
    n421,
    n280,
    n425
  );


  xor
  g478
  (
    n449,
    n417,
    n295,
    n291,
    n277
  );


  or
  g479
  (
    n527,
    n156,
    n414,
    n418,
    n301
  );


  and
  g480
  (
    n441,
    n402,
    n234,
    n295,
    n292
  );


  nor
  g481
  (
    n471,
    n167,
    n238,
    n145,
    n307
  );


  xor
  g482
  (
    n525,
    n424,
    n267,
    n281,
    n402
  );


  xor
  g483
  (
    n486,
    n304,
    n403,
    n152,
    n247
  );


  or
  g484
  (
    n460,
    n289,
    n416,
    n410,
    n309
  );


  or
  g485
  (
    n432,
    n231,
    n279,
    n301,
    n298
  );


  xor
  g486
  (
    n493,
    n274,
    n306,
    n273,
    n165
  );


  nand
  g487
  (
    n477,
    n219,
    n294,
    n126,
    n277
  );


  nor
  g488
  (
    n466,
    n170,
    n281,
    n190,
    n408
  );


  xor
  g489
  (
    n524,
    n419,
    n237,
    n288,
    n213
  );


  nand
  g490
  (
    n510,
    n419,
    n416,
    n272,
    n418
  );


  xor
  g491
  (
    n489,
    n293,
    n296,
    n291,
    n286
  );


  and
  g492
  (
    KeyWire_0_39,
    n276,
    n310,
    n242,
    n283
  );


  nor
  g493
  (
    n499,
    n419,
    n309,
    n278,
    n300
  );


  xor
  g494
  (
    KeyWire_0_36,
    n297,
    n143,
    n226,
    n423
  );


  nand
  g495
  (
    KeyWire_0_11,
    n300,
    n406,
    n212,
    n424
  );


  nand
  g496
  (
    n485,
    n415,
    n307,
    n411,
    n251
  );


  xnor
  g497
  (
    n446,
    n284,
    n423,
    n417,
    n288
  );


  xor
  g498
  (
    n473,
    n294,
    n149,
    n177,
    n195
  );


  xor
  g499
  (
    n526,
    n414,
    n260,
    n180,
    n178
  );


  and
  g500
  (
    n452,
    n403,
    n147,
    n310,
    n189
  );


  nand
  g501
  (
    n520,
    n198,
    n420,
    n414,
    n266
  );


  nand
  g502
  (
    KeyWire_0_24,
    n124,
    n245,
    n288,
    n400
  );


  xnor
  g503
  (
    KeyWire_0_2,
    n412,
    n290,
    n297,
    n425
  );


  and
  g504
  (
    n451,
    n306,
    n150,
    n418,
    n232
  );


  xnor
  g505
  (
    KeyWire_0_42,
    n159,
    n295,
    n274,
    n220
  );


  or
  g506
  (
    n503,
    n214,
    n179,
    n283,
    n176
  );


  and
  g507
  (
    n529,
    n224,
    n196,
    n207,
    n148
  );


  and
  g508
  (
    n501,
    n276,
    n422,
    n284,
    n297
  );


  or
  g509
  (
    n507,
    n290,
    n146,
    n277,
    n225
  );


  not
  g510
  (
    n539,
    n440
  );


  not
  g511
  (
    n533,
    n437
  );


  not
  g512
  (
    n549,
    n434
  );


  not
  g513
  (
    n536,
    n430
  );


  not
  g514
  (
    n544,
    n427
  );


  buf
  g515
  (
    n548,
    n444
  );


  not
  g516
  (
    n540,
    n432
  );


  not
  g517
  (
    n547,
    n445
  );


  not
  g518
  (
    n534,
    n429
  );


  not
  g519
  (
    KeyWire_0_17,
    n438
  );


  buf
  g520
  (
    n532,
    n428
  );


  not
  g521
  (
    KeyWire_0_3,
    n446
  );


  buf
  g522
  (
    n550,
    n436
  );


  buf
  g523
  (
    n537,
    n431
  );


  buf
  g524
  (
    KeyWire_0_33,
    n439
  );


  buf
  g525
  (
    n542,
    n441
  );


  not
  g526
  (
    KeyWire_0_20,
    n435
  );


  buf
  g527
  (
    n531,
    n426
  );


  buf
  g528
  (
    n546,
    n433
  );


  not
  g529
  (
    n545,
    n443
  );


  buf
  g530
  (
    n543,
    n442
  );


  not
  g531
  (
    n535,
    n447
  );


  nand
  g532
  (
    n579,
    n375,
    n545,
    n368,
    n345
  );


  xnor
  g533
  (
    KeyWire_0_57,
    n322,
    n342,
    n375,
    n534
  );


  nand
  g534
  (
    n617,
    n313,
    n318,
    n368,
    n531
  );


  and
  g535
  (
    KeyWire_0_49,
    n537,
    n548,
    n350,
    n339
  );


  xor
  g536
  (
    n616,
    n360,
    n358,
    n366,
    n349
  );


  nand
  g537
  (
    n587,
    n541,
    n324,
    n355,
    n330
  );


  or
  g538
  (
    n602,
    n363,
    n338,
    n334,
    n549
  );


  nand
  g539
  (
    n614,
    n367,
    n336,
    n318,
    n348
  );


  nand
  g540
  (
    n583,
    n547,
    n374,
    n337,
    n369
  );


  xnor
  g541
  (
    KeyWire_0_61,
    n352,
    n332,
    n327,
    n334
  );


  and
  g542
  (
    n637,
    n539,
    n362,
    n544,
    n549
  );


  or
  g543
  (
    n606,
    n341,
    n353,
    n330,
    n359
  );


  or
  g544
  (
    n597,
    n327,
    n359,
    n339,
    n364
  );


  or
  g545
  (
    n611,
    n544,
    n544,
    n342,
    n537
  );


  xor
  g546
  (
    n553,
    n343,
    n365,
    n356,
    n545
  );


  xnor
  g547
  (
    n556,
    n328,
    n322,
    n354,
    n351
  );


  and
  g548
  (
    n568,
    n550,
    n368,
    n535,
    n325
  );


  or
  g549
  (
    n608,
    n312,
    n355,
    n337,
    n361
  );


  nor
  g550
  (
    n559,
    n534,
    n344,
    n373,
    n316
  );


  or
  g551
  (
    n585,
    n542,
    n362,
    n336,
    n546
  );


  and
  g552
  (
    n627,
    n539,
    n348,
    n340,
    n352
  );


  nand
  g553
  (
    n601,
    n329,
    n371,
    n538,
    n375
  );


  and
  g554
  (
    n558,
    n372,
    n326,
    n551,
    n366
  );


  xor
  g555
  (
    n565,
    n534,
    n549,
    n363,
    n323
  );


  nand
  g556
  (
    n610,
    n322,
    n317,
    n319,
    n316
  );


  nor
  g557
  (
    n599,
    n548,
    n364,
    n543,
    n329
  );


  or
  g558
  (
    n612,
    n546,
    n370,
    n371,
    n327
  );


  and
  g559
  (
    n563,
    n534,
    n348,
    n325,
    n344
  );


  nor
  g560
  (
    n630,
    n321,
    n321,
    n541,
    n344
  );


  nor
  g561
  (
    n605,
    n539,
    n339,
    n314,
    n333
  );


  xor
  g562
  (
    n596,
    n335,
    n337,
    n369,
    n550
  );


  nor
  g563
  (
    n586,
    n321,
    n315,
    n338,
    n312
  );


  xnor
  g564
  (
    n581,
    n533,
    n329,
    n320,
    n351
  );


  and
  g565
  (
    n623,
    n530,
    n535,
    n312
  );


  xor
  g566
  (
    n625,
    n348,
    n361,
    n363
  );


  nand
  g567
  (
    n632,
    n547,
    n541,
    n343,
    n326
  );


  nor
  g568
  (
    KeyWire_0_18,
    n361,
    n341,
    n342,
    n547
  );


  and
  g569
  (
    n621,
    n542,
    n347,
    n346,
    n355
  );


  xnor
  g570
  (
    n580,
    n349,
    n314,
    n326,
    n319
  );


  xnor
  g571
  (
    n584,
    n320,
    n533,
    n346,
    n312
  );


  xor
  g572
  (
    n569,
    n345,
    n350,
    n341,
    n548
  );


  xor
  g573
  (
    n577,
    n372,
    n550,
    n365,
    n539
  );


  xnor
  g574
  (
    n600,
    n363,
    n365,
    n356,
    n359
  );


  xnor
  g575
  (
    n560,
    n341,
    n338,
    n328,
    n374
  );


  and
  g576
  (
    n572,
    n547,
    n376,
    n373,
    n317
  );


  or
  g577
  (
    n635,
    n358,
    n340,
    n537,
    n342
  );


  nand
  g578
  (
    n620,
    n335,
    n364,
    n365,
    n336
  );


  nand
  g579
  (
    n590,
    n330,
    n543,
    n332,
    n360
  );


  and
  g580
  (
    n615,
    n357,
    n347,
    n549
  );


  nor
  g581
  (
    n589,
    n357,
    n538,
    n325,
    n374
  );


  nand
  g582
  (
    n613,
    n343,
    n354,
    n331,
    n340
  );


  nor
  g583
  (
    KeyWire_0_4,
    n545,
    n332,
    n347,
    n366
  );


  nand
  g584
  (
    n636,
    n338,
    n370,
    n548,
    n536
  );


  nand
  g585
  (
    n626,
    n315,
    n339,
    n335,
    n328
  );


  xnor
  g586
  (
    n566,
    n354,
    n536,
    n311,
    n367
  );


  xnor
  g587
  (
    n562,
    n349,
    n531,
    n533
  );


  and
  g588
  (
    n598,
    n331,
    n540,
    n542,
    n353
  );


  and
  g589
  (
    n618,
    n375,
    n536,
    n360,
    n543
  );


  or
  g590
  (
    n552,
    n318,
    n343,
    n537,
    n535
  );


  nor
  g591
  (
    n588,
    n315,
    n356,
    n536,
    n340
  );


  or
  g592
  (
    KeyWire_0_51,
    n324,
    n333,
    n326,
    n321
  );


  nor
  g593
  (
    n582,
    n369,
    n316,
    n351,
    n333
  );


  xor
  g594
  (
    n593,
    n344,
    n355,
    n333,
    n550
  );


  and
  g595
  (
    KeyWire_0_40,
    n334,
    n315,
    n328,
    n353
  );


  xor
  g596
  (
    KeyWire_0_60,
    n327,
    n317,
    n551
  );


  nor
  g597
  (
    n561,
    n371,
    n357,
    n362,
    n551
  );


  xor
  g598
  (
    n570,
    n357,
    n356,
    n532,
    n543
  );


  xnor
  g599
  (
    n619,
    n372,
    n352,
    n532,
    n335
  );


  nor
  g600
  (
    n595,
    n367,
    n334,
    n370,
    n358
  );


  or
  g601
  (
    n607,
    n352,
    n370,
    n373,
    n350
  );


  xnor
  g602
  (
    n624,
    n362,
    n530,
    n314,
    n313
  );


  and
  g603
  (
    n557,
    n371,
    n313,
    n346,
    n324
  );


  or
  g604
  (
    n576,
    n331,
    n325,
    n531,
    n532
  );


  or
  g605
  (
    n564,
    n345,
    n329,
    n351,
    n322
  );


  nand
  g606
  (
    n603,
    n319,
    n366,
    n368,
    n323
  );


  nand
  g607
  (
    n573,
    n540,
    n372,
    n337,
    n546
  );


  nand
  g608
  (
    n604,
    n364,
    n353,
    n358,
    n545
  );


  xor
  g609
  (
    n567,
    n540,
    n354,
    n320,
    n533
  );


  or
  g610
  (
    n592,
    n332,
    n313,
    n350,
    n532
  );


  nor
  g611
  (
    n571,
    n319,
    n541,
    n367,
    n374
  );


  nor
  g612
  (
    n633,
    n324,
    n538,
    n316,
    n323
  );


  xnor
  g613
  (
    KeyWire_0_63,
    n331,
    n314,
    n359,
    n542
  );


  xor
  g614
  (
    n555,
    n540,
    n544,
    n318,
    n538
  );


  and
  g615
  (
    n554,
    n317,
    n373,
    n320,
    n336
  );


  nor
  g616
  (
    n631,
    n346,
    n323,
    n349,
    n360
  );


  nor
  g617
  (
    n622,
    n330,
    n546,
    n369,
    n345
  );


  xor
  g618
  (
    n661,
    n377,
    n388,
    n379,
    n378
  );


  and
  g619
  (
    n658,
    n386,
    n388,
    n393,
    n383
  );


  xnor
  g620
  (
    KeyWire_0_56,
    n394,
    n386,
    n392
  );


  nor
  g621
  (
    n655,
    n575,
    n568,
    n387,
    n560
  );


  or
  g622
  (
    n652,
    n385,
    n555,
    n381,
    n382
  );


  or
  g623
  (
    n643,
    n566,
    n381,
    n388,
    n552
  );


  xor
  g624
  (
    n662,
    n384,
    n379,
    n564,
    n385
  );


  and
  g625
  (
    KeyWire_0_29,
    n384,
    n387,
    n576,
    n385
  );


  xnor
  g626
  (
    n639,
    n573,
    n380,
    n553,
    n377
  );


  xor
  g627
  (
    n638,
    n569,
    n380,
    n383,
    n385
  );


  xor
  g628
  (
    n641,
    n384,
    n578,
    n392,
    n559
  );


  nor
  g629
  (
    n660,
    n391,
    n574,
    n381,
    n380
  );


  xnor
  g630
  (
    KeyWire_0_15,
    n563,
    n376,
    n383,
    n378
  );


  xnor
  g631
  (
    KeyWire_0_32,
    n567,
    n394,
    n388,
    n392
  );


  xor
  g632
  (
    n656,
    n554,
    n389,
    n390,
    n377
  );


  xnor
  g633
  (
    n645,
    n380,
    n386,
    n394,
    n382
  );


  xnor
  g634
  (
    KeyWire_0_31,
    n561,
    n390,
    n389,
    n577
  );


  xnor
  g635
  (
    n644,
    n558,
    n379,
    n384,
    n390
  );


  or
  g636
  (
    n649,
    n387,
    n392,
    n572,
    n393
  );


  nand
  g637
  (
    n648,
    n383,
    n382,
    n389,
    n394
  );


  nor
  g638
  (
    n642,
    n376,
    n378,
    n390,
    n382
  );


  xor
  g639
  (
    n651,
    n565,
    n389,
    n381,
    n379
  );


  or
  g640
  (
    n653,
    n556,
    n378,
    n393,
    n391
  );


  and
  g641
  (
    n657,
    n571,
    n562,
    n395
  );


  or
  g642
  (
    n647,
    n376,
    n391,
    n557
  );


  nand
  g643
  (
    n654,
    n570,
    n393,
    n377,
    n387
  );


  and
  g644
  (
    n668,
    n639,
    n597,
    n468,
    n588
  );


  xor
  g645
  (
    n675,
    n591,
    n654,
    n587,
    n464
  );


  nor
  g646
  (
    n671,
    n604,
    n644,
    n661,
    n638
  );


  xnor
  g647
  (
    n667,
    n618,
    n602,
    n583,
    n624
  );


  or
  g648
  (
    n687,
    n585,
    n647,
    n615,
    n601
  );


  nor
  g649
  (
    n684,
    n617,
    n593,
    n449,
    n579
  );


  nor
  g650
  (
    n679,
    n450,
    n456,
    n610,
    n599
  );


  and
  g651
  (
    KeyWire_0_10,
    n590,
    n596,
    n613,
    n607
  );


  or
  g652
  (
    n686,
    n660,
    n622,
    n470,
    n651
  );


  nand
  g653
  (
    n665,
    n603,
    n642,
    n467,
    n471
  );


  nor
  g654
  (
    n669,
    n625,
    n581,
    n472,
    n649
  );


  or
  g655
  (
    n666,
    n620,
    n606,
    n452,
    n463
  );


  nand
  g656
  (
    n673,
    n457,
    n612,
    n655,
    n592
  );


  xnor
  g657
  (
    n674,
    n646,
    n458,
    n460,
    n448
  );


  xnor
  g658
  (
    n680,
    n461,
    n451,
    n641,
    n598
  );


  or
  g659
  (
    n664,
    n658,
    n584,
    n459,
    n648
  );


  nor
  g660
  (
    n677,
    n627,
    n623,
    n594,
    n453
  );


  or
  g661
  (
    n670,
    n656,
    n454,
    n650,
    n652
  );


  or
  g662
  (
    n688,
    n659,
    n662,
    n643,
    n466
  );


  and
  g663
  (
    n672,
    n614,
    n605,
    n645,
    n640
  );


  xor
  g664
  (
    n681,
    n657,
    n589,
    n462,
    n619
  );


  nor
  g665
  (
    n676,
    n626,
    n469,
    n455,
    n621
  );


  or
  g666
  (
    n682,
    n608,
    n628,
    n653,
    n465
  );


  or
  g667
  (
    n685,
    n611,
    n616,
    n586,
    n609
  );


  or
  g668
  (
    n678,
    n582,
    n580,
    n595,
    n600
  );


  or
  g669
  (
    n723,
    n527,
    n507,
    n491,
    n396
  );


  and
  g670
  (
    n721,
    n509,
    n479,
    n514
  );


  nand
  g671
  (
    n725,
    n493,
    n517,
    n527,
    n498
  );


  nor
  g672
  (
    n698,
    n514,
    n485,
    n526,
    n666
  );


  xnor
  g673
  (
    n719,
    n396,
    n688,
    n474,
    n397
  );


  xor
  g674
  (
    n720,
    n523,
    n516,
    n477,
    n686
  );


  nor
  g675
  (
    n691,
    n499,
    n500,
    n503,
    n675
  );


  or
  g676
  (
    n730,
    n511,
    n398,
    n517,
    n515
  );


  or
  g677
  (
    n703,
    n667,
    n478,
    n529,
    n528
  );


  nor
  g678
  (
    n704,
    n668,
    n524,
    n492,
    n515
  );


  nand
  g679
  (
    n729,
    n512,
    n670,
    n520,
    n523
  );


  and
  g680
  (
    n708,
    n669,
    n520,
    n686,
    n665
  );


  nand
  g681
  (
    n713,
    n519,
    n522,
    n686,
    n398
  );


  and
  g682
  (
    n692,
    n671,
    n688,
    n686,
    n677
  );


  xnor
  g683
  (
    n715,
    n522,
    n684,
    n529,
    n395
  );


  or
  g684
  (
    n728,
    n396,
    n504,
    n672,
    n496
  );


  xnor
  g685
  (
    n718,
    n683,
    n688,
    n399,
    n528
  );


  xnor
  g686
  (
    n717,
    n682,
    n508,
    n664,
    n521
  );


  or
  g687
  (
    n701,
    n473,
    n524,
    n521,
    n687
  );


  xnor
  g688
  (
    n707,
    n501,
    n688,
    n684,
    n399
  );


  and
  g689
  (
    n709,
    n519,
    n517,
    n528,
    n397
  );


  nand
  g690
  (
    n695,
    n687,
    n685,
    n680,
    n525
  );


  nand
  g691
  (
    n711,
    n683,
    n480,
    n481,
    n522
  );


  nand
  g692
  (
    n689,
    n516,
    n678,
    n475,
    n513
  );


  or
  g693
  (
    n697,
    n521,
    n487,
    n510,
    n524
  );


  and
  g694
  (
    n712,
    n529,
    n513,
    n685,
    n519
  );


  nand
  g695
  (
    n726,
    n513,
    n505,
    n523,
    n522
  );


  nand
  g696
  (
    n710,
    n518,
    n525,
    n516
  );


  and
  g697
  (
    n716,
    n506,
    n673,
    n515,
    n687
  );


  nor
  g698
  (
    n693,
    n685,
    n513,
    n476,
    n515
  );


  nor
  g699
  (
    n702,
    n526,
    n527,
    n483,
    n518
  );


  xnor
  g700
  (
    n727,
    n486,
    n679,
    n489,
    n681
  );


  and
  g701
  (
    n724,
    n488,
    n399,
    n495,
    n490
  );


  xnor
  g702
  (
    n714,
    n502,
    n523,
    n687,
    n395
  );


  xor
  g703
  (
    n700,
    n684,
    n529,
    n521,
    n674
  );


  xnor
  g704
  (
    n690,
    n520,
    n676,
    n517,
    n398
  );


  and
  g705
  (
    n722,
    n397,
    n518,
    n494,
    n685
  );


  nand
  g706
  (
    n706,
    n520,
    n497,
    n396,
    n518
  );


  xor
  g707
  (
    n696,
    n528,
    n524,
    n527,
    n399
  );


  xor
  g708
  (
    n705,
    n482,
    n484,
    n514,
    n519
  );


  and
  g709
  (
    n699,
    n682,
    n525,
    n397,
    n516
  );


  xnor
  g710
  (
    n694,
    n684,
    n398,
    n526
  );


  buf
  g711
  (
    n786,
    n730
  );


  buf
  g712
  (
    n770,
    n722
  );


  not
  g713
  (
    n753,
    n719
  );


  not
  g714
  (
    n748,
    n723
  );


  not
  g715
  (
    n731,
    n726
  );


  not
  g716
  (
    n762,
    n629
  );


  buf
  g717
  (
    n788,
    n712
  );


  not
  g718
  (
    n775,
    n730
  );


  not
  g719
  (
    n732,
    n727
  );


  not
  g720
  (
    n756,
    n699
  );


  not
  g721
  (
    n735,
    n631
  );


  buf
  g722
  (
    n768,
    n705
  );


  not
  g723
  (
    n736,
    n727
  );


  buf
  g724
  (
    n789,
    n633
  );


  buf
  g725
  (
    n777,
    n703
  );


  buf
  g726
  (
    n744,
    n690
  );


  not
  g727
  (
    n769,
    n729
  );


  not
  g728
  (
    KeyWire_0_30,
    n713
  );


  buf
  g729
  (
    n764,
    n726
  );


  buf
  g730
  (
    KeyWire_0_62,
    n730
  );


  not
  g731
  (
    n759,
    n716
  );


  not
  g732
  (
    n785,
    n729
  );


  buf
  g733
  (
    n780,
    n724
  );


  buf
  g734
  (
    n743,
    n702
  );


  buf
  g735
  (
    n761,
    n691
  );


  not
  g736
  (
    n790,
    n727
  );


  not
  g737
  (
    n779,
    n718
  );


  not
  g738
  (
    n749,
    n729
  );


  buf
  g739
  (
    n747,
    n698
  );


  not
  g740
  (
    n752,
    n692
  );


  not
  g741
  (
    KeyWire_0_48,
    n715
  );


  not
  g742
  (
    n763,
    n730
  );


  not
  g743
  (
    n755,
    n720
  );


  not
  g744
  (
    n757,
    n709
  );


  not
  g745
  (
    n734,
    n701
  );


  not
  g746
  (
    n733,
    n717
  );


  not
  g747
  (
    n773,
    n728
  );


  not
  g748
  (
    n737,
    n721
  );


  buf
  g749
  (
    n750,
    n696
  );


  buf
  g750
  (
    n760,
    n689
  );


  buf
  g751
  (
    n738,
    n700
  );


  not
  g752
  (
    n792,
    n724
  );


  buf
  g753
  (
    n739,
    n726
  );


  not
  g754
  (
    n765,
    n724
  );


  not
  g755
  (
    n778,
    n725
  );


  not
  g756
  (
    KeyWire_0_37,
    n697
  );


  not
  g757
  (
    n741,
    n725
  );


  buf
  g758
  (
    n758,
    n708
  );


  buf
  g759
  (
    n754,
    n707
  );


  not
  g760
  (
    n787,
    n714
  );


  not
  g761
  (
    n781,
    n726
  );


  not
  g762
  (
    n784,
    n632
  );


  buf
  g763
  (
    n774,
    n630
  );


  buf
  g764
  (
    n767,
    n706
  );


  buf
  g765
  (
    n776,
    n728
  );


  buf
  g766
  (
    n740,
    n729
  );


  buf
  g767
  (
    n791,
    n724
  );


  not
  g768
  (
    n742,
    n725
  );


  buf
  g769
  (
    n793,
    n711
  );


  not
  g770
  (
    KeyWire_0_50,
    n728
  );


  not
  g771
  (
    n746,
    n693
  );


  and
  g772
  (
    n782,
    n695,
    n710,
    n725
  );


  xor
  g773
  (
    n772,
    n704,
    n727,
    n728,
    n694
  );


  nor
  g774
  (
    n803,
    n747,
    n789,
    n637,
    n749
  );


  nand
  g775
  (
    n800,
    n772,
    n741,
    n742,
    n737
  );


  or
  g776
  (
    n799,
    n771,
    n752,
    n738,
    n774
  );


  nor
  g777
  (
    n810,
    n783,
    n760,
    n635,
    n663
  );


  nand
  g778
  (
    n805,
    n731,
    n782,
    n756,
    n751
  );


  nor
  g779
  (
    n809,
    n745,
    n777,
    n765,
    n732
  );


  xnor
  g780
  (
    n797,
    n634,
    n768,
    n761,
    n735
  );


  xnor
  g781
  (
    n796,
    n781,
    n788,
    n750,
    n769
  );


  or
  g782
  (
    n794,
    n753,
    n778,
    n762,
    n757
  );


  or
  g783
  (
    n795,
    n734,
    n766,
    n733,
    n779
  );


  and
  g784
  (
    n801,
    n764,
    n758,
    n787,
    n785
  );


  nor
  g785
  (
    n798,
    n740,
    n767,
    n791,
    n773
  );


  and
  g786
  (
    n807,
    n763,
    n775,
    n744,
    n770
  );


  xnor
  g787
  (
    n808,
    n790,
    n636,
    n755,
    n754
  );


  nor
  g788
  (
    n802,
    n784,
    n776,
    n746,
    n759
  );


  xor
  g789
  (
    n804,
    n780,
    n736,
    n743,
    n786
  );


  or
  g790
  (
    n806,
    n748,
    n739,
    n793,
    n792
  );


  xnor
  KeyGate_0_0
  (
    n55,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n58,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n521,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n541,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n594,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n258,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n320,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n75,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n301,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n364,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n683,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n445,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n231,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n394,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n387,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n646,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n470,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n530,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n628,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n24,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n551,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n468,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n31,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n110,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n461,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n382,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n436,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n313,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n201,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n663,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n783,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n640,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n659,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n538,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n223,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n114,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n464,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n745,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n504,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n444,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n634,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n456,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n440,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n453,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n399,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n178,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n109,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n358,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n751,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n609,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n766,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n591,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n36,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n331,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n380,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n462,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n650,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n575,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n392,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n170,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n578,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n629,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n771,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n574,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

