// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_156 written by SynthGen on 2021/04/05 11:08:35
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_156 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1023, n1025, n1006, n1013, n1030, n1002, n1016, n1011,
 n1022, n1014, n1027, n1019, n1018, n1004, n1028, n1005,
 n1008, n1026, n1001, n1021, n1029, n1012, n1032, n1031,
 n1003, n1017, n1010, n1007, n1024, n1015, n1009, n1020);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1023, n1025, n1006, n1013, n1030, n1002, n1016, n1011,
 n1022, n1014, n1027, n1019, n1018, n1004, n1028, n1005,
 n1008, n1026, n1001, n1021, n1029, n1012, n1032, n1031,
 n1003, n1017, n1010, n1007, n1024, n1015, n1009, n1020;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000;

not  g0 (n68, n1);
not  g1 (n109, n4);
not  g2 (n95, n8);
not  g3 (n89, n17);
buf  g4 (n111, n13);
not  g5 (n74, n18);
not  g6 (n110, n18);
not  g7 (n49, n13);
not  g8 (n57, n16);
buf  g9 (n54, n7);
not  g10 (n35, n24);
buf  g11 (n102, n5);
not  g12 (n71, n4);
buf  g13 (n59, n20);
not  g14 (n77, n16);
not  g15 (n56, n23);
not  g16 (n86, n26);
not  g17 (n70, n7);
not  g18 (n94, n10);
buf  g19 (n48, n8);
not  g20 (n63, n12);
not  g21 (n60, n6);
buf  g22 (n55, n4);
buf  g23 (n88, n3);
buf  g24 (n38, n13);
not  g25 (n87, n9);
not  g26 (n66, n26);
not  g27 (n42, n11);
buf  g28 (n84, n4);
not  g29 (n79, n8);
not  g30 (n81, n25);
buf  g31 (n46, n9);
buf  g32 (n58, n1);
not  g33 (n34, n24);
buf  g34 (n96, n18);
buf  g35 (n33, n25);
not  g36 (n51, n14);
not  g37 (n104, n3);
buf  g38 (n98, n12);
buf  g39 (n40, n24);
buf  g40 (n52, n16);
not  g41 (n80, n11);
not  g42 (n108, n25);
buf  g43 (n75, n15);
buf  g44 (n103, n6);
buf  g45 (n39, n15);
buf  g46 (n72, n26);
not  g47 (n61, n7);
buf  g48 (n100, n19);
buf  g49 (n36, n16);
buf  g50 (n83, n20);
buf  g51 (n97, n21);
buf  g52 (n90, n17);
buf  g53 (n99, n22);
not  g54 (n45, n13);
buf  g55 (n44, n22);
buf  g56 (n43, n27);
buf  g57 (n64, n12);
buf  g58 (n41, n12);
not  g59 (n93, n6);
buf  g60 (n47, n6);
not  g61 (n53, n23);
not  g62 (n106, n9);
not  g63 (n91, n5);
buf  g64 (n76, n1);
not  g65 (n85, n3);
not  g66 (n73, n2);
buf  g67 (n37, n11);
buf  g68 (n62, n9);
buf  g69 (n78, n3);
not  g70 (n65, n24);
xnor g71 (n107, n1, n23, n11);
and  g72 (n101, n5, n15, n23);
nor  g73 (n105, n21, n27, n19);
or   g74 (n67, n21, n8, n10, n14);
xnor g75 (n82, n25, n20, n14, n17);
xor  g76 (n50, n10, n18, n2, n21);
or   g77 (n92, n19, n26, n14, n22);
xor  g78 (n69, n2, n10, n5, n17);
xor  g79 (n112, n22, n2, n20, n7);
buf  g80 (n238, n48);
not  g81 (n161, n68);
buf  g82 (n145, n37);
buf  g83 (n226, n93);
not  g84 (n119, n107);
not  g85 (n183, n53);
buf  g86 (n160, n56);
buf  g87 (n202, n95);
buf  g88 (n115, n51);
buf  g89 (n212, n38);
not  g90 (n125, n104);
not  g91 (n219, n85);
buf  g92 (n193, n41);
not  g93 (n120, n33);
buf  g94 (n234, n104);
not  g95 (n171, n76);
buf  g96 (n124, n94);
buf  g97 (n213, n87);
not  g98 (n140, n49);
not  g99 (n233, n110);
buf  g100 (n116, n62);
buf  g101 (n200, n54);
not  g102 (n228, n47);
buf  g103 (n205, n75);
buf  g104 (n242, n102);
buf  g105 (n169, n78);
buf  g106 (n209, n96);
buf  g107 (n184, n52);
buf  g108 (n144, n89);
buf  g109 (n166, n109);
buf  g110 (n173, n47);
buf  g111 (n240, n65);
buf  g112 (n231, n73);
not  g113 (n186, n40);
not  g114 (n117, n51);
buf  g115 (n187, n76);
not  g116 (n154, n95);
buf  g117 (n182, n64);
not  g118 (n135, n87);
buf  g119 (n156, n56);
nor  g120 (n235, n35, n106, n100);
xor  g121 (n153, n39, n86, n105);
nor  g122 (n129, n59, n35, n60);
xnor g123 (n151, n72, n85, n74);
nor  g124 (n114, n41, n35, n79);
xnor g125 (n163, n78, n52, n90);
xor  g126 (n195, n60, n44, n103);
nor  g127 (n147, n51, n101, n34);
or   g128 (n152, n47, n105, n101);
nor  g129 (n241, n58, n65, n92);
nand g130 (n201, n98, n108, n45);
xnor g131 (n220, n59, n80, n108);
nand g132 (n211, n54, n61, n83);
and  g133 (n198, n58, n111, n63);
and  g134 (n139, n97, n109, n53);
nor  g135 (n142, n81, n73, n76);
and  g136 (n168, n46, n52, n77);
nor  g137 (n199, n84, n91, n72);
nor  g138 (n237, n94, n83, n79);
nand g139 (n218, n55, n94, n44);
nor  g140 (n123, n55, n99, n41);
nand g141 (n143, n80, n49, n33);
and  g142 (n207, n71, n43, n35);
or   g143 (n131, n60, n107, n98);
nor  g144 (n172, n86, n68, n56);
and  g145 (n224, n42, n98, n78);
nand g146 (n197, n81, n101, n69);
nand g147 (n146, n90, n105, n38);
xnor g148 (n157, n72, n99, n50);
nor  g149 (n179, n57, n43, n91);
nor  g150 (n150, n40, n75, n87);
nor  g151 (n138, n82, n106, n54);
nand g152 (n158, n93, n81, n94);
xor  g153 (n221, n103, n71, n72);
xor  g154 (n181, n38, n89, n85);
nor  g155 (n164, n65, n89, n109);
or   g156 (n127, n62, n46, n42);
or   g157 (n128, n33, n63, n40);
nor  g158 (n149, n97, n39, n106);
nor  g159 (n180, n66, n75, n83);
and  g160 (n177, n62, n49, n45);
nand g161 (n133, n45, n100, n54);
xnor g162 (n239, n61, n36, n58);
xor  g163 (n203, n55, n57, n41);
xnor g164 (n136, n104, n82, n101);
nand g165 (n204, n82, n80);
xor  g166 (n122, n88, n40, n104);
xnor g167 (n196, n36, n34, n52);
xor  g168 (n194, n76, n93);
xor  g169 (n191, n62, n86, n49);
nand g170 (n225, n55, n64, n84);
xnor g171 (n165, n78, n77, n84);
and  g172 (n227, n66, n88, n64);
xnor g173 (n132, n88, n71, n39);
nand g174 (n190, n60, n43, n103);
nor  g175 (n170, n58, n33, n57);
or   g176 (n230, n46, n103, n96);
nand g177 (n236, n57, n96, n48);
xor  g178 (n175, n108, n107, n84);
xor  g179 (n223, n81, n91, n70);
xor  g180 (n141, n97, n110, n108);
and  g181 (n134, n50, n102, n74);
nor  g182 (n188, n53, n90, n64);
nor  g183 (n206, n110, n96, n107);
xor  g184 (n214, n39, n36, n67);
nand g185 (n118, n100, n51, n38);
xnor g186 (n189, n44, n110, n65);
nand g187 (n232, n66, n70, n73);
or   g188 (n229, n53, n46, n61);
xnor g189 (n210, n36, n42, n69);
and  g190 (n137, n92, n45, n88);
nor  g191 (n243, n82, n86, n100);
and  g192 (n222, n98, n77);
xnor g193 (n148, n67, n37, n63);
nand g194 (n217, n90, n70, n47);
or   g195 (n121, n95, n105, n92);
xor  g196 (n215, n102, n42, n106);
xnor g197 (n174, n75, n79, n85);
and  g198 (n126, n59, n67);
xor  g199 (n216, n56, n73, n66);
nand g200 (n167, n43, n63, n102);
xor  g201 (n185, n48, n79, n71);
or   g202 (n113, n99, n61, n74);
nand g203 (n192, n70, n95, n69);
nand g204 (n130, n92, n68, n34);
xor  g205 (n178, n69, n50);
nand g206 (n176, n34, n59, n91);
and  g207 (n162, n87, n37, n48);
nand g208 (n208, n68, n89, n99);
xnor g209 (n155, n83, n74, n97);
nand g210 (n159, n37, n44, n109);
not  g211 (n300, n127);
buf  g212 (n339, n113);
buf  g213 (n315, n127);
not  g214 (n245, n125);
buf  g215 (n348, n115);
buf  g216 (n316, n123);
not  g217 (n354, n128);
not  g218 (n318, n142);
buf  g219 (n351, n123);
buf  g220 (n273, n120);
not  g221 (n319, n120);
not  g222 (n272, n121);
not  g223 (n337, n121);
not  g224 (n249, n141);
not  g225 (n342, n133);
not  g226 (n280, n126);
buf  g227 (n266, n133);
buf  g228 (n358, n115);
not  g229 (n327, n118);
not  g230 (n289, n125);
not  g231 (n331, n117);
not  g232 (n244, n135);
buf  g233 (n290, n135);
buf  g234 (n279, n129);
buf  g235 (n341, n130);
not  g236 (n326, n114);
not  g237 (n284, n138);
not  g238 (n323, n127);
buf  g239 (n340, n127);
not  g240 (n302, n130);
not  g241 (n260, n141);
buf  g242 (n322, n115);
buf  g243 (n275, n132);
not  g244 (n285, n123);
buf  g245 (n254, n126);
not  g246 (n291, n139);
buf  g247 (n248, n128);
not  g248 (n335, n119);
buf  g249 (n287, n134);
not  g250 (n252, n132);
buf  g251 (n309, n131);
not  g252 (n265, n118);
not  g253 (n256, n117);
not  g254 (n262, n128);
not  g255 (n310, n137);
buf  g256 (n277, n130);
not  g257 (n333, n119);
buf  g258 (n283, n137);
buf  g259 (n274, n129);
buf  g260 (n336, n134);
not  g261 (n301, n136);
not  g262 (n347, n121);
buf  g263 (n320, n119);
not  g264 (n250, n131);
not  g265 (n294, n119);
not  g266 (n356, n136);
not  g267 (n346, n122);
buf  g268 (n355, n138);
buf  g269 (n324, n133);
buf  g270 (n271, n124);
not  g271 (n267, n139);
not  g272 (n314, n117);
buf  g273 (n334, n139);
buf  g274 (n286, n123);
not  g275 (n247, n125);
buf  g276 (n345, n114);
not  g277 (n352, n135);
not  g278 (n292, n124);
not  g279 (n312, n120);
not  g280 (n255, n114);
buf  g281 (n305, n122);
buf  g282 (n321, n117);
not  g283 (n353, n140);
not  g284 (n257, n128);
buf  g285 (n343, n129);
buf  g286 (n357, n118);
not  g287 (n264, n140);
not  g288 (n303, n131);
not  g289 (n278, n137);
buf  g290 (n253, n124);
buf  g291 (n270, n130);
not  g292 (n295, n116);
not  g293 (n293, n132);
buf  g294 (n299, n138);
buf  g295 (n344, n138);
buf  g296 (n311, n121);
buf  g297 (n308, n126);
not  g298 (n349, n120);
not  g299 (n251, n134);
not  g300 (n269, n113);
buf  g301 (n329, n140);
not  g302 (n261, n139);
buf  g303 (n328, n142);
buf  g304 (n313, n113);
buf  g305 (n282, n125);
not  g306 (n276, n124);
not  g307 (n258, n141);
buf  g308 (n246, n122);
buf  g309 (n268, n131);
buf  g310 (n317, n115);
buf  g311 (n263, n140);
buf  g312 (n281, n135);
not  g313 (n259, n116);
buf  g314 (n338, n137);
not  g315 (n296, n136);
buf  g316 (n298, n134);
buf  g317 (n332, n126);
buf  g318 (n304, n136);
buf  g319 (n325, n113);
buf  g320 (n350, n114);
buf  g321 (n288, n141);
buf  g322 (n297, n129);
buf  g323 (n330, n118);
buf  g324 (n306, n122);
nand g325 (n307, n116, n116, n133, n132);
buf  g326 (n365, n320);
buf  g327 (n441, n152);
buf  g328 (n436, n156);
not  g329 (n407, n150);
not  g330 (n375, n142);
not  g331 (n404, n255);
buf  g332 (n382, n307);
buf  g333 (n389, n152);
buf  g334 (n438, n144);
not  g335 (n414, n111);
not  g336 (n384, n276);
buf  g337 (n437, n315);
buf  g338 (n403, n295);
buf  g339 (n413, n149);
buf  g340 (n385, n287);
buf  g341 (n387, n259);
buf  g342 (n439, n149);
not  g343 (n425, n155);
buf  g344 (n405, n291);
buf  g345 (n372, n286);
buf  g346 (n399, n268);
not  g347 (n411, n278);
not  g348 (n377, n152);
not  g349 (n381, n153);
not  g350 (n431, n145);
buf  g351 (n435, n252);
buf  g352 (n363, n303);
buf  g353 (n434, n287);
buf  g354 (n364, n112);
not  g355 (n417, n151);
not  g356 (n400, n270);
not  g357 (n402, n313);
not  g358 (n374, n312);
not  g359 (n409, n301);
buf  g360 (n392, n265);
not  g361 (n420, n146);
not  g362 (n408, n260);
buf  g363 (n433, n245);
not  g364 (n360, n294);
buf  g365 (n366, n154);
buf  g366 (n376, n253);
buf  g367 (n398, n300);
not  g368 (n421, n157);
not  g369 (n371, n294);
nor  g370 (n361, n289, n276, n302, n292);
nor  g371 (n370, n248, n144, n151, n282);
and  g372 (n419, n302, n151, n305, n268);
and  g373 (n367, n152, n295, n111, n246);
or   g374 (n390, n149, n275, n254, n306);
xnor g375 (n388, n278, n310, n155);
xnor g376 (n396, n272, n156, n308, n304);
nand g377 (n380, n281, n313, n298, n150);
xor  g378 (n429, n153, n301, n154, n277);
nor  g379 (n394, n311, n112, n269, n148);
nand g380 (n418, n290, n147, n143, n251);
xnor g381 (n415, n285, n284, n257, n308);
nand g382 (n359, n155, n27, n320, n280);
xor  g383 (n424, n305, n304, n286, n150);
xor  g384 (n410, n153, n307, n275, n266);
nand g385 (n426, n296, n154, n146, n148);
nor  g386 (n373, n145, n279, n281, n288);
nor  g387 (n427, n146, n144, n317, n258);
and  g388 (n369, n277, n309, n315, n297);
nor  g389 (n379, n292, n155, n148, n143);
nor  g390 (n395, n145, n306, n314, n267);
nor  g391 (n391, n273, n290, n112, n144);
xor  g392 (n386, n291, n256, n269, n264);
xnor g393 (n378, n319, n293, n303, n148);
xor  g394 (n401, n271, n274, n316, n288);
and  g395 (n406, n143, n311, n314, n284);
and  g396 (n393, n282, n147, n289, n299);
xnor g397 (n397, n147, n111, n280, n142);
or   g398 (n432, n312, n293, n154, n271);
and  g399 (n412, n262, n272, n298, n299);
xor  g400 (n362, n244, n151, n112, n285);
or   g401 (n416, n318, n267, n27, n283);
and  g402 (n422, n274, n143, n283, n146);
nor  g403 (n428, n156, n249, n296, n316);
and  g404 (n368, n270, n317, n263, n319);
or   g405 (n430, n145, n318, n273, n149);
and  g406 (n440, n153, n266, n147, n156);
and  g407 (n383, n279, n309, n247, n250);
xnor g408 (n423, n300, n150, n297, n261);
xnor g409 (n445, n362, n364, n363);
xnor g410 (n448, n364, n360);
and  g411 (n447, n361, n360, n363);
or   g412 (n444, n360, n361, n366, n362);
xnor g413 (n442, n362, n361, n366, n364);
xnor g414 (n443, n362, n366, n365);
nor  g415 (n446, n364, n365);
xnor g416 (n449, n359, n363, n361, n367);
nor  g417 (n452, n157, n28, n158);
xnor g418 (n451, n443, n445, n157, n29);
nand g419 (n450, n28, n158, n157);
xor  g420 (n453, n158, n28, n444, n442);
nor  g421 (n463, n450, n369, n453, n373);
or   g422 (n461, n371, n372, n367);
nor  g423 (n456, n370, n373, n368);
nand g424 (n460, n374, n371, n452, n369);
nand g425 (n458, n370, n369, n452);
nor  g426 (n454, n453, n453, n374, n371);
or   g427 (n455, n368, n372, n451, n369);
xnor g428 (n457, n368, n453, n372, n367);
or   g429 (n462, n370, n372, n373, n374);
nand g430 (n459, n452, n370, n373, n371);
or   g431 (n497, n160, n463, n383, n461);
xnor g432 (n498, n167, n159, n171, n166);
xor  g433 (n489, n160, n164, n460, n457);
xor  g434 (n483, n381, n170, n456, n175);
xnor g435 (n468, n384, n177, n168, n383);
and  g436 (n492, n459, n163, n171, n461);
xnor g437 (n501, n159, n457, n379, n177);
nand g438 (n465, n164, n383, n173, n163);
nand g439 (n485, n164, n456, n378, n376);
xnor g440 (n477, n178, n457, n162);
nand g441 (n491, n379, n173, n459, n381);
nand g442 (n499, n455, n174, n159, n171);
or   g443 (n480, n461, n455, n462, n169);
and  g444 (n500, n455, n177, n174);
nand g445 (n478, n161, n461, n380, n383);
nor  g446 (n479, n378, n379, n377, n165);
xor  g447 (n503, n460, n160, n169, n378);
xor  g448 (n482, n172, n169, n375, n161);
xor  g449 (n487, n172, n169, n380, n170);
nand g450 (n502, n454, n382, n168, n375);
and  g451 (n488, n175, n454, n163, n166);
nor  g452 (n495, n160, n377, n176, n167);
nor  g453 (n496, n176, n458, n384, n382);
and  g454 (n466, n455, n172, n457, n463);
nor  g455 (n486, n379, n175, n459, n162);
or   g456 (n494, n463, n376, n176, n166);
nor  g457 (n472, n460, n165, n458, n175);
nand g458 (n470, n458, n170, n163, n167);
nor  g459 (n471, n172, n381, n173, n376);
xnor g460 (n481, n456, n384, n377, n176);
and  g461 (n490, n382, n380, n454, n462);
xor  g462 (n469, n374, n178, n168, n161);
xnor g463 (n484, n463, n159, n460, n173);
or   g464 (n467, n165, n462, n381, n161);
xnor g465 (n475, n384, n166, n459, n375);
or   g466 (n473, n454, n382, n168, n380);
xnor g467 (n476, n376, n378, n462, n174);
xnor g468 (n474, n377, n170, n456, n177);
nand g469 (n464, n162, n375, n171, n164);
or   g470 (n493, n167, n458, n165, n178);
and  g471 (n554, n343, n345, n391, n470);
xnor g472 (n551, n399, n397, n343, n478);
nand g473 (n530, n332, n350, n487, n347);
nor  g474 (n574, n467, n396, n464, n332);
xor  g475 (n508, n346, n358, n405, n487);
xnor g476 (n525, n349, n350, n386, n329);
nand g477 (n571, n483, n390, n485, n400);
xnor g478 (n548, n339, n327, n335, n386);
nor  g479 (n519, n397, n486, n475, n471);
xnor g480 (n512, n474, n393, n466, n355);
xnor g481 (n547, n487, n331, n330);
nor  g482 (n568, n354, n336, n346, n491);
xnor g483 (n572, n343, n345, n327, n349);
or   g484 (n529, n480, n355, n392, n485);
xor  g485 (n523, n355, n336, n348, n393);
or   g486 (n544, n321, n326, n332, n395);
xor  g487 (n567, n489, n404, n399, n391);
xor  g488 (n520, n385, n398, n395, n490);
xnor g489 (n504, n325, n388, n394, n341);
nand g490 (n536, n484, n488, n340, n321);
xor  g491 (n560, n484, n337, n396, n467);
or   g492 (n531, n400, n334, n335, n491);
xor  g493 (n527, n404, n348, n351, n388);
xor  g494 (n553, n482, n339, n328, n485);
xnor g495 (n555, n474, n336, n397, n485);
xnor g496 (n521, n401, n396, n358, n354);
xnor g497 (n549, n352, n387, n326, n338);
nand g498 (n558, n490, n489, n400, n335);
xor  g499 (n522, n357, n352, n472, n405);
or   g500 (n576, n464, n338, n337, n331);
and  g501 (n524, n338, n332, n385, n478);
nor  g502 (n575, n394, n352, n339, n403);
or   g503 (n557, n334, n385, n386, n477);
or   g504 (n569, n395, n353, n484, n487);
nand g505 (n528, n401, n390, n354, n490);
or   g506 (n518, n393, n483, n336, n356);
or   g507 (n507, n347, n340, n398, n472);
nand g508 (n566, n347, n339, n351, n398);
nor  g509 (n517, n356, n350, n387, n395);
xnor g510 (n573, n388, n324, n325, n391);
xor  g511 (n526, n335, n387, n340, n483);
nand g512 (n511, n466, n329, n405, n354);
nand g513 (n564, n473, n386, n398, n404);
xor  g514 (n546, n469, n331, n403, n481);
xor  g515 (n514, n337, n396, n394, n352);
nor  g516 (n539, n341, n390, n323, n322);
xor  g517 (n545, n402, n480, n330, n353);
xor  g518 (n550, n490, n402, n477, n355);
or   g519 (n542, n349, n330, n333, n358);
and  g520 (n537, n406, n337, n402, n342);
xor  g521 (n505, n473, n479, n322, n393);
nor  g522 (n562, n471, n402, n397, n481);
and  g523 (n535, n476, n333, n389, n486);
nor  g524 (n552, n331, n345, n399, n357);
nand g525 (n540, n479, n358, n392, n356);
xor  g526 (n509, n491, n344, n399, n400);
xor  g527 (n515, n324, n343, n338, n357);
and  g528 (n563, n465, n385, n486, n341);
nor  g529 (n559, n488, n475, n389, n333);
or   g530 (n543, n347, n353, n392, n334);
nand g531 (n534, n488, n345, n391, n390);
and  g532 (n570, n488, n340, n482, n468);
xor  g533 (n533, n489, n470, n476, n348);
nand g534 (n565, n394, n344, n349, n401);
xnor g535 (n516, n333, n484, n323, n357);
nand g536 (n532, n465, n403, n344, n405);
xor  g537 (n506, n334, n483, n401, n351);
or   g538 (n541, n342, n328, n387, n348);
nand g539 (n538, n342, n342, n350, n344);
nor  g540 (n561, n351, n468, n469, n403);
nor  g541 (n513, n486, n341, n392, n346);
or   g542 (n556, n404, n353, n389);
xnor g543 (n510, n388, n346, n489, n356);
xor  g544 (n584, n407, n510);
nor  g545 (n580, n406, n508);
nand g546 (n579, n504, n506);
xor  g547 (n582, n507, n505);
and  g548 (n578, n511, n408);
or   g549 (n583, n509, n406);
not  g550 (n581, n407);
xnor g551 (n577, n407, n406);
xnor g552 (n608, n411, n522, n448, n180);
xnor g553 (n603, n183, n583, n521, n578);
xnor g554 (n606, n409, n409, n551, n579);
and  g555 (n595, n525, n584, n526, n181);
or   g556 (n602, n183, n577, n181, n411);
and  g557 (n613, n578, n512, n534, n543);
nor  g558 (n607, n582, n180, n181, n579);
or   g559 (n612, n181, n179, n581);
nand g560 (n611, n449, n179, n580, n531);
nand g561 (n610, n532, n178, n411, n582);
xnor g562 (n609, n514, n446, n538, n410);
xnor g563 (n596, n180, n516, n581, n527);
nor  g564 (n592, n580, n523, n518, n515);
or   g565 (n588, n179, n408, n579, n183);
nor  g566 (n591, n546, n182, n410, n582);
xnor g567 (n587, n579, n547, n541, n580);
nand g568 (n604, n409, n550, n583, n517);
or   g569 (n593, n540, n533, n548, n182);
nand g570 (n599, n539, n583, n182, n584);
xnor g571 (n601, n410, n448, n449);
nand g572 (n594, n513, n583, n447, n520);
nand g573 (n600, n578, n524, n580, n544);
and  g574 (n589, n449, n581, n549);
or   g575 (n605, n447, n182, n578, n446);
nand g576 (n598, n582, n584, n408, n535);
and  g577 (n586, n584, n448, n491, n537);
xnor g578 (n597, n545, n409, n529, n542);
or   g579 (n585, n449, n536, n519, n180);
or   g580 (n590, n408, n528, n530, n410);
not  g581 (n658, n429);
buf  g582 (n665, n608);
not  g583 (n638, n610);
not  g584 (n620, n593);
not  g585 (n625, n596);
buf  g586 (n656, n592);
buf  g587 (n621, n594);
buf  g588 (n701, n590);
buf  g589 (n615, n594);
buf  g590 (n671, n599);
buf  g591 (n618, n591);
buf  g592 (n691, n418);
not  g593 (n666, n593);
not  g594 (n630, n603);
buf  g595 (n708, n613);
buf  g596 (n676, n417);
buf  g597 (n644, n589);
buf  g598 (n640, n595);
not  g599 (n672, n603);
buf  g600 (n633, n418);
not  g601 (n704, n606);
buf  g602 (n702, n608);
not  g603 (n614, n606);
not  g604 (n646, n590);
buf  g605 (n634, n604);
buf  g606 (n693, n600);
not  g607 (n684, n421);
not  g608 (n668, n598);
buf  g609 (n639, n564);
buf  g610 (n631, n432);
buf  g611 (n685, n436);
not  g612 (n653, n596);
not  g613 (n632, n613);
buf  g614 (n663, n593);
not  g615 (n675, n422);
buf  g616 (n679, n596);
not  g617 (n689, n607);
not  g618 (n623, n595);
not  g619 (n682, n604);
buf  g620 (n619, n594);
not  g621 (n698, n586);
not  g622 (n700, n554);
buf  g623 (n617, n592);
buf  g624 (n686, n415);
not  g625 (n648, n589);
buf  g626 (n664, n417);
buf  g627 (n667, n597);
not  g628 (n699, n607);
not  g629 (n641, n612);
xnor g630 (n705, n421, n493, n604);
nand g631 (n624, n420, n413, n434, n585);
nand g632 (n627, n420, n563, n492, n428);
nor  g633 (n637, n607, n426, n430, n417);
nor  g634 (n695, n587, n425, n424, n599);
xor  g635 (n661, n592, n426, n585, n588);
and  g636 (n696, n588, n428, n604, n559);
xor  g637 (n669, n412, n589, n429, n601);
xor  g638 (n642, n414, n435, n597, n436);
nand g639 (n655, n608, n595, n601, n416);
and  g640 (n673, n422, n594, n418, n600);
xnor g641 (n659, n424, n419, n602, n586);
and  g642 (n654, n601, n419, n608, n416);
nand g643 (n680, n609, n605, n420);
xnor g644 (n662, n427, n603, n426, n434);
xor  g645 (n690, n431, n599, n412, n585);
or   g646 (n687, n586, n427, n428, n588);
nor  g647 (n692, n597, n427, n416, n561);
nor  g648 (n651, n610, n613, n612, n598);
and  g649 (n706, n553, n432, n611, n590);
nand g650 (n626, n431, n415, n423);
xor  g651 (n678, n434, n492, n600, n423);
and  g652 (n703, n432, n421, n605, n593);
xor  g653 (n652, n430, n599, n421, n436);
nor  g654 (n694, n585, n592, n417, n425);
and  g655 (n709, n595, n414, n412, n424);
or   g656 (n677, n436, n590, n610, n557);
or   g657 (n636, n610, n435, n430, n429);
and  g658 (n616, n611, n596, n492, n430);
nor  g659 (n649, n415, n419, n432);
nor  g660 (n657, n612, n435, n414, n420);
or   g661 (n628, n556, n598, n413, n424);
or   g662 (n629, n586, n434, n611, n603);
xnor g663 (n660, n492, n598, n602, n425);
nor  g664 (n683, n429, n413, n613, n411);
and  g665 (n647, n428, n607, n609, n422);
nand g666 (n697, n431, n558, n433, n435);
or   g667 (n707, n560, n588, n605, n426);
nor  g668 (n674, n433, n587, n611, n600);
and  g669 (n645, n437, n602, n606, n601);
and  g670 (n670, n425, n589, n418, n609);
nor  g671 (n688, n552, n609, n591, n423);
nand g672 (n643, n597, n612, n427, n433);
nor  g673 (n681, n422, n555, n416, n602);
xnor g674 (n650, n414, n591, n413, n412);
and  g675 (n635, n606, n591, n587, n415);
xnor g676 (n622, n562, n587, n431, n433);
xor  g677 (n769, n184, n225, n706, n238);
nand g678 (n778, n198, n570, n188, n201);
nand g679 (n741, n617, n625, n643, n187);
nand g680 (n714, n189, n665, n623, n199);
xnor g681 (n755, n664, n672, n197, n627);
nor  g682 (n798, n681, n651, n668, n623);
or   g683 (n760, n686, n202, n661, n230);
or   g684 (n870, n238, n232, n672, n660);
and  g685 (n869, n241, n202, n679, n628);
or   g686 (n810, n688, n183, n208, n684);
and  g687 (n752, n690, n669, n682, n200);
nor  g688 (n751, n662, n663, n231, n614);
and  g689 (n802, n239, n186, n222, n194);
xor  g690 (n759, n217, n666, n243, n657);
and  g691 (n816, n619, n661, n683, n185);
nor  g692 (n844, n650, n683, n208, n673);
xnor g693 (n849, n677, n630, n642, n676);
or   g694 (n744, n224, n698, n628, n208);
xnor g695 (n713, n695, n635, n234, n216);
xor  g696 (n806, n196, n29, n630, n658);
nor  g697 (n753, n692, n617, n651, n622);
or   g698 (n850, n619, n203, n236, n211);
nand g699 (n848, n692, n237, n645, n243);
nand g700 (n818, n615, n235, n32, n625);
or   g701 (n854, n224, n646, n621, n620);
xnor g702 (n780, n653, n665, n631, n614);
xor  g703 (n735, n186, n209, n31, n236);
xnor g704 (n772, n701, n188, n689, n695);
xnor g705 (n811, n32, n232, n229, n646);
nand g706 (n716, n238, n654, n636, n632);
or   g707 (n732, n619, n666, n199, n639);
xor  g708 (n862, n659, n239, n706, n648);
nand g709 (n825, n659, n624, n184, n206);
xnor g710 (n787, n615, n652, n677, n223);
xnor g711 (n842, n694, n631, n30, n681);
nor  g712 (n796, n685, n187, n200, n680);
nand g713 (n710, n690, n650, n32, n693);
or   g714 (n853, n678, n702, n687, n654);
nand g715 (n805, n229, n228, n668, n618);
xor  g716 (n717, n184, n697, n632, n676);
nand g717 (n828, n214, n687, n194, n235);
and  g718 (n726, n653, n692, n626, n651);
or   g719 (n777, n213, n657, n696, n214);
and  g720 (n747, n226, n681, n682, n204);
nand g721 (n843, n635, n650, n693, n653);
and  g722 (n739, n189, n660, n215);
xnor g723 (n773, n218, n198, n695, n615);
and  g724 (n761, n703, n630, n203, n657);
xnor g725 (n856, n674, n677, n649, n234);
and  g726 (n768, n220, n678, n701, n615);
and  g727 (n738, n700, n185, n216, n637);
nor  g728 (n799, n237, n664, n201, n658);
nor  g729 (n861, n29, n231, n640, n652);
or   g730 (n840, n207, n184, n705, n627);
nor  g731 (n823, n239, n637, n221, n231);
or   g732 (n779, n617, n229, n678, n675);
xnor g733 (n871, n31, n618, n709, n191);
xnor g734 (n785, n699, n192, n220, n189);
or   g735 (n792, n201, n207, n645, n668);
xor  g736 (n794, n656, n679, n708, n698);
nor  g737 (n724, n669, n199, n639, n242);
or   g738 (n764, n225, n210, n204, n205);
xnor g739 (n733, n567, n193, n212, n655);
and  g740 (n743, n684, n190, n680, n212);
nor  g741 (n809, n650, n654, n236, n234);
nand g742 (n784, n242, n230, n31, n685);
or   g743 (n866, n235, n640, n656, n694);
xor  g744 (n837, n571, n689, n697, n645);
nor  g745 (n841, n206, n672, n212, n691);
or   g746 (n770, n675, n621, n620, n667);
or   g747 (n774, n572, n209, n236, n219);
xor  g748 (n807, n223, n233, n195, n621);
nand g749 (n725, n680, n696, n668, n624);
nand g750 (n762, n679, n639, n673, n235);
xnor g751 (n728, n691, n622, n687, n631);
or   g752 (n852, n654, n699, n671, n709);
nor  g753 (n833, n243, n689, n634, n209);
nand g754 (n808, n658, n662, n664, n240);
xor  g755 (n771, n200, n633, n241, n217);
xor  g756 (n832, n237, n706, n691, n651);
nor  g757 (n788, n194, n225, n709, n704);
or   g758 (n789, n704, n222, n210, n241);
nor  g759 (n863, n228, n189, n227, n637);
xor  g760 (n839, n217, n30, n240, n196);
xor  g761 (n814, n242, n221, n645, n614);
and  g762 (n845, n197, n697, n662, n660);
or   g763 (n864, n617, n618, n671, n679);
and  g764 (n781, n192, n633, n675, n569);
xor  g765 (n765, n202, n205, n627, n223);
and  g766 (n775, n216, n622, n638, n620);
nand g767 (n859, n694, n211, n648, n616);
nand g768 (n829, n206, n683, n700, n669);
nand g769 (n855, n641, n191, n672);
and  g770 (n860, n663, n685, n652, n618);
nor  g771 (n748, n698, n195, n691, n207);
and  g772 (n718, n629, n655, n215, n692);
or   g773 (n783, n662, n671, n218, n211);
xnor g774 (n750, n210, n212, n648, n702);
nand g775 (n820, n628, n242, n185, n674);
xnor g776 (n793, n690, n186, n667, n657);
nand g777 (n812, n576, n203, n688, n638);
xor  g778 (n831, n193, n211, n705, n641);
nand g779 (n786, n209, n226, n217, n31);
xnor g780 (n819, n222, n203, n221, n202);
and  g781 (n737, n233, n670, n683, n197);
nor  g782 (n740, n630, n204, n636, n656);
nor  g783 (n867, n634, n663, n701, n647);
or   g784 (n817, n685, n702, n616, n629);
nand g785 (n711, n195, n625, n640, n226);
and  g786 (n746, n695, n661, n636, n233);
xor  g787 (n797, n207, n208, n190);
nor  g788 (n834, n677, n638, n637, n204);
xnor g789 (n804, n642, n218, n641, n188);
or   g790 (n846, n214, n199, n633, n213);
nor  g791 (n721, n619, n644, n675, n655);
nor  g792 (n835, n648, n231, n193, n232);
nand g793 (n865, n703, n693, n700, n225);
xor  g794 (n715, n661, n214, n680, n684);
nand g795 (n857, n708, n671, n240, n647);
nand g796 (n749, n638, n227, n215, n224);
or   g797 (n754, n626, n566, n565, n240);
xor  g798 (n868, n674, n646, n206, n219);
and  g799 (n830, n660, n643, n190, n658);
nor  g800 (n791, n201, n699, n674, n633);
xor  g801 (n722, n186, n187, n655);
nor  g802 (n790, n29, n640, n621, n670);
or   g803 (n763, n676, n690, n688, n639);
nor  g804 (n742, n652, n686, n193, n626);
xor  g805 (n782, n620, n205, n644, n32);
and  g806 (n824, n684, n643, n234, n649);
xor  g807 (n858, n665, n229, n624, n641);
xnor g808 (n821, n699, n625, n669, n632);
and  g809 (n734, n227, n205, n707, n197);
xnor g810 (n723, n697, n708, n649, n30);
or   g811 (n801, n702, n696, n230, n653);
nor  g812 (n827, n705, n200, n701, n673);
and  g813 (n730, n647, n659, n670, n693);
xnor g814 (n712, n227, n196, n213, n707);
or   g815 (n795, n614, n195, n629, n704);
xor  g816 (n776, n664, n241, n646, n673);
nor  g817 (n847, n222, n676, n624, n686);
xnor g818 (n822, n192, n682, n191, n196);
xor  g819 (n758, n623, n221, n243, n696);
or   g820 (n836, n228, n198, n659, n213);
xnor g821 (n736, n670, n681, n708, n642);
or   g822 (n803, n705, n686, n706, n574);
xor  g823 (n800, n698, n220, n30, n623);
or   g824 (n851, n223, n704, n228, n649);
xor  g825 (n767, n634, n636, n707, n666);
nand g826 (n766, n682, n628, n631, n629);
and  g827 (n756, n687, n573, n233, n689);
nand g828 (n719, n627, n194, n703, n666);
nand g829 (n727, n694, n220, n622, n568);
xnor g830 (n720, n575, n700, n626, n678);
xnor g831 (n838, n616, n219, n218, n188);
nand g832 (n731, n667, n198, n185, n665);
xnor g833 (n745, n239, n709, n667, n226);
xnor g834 (n872, n688, n656, n644, n237);
xor  g835 (n826, n230, n224, n232, n703);
and  g836 (n813, n644, n219, n238, n616);
and  g837 (n757, n643, n192, n647, n635);
or   g838 (n729, n216, n635, n634, n632);
nand g839 (n815, n663, n642, n707, n210);
nand g840 (n873, n840, n813, n499, n860);
xnor g841 (n874, n754, n846, n815, n729);
xor  g842 (n907, n744, n755, n772, n831);
xor  g843 (n994, n503, n813, n869, n860);
xor  g844 (n990, n500, n867, n857, n777);
nor  g845 (n977, n712, n720, n779, n732);
or   g846 (n922, n765, n501, n819, n759);
or   g847 (n902, n791, n839, n726, n725);
nand g848 (n976, n749, n719, n751, n780);
and  g849 (n894, n748, n845, n820, n730);
xnor g850 (n941, n735, n764, n852, n503);
xnor g851 (n964, n843, n771, n441, n830);
nand g852 (n933, n827, n715, n870, n844);
nor  g853 (n958, n502, n822, n838, n438);
nor  g854 (n961, n821, n824, n865, n807);
or   g855 (n997, n857, n716, n765, n757);
nand g856 (n978, n762, n864, n816, n739);
and  g857 (n885, n734, n745, n728, n768);
xor  g858 (n955, n871, n828, n439, n494);
xor  g859 (n896, n499, n819, n835, n501);
nor  g860 (n965, n837, n806, n860, n856);
or   g861 (n995, n764, n761, n782, n824);
xor  g862 (n884, n800, n857, n774, n799);
or   g863 (n917, n835, n809, n743, n758);
xor  g864 (n932, n830, n864, n797, n847);
nor  g865 (n929, n718, n859, n823, n867);
and  g866 (n935, n752, n866, n857, n724);
xnor g867 (n892, n803, n786, n750, n837);
and  g868 (n943, n439, n803, n870, n817);
nand g869 (n887, n737, n871, n805, n786);
xnor g870 (n938, n727, n866, n710, n844);
xor  g871 (n942, n785, n806, n822, n790);
and  g872 (n973, n872, n823, n438, n862);
xnor g873 (n970, n828, n869, n836, n816);
xnor g874 (n881, n812, n805, n712, n822);
xor  g875 (n975, n866, n868, n842, n858);
xor  g876 (n918, n710, n812, n498, n865);
nand g877 (n927, n851, n494, n835, n804);
xnor g878 (n882, n437, n821, n841, n767);
or   g879 (n948, n830, n787, n441, n789);
nor  g880 (n987, n838, n440, n758, n794);
nand g881 (n969, n772, n747, n727, n501);
nand g882 (n924, n716, n856, n865, n736);
and  g883 (n891, n811, n755, n812, n852);
nor  g884 (n951, n776, n843, n761, n852);
and  g885 (n899, n719, n859, n814, n834);
xor  g886 (n993, n840, n869, n827, n731);
nand g887 (n926, n815, n833, n808, n438);
xor  g888 (n998, n815, n863, n853, n725);
xor  g889 (n963, n437, n802, n729, n438);
and  g890 (n999, n818, n849, n836, n824);
nand g891 (n931, n773, n868, n778, n825);
xnor g892 (n984, n770, n739, n763, n734);
xor  g893 (n880, n868, n793, n816, n503);
or   g894 (n986, n497, n495, n503, n861);
xnor g895 (n879, n846, n809, n850, n751);
nor  g896 (n979, n826, n733, n834, n441);
xnor g897 (n903, n826, n831, n847, n759);
and  g898 (n966, n849, n831, n722, n795);
or   g899 (n962, n753, n863, n495, n829);
xnor g900 (n991, n810, n818, n717, n842);
nand g901 (n901, n860, n837, n717, n825);
nor  g902 (n906, n754, n730, n791, n781);
nand g903 (n960, n796, n437, n836, n841);
xnor g904 (n928, n867, n496, n820, n846);
nand g905 (n980, n817, n845, n784, n833);
nand g906 (n919, n798, n496, n840, n807);
nor  g907 (n972, n748, n861, n817, n823);
xor  g908 (n936, n778, n871, n851, n753);
xnor g909 (n920, n866, n854, n711, n439);
or   g910 (n953, n721, n827, n845, n499);
nor  g911 (n944, n811, n855, n835, n856);
xnor g912 (n921, n850, n752, n496, n771);
nand g913 (n949, n819, n830, n840, n861);
xor  g914 (n908, n826, n818, n870, n781);
and  g915 (n952, n841, n834, n728, n863);
nand g916 (n1000, n726, n847, n797, n826);
and  g917 (n945, n747, n494, n824, n838);
or   g918 (n915, n849, n777, n762, n838);
nor  g919 (n897, n812, n832, n766, n825);
nand g920 (n946, n837, n774, n839, n871);
nand g921 (n937, n740, n862, n813, n497);
xor  g922 (n959, n832, n502, n831, n796);
xor  g923 (n895, n861, n802, n746, n864);
xnor g924 (n940, n440, n801, n843, n821);
or   g925 (n878, n800, n783, n855, n769);
or   g926 (n883, n849, n844, n848, n845);
nor  g927 (n890, n848, n767, n850, n822);
xnor g928 (n898, n779, n872, n495, n783);
nor  g929 (n983, n500, n869, n713, n497);
xnor g930 (n981, n742, n868, n821, n862);
xor  g931 (n914, n780, n763, n801, n858);
nand g932 (n925, n834, n808, n851, n493);
xor  g933 (n947, n863, n833, n740, n746);
and  g934 (n886, n804, n832, n792, n776);
xnor g935 (n877, n789, n718, n501, n724);
nor  g936 (n889, n735, n440, n496, n741);
nand g937 (n888, n825, n768, n766, n815);
xnor g938 (n909, n757, n814, n775, n817);
or   g939 (n996, n723, n811, n502, n848);
xor  g940 (n930, n798, n738, n852, n745);
or   g941 (n971, n441, n782, n714, n721);
and  g942 (n934, n722, n744, n858, n788);
and  g943 (n904, n720, n736, n827, n829);
or   g944 (n893, n864, n855, n499, n738);
and  g945 (n985, n823, n500, n756, n819);
nor  g946 (n900, n836, n498, n872, n795);
or   g947 (n875, n829, n775, n498, n847);
xnor g948 (n967, n853, n816, n750, n713);
xnor g949 (n905, n440, n756, n493, n799);
xor  g950 (n956, n813, n714, n853, n787);
and  g951 (n968, n867, n773, n865, n828);
nand g952 (n923, n832, n493, n870, n502);
and  g953 (n910, n810, n732, n770, n829);
xnor g954 (n950, n828, n731, n737, n858);
and  g955 (n954, n872, n498, n814, n497);
nor  g956 (n916, n794, n842, n741, n495);
nor  g957 (n939, n859, n711, n855, n833);
and  g958 (n989, n818, n844, n839, n854);
nor  g959 (n913, n792, n854, n760, n715);
nor  g960 (n992, n851, n856, n788, n500);
nor  g961 (n911, n793, n841, n846, n814);
or   g962 (n982, n843, n862, n854, n784);
or   g963 (n974, n743, n494, n853, n439);
or   g964 (n912, n760, n769, n842, n820);
nand g965 (n876, n749, n848, n790, n742);
nand g966 (n988, n811, n850, n733, n820);
nor  g967 (n957, n785, n859, n839, n723);
xnor g968 (n1004, n878, n920, n958, n953);
nor  g969 (n1008, n996, n905, n992, n933);
or   g970 (n1021, n894, n909, n961, n918);
nand g971 (n1012, n881, n998, n934, n962);
xnor g972 (n1005, n883, n923, n874, n989);
nor  g973 (n1029, n939, n899, n926, n1000);
xor  g974 (n1023, n877, n959, n990, n936);
or   g975 (n1003, n982, n978, n882, n980);
nor  g976 (n1026, n949, n965, n979, n976);
nand g977 (n1013, n937, n960, n928, n999);
and  g978 (n1025, n985, n925, n890, n993);
and  g979 (n1010, n893, n900, n930, n895);
xor  g980 (n1011, n947, n903, n889, n946);
xnor g981 (n1015, n885, n897, n932, n983);
and  g982 (n1018, n986, n921, n951, n945);
xor  g983 (n1019, n964, n922, n896, n944);
nand g984 (n1027, n876, n888, n913, n910);
xnor g985 (n1009, n919, n972, n943, n935);
xnor g986 (n1028, n908, n954, n955, n880);
and  g987 (n1017, n940, n884, n929, n892);
xor  g988 (n1024, n995, n912, n991, n963);
nand g989 (n1030, n974, n952, n956, n970);
nor  g990 (n1016, n975, n948, n994, n927);
nand g991 (n1032, n906, n988, n931, n969);
xnor g992 (n1014, n981, n917, n987, n967);
nor  g993 (n1002, n957, n941, n875, n942);
xnor g994 (n1020, n911, n916, n887, n915);
xnor g995 (n1007, n977, n886, n966, n984);
nor  g996 (n1006, n898, n907, n971, n968);
and  g997 (n1022, n873, n904, n902, n924);
xor  g998 (n1001, n938, n950, n891, n914);
nand g999 (n1031, n997, n901, n973, n879);
endmodule
