

module Stat_100_47
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n110,
  n132,
  n126,
  n125,
  n102,
  n121,
  n127,
  n112,
  n115,
  n129,
  n119,
  n109,
  n107,
  n108,
  n128,
  n131,
  n114,
  n103,
  n104,
  n113,
  n111,
  n122,
  n105,
  n117,
  n118,
  n124,
  n101,
  n120,
  n116,
  n123,
  n106,
  n130
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n110;output n132;output n126;output n125;output n102;output n121;output n127;output n112;output n115;output n129;output n119;output n109;output n107;output n108;output n128;output n131;output n114;output n103;output n104;output n113;output n111;output n122;output n105;output n117;output n118;output n124;output n101;output n120;output n116;output n123;output n106;output n130;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    KeyWire_0_16,
    n1
  );


  buf
  g1
  (
    n37,
    n1
  );


  buf
  g2
  (
    n34,
    n1
  );


  not
  g3
  (
    n36,
    n2
  );


  not
  g4
  (
    KeyWire_0_44,
    n1
  );


  buf
  g5
  (
    n45,
    n34
  );


  buf
  g6
  (
    n46,
    n35
  );


  not
  g7
  (
    KeyWire_0_4,
    n34
  );


  buf
  g8
  (
    KeyWire_0_29,
    n34
  );


  buf
  g9
  (
    KeyWire_0_3,
    n33
  );


  buf
  g10
  (
    n42,
    n35
  );


  buf
  g11
  (
    KeyWire_0_12,
    n33
  );


  not
  g12
  (
    n44,
    n37
  );


  buf
  g13
  (
    n47,
    n36
  );


  buf
  g14
  (
    KeyWire_0_9,
    n33
  );


  buf
  g15
  (
    n38,
    n34
  );


  buf
  g16
  (
    n41,
    n37
  );


  buf
  g17
  (
    KeyWire_0_6,
    n36
  );


  not
  g18
  (
    KeyWire_0_5,
    n37
  );


  buf
  g19
  (
    n43,
    n33
  );


  buf
  g20
  (
    KeyWire_0_40,
    n36
  );


  buf
  g21
  (
    n51,
    n35
  );


  not
  g22
  (
    KeyWire_0_26,
    n35
  );


  buf
  g23
  (
    n39,
    n36
  );


  not
  g24
  (
    n79,
    n28
  );


  buf
  g25
  (
    KeyWire_0_56,
    n9
  );


  and
  g26
  (
    KeyWire_0_23,
    n47,
    n18,
    n8,
    n29
  );


  nor
  g27
  (
    KeyWire_0_52,
    n26,
    n8,
    n55,
    n20
  );


  or
  g28
  (
    KeyWire_0_25,
    n48,
    n11,
    n56,
    n6
  );


  xnor
  g29
  (
    KeyWire_0_0,
    n31,
    n42,
    n45,
    n29
  );


  xor
  g30
  (
    KeyWire_0_57,
    n7,
    n2,
    n50
  );


  xnor
  g31
  (
    n78,
    n22,
    n25,
    n13,
    n26
  );


  xor
  g32
  (
    KeyWire_0_39,
    n52,
    n5,
    n7,
    n40
  );


  nand
  g33
  (
    KeyWire_0_42,
    n52,
    n10,
    n7,
    n21
  );


  nor
  g34
  (
    KeyWire_0_63,
    n14,
    n11,
    n32,
    n21
  );


  or
  g35
  (
    KeyWire_0_60,
    n12,
    n17,
    n28,
    n21
  );


  nor
  g36
  (
    KeyWire_0_62,
    n6,
    n48,
    n41,
    n4
  );


  xor
  g37
  (
    KeyWire_0_13,
    n30,
    n16,
    n51,
    n27
  );


  nand
  g38
  (
    n71,
    n12,
    n4,
    n31,
    n27
  );


  nor
  g39
  (
    KeyWire_0_22,
    n53,
    n14,
    n17,
    n23
  );


  nor
  g40
  (
    KeyWire_0_48,
    n11,
    n15,
    n4,
    n25
  );


  or
  g41
  (
    KeyWire_0_10,
    n54,
    n26,
    n25,
    n3
  );


  and
  g42
  (
    n72,
    n24,
    n31,
    n9,
    n18
  );


  or
  g43
  (
    n97,
    n27,
    n22,
    n6,
    n24
  );


  or
  g44
  (
    KeyWire_0_21,
    n49,
    n43,
    n56,
    n39
  );


  and
  g45
  (
    KeyWire_0_53,
    n12,
    n52,
    n23,
    n51
  );


  nand
  g46
  (
    n61,
    n19,
    n50,
    n9
  );


  and
  g47
  (
    KeyWire_0_31,
    n22,
    n56,
    n28,
    n20
  );


  or
  g48
  (
    n84,
    n15,
    n19,
    n17,
    n47
  );


  xnor
  g49
  (
    KeyWire_0_45,
    n14,
    n19,
    n54,
    n16
  );


  or
  g50
  (
    KeyWire_0_33,
    n10,
    n13,
    n52,
    n51
  );


  xnor
  g51
  (
    n57,
    n46,
    n55,
    n18,
    n38
  );


  or
  g52
  (
    KeyWire_0_55,
    n29,
    n6,
    n48,
    n54
  );


  nand
  g53
  (
    KeyWire_0_46,
    n16,
    n15,
    n12,
    n14
  );


  and
  g54
  (
    n88,
    n51,
    n23,
    n47,
    n3
  );


  xor
  g55
  (
    KeyWire_0_14,
    n19,
    n30,
    n56,
    n47
  );


  or
  g56
  (
    n86,
    n3,
    n55,
    n15,
    n18
  );


  nor
  g57
  (
    KeyWire_0_34,
    n2,
    n13,
    n5,
    n10
  );


  and
  g58
  (
    KeyWire_0_2,
    n13,
    n32,
    n48,
    n11
  );


  and
  g59
  (
    n80,
    n23,
    n44,
    n7,
    n55
  );


  nor
  g60
  (
    KeyWire_0_38,
    n49,
    n20,
    n5,
    n54
  );


  or
  g61
  (
    KeyWire_0_37,
    n10,
    n8,
    n28,
    n26
  );


  or
  g62
  (
    n87,
    n17,
    n20,
    n2,
    n5
  );


  and
  g63
  (
    KeyWire_0_28,
    n4,
    n53,
    n49,
    n3
  );


  xnor
  g64
  (
    KeyWire_0_54,
    n31,
    n24,
    n27
  );


  xnor
  g65
  (
    KeyWire_0_24,
    n16,
    n29,
    n22,
    n50
  );


  xor
  g66
  (
    n96,
    n49,
    n53,
    n8
  );


  xnor
  g67
  (
    n90,
    n21,
    n30,
    n25
  );


  nor
  g68
  (
    n119,
    n79,
    n94,
    n64,
    n58
  );


  xor
  g69
  (
    KeyWire_0_30,
    n100,
    n79,
    n81,
    n87
  );


  xnor
  g70
  (
    KeyWire_0_35,
    n85,
    n98,
    n92,
    n91
  );


  nand
  g71
  (
    KeyWire_0_36,
    n78,
    n76,
    n95,
    n83
  );


  or
  g72
  (
    KeyWire_0_51,
    n67,
    n76,
    n92,
    n77
  );


  or
  g73
  (
    n105,
    n92,
    n95,
    n79,
    n68
  );


  nor
  g74
  (
    KeyWire_0_1,
    n95,
    n93,
    n80,
    n79
  );


  xor
  g75
  (
    KeyWire_0_47,
    n94,
    n94,
    n81,
    n90
  );


  xnor
  g76
  (
    KeyWire_0_32,
    n61,
    n77,
    n87,
    n82
  );


  and
  g77
  (
    KeyWire_0_41,
    n63,
    n72,
    n87,
    n78
  );


  or
  g78
  (
    KeyWire_0_11,
    n73,
    n96,
    n84,
    n80
  );


  xnor
  g79
  (
    KeyWire_0_20,
    n96,
    n97,
    n81,
    n74
  );


  and
  g80
  (
    KeyWire_0_27,
    n84,
    n96,
    n71,
    n83
  );


  nor
  g81
  (
    KeyWire_0_58,
    n85,
    n88,
    n84,
    n98
  );


  and
  g82
  (
    n111,
    n65,
    n100,
    n97,
    n94
  );


  and
  g83
  (
    KeyWire_0_59,
    n88,
    n59,
    n76,
    n99
  );


  or
  g84
  (
    KeyWire_0_43,
    n75,
    n60,
    n97,
    n57
  );


  or
  g85
  (
    KeyWire_0_19,
    n74,
    n66,
    n77,
    n93
  );


  xor
  g86
  (
    KeyWire_0_17,
    n77,
    n99,
    n93,
    n74
  );


  xor
  g87
  (
    n102,
    n89,
    n86,
    n90,
    n82
  );


  nor
  g88
  (
    KeyWire_0_15,
    n82,
    n90,
    n76,
    n78
  );


  nor
  g89
  (
    KeyWire_0_18,
    n89,
    n82,
    n88,
    n100
  );


  xor
  g90
  (
    n120,
    n83,
    n88,
    n86,
    n91
  );


  nand
  g91
  (
    n125,
    n100,
    n99,
    n32,
    n75
  );


  xor
  g92
  (
    KeyWire_0_7,
    n93,
    n92,
    n74,
    n98
  );


  xnor
  g93
  (
    n106,
    n99,
    n70,
    n80
  );


  or
  g94
  (
    KeyWire_0_49,
    n90,
    n87,
    n91,
    n69
  );


  xnor
  g95
  (
    KeyWire_0_50,
    n86,
    n78,
    n98,
    n83
  );


  and
  g96
  (
    n126,
    n95,
    n62,
    n85,
    n89
  );


  xor
  g97
  (
    KeyWire_0_8,
    n84,
    n37,
    n91,
    n97
  );


  and
  g98
  (
    KeyWire_0_61,
    n86,
    n85,
    n75
  );


  and
  g99
  (
    n107,
    n32,
    n89,
    n81,
    n96
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n63,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n108,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n68,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n56,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n40,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n54,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n55,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n103,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n117,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n52,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n89,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n131,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n53,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n58,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n74,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n113,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n33,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n109,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n122,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n112,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n127,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n83,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n93,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n65,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n95,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n91,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n49,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n116,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n99,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n48,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n115,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n73,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n128,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n81,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n76,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n123,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n132,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n59,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n64,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n92,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n50,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n121,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n67,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n130,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n35,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n100,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n62,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n118,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n66,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n114,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n104,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n101,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n70,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n98,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n77,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n69,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n75,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n82,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n129,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n124,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n60,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n110,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n85,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n94,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


