// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_392_937 written by SynthGen on 2021/05/24 19:47:35
module Stat_392_937( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23,
 n399, n403, n395, n396, n408, n397, n414, n405,
 n410, n398, n411, n413, n407, n400, n393, n409,
 n402, n415, n404, n401, n394, n412, n406);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23;

output n399, n403, n395, n396, n408, n397, n414, n405,
 n410, n398, n411, n413, n407, n400, n393, n409,
 n402, n415, n404, n401, n394, n412, n406;

wire n24, n25, n26, n27, n28, n29, n30, n31,
 n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392;

not  g0 (n24, n1);
not  g1 (n37, n4);
not  g2 (n29, n2);
not  g3 (n33, n2);
buf  g4 (n25, n1);
not  g5 (n30, n1);
not  g6 (n36, n3);
not  g7 (n26, n3);
not  g8 (n32, n2);
buf  g9 (n35, n4);
buf  g10 (n34, n1);
buf  g11 (n31, n3);
buf  g12 (n27, n2);
not  g13 (n28, n3);
not  g14 (n50, n24);
buf  g15 (n41, n29);
buf  g16 (n59, n28);
buf  g17 (n55, n27);
buf  g18 (n42, n26);
buf  g19 (n43, n25);
buf  g20 (n48, n26);
not  g21 (n58, n24);
buf  g22 (n52, n29);
buf  g23 (n57, n27);
buf  g24 (n39, n24);
buf  g25 (n46, n27);
not  g26 (n44, n25);
buf  g27 (n40, n24);
buf  g28 (n45, n30);
not  g29 (n38, n27);
not  g30 (n53, n26);
buf  g31 (n60, n25);
buf  g32 (n56, n28);
buf  g33 (n51, n29);
not  g34 (n54, n26);
not  g35 (n47, n28);
buf  g36 (n61, n28);
not  g37 (n62, n25);
not  g38 (n49, n29);
not  g39 (n75, n39);
buf  g40 (n68, n45);
not  g41 (n83, n40);
not  g42 (n78, n41);
buf  g43 (n73, n42);
buf  g44 (n79, n46);
buf  g45 (n66, n39);
buf  g46 (n65, n38);
not  g47 (n80, n42);
buf  g48 (n76, n48);
not  g49 (n64, n47);
not  g50 (n71, n46);
buf  g51 (n77, n45);
not  g52 (n69, n43);
not  g53 (n72, n43);
buf  g54 (n70, n41);
not  g55 (n82, n47);
buf  g56 (n67, n44);
buf  g57 (n74, n44);
buf  g58 (n81, n48);
not  g59 (n63, n40);
buf  g60 (n105, n71);
buf  g61 (n136, n63);
not  g62 (n107, n70);
buf  g63 (n93, n65);
buf  g64 (n91, n63);
buf  g65 (n114, n75);
not  g66 (n87, n76);
buf  g67 (n96, n69);
not  g68 (n89, n68);
not  g69 (n110, n68);
not  g70 (n137, n71);
not  g71 (n104, n74);
not  g72 (n102, n64);
not  g73 (n113, n65);
buf  g74 (n116, n73);
buf  g75 (n126, n66);
not  g76 (n106, n67);
not  g77 (n88, n70);
buf  g78 (n123, n75);
buf  g79 (n86, n70);
buf  g80 (n98, n69);
buf  g81 (n109, n74);
not  g82 (n131, n69);
buf  g83 (n128, n66);
not  g84 (n135, n75);
not  g85 (n118, n63);
not  g86 (n108, n72);
buf  g87 (n115, n72);
not  g88 (n85, n74);
buf  g89 (n99, n74);
not  g90 (n133, n64);
not  g91 (n117, n63);
not  g92 (n125, n76);
not  g93 (n132, n72);
buf  g94 (n122, n69);
buf  g95 (n95, n72);
not  g96 (n134, n73);
buf  g97 (n121, n75);
buf  g98 (n97, n67);
not  g99 (n101, n70);
not  g100 (n90, n71);
buf  g101 (n103, n67);
buf  g102 (n130, n76);
not  g103 (n111, n68);
buf  g104 (n139, n65);
buf  g105 (n129, n67);
not  g106 (n127, n73);
not  g107 (n120, n71);
buf  g108 (n84, n68);
not  g109 (n92, n73);
buf  g110 (n119, n66);
not  g111 (n112, n66);
not  g112 (n94, n76);
not  g113 (n100, n65);
not  g114 (n138, n64);
buf  g115 (n124, n64);
not  g116 (n199, n116);
not  g117 (n183, n96);
not  g118 (n181, n111);
not  g119 (n155, n22);
not  g120 (n141, n84);
buf  g121 (n158, n125);
buf  g122 (n178, n86);
not  g123 (n184, n101);
not  g124 (n210, n5);
not  g125 (n145, n112);
not  g126 (n186, n100);
buf  g127 (n177, n118);
not  g128 (n148, n90);
not  g129 (n195, n115);
and  g130 (n176, n95, n112, n11, n86);
nor  g131 (n206, n120, n22, n121, n92);
nor  g132 (n157, n110, n116, n106, n92);
xnor g133 (n191, n84, n14, n113, n115);
nor  g134 (n179, n85, n113, n104, n110);
nor  g135 (n156, n12, n120, n18, n104);
nor  g136 (n162, n115, n10, n12, n101);
nand g137 (n147, n119, n93, n90, n100);
nand g138 (n182, n102, n21, n119, n118);
xnor g139 (n154, n125, n114, n5, n97);
xor  g140 (n149, n15, n113, n122, n21);
nand g141 (n205, n10, n12, n7, n95);
xnor g142 (n173, n87, n10, n19, n14);
xnor g143 (n172, n98, n86, n18, n95);
xnor g144 (n152, n85, n102, n98, n124);
or   g145 (n194, n93, n20, n13, n89);
xnor g146 (n207, n5, n94, n95, n86);
nand g147 (n203, n123, n14, n104, n119);
xor  g148 (n165, n11, n122, n124, n109);
xor  g149 (n200, n8, n104, n22, n93);
nor  g150 (n174, n90, n119, n109, n107);
nor  g151 (n167, n121, n85, n108, n4);
xor  g152 (n202, n106, n102, n96, n89);
or   g153 (n185, n6, n17, n124, n111);
xnor g154 (n159, n114, n102, n92, n108);
or   g155 (n196, n121, n84, n93, n17);
nor  g156 (n198, n21, n18, n94, n88);
xor  g157 (n169, n117, n112, n6, n22);
nand g158 (n146, n8, n88, n106, n107);
nor  g159 (n144, n105, n96, n111, n13);
xnor g160 (n201, n88, n15, n87, n97);
xor  g161 (n175, n113, n120, n122, n16);
nand g162 (n142, n108, n8, n7, n18);
xnor g163 (n153, n111, n94, n96, n91);
and  g164 (n190, n13, n7, n100, n9);
nor  g165 (n150, n84, n109, n6, n100);
xnor g166 (n197, n91, n5, n121, n17);
and  g167 (n192, n123, n99, n98, n21);
or   g168 (n168, n124, n15, n103, n90);
nor  g169 (n204, n8, n108, n16, n103);
and  g170 (n143, n15, n20, n13, n114);
nand g171 (n160, n20, n94, n19, n120);
nand g172 (n193, n91, n11, n110, n17);
xor  g173 (n208, n122, n16, n106, n9);
xnor g174 (n189, n107, n97, n12, n89);
nor  g175 (n166, n101, n99, n23, n16);
or   g176 (n171, n117, n9, n116, n92);
or   g177 (n161, n114, n123, n101, n105);
and  g178 (n151, n19, n118, n105, n112);
and  g179 (n163, n103, n118, n9, n14);
nand g180 (n209, n117, n116, n19, n87);
xnor g181 (n187, n110, n88, n91, n87);
nor  g182 (n180, n10, n89, n7, n6);
xnor g183 (n170, n109, n23, n115, n117);
or   g184 (n188, n11, n103, n99, n20);
nor  g185 (n140, n98, n85, n97, n107);
xor  g186 (n164, n105, n123, n4, n99);
buf  g187 (n259, n162);
not  g188 (n223, n158);
buf  g189 (n219, n156);
not  g190 (n231, n153);
not  g191 (n220, n166);
not  g192 (n255, n153);
not  g193 (n243, n164);
buf  g194 (n237, n156);
not  g195 (n236, n165);
not  g196 (n214, n151);
not  g197 (n215, n163);
not  g198 (n252, n144);
buf  g199 (n249, n171);
buf  g200 (n253, n174);
buf  g201 (n212, n167);
not  g202 (n230, n168);
buf  g203 (n225, n150);
buf  g204 (n216, n172);
buf  g205 (n261, n157);
not  g206 (n222, n162);
buf  g207 (n227, n152);
not  g208 (n257, n164);
not  g209 (n256, n155);
buf  g210 (n260, n166);
buf  g211 (n244, n170);
buf  g212 (n213, n168);
buf  g213 (n238, n165);
buf  g214 (n258, n163);
not  g215 (n226, n167);
not  g216 (n228, n150);
not  g217 (n248, n157);
not  g218 (n232, n161);
buf  g219 (n239, n148);
buf  g220 (n240, n155);
buf  g221 (n224, n149);
buf  g222 (n221, n154);
buf  g223 (n241, n175);
buf  g224 (n229, n151);
not  g225 (n235, n175);
not  g226 (n211, n170);
buf  g227 (n246, n176);
buf  g228 (n254, n141);
buf  g229 (n217, n158);
buf  g230 (n262, n143);
buf  g231 (n247, n172);
not  g232 (n251, n173);
not  g233 (n245, n146);
buf  g234 (n242, n173);
xnor g235 (n233, n174, n159, n169, n161);
xor  g236 (n218, n160, n149, n159, n169);
and  g237 (n250, n160, n154, n147, n142);
nor  g238 (n234, n145, n152, n140, n171);
or   g239 (n315, n208, n202, n225, n199);
nand g240 (n299, n229, n227, n197, n177);
and  g241 (n331, n204, n201, n254, n229);
or   g242 (n302, n204, n240, n202, n255);
nand g243 (n274, n207, n260, n252, n190);
nand g244 (n319, n218, n230, n236, n256);
nor  g245 (n291, n183, n241, n255, n246);
nor  g246 (n306, n199, n215, n252, n253);
xor  g247 (n280, n194, n206, n259, n180);
or   g248 (n344, n33, n182, n200, n219);
and  g249 (n263, n228, n185, n243, n180);
nand g250 (n296, n254, n254, n49, n196);
or   g251 (n316, n225, n258, n213, n256);
nor  g252 (n339, n203, n58, n222, n259);
xor  g253 (n286, n235, n217, n176, n224);
nand g254 (n295, n230, n233, n262, n208);
xor  g255 (n334, n223, n216, n183, n227);
xnor g256 (n325, n209, n210, n187, n217);
or   g257 (n345, n247, n205, n34, n202);
or   g258 (n271, n236, n52, n228, n50);
nand g259 (n355, n238, n185, n226, n178);
xor  g260 (n288, n232, n57, n33, n240);
nand g261 (n273, n213, n216, n234, n30);
nor  g262 (n303, n245, n178, n181, n220);
nor  g263 (n323, n230, n195, n248, n228);
nor  g264 (n298, n62, n246, n60, n204);
xor  g265 (n264, n203, n221, n248, n179);
xnor g266 (n292, n196, n198, n257, n237);
and  g267 (n324, n257, n195, n53, n238);
xnor g268 (n279, n211, n198, n53, n260);
and  g269 (n352, n190, n198, n33, n32);
xor  g270 (n276, n249, n258, n219, n177);
xnor g271 (n275, n251, n258, n32, n252);
nand g272 (n332, n193, n210, n239, n214);
and  g273 (n343, n237, n193, n52, n31);
xnor g274 (n349, n199, n214, n207, n210);
and  g275 (n267, n184, n259, n215, n261);
nor  g276 (n317, n197, n30, n227, n242);
or   g277 (n353, n250, n222, n229, n232);
xnor g278 (n328, n59, n235, n221, n191);
nor  g279 (n351, n187, n215, n186, n238);
nand g280 (n341, n54, n250, n242, n193);
and  g281 (n300, n225, n247, n233, n198);
and  g282 (n333, n219, n251, n246, n248);
nand g283 (n304, n245, n243, n261, n31);
nor  g284 (n294, n182, n34, n197, n212);
or   g285 (n322, n234, n236, n190, n215);
nor  g286 (n283, n253, n35, n61, n216);
or   g287 (n270, n184, n209, n260, n186);
or   g288 (n312, n192, n234, n194, n23);
nand g289 (n301, n235, n207, n241, n210);
xnor g290 (n313, n254, n194, n196, n244);
xor  g291 (n342, n245, n230, n229, n255);
xor  g292 (n284, n239, n214, n244, n192);
and  g293 (n268, n257, n208, n255, n233);
or   g294 (n307, n189, n189, n219, n221);
nand g295 (n277, n61, n227, n197, n261);
xnor g296 (n290, n231, n200, n220, n30);
xnor g297 (n348, n221, n202, n231, n56);
xnor g298 (n272, n32, n31, n238, n239);
and  g299 (n326, n54, n223, n182, n257);
nor  g300 (n356, n192, n256, n232, n199);
nand g301 (n338, n188, n249, n204, n245);
nand g302 (n309, n212, n201, n49, n250);
xor  g303 (n269, n50, n212, n183, n251);
xnor g304 (n327, n185, n187, n188, n205);
or   g305 (n311, n253, n222, n191, n205);
and  g306 (n285, n218, n225, n224, n188);
or   g307 (n308, n195, n243, n59, n248);
and  g308 (n310, n240, n247, n193, n218);
and  g309 (n337, n251, n182, n207, n208);
nand g310 (n318, n241, n226, n234, n224);
and  g311 (n346, n31, n55, n214, n216);
nor  g312 (n314, n223, n190, n256, n262);
nand g313 (n329, n247, n51, n60, n261);
or   g314 (n297, n184, n262, n236, n200);
xor  g315 (n320, n258, n181, n253, n239);
and  g316 (n278, n246, n189, n58, n213);
xor  g317 (n350, n185, n220, n206, n188);
xnor g318 (n335, n206, n241, n209, n203);
and  g319 (n357, n194, n212, n237, n235);
nor  g320 (n347, n183, n217, n213);
xnor g321 (n266, n203, n243, n201, n244);
and  g322 (n293, n262, n226, n55, n231);
nor  g323 (n358, n201, n249, n244, n224);
nor  g324 (n282, n191, n220, n249, n184);
xnor g325 (n336, n192, n260, n237, n196);
xor  g326 (n265, n242, n223, n179, n189);
nor  g327 (n281, n259, n205, n51, n186);
and  g328 (n330, n57, n56, n250, n195);
nor  g329 (n340, n187, n206, n232, n222);
and  g330 (n321, n209, n211, n33, n34);
and  g331 (n354, n228, n181, n218, n32);
or   g332 (n287, n252, n200, n233, n23);
xor  g333 (n305, n242, n186, n191, n240);
nand g334 (n289, n181, n231, n34, n226);
nor  g335 (n380, n355, n340, n290, n62);
nand g336 (n373, n281, n83, n351, n36);
or   g337 (n364, n343, n319, n317, n35);
nor  g338 (n377, n273, n282, n287, n35);
xor  g339 (n367, n350, n323, n306, n81);
xor  g340 (n387, n325, n302, n283, n295);
nand g341 (n362, n298, n313, n336, n288);
xnor g342 (n389, n324, n307, n81, n82);
or   g343 (n375, n80, n83, n267, n345);
nor  g344 (n392, n321, n37, n286, n263);
xnor g345 (n388, n80, n320, n266, n277);
nand g346 (n383, n356, n301, n357, n82);
xor  g347 (n363, n352, n304, n312, n293);
nor  g348 (n365, n272, n36, n309, n78);
xor  g349 (n374, n82, n81, n303, n326);
and  g350 (n390, n308, n331, n83, n285);
xnor g351 (n384, n289, n344, n314, n341);
nor  g352 (n391, n280, n354, n318, n347);
and  g353 (n376, n316, n268, n78, n264);
or   g354 (n368, n77, n333, n353, n327);
and  g355 (n359, n346, n77, n274, n35);
xor  g356 (n360, n37, n339, n292, n80);
nand g357 (n382, n335, n279, n77, n278);
nand g358 (n371, n83, n322, n358, n79);
nand g359 (n370, n79, n37, n299, n82);
xnor g360 (n372, n300, n276, n37, n275);
or   g361 (n385, n349, n310, n315, n338);
xor  g362 (n379, n328, n305, n79, n78);
and  g363 (n381, n296, n79, n311, n80);
nand g364 (n369, n297, n36, n77, n348);
nor  g365 (n366, n337, n294, n270, n265);
or   g366 (n361, n269, n291, n81, n334);
or   g367 (n386, n332, n78, n36, n271);
and  g368 (n378, n342, n330, n284, n329);
and  g369 (n411, n129, n132, n374);
nor  g370 (n399, n377, n133, n130, n135);
xnor g371 (n415, n371, n130, n135, n139);
or   g372 (n397, n128, n131, n137);
nor  g373 (n414, n135, n375, n360, n385);
or   g374 (n405, n128, n128, n138, n129);
xnor g375 (n398, n132, n362, n134, n126);
nor  g376 (n408, n384, n380, n369, n129);
nand g377 (n401, n364, n390, n135, n139);
nand g378 (n407, n359, n368, n125, n131);
nand g379 (n400, n125, n373, n131, n138);
or   g380 (n394, n379, n386, n365, n367);
xor  g381 (n413, n134, n137, n361, n139);
xnor g382 (n403, n127, n370, n388, n392);
or   g383 (n406, n139, n126, n382, n137);
nor  g384 (n409, n391, n133, n387, n372);
xnor g385 (n410, n126, n127, n133, n130);
xnor g386 (n395, n136, n378, n130, n138);
xor  g387 (n412, n389, n134, n127);
and  g388 (n393, n366, n128, n127, n136);
nand g389 (n402, n126, n133, n137, n138);
xor  g390 (n404, n383, n132, n363, n136);
xor  g391 (n396, n376, n129, n381, n136);
endmodule
