// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_222 written by SynthGen on 2021/04/05 11:23:25
module Stat_2000_222( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n83, n289, n339, n998, n831, n1002, n1072, n876,
 n1097, n967, n1087, n1064, n1039, n955, n978, n1093,
 n871, n965, n870, n1871, n1883, n2027, n2022, n2026,
 n2024, n2030, n2032, n2029, n2028, n2025, n2031, n2023);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n83, n289, n339, n998, n831, n1002, n1072, n876,
 n1097, n967, n1087, n1064, n1039, n955, n978, n1093,
 n871, n965, n870, n1871, n1883, n2027, n2022, n2026,
 n2024, n2030, n2032, n2029, n2028, n2025, n2031, n2023;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n340, n341, n342, n343, n344, n345, n346, n347,
 n348, n349, n350, n351, n352, n353, n354, n355,
 n356, n357, n358, n359, n360, n361, n362, n363,
 n364, n365, n366, n367, n368, n369, n370, n371,
 n372, n373, n374, n375, n376, n377, n378, n379,
 n380, n381, n382, n383, n384, n385, n386, n387,
 n388, n389, n390, n391, n392, n393, n394, n395,
 n396, n397, n398, n399, n400, n401, n402, n403,
 n404, n405, n406, n407, n408, n409, n410, n411,
 n412, n413, n414, n415, n416, n417, n418, n419,
 n420, n421, n422, n423, n424, n425, n426, n427,
 n428, n429, n430, n431, n432, n433, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n634, n635,
 n636, n637, n638, n639, n640, n641, n642, n643,
 n644, n645, n646, n647, n648, n649, n650, n651,
 n652, n653, n654, n655, n656, n657, n658, n659,
 n660, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685, n686, n687, n688, n689, n690, n691,
 n692, n693, n694, n695, n696, n697, n698, n699,
 n700, n701, n702, n703, n704, n705, n706, n707,
 n708, n709, n710, n711, n712, n713, n714, n715,
 n716, n717, n718, n719, n720, n721, n722, n723,
 n724, n725, n726, n727, n728, n729, n730, n731,
 n732, n733, n734, n735, n736, n737, n738, n739,
 n740, n741, n742, n743, n744, n745, n746, n747,
 n748, n749, n750, n751, n752, n753, n754, n755,
 n756, n757, n758, n759, n760, n761, n762, n763,
 n764, n765, n766, n767, n768, n769, n770, n771,
 n772, n773, n774, n775, n776, n777, n778, n779,
 n780, n781, n782, n783, n784, n785, n786, n787,
 n788, n789, n790, n791, n792, n793, n794, n795,
 n796, n797, n798, n799, n800, n801, n802, n803,
 n804, n805, n806, n807, n808, n809, n810, n811,
 n812, n813, n814, n815, n816, n817, n818, n819,
 n820, n821, n822, n823, n824, n825, n826, n827,
 n828, n829, n830, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n865, n866, n867, n868,
 n869, n872, n873, n874, n875, n877, n878, n879,
 n880, n881, n882, n883, n884, n885, n886, n887,
 n888, n889, n890, n891, n892, n893, n894, n895,
 n896, n897, n898, n899, n900, n901, n902, n903,
 n904, n905, n906, n907, n908, n909, n910, n911,
 n912, n913, n914, n915, n916, n917, n918, n919,
 n920, n921, n922, n923, n924, n925, n926, n927,
 n928, n929, n930, n931, n932, n933, n934, n935,
 n936, n937, n938, n939, n940, n941, n942, n943,
 n944, n945, n946, n947, n948, n949, n950, n951,
 n952, n953, n954, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n966, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n979,
 n980, n981, n982, n983, n984, n985, n986, n987,
 n988, n989, n990, n991, n992, n993, n994, n995,
 n996, n997, n999, n1000, n1001, n1003, n1004, n1005,
 n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
 n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
 n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
 n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
 n1038, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
 n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
 n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
 n1063, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1088, n1089,
 n1090, n1091, n1092, n1094, n1095, n1096, n1098, n1099,
 n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
 n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
 n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
 n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
 n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
 n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
 n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
 n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
 n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
 n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
 n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
 n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
 n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
 n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
 n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
 n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
 n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
 n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
 n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
 n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
 n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
 n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
 n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
 n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
 n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
 n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
 n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
 n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
 n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
 n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
 n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
 n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
 n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
 n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
 n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
 n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
 n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
 n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
 n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
 n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
 n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
 n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
 n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
 n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
 n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
 n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
 n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
 n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
 n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
 n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
 n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
 n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
 n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
 n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
 n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
 n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
 n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
 n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
 n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
 n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
 n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
 n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
 n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
 n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
 n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
 n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
 n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
 n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
 n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
 n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
 n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
 n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
 n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
 n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
 n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
 n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
 n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
 n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
 n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
 n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
 n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
 n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
 n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
 n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
 n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
 n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
 n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
 n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
 n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
 n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
 n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
 n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
 n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
 n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
 n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
 n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
 n1868, n1869, n1870, n1872, n1873, n1874, n1875, n1876,
 n1877, n1878, n1879, n1880, n1881, n1882, n1884, n1885,
 n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
 n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
 n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
 n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
 n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
 n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
 n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
 n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
 n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
 n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
 n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
 n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
 n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
 n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
 n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
 n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
 n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021;

buf  g0 (n47, n7);
buf  g1 (n34, n3);
not  g2 (n40, n6);
not  g3 (n60, n6);
not  g4 (n37, n7);
not  g5 (n38, n2);
buf  g6 (n33, n7);
buf  g7 (n54, n4);
buf  g8 (n49, n1);
not  g9 (n59, n2);
buf  g10 (n62, n8);
buf  g11 (n57, n5);
buf  g12 (n52, n5);
buf  g13 (n61, n8);
buf  g14 (n55, n1);
buf  g15 (n58, n7);
not  g16 (n53, n2);
buf  g17 (n43, n4);
buf  g18 (n44, n5);
buf  g19 (n46, n2);
buf  g20 (n56, n1);
not  g21 (n63, n3);
not  g22 (n39, n3);
buf  g23 (n51, n3);
not  g24 (n50, n4);
buf  g25 (n48, n6);
buf  g26 (n35, n8);
not  g27 (n45, n6);
not  g28 (n36, n1);
buf  g29 (n42, n4);
buf  g30 (n41, n5);
not  g31 (n121, n59);
buf  g32 (n181, n58);
not  g33 (n81, n60);
not  g34 (n139, n41);
not  g35 (n128, n49);
buf  g36 (n103, n37);
buf  g37 (n64, n54);
buf  g38 (n100, n44);
not  g39 (n158, n63);
not  g40 (n115, n58);
buf  g41 (n71, n59);
not  g42 (n177, n36);
buf  g43 (n160, n41);
buf  g44 (n68, n37);
not  g45 (n92, n52);
not  g46 (n186, n43);
buf  g47 (n164, n39);
not  g48 (n79, n54);
not  g49 (n182, n60);
not  g50 (n110, n34);
buf  g51 (n108, n48);
buf  g52 (n73, n52);
not  g53 (n78, n63);
not  g54 (n159, n58);
not  g55 (n83, n62);
buf  g56 (n187, n39);
buf  g57 (n173, n49);
not  g58 (n118, n48);
not  g59 (n113, n63);
not  g60 (n133, n53);
buf  g61 (n141, n42);
not  g62 (n179, n50);
not  g63 (n114, n57);
not  g64 (n180, n57);
buf  g65 (n161, n56);
buf  g66 (n163, n34);
buf  g67 (n87, n45);
not  g68 (n126, n46);
not  g69 (n104, n47);
not  g70 (n174, n35);
not  g71 (n96, n55);
not  g72 (n109, n33);
not  g73 (n91, n55);
buf  g74 (n152, n51);
not  g75 (n76, n35);
buf  g76 (n99, n62);
buf  g77 (n144, n48);
buf  g78 (n112, n46);
buf  g79 (n137, n33);
buf  g80 (n138, n60);
not  g81 (n67, n41);
buf  g82 (n65, n61);
not  g83 (n129, n60);
buf  g84 (n172, n37);
not  g85 (n165, n57);
not  g86 (n125, n41);
not  g87 (n127, n62);
buf  g88 (n148, n47);
buf  g89 (n82, n33);
buf  g90 (n157, n50);
buf  g91 (n135, n54);
buf  g92 (n106, n34);
buf  g93 (n124, n42);
not  g94 (n117, n45);
not  g95 (n88, n45);
not  g96 (n151, n56);
buf  g97 (n156, n53);
not  g98 (n105, n57);
buf  g99 (n131, n34);
buf  g100 (n145, n47);
not  g101 (n169, n39);
not  g102 (n97, n42);
not  g103 (n74, n55);
not  g104 (n143, n58);
buf  g105 (n175, n56);
not  g106 (n154, n40);
buf  g107 (n116, n46);
buf  g108 (n80, n44);
not  g109 (n72, n59);
not  g110 (n94, n59);
buf  g111 (n66, n61);
buf  g112 (n155, n50);
not  g113 (n146, n51);
buf  g114 (n90, n62);
buf  g115 (n132, n51);
buf  g116 (n147, n63);
not  g117 (n107, n43);
not  g118 (n101, n51);
buf  g119 (n77, n35);
buf  g120 (n85, n36);
not  g121 (n167, n40);
not  g122 (n178, n52);
buf  g123 (n119, n38);
buf  g124 (n122, n40);
not  g125 (n176, n53);
buf  g126 (n166, n47);
buf  g127 (n168, n43);
not  g128 (n134, n43);
buf  g129 (n140, n55);
not  g130 (n170, n38);
not  g131 (n98, n61);
buf  g132 (n111, n46);
buf  g133 (n123, n54);
buf  g134 (n130, n39);
not  g135 (n183, n38);
buf  g136 (n70, n48);
not  g137 (n93, n56);
buf  g138 (n150, n35);
buf  g139 (n136, n61);
not  g140 (n69, n36);
buf  g141 (n171, n52);
not  g142 (n86, n49);
not  g143 (n162, n37);
not  g144 (n95, n44);
not  g145 (n102, n33);
not  g146 (n75, n50);
buf  g147 (n184, n38);
buf  g148 (n153, n49);
buf  g149 (n142, n45);
buf  g150 (n89, n40);
not  g151 (n84, n44);
buf  g152 (n185, n42);
not  g153 (n149, n36);
not  g154 (n120, n53);
buf  g155 (n433, n65);
buf  g156 (n313, n96);
buf  g157 (n192, n135);
not  g158 (n398, n102);
not  g159 (n269, n79);
buf  g160 (n213, n131);
buf  g161 (n263, n80);
buf  g162 (n209, n119);
buf  g163 (n397, n96);
not  g164 (n326, n137);
not  g165 (n412, n130);
not  g166 (n280, n141);
buf  g167 (n310, n97);
not  g168 (n282, n119);
not  g169 (n381, n116);
not  g170 (n416, n84);
not  g171 (n320, n105);
not  g172 (n427, n136);
not  g173 (n242, n133);
buf  g174 (n262, n115);
not  g175 (n333, n125);
not  g176 (n402, n88);
not  g177 (n226, n121);
not  g178 (n272, n85);
buf  g179 (n250, n84);
buf  g180 (n220, n95);
not  g181 (n383, n104);
not  g182 (n434, n112);
buf  g183 (n240, n129);
not  g184 (n445, n97);
not  g185 (n329, n85);
buf  g186 (n404, n73);
buf  g187 (n254, n142);
buf  g188 (n447, n89);
buf  g189 (n258, n103);
buf  g190 (n260, n66);
buf  g191 (n345, n82);
buf  g192 (n222, n94);
buf  g193 (n439, n126);
not  g194 (n230, n117);
buf  g195 (n432, n83);
not  g196 (n219, n99);
buf  g197 (n245, n138);
not  g198 (n335, n67);
not  g199 (n443, n70);
not  g200 (n415, n88);
not  g201 (n444, n143);
not  g202 (n207, n132);
buf  g203 (n261, n134);
not  g204 (n348, n92);
not  g205 (n462, n134);
not  g206 (n373, n87);
not  g207 (n248, n82);
buf  g208 (n198, n90);
not  g209 (n399, n65);
buf  g210 (n332, n117);
not  g211 (n237, n103);
buf  g212 (n425, n140);
not  g213 (n300, n100);
not  g214 (n211, n117);
buf  g215 (n372, n109);
not  g216 (n252, n107);
buf  g217 (n291, n132);
not  g218 (n243, n81);
not  g219 (n442, n129);
not  g220 (n461, n118);
not  g221 (n297, n88);
buf  g222 (n351, n74);
not  g223 (n414, n144);
buf  g224 (n359, n71);
buf  g225 (n403, n101);
not  g226 (n380, n113);
not  g227 (n370, n122);
buf  g228 (n441, n77);
buf  g229 (n301, n83);
buf  g230 (n321, n120);
buf  g231 (n424, n140);
not  g232 (n318, n80);
not  g233 (n188, n125);
buf  g234 (n354, n143);
not  g235 (n435, n87);
not  g236 (n361, n137);
buf  g237 (n456, n113);
buf  g238 (n305, n64);
buf  g239 (n277, n123);
not  g240 (n306, n95);
buf  g241 (n457, n124);
buf  g242 (n249, n130);
not  g243 (n239, n86);
buf  g244 (n406, n132);
buf  g245 (n355, n88);
buf  g246 (n307, n109);
not  g247 (n448, n96);
buf  g248 (n256, n87);
not  g249 (n394, n94);
buf  g250 (n460, n109);
not  g251 (n322, n138);
buf  g252 (n386, n95);
buf  g253 (n289, n133);
buf  g254 (n304, n141);
not  g255 (n193, n139);
not  g256 (n238, n72);
buf  g257 (n257, n107);
not  g258 (n266, n117);
not  g259 (n377, n132);
buf  g260 (n431, n102);
not  g261 (n452, n122);
buf  g262 (n411, n140);
not  g263 (n352, n116);
not  g264 (n255, n138);
buf  g265 (n276, n82);
buf  g266 (n421, n89);
not  g267 (n270, n90);
buf  g268 (n298, n111);
not  g269 (n204, n86);
buf  g270 (n367, n119);
buf  g271 (n410, n74);
not  g272 (n206, n99);
not  g273 (n316, n128);
not  g274 (n196, n91);
buf  g275 (n217, n85);
buf  g276 (n283, n108);
buf  g277 (n311, n86);
buf  g278 (n393, n121);
not  g279 (n303, n105);
buf  g280 (n340, n115);
buf  g281 (n227, n94);
buf  g282 (n287, n84);
not  g283 (n286, n92);
buf  g284 (n293, n104);
not  g285 (n374, n94);
buf  g286 (n378, n114);
not  g287 (n194, n112);
buf  g288 (n247, n83);
not  g289 (n224, n81);
buf  g290 (n376, n108);
buf  g291 (n360, n106);
buf  g292 (n234, n119);
not  g293 (n218, n101);
not  g294 (n265, n75);
buf  g295 (n429, n145);
not  g296 (n323, n103);
buf  g297 (n195, n133);
buf  g298 (n387, n118);
buf  g299 (n274, n139);
buf  g300 (n459, n69);
buf  g301 (n317, n64);
not  g302 (n437, n128);
not  g303 (n401, n105);
not  g304 (n369, n122);
buf  g305 (n395, n145);
not  g306 (n210, n74);
not  g307 (n446, n140);
not  g308 (n338, n93);
not  g309 (n407, n93);
buf  g310 (n251, n137);
buf  g311 (n353, n144);
not  g312 (n396, n92);
buf  g313 (n454, n71);
buf  g314 (n229, n84);
buf  g315 (n418, n121);
buf  g316 (n392, n116);
buf  g317 (n357, n126);
buf  g318 (n267, n141);
buf  g319 (n236, n100);
buf  g320 (n365, n130);
buf  g321 (n228, n134);
not  g322 (n190, n113);
buf  g323 (n408, n85);
not  g324 (n319, n89);
buf  g325 (n356, n78);
not  g326 (n212, n112);
buf  g327 (n391, n116);
not  g328 (n290, n114);
buf  g329 (n232, n110);
buf  g330 (n241, n66);
buf  g331 (n314, n115);
buf  g332 (n349, n92);
not  g333 (n233, n124);
buf  g334 (n388, n127);
not  g335 (n341, n138);
not  g336 (n201, n76);
buf  g337 (n324, n125);
not  g338 (n302, n89);
buf  g339 (n273, n136);
buf  g340 (n264, n75);
buf  g341 (n390, n93);
not  g342 (n366, n81);
buf  g343 (n191, n130);
not  g344 (n288, n80);
buf  g345 (n450, n128);
not  g346 (n231, n74);
not  g347 (n244, n76);
not  g348 (n363, n86);
buf  g349 (n405, n98);
buf  g350 (n271, n79);
not  g351 (n455, n111);
buf  g352 (n202, n70);
not  g353 (n284, n97);
buf  g354 (n253, n142);
not  g355 (n400, n82);
buf  g356 (n309, n123);
not  g357 (n458, n90);
not  g358 (n344, n123);
buf  g359 (n451, n102);
buf  g360 (n423, n68);
buf  g361 (n368, n134);
not  g362 (n214, n73);
buf  g363 (n337, n98);
not  g364 (n440, n125);
buf  g365 (n312, n126);
not  g366 (n328, n127);
not  g367 (n268, n131);
not  g368 (n325, n139);
not  g369 (n205, n101);
buf  g370 (n278, n142);
buf  g371 (n197, n107);
buf  g372 (n294, n123);
not  g373 (n189, n76);
not  g374 (n417, n83);
not  g375 (n426, n87);
buf  g376 (n409, n75);
not  g377 (n275, n145);
buf  g378 (n334, n101);
buf  g379 (n347, n79);
buf  g380 (n331, n111);
buf  g381 (n295, n104);
buf  g382 (n299, n106);
buf  g383 (n279, n100);
not  g384 (n327, n95);
not  g385 (n375, n78);
not  g386 (n225, n99);
not  g387 (n285, n102);
buf  g388 (n342, n114);
buf  g389 (n384, n80);
not  g390 (n436, n109);
not  g391 (n199, n68);
not  g392 (n259, n122);
buf  g393 (n292, n77);
not  g394 (n364, n77);
not  g395 (n315, n126);
not  g396 (n382, n118);
not  g397 (n281, n136);
buf  g398 (n389, n141);
not  g399 (n438, n105);
buf  g400 (n235, n144);
not  g401 (n208, n78);
buf  g402 (n430, n124);
not  g403 (n413, n67);
not  g404 (n221, n96);
not  g405 (n330, n133);
not  g406 (n215, n135);
buf  g407 (n428, n131);
not  g408 (n346, n79);
not  g409 (n379, n77);
buf  g410 (n422, n106);
not  g411 (n246, n110);
buf  g412 (n308, n131);
buf  g413 (n385, n135);
buf  g414 (n350, n127);
not  g415 (n343, n120);
not  g416 (n223, n104);
not  g417 (n371, n128);
buf  g418 (n216, n121);
or   g419 (n296, n127, n76, n90, n72);
xor  g420 (n339, n78, n144, n129, n120);
xor  g421 (n449, n115, n100, n106, n136);
nand g422 (n419, n113, n97, n110, n69);
and  g423 (n336, n98, n129, n118, n111);
and  g424 (n203, n108, n99, n107, n112);
xnor g425 (n358, n137, n75, n135, n145);
nor  g426 (n420, n81, n91, n120, n124);
or   g427 (n362, n143, n108, n142, n139);
nand g428 (n453, n143, n91, n98);
xor  g429 (n200, n110, n114, n103, n93);
not  g430 (n463, n190);
buf  g431 (n464, n191);
buf  g432 (n466, n463);
buf  g433 (n465, n463);
and  g434 (n472, n196, n147, n197);
xnor g435 (n473, n195, n149, n199, n146);
xnor g436 (n471, n146, n466, n148, n465);
or   g437 (n468, n201, n146, n465);
xor  g438 (n474, n466, n148, n147);
nand g439 (n470, n148, n200, n192, n466);
xor  g440 (n467, n193, n194, n465, n466);
xor  g441 (n469, n148, n149, n465, n198);
buf  g442 (n502, n468);
not  g443 (n475, n472);
buf  g444 (n499, n467);
buf  g445 (n500, n473);
not  g446 (n497, n474);
not  g447 (n504, n471);
buf  g448 (n484, n469);
not  g449 (n486, n468);
buf  g450 (n506, n473);
buf  g451 (n498, n470);
buf  g452 (n505, n467);
buf  g453 (n492, n471);
buf  g454 (n478, n472);
not  g455 (n479, n469);
buf  g456 (n477, n469);
buf  g457 (n487, n471);
not  g458 (n485, n472);
buf  g459 (n493, n473);
buf  g460 (n496, n468);
buf  g461 (n480, n474);
not  g462 (n489, n470);
buf  g463 (n491, n472);
not  g464 (n503, n469);
not  g465 (n483, n474);
not  g466 (n490, n467);
not  g467 (n476, n467);
not  g468 (n501, n470);
not  g469 (n495, n471);
not  g470 (n482, n468);
not  g471 (n481, n473);
not  g472 (n494, n470);
buf  g473 (n488, n474);
not  g474 (n554, n480);
not  g475 (n540, n495);
buf  g476 (n525, n490);
buf  g477 (n544, n494);
buf  g478 (n509, n495);
buf  g479 (n543, n491);
buf  g480 (n515, n487);
not  g481 (n570, n481);
not  g482 (n572, n492);
not  g483 (n580, n500);
buf  g484 (n533, n488);
not  g485 (n508, n499);
not  g486 (n581, n489);
not  g487 (n567, n475);
not  g488 (n552, n502);
not  g489 (n542, n479);
buf  g490 (n557, n499);
buf  g491 (n568, n493);
buf  g492 (n573, n494);
buf  g493 (n583, n498);
buf  g494 (n553, n502);
buf  g495 (n527, n486);
buf  g496 (n546, n500);
not  g497 (n561, n500);
buf  g498 (n551, n482);
not  g499 (n518, n497);
buf  g500 (n526, n484);
buf  g501 (n584, n485);
buf  g502 (n585, n484);
not  g503 (n510, n478);
not  g504 (n556, n488);
buf  g505 (n530, n496);
not  g506 (n535, n496);
buf  g507 (n507, n501);
buf  g508 (n531, n494);
not  g509 (n582, n498);
buf  g510 (n569, n501);
buf  g511 (n548, n483);
buf  g512 (n511, n493);
not  g513 (n576, n497);
not  g514 (n545, n497);
buf  g515 (n516, n497);
buf  g516 (n555, n487);
buf  g517 (n547, n475);
buf  g518 (n528, n485);
buf  g519 (n566, n499);
not  g520 (n522, n493);
buf  g521 (n550, n496);
not  g522 (n523, n498);
not  g523 (n562, n494);
buf  g524 (n560, n491);
not  g525 (n559, n486);
buf  g526 (n575, n492);
buf  g527 (n517, n491);
buf  g528 (n565, n491);
not  g529 (n524, n490);
not  g530 (n574, n495);
not  g531 (n532, n480);
buf  g532 (n578, n483);
not  g533 (n538, n479);
not  g534 (n586, n499);
buf  g535 (n512, n477);
buf  g536 (n564, n501);
not  g537 (n537, n500);
buf  g538 (n514, n476);
not  g539 (n519, n501);
buf  g540 (n571, n489);
not  g541 (n558, n498);
buf  g542 (n539, n490);
not  g543 (n579, n490);
buf  g544 (n521, n477);
buf  g545 (n534, n482);
buf  g546 (n549, n496);
not  g547 (n536, n481);
not  g548 (n541, n476);
not  g549 (n529, n478);
not  g550 (n520, n495);
buf  g551 (n513, n492);
buf  g552 (n577, n493);
buf  g553 (n563, n492);
not  g554 (n597, n513);
not  g555 (n610, n510);
buf  g556 (n601, n513);
not  g557 (n594, n509);
not  g558 (n609, n512);
not  g559 (n603, n507);
buf  g560 (n605, n509);
not  g561 (n589, n510);
buf  g562 (n592, n514);
not  g563 (n604, n508);
buf  g564 (n611, n513);
not  g565 (n593, n507);
buf  g566 (n599, n511);
not  g567 (n607, n507);
buf  g568 (n608, n512);
buf  g569 (n590, n514);
not  g570 (n595, n511);
not  g571 (n606, n512);
buf  g572 (n588, n510);
buf  g573 (n596, n514);
buf  g574 (n587, n511);
buf  g575 (n600, n508);
or   g576 (n598, n507, n509);
xor  g577 (n591, n513, n508, n514);
nor  g578 (n602, n510, n511, n509, n512);
xnor g579 (n626, n588, n15, n610);
or   g580 (n637, n609, n589, n18);
and  g581 (n614, n14, n12, n595);
or   g582 (n615, n9, n19, n21);
or   g583 (n628, n13, n590, n15);
xor  g584 (n632, n20, n9, n18);
nand g585 (n621, n603, n18, n12);
nor  g586 (n624, n600, n13, n611);
nor  g587 (n627, n605, n606, n14);
nand g588 (n635, n13, n9, n16);
or   g589 (n619, n21, n12, n20);
xor  g590 (n612, n14, n16, n17);
nand g591 (n623, n16, n602, n21);
xnor g592 (n630, n8, n10, n15);
nor  g593 (n634, n596, n12, n597);
or   g594 (n618, n598, n18, n593);
xnor g595 (n633, n609, n17, n9);
xor  g596 (n616, n19, n592, n11);
nor  g597 (n620, n14, n587, n604);
xnor g598 (n617, n16, n11);
nor  g599 (n625, n10, n611, n17);
nand g600 (n622, n11, n10);
nand g601 (n613, n608, n607, n17);
and  g602 (n629, n13, n591, n610);
and  g603 (n636, n601, n20, n594);
xor  g604 (n631, n15, n19, n599);
buf  g605 (n643, n522);
buf  g606 (n684, n550);
not  g607 (n708, n618);
buf  g608 (n674, n542);
not  g609 (n710, n520);
and  g610 (n660, n26, n544, n519, n554);
nor  g611 (n707, n515, n536, n631, n503);
or   g612 (n661, n503, n551, n636);
xnor g613 (n658, n519, n27, n560, n522);
nor  g614 (n687, n620, n546, n619, n615);
and  g615 (n666, n629, n550, n517, n529);
xnor g616 (n662, n530, n539, n634, n624);
xor  g617 (n655, n620, n534, n205, n537);
xor  g618 (n668, n615, n522, n627, n637);
xor  g619 (n688, n618, n526, n544, n635);
and  g620 (n725, n505, n636, n540, n522);
nand g621 (n716, n545, n532, n527);
nor  g622 (n648, n543, n619, n612, n553);
or   g623 (n673, n553, n634, n502, n627);
and  g624 (n719, n24, n621, n551, n561);
xor  g625 (n652, n547, n534, n562, n520);
and  g626 (n646, n614, n560, n622, n628);
or   g627 (n709, n25, n503, n22, n621);
xnor g628 (n715, n540, n626, n539, n549);
or   g629 (n657, n618, n519, n633, n553);
xor  g630 (n650, n534, n516, n530, n622);
xnor g631 (n703, n526, n615, n516, n559);
xor  g632 (n690, n26, n543, n539, n23);
and  g633 (n711, n627, n526, n558, n534);
xor  g634 (n689, n535, n533, n24);
nand g635 (n726, n612, n549, n558, n547);
xor  g636 (n691, n26, n525, n540);
or   g637 (n718, n517, n202, n633, n532);
nand g638 (n683, n553, n531, n622, n617);
xnor g639 (n685, n515, n554, n630, n632);
and  g640 (n677, n541, n24, n525, n518);
xor  g641 (n695, n535, n623, n556, n629);
xor  g642 (n638, n204, n538, n530, n556);
nor  g643 (n681, n631, n22, n555, n623);
xor  g644 (n705, n614, n525, n552, n632);
nand g645 (n675, n545, n521, n555, n619);
xor  g646 (n713, n517, n632, n519, n525);
xor  g647 (n671, n615, n537, n622, n506);
or   g648 (n639, n22, n503, n547, n633);
xnor g649 (n680, n541, n555, n21, n504);
and  g650 (n679, n551, n618, n528, n504);
nor  g651 (n697, n535, n635, n27, n557);
and  g652 (n698, n631, n557, n25, n613);
or   g653 (n712, n546, n515, n536, n614);
nand g654 (n669, n628, n533, n541, n613);
or   g655 (n682, n626, n531, n23, n518);
xnor g656 (n699, n203, n523, n504, n520);
nand g657 (n642, n554, n637, n625, n505);
xor  g658 (n656, n26, n561, n616, n549);
nand g659 (n692, n505, n558, n523, n625);
xor  g660 (n720, n531, n559, n527, n504);
nand g661 (n696, n544, n526, n548, n624);
or   g662 (n694, n558, n537, n532, n531);
nand g663 (n653, n556, n520, n27, n560);
and  g664 (n654, n523, n627, n517, n541);
nor  g665 (n723, n635, n552, n521, n557);
xnor g666 (n651, n559, n620, n530, n630);
nor  g667 (n659, n628, n632, n551, n626);
and  g668 (n701, n515, n560, n613, n554);
and  g669 (n706, n516, n634, n506, n617);
nor  g670 (n645, n614, n542, n538, n613);
xnor g671 (n641, n624, n617, n625, n549);
nand g672 (n704, n527, n550, n633, n529);
nand g673 (n672, n556, n521, n524, n542);
nor  g674 (n722, n529, n628, n626, n543);
xor  g675 (n647, n542, n637, n546, n544);
nor  g676 (n724, n612, n535, n624, n634);
and  g677 (n676, n548, n555, n621, n543);
or   g678 (n640, n518, n616, n506);
xor  g679 (n649, n616, n636, n502, n537);
xnor g680 (n717, n545, n529, n518, n562);
xor  g681 (n665, n516, n629, n623, n635);
xnor g682 (n686, n528, n25, n557, n539);
nand g683 (n721, n548, n548, n524, n532);
xor  g684 (n667, n552, n25, n612, n545);
nor  g685 (n700, n521, n561, n505, n552);
and  g686 (n678, n623, n617, n528, n538);
xor  g687 (n663, n23, n23, n620, n506);
nand g688 (n644, n625, n637, n528, n630);
and  g689 (n670, n547, n24, n550, n524);
xor  g690 (n664, n536, n559, n631, n629);
xor  g691 (n702, n619, n630, n533, n206);
nand g692 (n714, n524, n561, n538, n621);
and  g693 (n693, n523, n546, n536, n22);
not  g694 (n752, n652);
buf  g695 (n766, n179);
or   g696 (n764, n714, n643, n716, n221);
and  g697 (n777, n646, n183, n219, n564);
nor  g698 (n733, n173, n571, n149, n187);
or   g699 (n739, n151, n579, n155, n691);
nor  g700 (n744, n187, n581, n582, n573);
or   g701 (n798, n574, n572, n648, n693);
nand g702 (n793, n686, n583, n164);
nor  g703 (n768, n584, n668, n153, n657);
nor  g704 (n758, n723, n573, n162, n656);
nand g705 (n735, n567, n164, n681, n577);
nand g706 (n771, n162, n154, n661, n573);
or   g707 (n807, n564, n697, n692, n173);
nor  g708 (n815, n161, n159, n181, n180);
xnor g709 (n776, n570, n574, n176, n150);
nor  g710 (n727, n161, n678, n186, n212);
xnor g711 (n792, n694, n651, n575, n184);
nor  g712 (n789, n176, n169, n168);
or   g713 (n746, n568, n567, n170, n159);
nor  g714 (n791, n582, n169, n163, n181);
and  g715 (n809, n181, n572, n563, n578);
and  g716 (n782, n178, n165, n179, n183);
or   g717 (n737, n665, n168, n184, n707);
nand g718 (n743, n564, n169, n684, n719);
and  g719 (n800, n172, n161, n580, n177);
xnor g720 (n749, n208, n185, n577, n677);
xor  g721 (n738, n569, n573, n701, n562);
nor  g722 (n772, n674, n669, n171, n214);
xnor g723 (n781, n210, n175, n163, n577);
xor  g724 (n759, n169, n569, n584, n695);
and  g725 (n750, n152, n182, n172, n168);
and  g726 (n794, n569, n154, n185, n563);
nand g727 (n805, n164, n162, n181, n579);
xnor g728 (n761, n151, n578, n654, n175);
nor  g729 (n765, n163, n726, n722, n207);
xor  g730 (n799, n584, n645, n567, n581);
nand g731 (n757, n28, n151, n568, n27);
xor  g732 (n741, n670, n171, n155, n160);
and  g733 (n797, n690, n178, n700, n167);
and  g734 (n783, n566, n662, n562, n178);
and  g735 (n754, n698, n182, n174, n580);
xnor g736 (n773, n577, n564, n179, n463);
xnor g737 (n796, n176, n647, n655, n712);
xnor g738 (n779, n571, n166, n180, n704);
and  g739 (n748, n578, n213, n159);
and  g740 (n730, n574, n167, n566, n679);
or   g741 (n742, n570, n161, n571, n165);
xnor g742 (n767, n575, n158, n567, n150);
nor  g743 (n790, n580, n175, n582, n568);
xnor g744 (n745, n685, n152, n185, n184);
xor  g745 (n740, n725, n211, n177, n172);
or   g746 (n770, n565, n671, n157, n162);
nand g747 (n753, n724, n163, n170, n157);
xnor g748 (n810, n575, n154, n660, n572);
or   g749 (n780, n185, n582, n581, n153);
or   g750 (n762, n177, n166, n174, n157);
and  g751 (n804, n715, n720, n565, n170);
nor  g752 (n747, n160, n667, n570, n696);
xor  g753 (n731, n171, n150, n180, n676);
nand g754 (n786, n166, n644, n170, n569);
xnor g755 (n814, n566, n682, n718, n184);
or   g756 (n788, n689, n659, n180, n218);
nor  g757 (n736, n155, n176, n173, n642);
xor  g758 (n803, n699, n583, n179, n209);
xnor g759 (n801, n574, n156, n579, n167);
or   g760 (n806, n154, n702, n186, n653);
or   g761 (n778, n583, n708, n650, n666);
and  g762 (n811, n563, n165, n186, n153);
nor  g763 (n729, n706, n171, n158, n568);
nand g764 (n795, n153, n157, n710, n156);
nand g765 (n732, n673, n167, n182, n164);
and  g766 (n785, n158, n713, n658, n215);
or   g767 (n760, n580, n151, n177, n156);
and  g768 (n769, n217, n680, n641, n649);
or   g769 (n755, n703, n173, n672, n579);
and  g770 (n784, n174, n178, n576, n675);
nand g771 (n787, n220, n174, n571, n664);
and  g772 (n756, n687, n166, n663, n717);
nand g773 (n802, n575, n158, n705, n640);
xor  g774 (n774, n639, n576, n584, n638);
xnor g775 (n763, n565, n572, n152, n688);
nor  g776 (n751, n711, n152, n570, n563);
xor  g777 (n734, n576, n186, n172, n581);
nor  g778 (n813, n222, n565, n216, n160);
or   g779 (n775, n183, n709, n160, n156);
nand g780 (n808, n150, n576, n683, n149);
or   g781 (n728, n566, n183, n175, n165);
nor  g782 (n812, n721, n182, n155, n578);
not  g783 (n968, n434);
buf  g784 (n883, n737);
not  g785 (n1072, n771);
not  g786 (n1070, n766);
not  g787 (n919, n739);
buf  g788 (n928, n805);
buf  g789 (n1150, n745);
buf  g790 (n993, n350);
buf  g791 (n1047, n760);
not  g792 (n997, n765);
not  g793 (n895, n276);
buf  g794 (n1063, n397);
buf  g795 (n1033, n787);
not  g796 (n843, n731);
not  g797 (n1156, n774);
not  g798 (n956, n395);
not  g799 (n1034, n800);
buf  g800 (n835, n353);
not  g801 (n976, n305);
buf  g802 (n844, n420);
buf  g803 (n873, n396);
not  g804 (n1117, n403);
buf  g805 (n1028, n812);
not  g806 (n1018, n730);
buf  g807 (n1170, n746);
buf  g808 (n940, n386);
not  g809 (n1086, n738);
not  g810 (n1167, n752);
not  g811 (n861, n266);
not  g812 (n984, n811);
not  g813 (n1171, n273);
not  g814 (n995, n767);
not  g815 (n860, n777);
not  g816 (n897, n351);
buf  g817 (n1035, n813);
not  g818 (n1022, n287);
buf  g819 (n896, n734);
not  g820 (n890, n756);
not  g821 (n1134, n775);
buf  g822 (n948, n766);
buf  g823 (n1011, n807);
not  g824 (n977, n792);
buf  g825 (n937, n788);
buf  g826 (n961, n279);
not  g827 (n978, n763);
buf  g828 (n833, n762);
buf  g829 (n1073, n798);
buf  g830 (n899, n246);
buf  g831 (n971, n286);
not  g832 (n979, n257);
not  g833 (n945, n225);
buf  g834 (n885, n751);
not  g835 (n841, n442);
not  g836 (n1114, n363);
not  g837 (n1160, n732);
not  g838 (n982, n785);
not  g839 (n1030, n270);
buf  g840 (n1157, n763);
buf  g841 (n1082, n411);
not  g842 (n957, n759);
not  g843 (n966, n277);
not  g844 (n1109, n754);
buf  g845 (n1075, n740);
buf  g846 (n970, n727);
buf  g847 (n1040, n308);
not  g848 (n1162, n729);
not  g849 (n1087, n742);
not  g850 (n829, n756);
not  g851 (n1052, n388);
not  g852 (n1042, n318);
not  g853 (n1163, n771);
buf  g854 (n929, n789);
buf  g855 (n1068, n747);
not  g856 (n842, n748);
buf  g857 (n1020, n794);
buf  g858 (n973, n762);
buf  g859 (n852, n422);
buf  g860 (n1168, n373);
not  g861 (n974, n414);
buf  g862 (n1045, n416);
not  g863 (n1110, n783);
not  g864 (n1144, n746);
buf  g865 (n1085, n224);
not  g866 (n1126, n753);
not  g867 (n1107, n810);
not  g868 (n1000, n789);
not  g869 (n994, n773);
not  g870 (n851, n323);
not  g871 (n1089, n799);
buf  g872 (n969, n806);
not  g873 (n913, n809);
not  g874 (n869, n399);
not  g875 (n893, n242);
not  g876 (n942, n358);
not  g877 (n1146, n271);
buf  g878 (n1124, n755);
not  g879 (n1106, n333);
not  g880 (n891, n802);
buf  g881 (n820, n334);
buf  g882 (n911, n767);
not  g883 (n871, n437);
not  g884 (n906, n298);
not  g885 (n925, n743);
not  g886 (n1129, n766);
buf  g887 (n874, n325);
buf  g888 (n908, n243);
not  g889 (n838, n792);
not  g890 (n878, n247);
not  g891 (n858, n795);
buf  g892 (n1032, n762);
not  g893 (n923, n428);
buf  g894 (n1100, n789);
not  g895 (n1153, n736);
buf  g896 (n1002, n783);
not  g897 (n884, n274);
buf  g898 (n894, n387);
not  g899 (n1008, n744);
buf  g900 (n1001, n452);
not  g901 (n927, n359);
buf  g902 (n950, n750);
not  g903 (n1005, n757);
buf  g904 (n1061, n457);
buf  g905 (n1037, n776);
not  g906 (n931, n815);
buf  g907 (n830, n808);
not  g908 (n881, n784);
buf  g909 (n915, n748);
not  g910 (n868, n362);
buf  g911 (n826, n288);
buf  g912 (n1076, n779);
buf  g913 (n954, n187);
not  g914 (n932, n814);
not  g915 (n880, n790);
buf  g916 (n854, n430);
buf  g917 (n1029, n779);
buf  g918 (n1115, n311);
buf  g919 (n924, n769);
not  g920 (n1102, n393);
buf  g921 (n817, n253);
not  g922 (n1025, n417);
buf  g923 (n962, n354);
not  g924 (n1083, n309);
buf  g925 (n967, n728);
buf  g926 (n889, n407);
not  g927 (n920, n275);
buf  g928 (n1128, n753);
not  g929 (n863, n809);
buf  g930 (n986, n438);
buf  g931 (n898, n774);
not  g932 (n1069, n773);
not  g933 (n917, n789);
not  g934 (n1161, n295);
buf  g935 (n1125, n749);
not  g936 (n902, n767);
not  g937 (n1139, n775);
not  g938 (n845, n808);
not  g939 (n823, n729);
buf  g940 (n825, n239);
buf  g941 (n1036, n733);
buf  g942 (n990, n801);
not  g943 (n1155, n444);
buf  g944 (n1026, n806);
not  g945 (n938, n777);
not  g946 (n903, n813);
not  g947 (n1059, n365);
buf  g948 (n1053, n458);
buf  g949 (n939, n749);
buf  g950 (n850, n740);
buf  g951 (n828, n801);
buf  g952 (n946, n813);
buf  g953 (n1006, n733);
not  g954 (n1014, n327);
not  g955 (n1027, n228);
not  g956 (n1154, n302);
not  g957 (n992, n357);
not  g958 (n934, n262);
not  g959 (n892, n433);
not  g960 (n1091, n238);
buf  g961 (n963, n815);
buf  g962 (n1080, n368);
not  g963 (n1148, n223);
buf  g964 (n1130, n742);
buf  g965 (n1054, n768);
not  g966 (n983, n264);
not  g967 (n1031, n361);
buf  g968 (n955, n267);
buf  g969 (n933, n745);
not  g970 (n916, n782);
not  g971 (n901, n421);
buf  g972 (n910, n797);
not  g973 (n1133, n756);
not  g974 (n1169, n745);
not  g975 (n1140, n797);
not  g976 (n1090, n750);
buf  g977 (n996, n788);
not  g978 (n943, n765);
not  g979 (n853, n784);
buf  g980 (n1145, n376);
not  g981 (n988, n370);
buf  g982 (n1015, n381);
buf  g983 (n909, n347);
not  g984 (n1108, n377);
not  g985 (n1112, n768);
buf  g986 (n914, n296);
not  g987 (n947, n303);
not  g988 (n949, n764);
buf  g989 (n1098, n808);
buf  g990 (n1019, n432);
not  g991 (n1079, n380);
not  g992 (n855, n746);
not  g993 (n1135, n449);
not  g994 (n876, n348);
buf  g995 (n1119, n800);
buf  g996 (n1164, n418);
not  g997 (n1009, n797);
buf  g998 (n875, n794);
not  g999 (n827, n787);
not  g1000 (n1152, n770);
not  g1001 (n824, n811);
buf  g1002 (n1159, n383);
not  g1003 (n821, n774);
not  g1004 (n1105, n360);
buf  g1005 (n859, n291);
not  g1006 (n872, n732);
buf  g1007 (n1151, n769);
buf  g1008 (n818, n391);
not  g1009 (n1055, n810);
buf  g1010 (n1007, n743);
buf  g1011 (n964, n752);
not  g1012 (n921, n783);
buf  g1013 (n951, n755);
buf  g1014 (n1111, n366);
buf  g1015 (n972, n772);
not  g1016 (n1081, n235);
buf  g1017 (n864, n788);
buf  g1018 (n1060, n807);
not  g1019 (n1038, n342);
not  g1020 (n1127, n278);
not  g1021 (n936, n364);
buf  g1022 (n1048, n815);
not  g1023 (n1113, n770);
not  g1024 (n877, n772);
not  g1025 (n1013, n413);
not  g1026 (n867, n730);
buf  g1027 (n987, n751);
not  g1028 (n819, n328);
not  g1029 (n1149, n769);
buf  g1030 (n1067, n814);
buf  g1031 (n905, n423);
not  g1032 (n912, n732);
buf  g1033 (n989, n758);
buf  g1034 (n1093, n250);
not  g1035 (n839, n745);
not  g1036 (n840, n453);
not  g1037 (n952, n769);
not  g1038 (n1121, n755);
not  g1039 (n1123, n780);
not  g1040 (n1136, n321);
buf  g1041 (n1141, n786);
not  g1042 (n1021, n340);
buf  g1043 (n882, n258);
not  g1044 (n900, n747);
buf  g1045 (n1003, n390);
not  g1046 (n1137, n750);
buf  g1047 (n1074, n795);
buf  g1048 (n1065, n245);
buf  g1049 (n886, n229);
not  g1050 (n1039, n812);
buf  g1051 (n1120, n800);
not  g1052 (n980, n424);
buf  g1053 (n1101, n254);
not  g1054 (n998, n790);
not  g1055 (n1046, n284);
buf  g1056 (n1024, n252);
buf  g1057 (n1064, n734);
buf  g1058 (n862, n759);
and  g1059 (n837, n736, n792, n226, n728);
and  g1060 (n1057, n796, n796, n811, n777);
nor  g1061 (n1132, n748, n806, n742, n256);
nor  g1062 (n1088, n760, n751, n346, n289);
or   g1063 (n1094, n294, n753, n349, n802);
xor  g1064 (n1077, n731, n759, n737, n799);
and  g1065 (n1058, n255, n297, n332, n241);
or   g1066 (n1084, n763, n408, n793, n371);
or   g1067 (n1010, n786, n410, n272, n757);
xnor g1068 (n816, n727, n741, n744, n767);
xnor g1069 (n941, n419, n784, n736, n809);
xor  g1070 (n822, n251, n799, n236, n315);
or   g1071 (n1049, n791, n771, n441, n777);
nand g1072 (n865, n743, n740, n782, n356);
xor  g1073 (n1017, n234, n281, n394, n728);
or   g1074 (n1078, n259, n733, n770, n268);
or   g1075 (n922, n282, n743, n805, n324);
nand g1076 (n1016, n230, n786, n379, n764);
nor  g1077 (n1043, n747, n233, n730, n459);
or   g1078 (n981, n748, n436, n759, n765);
and  g1079 (n959, n802, n260, n741, n456);
xnor g1080 (n991, n780, n447, n446, n760);
or   g1081 (n1142, n392, n404, n736, n415);
nor  g1082 (n856, n749, n754, n797, n738);
nor  g1083 (n846, n727, n448, n755, n738);
xnor g1084 (n832, n782, n402, n739, n409);
and  g1085 (n1096, n772, n461, n785, n312);
xor  g1086 (n1138, n778, n780, n766, n269);
xor  g1087 (n907, n283, n426, n773, n369);
or   g1088 (n1131, n398, n310, n293, n319);
nand g1089 (n1050, n747, n749, n740, n753);
nand g1090 (n960, n385, n792, n355, n746);
nor  g1091 (n975, n778, n778, n754, n786);
xor  g1092 (n1118, n804, n344, n781);
nand g1093 (n1023, n782, n770, n375, n738);
xnor g1094 (n1071, n730, n809, n227, n244);
nand g1095 (n836, n737, n343, n799, n800);
and  g1096 (n918, n768, n313, n735, n378);
or   g1097 (n1004, n729, n773, n761, n460);
xor  g1098 (n958, n806, n815, n752, n248);
or   g1099 (n953, n427, n451, n454, n787);
xnor g1100 (n888, n322, n337, n790, n807);
or   g1101 (n831, n261, n320, n431, n285);
and  g1102 (n1092, n741, n810, n733, n808);
xor  g1103 (n904, n231, n791, n317, n754);
xor  g1104 (n847, n812, n425, n793, n795);
nand g1105 (n1147, n801, n739, n775, n735);
xor  g1106 (n1056, n791, n443, n810, n734);
xnor g1107 (n1103, n793, n445, n304, n300);
xnor g1108 (n887, n783, n751, n781, n455);
or   g1109 (n999, n729, n341, n280, n450);
and  g1110 (n849, n793, n232, n301, n237);
nor  g1111 (n1051, n316, n339, n771, n335);
xor  g1112 (n1012, n263, n814, n734, n741);
and  g1113 (n1062, n803, n744, n805, n768);
xor  g1114 (n965, n727, n763, n435, n735);
xnor g1115 (n930, n801, n249, n779, n401);
nor  g1116 (n879, n798, n802, n731, n336);
and  g1117 (n1097, n814, n776, n764, n372);
nor  g1118 (n1066, n440, n400, n778, n412);
or   g1119 (n1044, n761, n757, n811, n804);
xor  g1120 (n857, n299, n405, n240, n787);
xnor g1121 (n1104, n758, n804, n739, n757);
nand g1122 (n834, n774, n314, n790, n796);
or   g1123 (n1122, n794, n775, n785, n731);
xnor g1124 (n944, n784, n744, n798, n804);
and  g1125 (n848, n788, n389, n290, n756);
xor  g1126 (n1116, n791, n374, n429, n781);
or   g1127 (n1166, n785, n779, n742, n764);
xnor g1128 (n1143, n807, n367, n326, n331);
nor  g1129 (n935, n795, n338, n439, n758);
xnor g1130 (n1041, n758, n803, n406, n728);
nor  g1131 (n1158, n794, n803, n765, n780);
or   g1132 (n1165, n735, n384, n812, n776);
nor  g1133 (n870, n776, n382, n307, n752);
xnor g1134 (n1099, n329, n306, n762, n761);
or   g1135 (n866, n732, n737, n813, n798);
or   g1136 (n926, n760, n796, n352, n330);
or   g1137 (n1095, n803, n761, n805, n772);
xor  g1138 (n985, n265, n345, n750, n292);
not  g1139 (n1286, n907);
buf  g1140 (n1503, n1039);
buf  g1141 (n1618, n894);
not  g1142 (n1273, n831);
not  g1143 (n1421, n1136);
buf  g1144 (n1485, n1137);
not  g1145 (n1379, n1154);
not  g1146 (n1585, n1023);
not  g1147 (n1393, n1117);
not  g1148 (n1529, n1030);
buf  g1149 (n1659, n826);
not  g1150 (n1638, n1133);
buf  g1151 (n1268, n1035);
buf  g1152 (n1472, n902);
not  g1153 (n1470, n1086);
not  g1154 (n1207, n920);
not  g1155 (n1471, n1143);
buf  g1156 (n1222, n828);
buf  g1157 (n1604, n1029);
buf  g1158 (n1623, n906);
not  g1159 (n1336, n1103);
not  g1160 (n1329, n1077);
buf  g1161 (n1189, n1040);
buf  g1162 (n1647, n1066);
not  g1163 (n1317, n931);
not  g1164 (n1526, n1045);
not  g1165 (n1246, n1020);
not  g1166 (n1458, n1078);
buf  g1167 (n1274, n1113);
buf  g1168 (n1360, n1125);
not  g1169 (n1621, n1116);
buf  g1170 (n1474, n916);
buf  g1171 (n1247, n1123);
buf  g1172 (n1523, n911);
buf  g1173 (n1282, n1079);
not  g1174 (n1501, n1094);
buf  g1175 (n1365, n1049);
not  g1176 (n1578, n1168);
buf  g1177 (n1496, n1106);
buf  g1178 (n1567, n891);
buf  g1179 (n1557, n936);
buf  g1180 (n1257, n1041);
not  g1181 (n1518, n1148);
not  g1182 (n1413, n1004);
not  g1183 (n1616, n1171);
not  g1184 (n1548, n1133);
buf  g1185 (n1363, n1076);
not  g1186 (n1284, n1034);
not  g1187 (n1522, n860);
buf  g1188 (n1271, n839);
not  g1189 (n1532, n1058);
buf  g1190 (n1549, n1018);
buf  g1191 (n1198, n1072);
not  g1192 (n1188, n1038);
not  g1193 (n1303, n912);
buf  g1194 (n1179, n1168);
buf  g1195 (n1375, n1079);
not  g1196 (n1491, n1135);
not  g1197 (n1627, n1139);
buf  g1198 (n1202, n841);
buf  g1199 (n1452, n1080);
not  g1200 (n1617, n1016);
not  g1201 (n1597, n1124);
not  g1202 (n1519, n1060);
buf  g1203 (n1172, n1156);
not  g1204 (n1255, n1092);
not  g1205 (n1646, n942);
buf  g1206 (n1244, n1009);
buf  g1207 (n1592, n1161);
not  g1208 (n1463, n932);
buf  g1209 (n1542, n1043);
not  g1210 (n1309, n977);
not  g1211 (n1220, n926);
buf  g1212 (n1252, n871);
buf  g1213 (n1278, n934);
not  g1214 (n1376, n1150);
buf  g1215 (n1226, n1043);
buf  g1216 (n1346, n884);
not  g1217 (n1505, n988);
not  g1218 (n1615, n1151);
buf  g1219 (n1568, n1089);
buf  g1220 (n1287, n1063);
buf  g1221 (n1174, n1031);
buf  g1222 (n1398, n944);
not  g1223 (n1381, n991);
not  g1224 (n1429, n1081);
buf  g1225 (n1599, n824);
not  g1226 (n1575, n1166);
buf  g1227 (n1298, n1115);
buf  g1228 (n1353, n1088);
buf  g1229 (n1404, n1091);
buf  g1230 (n1301, n896);
buf  g1231 (n1279, n1051);
not  g1232 (n1307, n1052);
buf  g1233 (n1342, n827);
buf  g1234 (n1552, n917);
not  g1235 (n1612, n1134);
buf  g1236 (n1224, n1067);
buf  g1237 (n1639, n833);
not  g1238 (n1308, n1170);
buf  g1239 (n1643, n1116);
not  g1240 (n1281, n873);
buf  g1241 (n1658, n1167);
not  g1242 (n1311, n921);
not  g1243 (n1570, n1128);
not  g1244 (n1626, n1107);
buf  g1245 (n1454, n1071);
buf  g1246 (n1267, n967);
not  g1247 (n1242, n990);
buf  g1248 (n1664, n999);
buf  g1249 (n1359, n1061);
buf  g1250 (n1277, n866);
buf  g1251 (n1283, n835);
not  g1252 (n1370, n850);
not  g1253 (n1300, n1041);
buf  g1254 (n1602, n1010);
buf  g1255 (n1504, n930);
not  g1256 (n1251, n998);
not  g1257 (n1637, n1144);
buf  g1258 (n1324, n1064);
buf  g1259 (n1494, n1120);
not  g1260 (n1187, n1073);
not  g1261 (n1591, n957);
buf  g1262 (n1193, n970);
not  g1263 (n1673, n1047);
buf  g1264 (n1608, n1107);
buf  g1265 (n1313, n848);
buf  g1266 (n1624, n885);
not  g1267 (n1206, n1165);
not  g1268 (n1347, n1132);
not  g1269 (n1354, n1059);
not  g1270 (n1559, n1027);
not  g1271 (n1444, n1021);
not  g1272 (n1337, n1132);
buf  g1273 (n1331, n876);
not  g1274 (n1322, n847);
not  g1275 (n1306, n980);
not  g1276 (n1446, n929);
buf  g1277 (n1562, n1120);
not  g1278 (n1475, n1115);
not  g1279 (n1478, n1103);
buf  g1280 (n1237, n1024);
not  g1281 (n1424, n925);
buf  g1282 (n1304, n1129);
buf  g1283 (n1601, n1012);
not  g1284 (n1340, n845);
buf  g1285 (n1669, n1017);
buf  g1286 (n1565, n822);
buf  g1287 (n1238, n953);
not  g1288 (n1450, n1050);
not  g1289 (n1225, n898);
not  g1290 (n1356, n1036);
not  g1291 (n1316, n955);
buf  g1292 (n1514, n1137);
buf  g1293 (n1600, n1126);
buf  g1294 (n1479, n895);
buf  g1295 (n1590, n1162);
buf  g1296 (n1531, n837);
not  g1297 (n1345, n846);
buf  g1298 (n1293, n986);
buf  g1299 (n1481, n1150);
buf  g1300 (n1477, n1117);
not  g1301 (n1333, n886);
buf  g1302 (n1455, n1076);
buf  g1303 (n1314, n1139);
buf  g1304 (n1556, n820);
not  g1305 (n1199, n968);
not  g1306 (n1577, n1084);
buf  g1307 (n1217, n1138);
buf  g1308 (n1480, n1052);
buf  g1309 (n1425, n836);
not  g1310 (n1372, n825);
not  g1311 (n1482, n1068);
not  g1312 (n1405, n1002);
buf  g1313 (n1439, n961);
not  g1314 (n1266, n1037);
not  g1315 (n1371, n1031);
buf  g1316 (n1358, n1011);
buf  g1317 (n1228, n888);
not  g1318 (n1332, n950);
not  g1319 (n1384, n1071);
not  g1320 (n1232, n1087);
buf  g1321 (n1418, n995);
buf  g1322 (n1441, n1077);
not  g1323 (n1310, n1065);
not  g1324 (n1230, n868);
not  g1325 (n1392, n834);
buf  g1326 (n1364, n1040);
not  g1327 (n1609, n1085);
buf  g1328 (n1185, n913);
buf  g1329 (n1513, n1044);
buf  g1330 (n1334, n1099);
buf  g1331 (n1541, n1006);
not  g1332 (n1436, n877);
buf  g1333 (n1516, n1140);
not  g1334 (n1588, n857);
buf  g1335 (n1652, n1163);
not  g1336 (n1536, n1061);
not  g1337 (n1668, n865);
buf  g1338 (n1319, n1053);
buf  g1339 (n1378, n1109);
not  g1340 (n1512, n987);
buf  g1341 (n1305, n994);
not  g1342 (n1263, n1159);
not  g1343 (n1506, n1166);
buf  g1344 (n1390, n1149);
buf  g1345 (n1180, n946);
not  g1346 (n1666, n948);
not  g1347 (n1335, n1089);
not  g1348 (n1241, n849);
not  g1349 (n1619, n1083);
buf  g1350 (n1366, n1102);
not  g1351 (n1216, n855);
not  g1352 (n1665, n1057);
buf  g1353 (n1177, n973);
buf  g1354 (n1456, n1066);
buf  g1355 (n1508, n874);
not  g1356 (n1628, n949);
buf  g1357 (n1318, n1149);
not  g1358 (n1605, n962);
not  g1359 (n1606, n1112);
not  g1360 (n1396, n993);
buf  g1361 (n1330, n1090);
not  g1362 (n1640, n1112);
not  g1363 (n1598, n851);
buf  g1364 (n1248, n919);
buf  g1365 (n1631, n1088);
buf  g1366 (n1211, n1141);
buf  g1367 (n1397, n1068);
not  g1368 (n1419, n1095);
not  g1369 (n1476, n1171);
not  g1370 (n1484, n1074);
buf  g1371 (n1417, n960);
not  g1372 (n1649, n1145);
not  g1373 (n1488, n1058);
not  g1374 (n1321, n1055);
not  g1375 (n1576, n1160);
buf  g1376 (n1620, n889);
buf  g1377 (n1595, n933);
buf  g1378 (n1380, n963);
not  g1379 (n1383, n1145);
not  g1380 (n1409, n1032);
not  g1381 (n1195, n1148);
not  g1382 (n1462, n1063);
not  g1383 (n1483, n952);
buf  g1384 (n1350, n887);
buf  g1385 (n1593, n1001);
not  g1386 (n1495, n1101);
not  g1387 (n1447, n1160);
buf  g1388 (n1219, n1037);
buf  g1389 (n1490, n1169);
buf  g1390 (n1227, n829);
not  g1391 (n1655, n818);
buf  g1392 (n1367, n924);
buf  g1393 (n1190, n1104);
not  g1394 (n1539, n1026);
buf  g1395 (n1420, n1158);
buf  g1396 (n1465, n976);
buf  g1397 (n1569, n1057);
not  g1398 (n1415, n1070);
not  g1399 (n1181, n943);
not  g1400 (n1401, n1080);
not  g1401 (n1325, n947);
buf  g1402 (n1389, n1081);
not  g1403 (n1622, n1155);
buf  g1404 (n1412, n1114);
buf  g1405 (n1551, n821);
not  g1406 (n1355, n941);
buf  g1407 (n1408, n1073);
not  g1408 (n1660, n1101);
not  g1409 (n1427, n1140);
not  g1410 (n1486, n863);
buf  g1411 (n1528, n974);
buf  g1412 (n1262, n1108);
not  g1413 (n1521, n992);
not  g1414 (n1373, n890);
buf  g1415 (n1594, n1157);
buf  g1416 (n1250, n1067);
not  g1417 (n1579, n817);
buf  g1418 (n1611, n856);
not  g1419 (n1445, n1054);
not  g1420 (n1391, n1062);
buf  g1421 (n1289, n989);
buf  g1422 (n1201, n1059);
buf  g1423 (n1416, n1122);
buf  g1424 (n1527, n1097);
buf  g1425 (n1582, n1056);
not  g1426 (n1341, n1126);
not  g1427 (n1186, n1015);
not  g1428 (n1657, n1095);
not  g1429 (n1492, n838);
not  g1430 (n1196, n1106);
buf  g1431 (n1525, n893);
buf  g1432 (n1610, n1144);
not  g1433 (n1603, n1054);
not  g1434 (n1269, n1099);
buf  g1435 (n1339, n1042);
buf  g1436 (n1629, n1119);
not  g1437 (n1435, n853);
not  g1438 (n1614, n959);
buf  g1439 (n1368, n1086);
buf  g1440 (n1630, n1128);
not  g1441 (n1498, n914);
not  g1442 (n1208, n1028);
not  g1443 (n1641, n1046);
not  g1444 (n1254, n909);
buf  g1445 (n1328, n1027);
not  g1446 (n1583, n1154);
not  g1447 (n1607, n903);
not  g1448 (n1651, n1049);
not  g1449 (n1218, n1093);
buf  g1450 (n1402, n1124);
not  g1451 (n1497, n1094);
not  g1452 (n1352, n966);
buf  g1453 (n1385, n1029);
not  g1454 (n1349, n975);
buf  g1455 (n1547, n1030);
not  g1456 (n1449, n1108);
not  g1457 (n1534, n852);
not  g1458 (n1432, n1131);
not  g1459 (n1502, n938);
not  g1460 (n1587, n901);
not  g1461 (n1538, n1110);
buf  g1462 (n1428, n854);
buf  g1463 (n1302, n1069);
buf  g1464 (n1410, n861);
buf  g1465 (n1291, n819);
buf  g1466 (n1361, n1075);
buf  g1467 (n1635, n1036);
buf  g1468 (n1414, n1127);
not  g1469 (n1369, n870);
buf  g1470 (n1192, n1048);
buf  g1471 (n1288, n1125);
buf  g1472 (n1558, n1046);
buf  g1473 (n1191, n1102);
buf  g1474 (n1400, n1096);
not  g1475 (n1243, n981);
not  g1476 (n1440, n844);
not  g1477 (n1468, n1135);
not  g1478 (n1442, n927);
buf  g1479 (n1434, n1118);
buf  g1480 (n1586, n1118);
buf  g1481 (n1249, n1113);
buf  g1482 (n1550, n1045);
not  g1483 (n1466, n1152);
buf  g1484 (n1203, n985);
buf  g1485 (n1221, n937);
not  g1486 (n1553, n1060);
not  g1487 (n1662, n1114);
not  g1488 (n1265, n1162);
not  g1489 (n1320, n1093);
not  g1490 (n1377, n965);
buf  g1491 (n1560, n869);
buf  g1492 (n1357, n1051);
not  g1493 (n1580, n859);
buf  g1494 (n1403, n1152);
not  g1495 (n1642, n1130);
buf  g1496 (n1259, n881);
buf  g1497 (n1633, n883);
buf  g1498 (n1387, n1070);
not  g1499 (n1566, n1111);
not  g1500 (n1178, n997);
not  g1501 (n1343, n1033);
not  g1502 (n1295, n1164);
buf  g1503 (n1323, n983);
not  g1504 (n1215, n1127);
buf  g1505 (n1173, n1083);
buf  g1506 (n1285, n1098);
buf  g1507 (n1453, n1169);
buf  g1508 (n1233, n958);
not  g1509 (n1194, n1005);
buf  g1510 (n1411, n875);
not  g1511 (n1388, n1129);
buf  g1512 (n1183, n935);
buf  g1513 (n1275, n1141);
buf  g1514 (n1636, n1082);
buf  g1515 (n1648, n972);
not  g1516 (n1571, n1003);
buf  g1517 (n1229, n956);
buf  g1518 (n1197, n922);
buf  g1519 (n1280, n1121);
not  g1520 (n1489, n1019);
not  g1521 (n1399, n1084);
buf  g1522 (n1661, n882);
buf  g1523 (n1653, n1121);
buf  g1524 (n1511, n979);
not  g1525 (n1625, n1164);
not  g1526 (n1184, n1014);
buf  g1527 (n1214, n897);
not  g1528 (n1239, n1111);
buf  g1529 (n1382, n867);
not  g1530 (n1543, n1143);
not  g1531 (n1299, n996);
buf  g1532 (n1656, n1050);
not  g1533 (n1563, n858);
buf  g1534 (n1672, n1092);
not  g1535 (n1423, n1082);
not  g1536 (n1264, n1136);
not  g1537 (n1644, n915);
buf  g1538 (n1327, n1074);
buf  g1539 (n1223, n1170);
buf  g1540 (n1584, n969);
not  g1541 (n1546, n823);
buf  g1542 (n1394, n1134);
buf  g1543 (n1431, n1034);
buf  g1544 (n1589, n1053);
buf  g1545 (n1312, n1069);
buf  g1546 (n1407, n1157);
buf  g1547 (n1437, n1085);
not  g1548 (n1362, n918);
not  g1549 (n1537, n1096);
buf  g1550 (n1294, n1109);
buf  g1551 (n1573, n978);
not  g1552 (n1175, n1158);
buf  g1553 (n1270, n1042);
not  g1554 (n1469, n1038);
buf  g1555 (n1272, n1091);
buf  g1556 (n1344, n864);
buf  g1557 (n1438, n879);
not  g1558 (n1260, n832);
not  g1559 (n1245, n971);
buf  g1560 (n1240, n1147);
buf  g1561 (n1654, n1104);
buf  g1562 (n1451, n880);
buf  g1563 (n1460, n964);
buf  g1564 (n1395, n984);
buf  g1565 (n1524, n892);
buf  g1566 (n1200, n1155);
buf  g1567 (n1459, n1007);
not  g1568 (n1315, n1142);
not  g1569 (n1457, n1039);
buf  g1570 (n1574, n954);
buf  g1571 (n1448, n940);
not  g1572 (n1540, n1048);
buf  g1573 (n1426, n1100);
not  g1574 (n1493, n1098);
not  g1575 (n1236, n923);
not  g1576 (n1234, n1156);
buf  g1577 (n1499, n1100);
not  g1578 (n1205, n1131);
not  g1579 (n1670, n1047);
buf  g1580 (n1613, n840);
not  g1581 (n1555, n908);
buf  g1582 (n1671, n939);
buf  g1583 (n1374, n1055);
buf  g1584 (n1209, n905);
buf  g1585 (n1430, n816);
not  g1586 (n1533, n1146);
not  g1587 (n1253, n1153);
buf  g1588 (n1487, n1025);
not  g1589 (n1663, n1013);
buf  g1590 (n1564, n1161);
buf  g1591 (n1596, n1110);
buf  g1592 (n1296, n1044);
buf  g1593 (n1338, n1138);
not  g1594 (n1348, n904);
buf  g1595 (n1210, n1123);
not  g1596 (n1473, n1151);
buf  g1597 (n1464, n928);
not  g1598 (n1182, n1026);
buf  g1599 (n1422, n1147);
buf  g1600 (n1500, n951);
buf  g1601 (n1461, n1159);
buf  g1602 (n1520, n842);
not  g1603 (n1545, n1078);
not  g1604 (n1572, n1032);
buf  g1605 (n1667, n1105);
buf  g1606 (n1645, n945);
not  g1607 (n1554, n862);
buf  g1608 (n1212, n899);
buf  g1609 (n1326, n1033);
buf  g1610 (n1443, n1072);
not  g1611 (n1581, n1022);
not  g1612 (n1213, n1000);
not  g1613 (n1386, n1035);
buf  g1614 (n1515, n843);
not  g1615 (n1510, n1064);
buf  g1616 (n1634, n910);
not  g1617 (n1176, n900);
buf  g1618 (n1406, n1167);
buf  g1619 (n1517, n1056);
buf  g1620 (n1258, n1075);
not  g1621 (n1231, n1008);
not  g1622 (n1235, n1163);
not  g1623 (n1351, n830);
not  g1624 (n1433, n1097);
not  g1625 (n1297, n982);
buf  g1626 (n1507, n1146);
buf  g1627 (n1256, n1119);
buf  g1628 (n1530, n1153);
not  g1629 (n1467, n1105);
buf  g1630 (n1509, n1065);
not  g1631 (n1204, n1130);
buf  g1632 (n1261, n1090);
buf  g1633 (n1544, n872);
buf  g1634 (n1650, n1142);
not  g1635 (n1632, n1062);
not  g1636 (n1561, n878);
buf  g1637 (n1276, n1028);
buf  g1638 (n1292, n1165);
not  g1639 (n1290, n1122);
buf  g1640 (n1535, n1087);
nor  g1641 (n1677, n1398, n1409, n1294, n1474);
nor  g1642 (n1854, n1202, n1595, n1230, n1626);
nor  g1643 (n1842, n1422, n1588, n1223, n1416);
nand g1644 (n1704, n1489, n1513, n1586, n1269);
or   g1645 (n1817, n1600, n1566, n1370, n1380);
nand g1646 (n1691, n1544, n1614, n1343, n1438);
xor  g1647 (n1818, n1606, n1514, n1497, n1596);
nor  g1648 (n1870, n1197, n1356, n1535, n1522);
xnor g1649 (n1770, n1330, n1569, n1289, n1409);
xnor g1650 (n1744, n1280, n1620, n1609, n1361);
nand g1651 (n1789, n1438, n1437, n1450, n1441);
and  g1652 (n1695, n1315, n1598, n1282, n1571);
or   g1653 (n1684, n1564, n1637, n1546, n1658);
xnor g1654 (n1805, n1417, n1576, n1428, n1559);
xor  g1655 (n1719, n1609, n1218, n1423, n1413);
and  g1656 (n1776, n1242, n1569, n1511, n1365);
or   g1657 (n1835, n1321, n1424, n1556, n1439);
nand g1658 (n1778, n1462, n1248, n1314, n1596);
xnor g1659 (n1806, n1585, n1394, n1436, n1526);
xor  g1660 (n1767, n1500, n1412, n1496, n1532);
xor  g1661 (n1836, n1564, n1404, n1493, n1542);
or   g1662 (n1846, n1515, n1599, n1204, n1527);
nand g1663 (n1742, n1369, n1581, n1465, n1429);
xnor g1664 (n1780, n1300, n1620, n1544, n1262);
nand g1665 (n1774, n1504, n1619, n1554, n1580);
nor  g1666 (n1861, n1534, n1452, n1236, n1389);
or   g1667 (n1699, n1509, n1471, n1489, n1541);
nor  g1668 (n1698, n1408, n1307, n1418, n1622);
xor  g1669 (n1843, n1196, n1344, n1348, n1266);
nand g1670 (n1771, n1427, n1618, n1577, n1368);
nor  g1671 (n1703, n1459, n1572, n1469, n1542);
nor  g1672 (n1718, n1525, n1540, n1408, n1422);
nor  g1673 (n1812, n1519, n1578, n1527, n1385);
nand g1674 (n1823, n1502, n1250, n1648, n1442);
and  g1675 (n1850, n1624, n1478, n1464, n1310);
xor  g1676 (n1747, n1411, n1507, n1560, n1547);
xor  g1677 (n1856, n1557, n1403, n1421, n1374);
nand g1678 (n1860, n1622, n1377, n1407, n1225);
xor  g1679 (n1775, n1256, n1653, n1481, n1425);
and  g1680 (n1735, n1654, n1529, n1631, n1499);
xnor g1681 (n1696, n1551, n1229, n1311, n1451);
nand g1682 (n1867, n1393, n1497, n1653, n1611);
xnor g1683 (n1755, n1550, n1377, n1477, n1479);
or   g1684 (n1847, n1574, n1610, n1652, n1659);
nor  g1685 (n1757, n1484, n1194, n1526, n1341);
xor  g1686 (n1716, n1440, n1301, n1628, n1444);
xnor g1687 (n1680, n1274, n1369, n1507, n1367);
and  g1688 (n1788, n1434, n1372, n1447, n1486);
nor  g1689 (n1781, n1320, n1513, n1428, n1302);
nor  g1690 (n1688, n1543, n1492, n1603, n1491);
nand g1691 (n1868, n1536, n1582, n1512, n1378);
or   g1692 (n1733, n1498, n1456, n1460, n1657);
and  g1693 (n1740, n1191, n1483, n1656, n1530);
or   g1694 (n1853, n1657, n1305, n1432, n1570);
and  g1695 (n1844, n1516, n1205, n1410);
xnor g1696 (n1675, n1487, n1543, n1354, n1187);
nand g1697 (n1804, n1501, n1648, n1328, n1630);
and  g1698 (n1679, n1453, n1538, n1560, n1433);
nor  g1699 (n1833, n1381, n1611, n1563);
or   g1700 (n1756, n1382, n1480, n1455, n1641);
or   g1701 (n1808, n1641, n1602, n1627, n1589);
xor  g1702 (n1768, n1368, n1631, n1467, n1608);
xnor g1703 (n1749, n1234, n1439, n1172, n1184);
and  g1704 (n1827, n1637, n1376, n1257, n1617);
or   g1705 (n1798, n1576, n1415, n1414, n1495);
xor  g1706 (n1869, n1496, n1470, n1258, n1384);
or   g1707 (n1711, n1499, n1295, n1567, n1616);
xnor g1708 (n1701, n1372, n1583, n1443, n1630);
and  g1709 (n1723, n1268, n1613, n1411, n1355);
nand g1710 (n1832, n1391, n1460, n1429, n1603);
nor  g1711 (n1813, n1226, n1207, n1283, n1284);
xnor g1712 (n1765, n1612, n1338, n1538, n1260);
xor  g1713 (n1810, n1469, n1592, n1627, n1500);
xor  g1714 (n1708, n1649, n1548, n1602, n1570);
nor  g1715 (n1731, n1480, n1402, n1566, n1493);
and  g1716 (n1840, n1625, n1209, n1435, n1655);
and  g1717 (n1790, n1550, n1643, n1340, n1203);
and  g1718 (n1687, n1523, n1491, n1178, n1649);
or   g1719 (n1766, n1233, n1216, n1299, n1359);
nor  g1720 (n1709, n1288, n1626, n1621, n1636);
xnor g1721 (n1859, n1173, n1634, n1474, n1510);
nor  g1722 (n1855, n1195, n1456, n1645, n1432);
nor  g1723 (n1779, n1519, n1647, n1201, n1575);
nor  g1724 (n1829, n1430, n1643, n1259, n1660);
xnor g1725 (n1700, n1317, n1632, n1222, n1593);
nand g1726 (n1786, n1579, n1190, n1612, n1431);
or   g1727 (n1732, n1463, n1616, n1575, n1539);
or   g1728 (n1692, n1552, n1365, n1624, n1179);
xnor g1729 (n1681, n1533, n1375, n1281, n1492);
xnor g1730 (n1816, n1390, n1503, n1451, n1436);
or   g1731 (n1801, n1578, n1582, n1373, n1235);
nor  g1732 (n1676, n1271, n1455, n1475, n1568);
nand g1733 (n1851, n1551, n1465, n1552, n1362);
nor  g1734 (n1683, n1445, n1594, n1387, n1598);
xnor g1735 (n1707, n1363, n1485, n1495, n1388);
nor  g1736 (n1821, n1249, n1593, n1220, n1437);
xnor g1737 (n1802, n1353, n1553, n1651, n1580);
nand g1738 (n1838, n1558, n1214, n1645, n1508);
and  g1739 (n1678, n1484, n1647, n1533, n1517);
and  g1740 (n1819, n1655, n1555, n1464, n1629);
and  g1741 (n1800, n1470, n1440, n1475, n1534);
nor  g1742 (n1752, n1567, n1450, n1403, n1388);
and  g1743 (n1824, n1448, n1419, n1264, n1515);
xnor g1744 (n1727, n1646, n1366, n1581, n1591);
and  g1745 (n1759, n1290, n1601, n1606, n1545);
xor  g1746 (n1841, n1350, n1514, n1524, n1420);
or   g1747 (n1725, n1399, n1397, n1594, n1595);
and  g1748 (n1685, n1607, n1312, n1441, n1459);
nand g1749 (n1694, n1419, n1521, n1434, n1556);
or   g1750 (n1748, n1378, n1406, n1349, n1633);
xnor g1751 (n1865, n1638, n1231, n1468, n1614);
or   g1752 (n1720, n1510, n1522, n1318, n1240);
nand g1753 (n1737, n1572, n1387, n1618, n1488);
xor  g1754 (n1724, n1363, n1654, n1177, n1477);
nand g1755 (n1845, n1490, n1394, n1273, n1454);
or   g1756 (n1762, n1476, n1345, n1568, n1386);
xor  g1757 (n1849, n1605, n1332, n1458, n1430);
nand g1758 (n1751, n1261, n1416, n1628, n1446);
nand g1759 (n1782, n1309, n1292, n1357, n1646);
xnor g1760 (n1803, n1211, n1185, n1393, n1640);
and  g1761 (n1745, n1639, n1574, n1454, n1461);
or   g1762 (n1773, n1186, n1400, n1447, n1633);
nand g1763 (n1784, n1478, n1431, n1293, n1296);
and  g1764 (n1797, n1584, n1613, n1390, n1287);
and  g1765 (n1783, n1597, n1379, n1585, n1382);
xnor g1766 (n1764, n1610, n1541, n1435, n1219);
nor  g1767 (n1857, n1254, n1243, n1562, n1498);
nor  g1768 (n1793, n1587, n1370, n1604, n1607);
xor  g1769 (n1753, n1488, n1241, n1506, n1535);
nor  g1770 (n1837, n1642, n1285, n1279, n1333);
or   g1771 (n1785, n1571, n1414, n1275, n1635);
xor  g1772 (n1769, n1418, n1392, n1659, n1494);
xor  g1773 (n1796, n1558, n1442, n1463, n1505);
xnor g1774 (n1761, n1175, n1413, n1335, n1181);
nor  g1775 (n1772, n1427, n1486, n1605, n1397);
nor  g1776 (n1794, n1650, n1263, n1505, n1481);
xnor g1777 (n1714, n1193, n1549, n1621, n1482);
xor  g1778 (n1795, n1358, n1506, n1265, n1401);
nand g1779 (n1831, n1426, n1188, n1656, n1482);
nor  g1780 (n1712, n1472, n1504, n1608, n1531);
nor  g1781 (n1746, n1402, n1217, n1373, n1351);
xnor g1782 (n1750, n1485, n1623, n1520, n1375);
nor  g1783 (n1852, n1371, n1457, n1466, n1587);
nor  g1784 (n1828, n1658, n1227, n1339, n1396);
and  g1785 (n1682, n1395, n1326, n1448, n1579);
or   g1786 (n1864, n1639, n1380, n1590, n1385);
and  g1787 (n1697, n1573, n1546, n1244, n1467);
or   g1788 (n1820, n1342, n1638, n1468, n1389);
nand g1789 (n1738, n1180, n1213, n1524, n1319);
xor  g1790 (n1792, n1642, n1278, n1245, n1453);
and  g1791 (n1689, n1400, n1520, n1529, n1530);
nand g1792 (n1693, n1276, n1379, n1415, n1334);
nand g1793 (n1807, n1208, n1597, n1200, n1395);
xnor g1794 (n1811, n1376, n1336, n1554, n1270);
and  g1795 (n1858, n1599, n1632, n1286, n1383);
xor  g1796 (n1743, n1635, n1421, n1215, n1325);
xor  g1797 (n1736, n1304, n1548, n1651, n1224);
xnor g1798 (n1763, n1228, n1617, n1396, n1423);
and  g1799 (n1863, n1246, n1425, n1583, n1518);
or   g1800 (n1760, n1640, n1650, n1532, n1267);
or   g1801 (n1722, n1462, n1199, n1619, n1444);
or   g1802 (n1826, n1210, n1360, n1629, n1277);
nor  g1803 (n1690, n1644, n1503, n1399, n1502);
xnor g1804 (n1822, n1509, n1424, n1392, n1324);
nor  g1805 (n1710, n1313, n1383, n1449, n1590);
or   g1806 (n1830, n1586, n1549, n1362, n1577);
nor  g1807 (n1734, n1573, n1545, n1457, n1523);
nand g1808 (n1741, n1366, n1297, n1471, n1537);
and  g1809 (n1809, n1405, n1255, n1625, n1555);
or   g1810 (n1705, n1604, n1511, n1206, n1557);
xor  g1811 (n1866, n1329, n1364, n1565, n1592);
and  g1812 (n1721, n1539, n1239, n1461, n1182);
xnor g1813 (n1848, n1238, n1251, n1487, n1600);
xor  g1814 (n1715, n1584, n1352, n1272, n1189);
xor  g1815 (n1702, n1174, n1561, n1623, n1406);
and  g1816 (n1726, n1636, n1508, n1443, n1323);
or   g1817 (n1706, n1384, n1212, n1536, n1391);
xnor g1818 (n1814, n1381, n1528, n1559, n1420);
and  g1819 (n1758, n1553, n1565, n1232, n1308);
xnor g1820 (n1839, n1521, n1404, n1652, n1252);
and  g1821 (n1739, n1449, n1407, n1322, n1426);
nand g1822 (n1729, n1361, n1634, n1528, n1483);
and  g1823 (n1730, n1472, n1364, n1562, n1452);
xnor g1824 (n1787, n1221, n1516, n1371, n1517);
xor  g1825 (n1825, n1291, n1306, n1615, n1445);
and  g1826 (n1791, n1525, n1473, n1331, n1367);
nand g1827 (n1815, n1588, n1494, n1591, n1417);
or   g1828 (n1754, n1303, n1537, n1531, n1473);
or   g1829 (n1674, n1298, n1547, n1512, n1253);
nand g1830 (n1713, n1183, n1466, n1644, n1198);
xnor g1831 (n1834, n1247, n1192, n1337, n1518);
nor  g1832 (n1686, n1374, n1479, n1405, n1316);
or   g1833 (n1728, n1458, n1589, n1490, n1540);
nor  g1834 (n1799, n1398, n1401, n1433, n1446);
nand g1835 (n1717, n1347, n1346, n1501, n1176);
and  g1836 (n1777, n1237, n1561, n1386, n1412);
nand g1837 (n1862, n1476, n1615, n1327, n1601);
nand g1838 (n1876, n1704, n1780, n1736, n1774);
nor  g1839 (n1877, n1694, n1778, n1767, n1787);
xor  g1840 (n1882, n1726, n1737, n1725, n1803);
nor  g1841 (n1888, n1749, n1784, n1788, n1684);
nand g1842 (n1872, n1768, n1791, n1748, n1722);
xnor g1843 (n1893, n1681, n1769, n1703, n1738);
and  g1844 (n1895, n1674, n1676, n1806, n1755);
nand g1845 (n1889, n1729, n1747, n1707, n1682);
or   g1846 (n1896, n1745, n1716, n1759, n1781);
nor  g1847 (n1890, n1809, n1798, n1782, n1779);
nor  g1848 (n1891, n1719, n1698, n1691, n1734);
and  g1849 (n1880, n1760, n1700, n1742, n1714);
xnor g1850 (n1894, n1706, n1772, n1757, n1804);
and  g1851 (n1873, n1705, n1740, n1802, n1730);
or   g1852 (n1898, n1708, n1689, n1688, n1786);
and  g1853 (n1875, n1686, n1796, n1690, n1765);
and  g1854 (n1884, n1812, n1711, n1785, n1801);
and  g1855 (n1881, n1728, n1800, n1741, n1766);
nand g1856 (n1883, n1721, n1754, n1699, n1697);
nand g1857 (n1900, n1761, n1743, n1763, n1713);
nand g1858 (n1892, n1756, n1770, n1687, n1685);
or   g1859 (n1879, n1762, n1678, n1753, n1795);
and  g1860 (n1904, n1783, n1744, n1773, n1777);
xor  g1861 (n1901, n1805, n1680, n1724, n1794);
xnor g1862 (n1878, n1797, n1776, n1731, n1807);
and  g1863 (n1903, n1746, n1712, n1808, n1750);
nand g1864 (n1902, n1709, n1732, n1813, n1710);
nor  g1865 (n1899, n1758, n1717, n1692, n1679);
and  g1866 (n1887, n1752, n1677, n1720, n1810);
xor  g1867 (n1886, n1702, n1683, n1715, n1789);
and  g1868 (n1871, n1733, n1811, n1793, n1751);
xnor g1869 (n1874, n1790, n1764, n1771, n1775);
xor  g1870 (n1905, n1723, n1799, n1695, n1727);
or   g1871 (n1885, n1693, n1701, n1675, n1696);
and  g1872 (n1897, n1792, n1718, n1735, n1739);
buf  g1873 (n1907, n1875);
not  g1874 (n1908, n1874);
xnor g1875 (n1906, n1876, n1660);
not  g1876 (n1914, n1908);
not  g1877 (n1913, n1906);
buf  g1878 (n1916, n1907);
buf  g1879 (n1915, n1906);
not  g1880 (n1910, n1907);
buf  g1881 (n1918, n1906);
buf  g1882 (n1911, n1907);
not  g1883 (n1909, n1907);
not  g1884 (n1912, n1908);
buf  g1885 (n1917, n1906);
not  g1886 (n1950, n1917);
not  g1887 (n1947, n1913);
not  g1888 (n1939, n1837);
not  g1889 (n1941, n1912);
buf  g1890 (n1946, n1840);
not  g1891 (n1937, n1911);
not  g1892 (n1923, n1842);
not  g1893 (n1949, n1916);
not  g1894 (n1942, n1914);
buf  g1895 (n1924, n1912);
not  g1896 (n1930, n1913);
not  g1897 (n1932, n1822);
not  g1898 (n1934, n1815);
buf  g1899 (n1920, n1820);
buf  g1900 (n1940, n1916);
buf  g1901 (n1922, n1829);
not  g1902 (n1925, n1913);
buf  g1903 (n1935, n1915);
not  g1904 (n1926, n1817);
buf  g1905 (n1948, n1828);
xnor g1906 (n1936, n1915, n1911);
xor  g1907 (n1928, n1917, n1912);
and  g1908 (n1927, n1913, n1827, n1823, n1835);
xor  g1909 (n1931, n1915, n1914, n1917, n1826);
nor  g1910 (n1919, n1844, n1832, n1845, n1909);
nand g1911 (n1921, n1918, n1918, n1910, n1816);
xor  g1912 (n1945, n1824, n1912, n1916, n1915);
xnor g1913 (n1944, n1821, n1909, n1819, n1914);
xnor g1914 (n1938, n1818, n1833, n1839, n1831);
xnor g1915 (n1929, n1834, n1814, n1838, n1836);
or   g1916 (n1943, n1830, n1843, n1910, n1917);
nand g1917 (n1933, n1825, n1841, n1914, n1916);
not  g1918 (n1972, n1908);
buf  g1919 (n1963, n1919);
xor  g1920 (n1953, n1905, n585, n1892, n1948);
and  g1921 (n1968, n1900, n1931, n1949, n1854);
xnor g1922 (n1951, n1856, n1937, n1883, n1897);
nand g1923 (n1961, n1887, n187, n1852, n1661);
or   g1924 (n1969, n1939, n1926, n464, n1866);
xnor g1925 (n1958, n1891, n1940, n1878, n1899);
or   g1926 (n1971, n1664, n585, n1663, n1847);
xnor g1927 (n1979, n1849, n463, n1853, n1867);
nor  g1928 (n1957, n1894, n1943, n1859, n586);
or   g1929 (n1974, n1855, n1935, n1934, n1862);
nand g1930 (n1967, n1663, n1941, n1858, n1902);
and  g1931 (n1970, n1932, n585, n1662, n1863);
nand g1932 (n1976, n1947, n586, n464, n1661);
and  g1933 (n1973, n1903, n1890, n1930, n1666);
and  g1934 (n1956, n1936, n1920, n1927, n1861);
nand g1935 (n1960, n1882, n464, n1860, n586);
and  g1936 (n1954, n1880, n1868, n1928, n1942);
and  g1937 (n1980, n1921, n586, n1945, n1946);
nand g1938 (n1965, n1901, n1893, n1667, n1851);
and  g1939 (n1964, n1846, n1857, n1662, n1888);
nor  g1940 (n1966, n1869, n1933, n585, n1898);
nor  g1941 (n1977, n1850, n1881, n1925, n1667);
and  g1942 (n1959, n1922, n1665, n1895, n1666);
and  g1943 (n1952, n1885, n1938, n1848, n1923);
and  g1944 (n1978, n1884, n1879, n1668, n1905);
and  g1945 (n1962, n1889, n1950, n1664, n464);
xnor g1946 (n1955, n1877, n1929, n1944, n1865);
nand g1947 (n1981, n1886, n462, n1864, n1665);
or   g1948 (n1975, n1908, n1896, n1904, n1924);
buf  g1949 (n2007, n1968);
not  g1950 (n2006, n1963);
buf  g1951 (n2013, n1964);
not  g1952 (n1992, n1951);
not  g1953 (n1991, n28);
not  g1954 (n2020, n1973);
buf  g1955 (n1996, n1954);
buf  g1956 (n2005, n1975);
not  g1957 (n2010, n1971);
not  g1958 (n2011, n29);
not  g1959 (n1986, n1965);
not  g1960 (n2000, n1965);
buf  g1961 (n2009, n29);
buf  g1962 (n2015, n1975);
not  g1963 (n1990, n1978);
buf  g1964 (n1993, n1670);
not  g1965 (n2002, n1972);
not  g1966 (n1999, n1967);
buf  g1967 (n1988, n1959);
not  g1968 (n2008, n1962);
buf  g1969 (n1985, n31);
buf  g1970 (n2001, n1970);
not  g1971 (n2004, n1971);
buf  g1972 (n2016, n1918);
buf  g1973 (n1998, n31);
buf  g1974 (n2003, n1972);
or   g1975 (n1989, n1966, n1981, n28);
and  g1976 (n1987, n30, n31, n1973, n1976);
and  g1977 (n1982, n1974, n1981, n29, n1979);
or   g1978 (n2018, n1960, n1918, n1963, n1977);
nand g1979 (n2019, n1957, n1961, n30, n1953);
nand g1980 (n1997, n1974, n29, n1955, n28);
xor  g1981 (n2021, n31, n1980, n32, n1966);
nor  g1982 (n1994, n1977, n1952, n1956, n1671);
nand g1983 (n2012, n1964, n1970, n1958, n1672);
nand g1984 (n2017, n1670, n1968, n1980, n1671);
and  g1985 (n2014, n30, n1668, n1976, n1967);
nand g1986 (n1983, n30, n1870, n1969, n1669);
nor  g1987 (n1984, n1672, n1961, n1978, n1979);
xnor g1988 (n1995, n1962, n1969, n1669, n1673);
or   g1989 (n2031, n2015, n2011, n1993, n2003);
or   g1990 (n2028, n32, n32, n1985, n2005);
xnor g1991 (n2032, n2008, n2018, n2000, n2014);
nand g1992 (n2022, n2007, n2017, n2010, n1992);
nand g1993 (n2024, n1987, n1988, n1983, n1995);
xnor g1994 (n2026, n2019, n1673, n2012, n2013);
or   g1995 (n2027, n1984, n1999, n2001, n1982);
xor  g1996 (n2023, n1991, n2016, n1996, n2020);
or   g1997 (n2025, n2002, n1986, n1989, n2021);
xor  g1998 (n2029, n1997, n2009, n1994, n1998);
xnor g1999 (n2030, n32, n1990, n2004, n2006);
endmodule
