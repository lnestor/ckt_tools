

module Stat_1343_29_11
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1000,
  n997,
  n1007,
  n1016,
  n1014,
  n1025,
  n1024,
  n1003,
  n1002,
  n1022,
  n1005,
  n996,
  n998,
  n1023,
  n1001,
  n1021,
  n1004,
  n1015,
  n1017,
  n1010,
  n1006,
  n1013,
  n999,
  n1009,
  n1011,
  n1008,
  n1094,
  n1089,
  n1092,
  n1096,
  n1100,
  n1098,
  n1097,
  n1375,
  n1373,
  n1372,
  n1371,
  n1370,
  n1374,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1000;
  output n997;
  output n1007;
  output n1016;
  output n1014;
  output n1025;
  output n1024;
  output n1003;
  output n1002;
  output n1022;
  output n1005;
  output n996;
  output n998;
  output n1023;
  output n1001;
  output n1021;
  output n1004;
  output n1015;
  output n1017;
  output n1010;
  output n1006;
  output n1013;
  output n999;
  output n1009;
  output n1011;
  output n1008;
  output n1094;
  output n1089;
  output n1092;
  output n1096;
  output n1100;
  output n1098;
  output n1097;
  output n1375;
  output n1373;
  output n1372;
  output n1371;
  output n1370;
  output n1374;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n1012;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1090;
  wire n1091;
  wire n1093;
  wire n1095;
  wire n1099;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n104,
    n31
  );


  buf
  g1
  (
    n97,
    n5
  );


  buf
  g2
  (
    n101,
    n7
  );


  not
  g3
  (
    n148,
    n5
  );


  buf
  g4
  (
    n35,
    n11
  );


  not
  g5
  (
    n125,
    n24
  );


  not
  g6
  (
    n61,
    n9
  );


  not
  g7
  (
    n139,
    n25
  );


  not
  g8
  (
    n149,
    n4
  );


  not
  g9
  (
    n128,
    n28
  );


  buf
  g10
  (
    n105,
    n28
  );


  not
  g11
  (
    n96,
    n24
  );


  buf
  g12
  (
    n89,
    n28
  );


  not
  g13
  (
    n67,
    n10
  );


  not
  g14
  (
    n45,
    n15
  );


  buf
  g15
  (
    n134,
    n2
  );


  not
  g16
  (
    n116,
    n29
  );


  buf
  g17
  (
    n133,
    n30
  );


  buf
  g18
  (
    n131,
    n19
  );


  buf
  g19
  (
    n43,
    n31
  );


  not
  g20
  (
    n159,
    n1
  );


  not
  g21
  (
    n106,
    n21
  );


  buf
  g22
  (
    n103,
    n22
  );


  not
  g23
  (
    n102,
    n12
  );


  not
  g24
  (
    n121,
    n27
  );


  not
  g25
  (
    n113,
    n27
  );


  buf
  g26
  (
    n68,
    n11
  );


  not
  g27
  (
    n123,
    n12
  );


  not
  g28
  (
    n79,
    n8
  );


  not
  g29
  (
    n76,
    n6
  );


  buf
  g30
  (
    n80,
    n28
  );


  not
  g31
  (
    n160,
    n10
  );


  not
  g32
  (
    n98,
    n22
  );


  buf
  g33
  (
    n95,
    n22
  );


  buf
  g34
  (
    n114,
    n26
  );


  buf
  g35
  (
    n120,
    n7
  );


  not
  g36
  (
    n60,
    n25
  );


  buf
  g37
  (
    n40,
    n15
  );


  buf
  g38
  (
    n47,
    n7
  );


  buf
  g39
  (
    n37,
    n16
  );


  not
  g40
  (
    n132,
    n6
  );


  not
  g41
  (
    n138,
    n30
  );


  buf
  g42
  (
    n74,
    n26
  );


  not
  g43
  (
    n115,
    n32
  );


  buf
  g44
  (
    n84,
    n9
  );


  not
  g45
  (
    n92,
    n5
  );


  not
  g46
  (
    n136,
    n2
  );


  buf
  g47
  (
    n65,
    n10
  );


  not
  g48
  (
    n34,
    n6
  );


  not
  g49
  (
    n143,
    n29
  );


  not
  g50
  (
    n151,
    n17
  );


  not
  g51
  (
    n81,
    n26
  );


  buf
  g52
  (
    n49,
    n16
  );


  not
  g53
  (
    n56,
    n32
  );


  not
  g54
  (
    n62,
    n24
  );


  buf
  g55
  (
    n155,
    n29
  );


  not
  g56
  (
    n150,
    n6
  );


  not
  g57
  (
    n145,
    n31
  );


  buf
  g58
  (
    n108,
    n14
  );


  buf
  g59
  (
    n156,
    n14
  );


  not
  g60
  (
    n75,
    n23
  );


  buf
  g61
  (
    n99,
    n9
  );


  buf
  g62
  (
    n83,
    n22
  );


  not
  g63
  (
    n54,
    n11
  );


  not
  g64
  (
    n82,
    n20
  );


  not
  g65
  (
    n88,
    n19
  );


  not
  g66
  (
    n158,
    n18
  );


  not
  g67
  (
    n73,
    n24
  );


  not
  g68
  (
    n129,
    n14
  );


  not
  g69
  (
    n146,
    n1
  );


  not
  g70
  (
    n107,
    n4
  );


  not
  g71
  (
    n87,
    n19
  );


  buf
  g72
  (
    n69,
    n13
  );


  not
  g73
  (
    n117,
    n23
  );


  not
  g74
  (
    n46,
    n13
  );


  buf
  g75
  (
    n126,
    n25
  );


  not
  g76
  (
    n86,
    n8
  );


  not
  g77
  (
    n90,
    n13
  );


  not
  g78
  (
    n110,
    n1
  );


  not
  g79
  (
    n42,
    n3
  );


  buf
  g80
  (
    n144,
    n14
  );


  buf
  g81
  (
    n109,
    n23
  );


  buf
  g82
  (
    n53,
    n20
  );


  not
  g83
  (
    KeyWire_0_0,
    n17
  );


  not
  g84
  (
    n33,
    n20
  );


  not
  g85
  (
    n36,
    n32
  );


  not
  g86
  (
    n127,
    n16
  );


  buf
  g87
  (
    n58,
    n3
  );


  not
  g88
  (
    n63,
    n13
  );


  buf
  g89
  (
    n64,
    n15
  );


  buf
  g90
  (
    n66,
    n5
  );


  buf
  g91
  (
    n78,
    n31
  );


  not
  g92
  (
    n94,
    n2
  );


  not
  g93
  (
    n51,
    n15
  );


  not
  g94
  (
    KeyWire_0_12,
    n9
  );


  not
  g95
  (
    n50,
    n23
  );


  buf
  g96
  (
    n112,
    n18
  );


  buf
  g97
  (
    n59,
    n2
  );


  not
  g98
  (
    n142,
    n8
  );


  not
  g99
  (
    n135,
    n21
  );


  buf
  g100
  (
    n154,
    n10
  );


  not
  g101
  (
    n157,
    n18
  );


  not
  g102
  (
    n72,
    n25
  );


  not
  g103
  (
    n57,
    n7
  );


  not
  g104
  (
    n140,
    n17
  );


  not
  g105
  (
    n147,
    n27
  );


  not
  g106
  (
    n118,
    n20
  );


  buf
  g107
  (
    n77,
    n29
  );


  not
  g108
  (
    n91,
    n30
  );


  not
  g109
  (
    n130,
    n4
  );


  not
  g110
  (
    n124,
    n3
  );


  not
  g111
  (
    n141,
    n3
  );


  not
  g112
  (
    n71,
    n21
  );


  buf
  g113
  (
    n137,
    n18
  );


  not
  g114
  (
    n48,
    n12
  );


  not
  g115
  (
    n52,
    n30
  );


  buf
  g116
  (
    n41,
    n11
  );


  buf
  g117
  (
    n122,
    n1
  );


  not
  g118
  (
    n85,
    n8
  );


  not
  g119
  (
    n152,
    n21
  );


  buf
  g120
  (
    n44,
    n12
  );


  buf
  g121
  (
    n153,
    n26
  );


  not
  g122
  (
    n111,
    n17
  );


  buf
  g123
  (
    n39,
    n4
  );


  buf
  g124
  (
    n119,
    n32
  );


  not
  g125
  (
    n100,
    n16
  );


  not
  g126
  (
    n70,
    n27
  );


  buf
  g127
  (
    n93,
    n19
  );


  not
  g128
  (
    n487,
    n110
  );


  not
  g129
  (
    n547,
    n81
  );


  buf
  g130
  (
    n604,
    n125
  );


  buf
  g131
  (
    n312,
    n71
  );


  buf
  g132
  (
    n376,
    n101
  );


  not
  g133
  (
    n372,
    n47
  );


  not
  g134
  (
    n586,
    n129
  );


  not
  g135
  (
    n526,
    n112
  );


  not
  g136
  (
    n433,
    n137
  );


  buf
  g137
  (
    n231,
    n87
  );


  buf
  g138
  (
    n582,
    n106
  );


  not
  g139
  (
    KeyWire_0_6,
    n96
  );


  buf
  g140
  (
    n406,
    n107
  );


  not
  g141
  (
    n248,
    n69
  );


  not
  g142
  (
    n218,
    n74
  );


  buf
  g143
  (
    n193,
    n97
  );


  buf
  g144
  (
    n513,
    n127
  );


  not
  g145
  (
    n198,
    n58
  );


  not
  g146
  (
    n332,
    n88
  );


  buf
  g147
  (
    n187,
    n132
  );


  buf
  g148
  (
    n352,
    n53
  );


  buf
  g149
  (
    n163,
    n112
  );


  not
  g150
  (
    n573,
    n117
  );


  buf
  g151
  (
    n359,
    n45
  );


  not
  g152
  (
    n466,
    n44
  );


  not
  g153
  (
    n316,
    n62
  );


  buf
  g154
  (
    n483,
    n76
  );


  not
  g155
  (
    n377,
    n79
  );


  not
  g156
  (
    n293,
    n86
  );


  buf
  g157
  (
    n562,
    n70
  );


  not
  g158
  (
    n400,
    n92
  );


  not
  g159
  (
    n486,
    n109
  );


  not
  g160
  (
    n253,
    n45
  );


  buf
  g161
  (
    n602,
    n120
  );


  not
  g162
  (
    n267,
    n83
  );


  not
  g163
  (
    n386,
    n126
  );


  buf
  g164
  (
    n226,
    n103
  );


  buf
  g165
  (
    n407,
    n91
  );


  not
  g166
  (
    n511,
    n86
  );


  not
  g167
  (
    n503,
    n70
  );


  not
  g168
  (
    n334,
    n122
  );


  buf
  g169
  (
    n328,
    n89
  );


  not
  g170
  (
    n369,
    n71
  );


  buf
  g171
  (
    n385,
    n55
  );


  buf
  g172
  (
    n257,
    n49
  );


  buf
  g173
  (
    n454,
    n116
  );


  not
  g174
  (
    n566,
    n105
  );


  buf
  g175
  (
    n393,
    n121
  );


  not
  g176
  (
    n176,
    n46
  );


  not
  g177
  (
    n202,
    n68
  );


  not
  g178
  (
    n571,
    n109
  );


  buf
  g179
  (
    n601,
    n52
  );


  buf
  g180
  (
    n476,
    n53
  );


  buf
  g181
  (
    n205,
    n117
  );


  not
  g182
  (
    n471,
    n128
  );


  buf
  g183
  (
    n296,
    n89
  );


  buf
  g184
  (
    n256,
    n41
  );


  buf
  g185
  (
    n451,
    n115
  );


  not
  g186
  (
    n525,
    n45
  );


  not
  g187
  (
    n184,
    n142
  );


  not
  g188
  (
    n335,
    n42
  );


  not
  g189
  (
    n264,
    n79
  );


  buf
  g190
  (
    n346,
    n118
  );


  not
  g191
  (
    n307,
    n131
  );


  not
  g192
  (
    n445,
    n37
  );


  not
  g193
  (
    n404,
    n98
  );


  buf
  g194
  (
    n188,
    n91
  );


  not
  g195
  (
    n214,
    n53
  );


  buf
  g196
  (
    n438,
    n82
  );


  not
  g197
  (
    n277,
    n77
  );


  not
  g198
  (
    n192,
    n99
  );


  buf
  g199
  (
    n431,
    n37
  );


  buf
  g200
  (
    n512,
    n69
  );


  not
  g201
  (
    n272,
    n112
  );


  not
  g202
  (
    n494,
    n114
  );


  buf
  g203
  (
    n380,
    n141
  );


  buf
  g204
  (
    n165,
    n99
  );


  not
  g205
  (
    n331,
    n64
  );


  buf
  g206
  (
    n230,
    n66
  );


  buf
  g207
  (
    n164,
    n133
  );


  buf
  g208
  (
    n429,
    n47
  );


  not
  g209
  (
    n458,
    n117
  );


  not
  g210
  (
    n572,
    n68
  );


  buf
  g211
  (
    n215,
    n87
  );


  not
  g212
  (
    n554,
    n49
  );


  not
  g213
  (
    n227,
    n80
  );


  buf
  g214
  (
    n373,
    n115
  );


  not
  g215
  (
    n489,
    n125
  );


  buf
  g216
  (
    n460,
    n113
  );


  not
  g217
  (
    n271,
    n142
  );


  buf
  g218
  (
    n500,
    n117
  );


  not
  g219
  (
    n200,
    n36
  );


  not
  g220
  (
    n493,
    n137
  );


  buf
  g221
  (
    n576,
    n58
  );


  not
  g222
  (
    n415,
    n83
  );


  buf
  g223
  (
    n375,
    n75
  );


  buf
  g224
  (
    n515,
    n78
  );


  not
  g225
  (
    n244,
    n133
  );


  buf
  g226
  (
    n242,
    n90
  );


  not
  g227
  (
    n565,
    n103
  );


  not
  g228
  (
    n261,
    n63
  );


  not
  g229
  (
    n358,
    n49
  );


  not
  g230
  (
    n574,
    n67
  );


  not
  g231
  (
    n343,
    n103
  );


  buf
  g232
  (
    n496,
    n88
  );


  buf
  g233
  (
    n440,
    n130
  );


  not
  g234
  (
    n491,
    n104
  );


  not
  g235
  (
    n599,
    n93
  );


  buf
  g236
  (
    n351,
    n61
  );


  not
  g237
  (
    n459,
    n131
  );


  not
  g238
  (
    n243,
    n110
  );


  not
  g239
  (
    n347,
    n135
  );


  buf
  g240
  (
    n546,
    n108
  );


  buf
  g241
  (
    n357,
    n80
  );


  not
  g242
  (
    n583,
    n79
  );


  not
  g243
  (
    n324,
    n94
  );


  not
  g244
  (
    n603,
    n113
  );


  not
  g245
  (
    n559,
    n79
  );


  buf
  g246
  (
    n366,
    n84
  );


  not
  g247
  (
    n502,
    n118
  );


  not
  g248
  (
    n402,
    n67
  );


  not
  g249
  (
    n298,
    n47
  );


  buf
  g250
  (
    n301,
    n81
  );


  buf
  g251
  (
    n234,
    n139
  );


  buf
  g252
  (
    n428,
    n43
  );


  not
  g253
  (
    n222,
    n68
  );


  buf
  g254
  (
    n306,
    n51
  );


  buf
  g255
  (
    n439,
    n95
  );


  not
  g256
  (
    n560,
    n57
  );


  buf
  g257
  (
    n474,
    n142
  );


  not
  g258
  (
    n521,
    n108
  );


  buf
  g259
  (
    n452,
    n93
  );


  not
  g260
  (
    n421,
    n136
  );


  not
  g261
  (
    n490,
    n102
  );


  not
  g262
  (
    n262,
    n63
  );


  buf
  g263
  (
    n172,
    n118
  );


  buf
  g264
  (
    n279,
    n34
  );


  buf
  g265
  (
    n555,
    n138
  );


  not
  g266
  (
    n178,
    n98
  );


  buf
  g267
  (
    n529,
    n95
  );


  not
  g268
  (
    n225,
    n135
  );


  not
  g269
  (
    n436,
    n52
  );


  not
  g270
  (
    n598,
    n95
  );


  buf
  g271
  (
    n553,
    n143
  );


  not
  g272
  (
    n223,
    n74
  );


  not
  g273
  (
    n191,
    n47
  );


  buf
  g274
  (
    n414,
    n40
  );


  buf
  g275
  (
    n396,
    n123
  );


  buf
  g276
  (
    n367,
    n138
  );


  buf
  g277
  (
    n287,
    n137
  );


  not
  g278
  (
    n542,
    n59
  );


  buf
  g279
  (
    n300,
    n111
  );


  buf
  g280
  (
    n520,
    n130
  );


  buf
  g281
  (
    n282,
    n137
  );


  buf
  g282
  (
    n238,
    n98
  );


  not
  g283
  (
    n561,
    n97
  );


  buf
  g284
  (
    n278,
    n121
  );


  not
  g285
  (
    n587,
    n41
  );


  buf
  g286
  (
    KeyWire_0_11,
    n140
  );


  buf
  g287
  (
    n390,
    n114
  );


  buf
  g288
  (
    n353,
    n65
  );


  not
  g289
  (
    n568,
    n69
  );


  not
  g290
  (
    n322,
    n91
  );


  buf
  g291
  (
    n302,
    n73
  );


  buf
  g292
  (
    n444,
    n119
  );


  buf
  g293
  (
    n528,
    n83
  );


  buf
  g294
  (
    n434,
    n33
  );


  not
  g295
  (
    n340,
    n124
  );


  not
  g296
  (
    n510,
    n80
  );


  buf
  g297
  (
    n391,
    n120
  );


  not
  g298
  (
    n548,
    n60
  );


  buf
  g299
  (
    n195,
    n105
  );


  not
  g300
  (
    n318,
    n128
  );


  not
  g301
  (
    n326,
    n120
  );


  buf
  g302
  (
    n240,
    n110
  );


  buf
  g303
  (
    n294,
    n124
  );


  not
  g304
  (
    n456,
    n85
  );


  buf
  g305
  (
    n285,
    n55
  );


  not
  g306
  (
    n299,
    n141
  );


  not
  g307
  (
    n442,
    n134
  );


  not
  g308
  (
    n311,
    n96
  );


  not
  g309
  (
    n484,
    n52
  );


  not
  g310
  (
    n167,
    n129
  );


  buf
  g311
  (
    n286,
    n48
  );


  not
  g312
  (
    n304,
    n81
  );


  not
  g313
  (
    n410,
    n124
  );


  not
  g314
  (
    n196,
    n102
  );


  not
  g315
  (
    n580,
    n126
  );


  not
  g316
  (
    n435,
    n134
  );


  buf
  g317
  (
    n585,
    n106
  );


  not
  g318
  (
    n541,
    n116
  );


  not
  g319
  (
    n501,
    n41
  );


  buf
  g320
  (
    n329,
    n122
  );


  buf
  g321
  (
    n535,
    n46
  );


  not
  g322
  (
    n310,
    n40
  );


  not
  g323
  (
    n588,
    n100
  );


  not
  g324
  (
    n563,
    n136
  );


  not
  g325
  (
    n464,
    n108
  );


  buf
  g326
  (
    n412,
    n97
  );


  buf
  g327
  (
    n250,
    n34
  );


  buf
  g328
  (
    n337,
    n114
  );


  not
  g329
  (
    n213,
    n54
  );


  not
  g330
  (
    n259,
    n62
  );


  buf
  g331
  (
    n177,
    n77
  );


  not
  g332
  (
    n246,
    n73
  );


  not
  g333
  (
    n170,
    n101
  );


  buf
  g334
  (
    n179,
    n71
  );


  buf
  g335
  (
    n488,
    n69
  );


  not
  g336
  (
    n325,
    n92
  );


  buf
  g337
  (
    n544,
    n78
  );


  not
  g338
  (
    n189,
    n107
  );


  buf
  g339
  (
    n185,
    n129
  );


  buf
  g340
  (
    n403,
    n130
  );


  not
  g341
  (
    n204,
    n66
  );


  not
  g342
  (
    n543,
    n54
  );


  buf
  g343
  (
    n537,
    n72
  );


  buf
  g344
  (
    n523,
    n135
  );


  buf
  g345
  (
    n216,
    n143
  );


  buf
  g346
  (
    n365,
    n115
  );


  not
  g347
  (
    n453,
    n134
  );


  buf
  g348
  (
    n449,
    n139
  );


  not
  g349
  (
    n345,
    n82
  );


  buf
  g350
  (
    n273,
    n55
  );


  not
  g351
  (
    n290,
    n127
  );


  not
  g352
  (
    n443,
    n57
  );


  not
  g353
  (
    n221,
    n40
  );


  buf
  g354
  (
    n239,
    n107
  );


  not
  g355
  (
    n382,
    n43
  );


  buf
  g356
  (
    n423,
    n95
  );


  not
  g357
  (
    KeyWire_0_3,
    n56
  );


  not
  g358
  (
    n288,
    n82
  );


  not
  g359
  (
    n245,
    n52
  );


  not
  g360
  (
    n505,
    n128
  );


  not
  g361
  (
    n263,
    n105
  );


  buf
  g362
  (
    n564,
    n64
  );


  not
  g363
  (
    n570,
    n86
  );


  buf
  g364
  (
    n397,
    n74
  );


  not
  g365
  (
    n190,
    n55
  );


  not
  g366
  (
    n508,
    n39
  );


  not
  g367
  (
    n274,
    n65
  );


  not
  g368
  (
    n409,
    n87
  );


  not
  g369
  (
    n379,
    n143
  );


  buf
  g370
  (
    n252,
    n67
  );


  buf
  g371
  (
    n203,
    n48
  );


  not
  g372
  (
    n219,
    n111
  );


  buf
  g373
  (
    n595,
    n99
  );


  buf
  g374
  (
    n197,
    n43
  );


  buf
  g375
  (
    n478,
    n71
  );


  not
  g376
  (
    n498,
    n132
  );


  not
  g377
  (
    n388,
    n113
  );


  buf
  g378
  (
    n507,
    n33
  );


  not
  g379
  (
    n249,
    n101
  );


  buf
  g380
  (
    n339,
    n48
  );


  not
  g381
  (
    n371,
    n141
  );


  buf
  g382
  (
    n364,
    n85
  );


  buf
  g383
  (
    n509,
    n60
  );


  not
  g384
  (
    n551,
    n36
  );


  buf
  g385
  (
    n519,
    n61
  );


  buf
  g386
  (
    n321,
    n135
  );


  buf
  g387
  (
    n284,
    n108
  );


  buf
  g388
  (
    n592,
    n59
  );


  buf
  g389
  (
    n527,
    n140
  );


  not
  g390
  (
    n208,
    n131
  );


  buf
  g391
  (
    n236,
    n62
  );


  buf
  g392
  (
    n534,
    n64
  );


  buf
  g393
  (
    n417,
    n100
  );


  buf
  g394
  (
    n480,
    n127
  );


  buf
  g395
  (
    n538,
    n54
  );


  buf
  g396
  (
    n465,
    n127
  );


  buf
  g397
  (
    n430,
    n142
  );


  buf
  g398
  (
    n292,
    n123
  );


  not
  g399
  (
    n497,
    n124
  );


  buf
  g400
  (
    n600,
    n38
  );


  not
  g401
  (
    n539,
    n63
  );


  buf
  g402
  (
    n405,
    n39
  );


  not
  g403
  (
    n360,
    n76
  );


  not
  g404
  (
    n427,
    n126
  );


  buf
  g405
  (
    n330,
    n50
  );


  buf
  g406
  (
    n295,
    n133
  );


  buf
  g407
  (
    n313,
    n56
  );


  buf
  g408
  (
    n420,
    n141
  );


  not
  g409
  (
    n462,
    n105
  );


  not
  g410
  (
    n395,
    n125
  );


  not
  g411
  (
    n171,
    n98
  );


  not
  g412
  (
    n408,
    n46
  );


  not
  g413
  (
    n597,
    n33
  );


  not
  g414
  (
    n199,
    n66
  );


  buf
  g415
  (
    n499,
    n96
  );


  not
  g416
  (
    n220,
    n139
  );


  buf
  g417
  (
    n556,
    n87
  );


  buf
  g418
  (
    n291,
    n78
  );


  buf
  g419
  (
    n550,
    n111
  );


  buf
  g420
  (
    n530,
    n90
  );


  not
  g421
  (
    n591,
    n61
  );


  buf
  g422
  (
    n461,
    n78
  );


  buf
  g423
  (
    n447,
    n94
  );


  not
  g424
  (
    n398,
    n44
  );


  not
  g425
  (
    n470,
    n109
  );


  not
  g426
  (
    n581,
    n133
  );


  not
  g427
  (
    n338,
    n46
  );


  buf
  g428
  (
    n206,
    n68
  );


  not
  g429
  (
    n348,
    n96
  );


  not
  g430
  (
    n174,
    n75
  );


  not
  g431
  (
    n342,
    n84
  );


  buf
  g432
  (
    n383,
    n50
  );


  buf
  g433
  (
    n211,
    n51
  );


  not
  g434
  (
    n590,
    n123
  );


  buf
  g435
  (
    n229,
    n104
  );


  not
  g436
  (
    n168,
    n140
  );


  not
  g437
  (
    n522,
    n104
  );


  not
  g438
  (
    n224,
    n50
  );


  not
  g439
  (
    n593,
    n51
  );


  not
  g440
  (
    n166,
    n60
  );


  not
  g441
  (
    n247,
    n66
  );


  not
  g442
  (
    n552,
    n35
  );


  buf
  g443
  (
    n514,
    n59
  );


  buf
  g444
  (
    n567,
    n70
  );


  not
  g445
  (
    n394,
    n128
  );


  buf
  g446
  (
    n210,
    n43
  );


  buf
  g447
  (
    n201,
    n33
  );


  not
  g448
  (
    n232,
    n94
  );


  buf
  g449
  (
    n241,
    n72
  );


  not
  g450
  (
    n477,
    n35
  );


  buf
  g451
  (
    n485,
    n140
  );


  buf
  g452
  (
    n584,
    n56
  );


  not
  g453
  (
    n536,
    n77
  );


  not
  g454
  (
    n255,
    n48
  );


  not
  g455
  (
    KeyWire_0_5,
    n85
  );


  not
  g456
  (
    n320,
    n44
  );


  buf
  g457
  (
    n579,
    n38
  );


  not
  g458
  (
    n549,
    n91
  );


  buf
  g459
  (
    n569,
    n63
  );


  buf
  g460
  (
    n381,
    n35
  );


  not
  g461
  (
    n557,
    n60
  );


  not
  g462
  (
    n186,
    n134
  );


  buf
  g463
  (
    n578,
    n122
  );


  buf
  g464
  (
    n289,
    n125
  );


  not
  g465
  (
    n419,
    n113
  );


  buf
  g466
  (
    n387,
    n38
  );


  buf
  g467
  (
    n506,
    n102
  );


  not
  g468
  (
    n162,
    n119
  );


  not
  g469
  (
    n441,
    n81
  );


  not
  g470
  (
    n424,
    n83
  );


  not
  g471
  (
    n319,
    n103
  );


  not
  g472
  (
    n275,
    n110
  );


  buf
  g473
  (
    n260,
    n106
  );


  not
  g474
  (
    n475,
    n89
  );


  not
  g475
  (
    n492,
    n131
  );


  buf
  g476
  (
    n309,
    n136
  );


  not
  g477
  (
    n297,
    n36
  );


  not
  g478
  (
    n182,
    n143
  );


  not
  g479
  (
    n370,
    n44
  );


  buf
  g480
  (
    n323,
    n57
  );


  buf
  g481
  (
    n384,
    n76
  );


  buf
  g482
  (
    n207,
    n107
  );


  not
  g483
  (
    n173,
    n73
  );


  not
  g484
  (
    n350,
    n54
  );


  buf
  g485
  (
    n180,
    n67
  );


  buf
  g486
  (
    n532,
    n129
  );


  not
  g487
  (
    n254,
    n109
  );


  buf
  g488
  (
    n266,
    n132
  );


  not
  g489
  (
    n596,
    n122
  );


  not
  g490
  (
    n378,
    n136
  );


  not
  g491
  (
    n268,
    n114
  );


  buf
  g492
  (
    n463,
    n92
  );


  buf
  g493
  (
    n577,
    n86
  );


  not
  g494
  (
    n235,
    n34
  );


  not
  g495
  (
    n399,
    n112
  );


  not
  g496
  (
    n411,
    n89
  );


  not
  g497
  (
    n349,
    n121
  );


  not
  g498
  (
    n516,
    n99
  );


  not
  g499
  (
    n265,
    n88
  );


  buf
  g500
  (
    n169,
    n88
  );


  not
  g501
  (
    n281,
    n35
  );


  not
  g502
  (
    n504,
    n36
  );


  buf
  g503
  (
    n479,
    n139
  );


  buf
  g504
  (
    n468,
    n53
  );


  not
  g505
  (
    n209,
    n94
  );


  buf
  g506
  (
    KeyWire_0_15,
    n93
  );


  not
  g507
  (
    n432,
    n37
  );


  not
  g508
  (
    n269,
    n74
  );


  not
  g509
  (
    n531,
    n90
  );


  not
  g510
  (
    n212,
    n106
  );


  buf
  g511
  (
    n540,
    n50
  );


  buf
  g512
  (
    n374,
    n119
  );


  not
  g513
  (
    n276,
    n42
  );


  buf
  g514
  (
    n258,
    n119
  );


  not
  g515
  (
    n315,
    n93
  );


  not
  g516
  (
    n341,
    n116
  );


  buf
  g517
  (
    n314,
    n42
  );


  buf
  g518
  (
    n413,
    n40
  );


  buf
  g519
  (
    n336,
    n104
  );


  not
  g520
  (
    n450,
    n37
  );


  buf
  g521
  (
    n495,
    n102
  );


  buf
  g522
  (
    n473,
    n76
  );


  buf
  g523
  (
    n270,
    n85
  );


  buf
  g524
  (
    n183,
    n82
  );


  buf
  g525
  (
    n448,
    n84
  );


  not
  g526
  (
    n482,
    n42
  );


  not
  g527
  (
    n354,
    n75
  );


  buf
  g528
  (
    n181,
    n123
  );


  buf
  g529
  (
    n533,
    n121
  );


  not
  g530
  (
    KeyWire_0_4,
    n75
  );


  not
  g531
  (
    n437,
    n130
  );


  not
  g532
  (
    n280,
    n59
  );


  buf
  g533
  (
    n389,
    n111
  );


  buf
  g534
  (
    n368,
    n118
  );


  not
  g535
  (
    n418,
    n100
  );


  not
  g536
  (
    n175,
    n64
  );


  buf
  g537
  (
    n362,
    n39
  );


  buf
  g538
  (
    n455,
    n49
  );


  not
  g539
  (
    n356,
    n100
  );


  buf
  g540
  (
    n457,
    n77
  );


  not
  g541
  (
    n481,
    n39
  );


  buf
  g542
  (
    n425,
    n72
  );


  not
  g543
  (
    n228,
    n62
  );


  not
  g544
  (
    n518,
    n92
  );


  not
  g545
  (
    n416,
    n58
  );


  buf
  g546
  (
    n558,
    n126
  );


  not
  g547
  (
    n472,
    n72
  );


  buf
  g548
  (
    n283,
    n116
  );


  not
  g549
  (
    n327,
    n115
  );


  buf
  g550
  (
    n305,
    n132
  );


  not
  g551
  (
    n517,
    n101
  );


  buf
  g552
  (
    n233,
    n70
  );


  buf
  g553
  (
    n422,
    n34
  );


  not
  g554
  (
    n303,
    n56
  );


  buf
  g555
  (
    n575,
    n58
  );


  not
  g556
  (
    n355,
    n41
  );


  not
  g557
  (
    n317,
    n38
  );


  not
  g558
  (
    n308,
    n90
  );


  not
  g559
  (
    n467,
    n120
  );


  buf
  g560
  (
    n524,
    n57
  );


  not
  g561
  (
    n344,
    n51
  );


  not
  g562
  (
    n161,
    n138
  );


  buf
  g563
  (
    n594,
    n97
  );


  buf
  g564
  (
    n469,
    n73
  );


  not
  g565
  (
    n426,
    n65
  );


  not
  g566
  (
    n361,
    n45
  );


  buf
  g567
  (
    n194,
    n65
  );


  not
  g568
  (
    n363,
    n84
  );


  not
  g569
  (
    n401,
    n80
  );


  buf
  g570
  (
    n589,
    n61
  );


  buf
  g571
  (
    n545,
    n138
  );


  or
  g572
  (
    n723,
    n429,
    n463,
    n301
  );


  nand
  g573
  (
    n657,
    n509,
    n435,
    n321,
    n394
  );


  nand
  g574
  (
    n648,
    n308,
    n425,
    n486,
    n402
  );


  or
  g575
  (
    n758,
    n306,
    n211,
    n491,
    n506
  );


  xor
  g576
  (
    n669,
    n173,
    n441,
    n397,
    n182
  );


  nor
  g577
  (
    n654,
    n373,
    n469,
    n482,
    n219
  );


  xor
  g578
  (
    n773,
    n443,
    n237,
    n435,
    n424
  );


  nand
  g579
  (
    n794,
    n292,
    n177,
    n496,
    n461
  );


  xor
  g580
  (
    n743,
    n244,
    n431,
    n473,
    n163
  );


  nor
  g581
  (
    n649,
    n456,
    n389,
    n439,
    n512
  );


  and
  g582
  (
    n746,
    n190,
    n481,
    n287,
    n386
  );


  xnor
  g583
  (
    n817,
    n269,
    n317,
    n283,
    n281
  );


  xor
  g584
  (
    n802,
    n283,
    n489,
    n192,
    n291
  );


  and
  g585
  (
    n719,
    n456,
    n462,
    n369,
    n227
  );


  xor
  g586
  (
    n781,
    n169,
    n466,
    n462,
    n473
  );


  nand
  g587
  (
    n697,
    n392,
    n360,
    n413,
    n340
  );


  and
  g588
  (
    n680,
    n377,
    n252,
    n502,
    n288
  );


  xnor
  g589
  (
    n606,
    n484,
    n490,
    n407,
    n355
  );


  nor
  g590
  (
    n608,
    n253,
    n313,
    n494,
    n183
  );


  xor
  g591
  (
    n644,
    n231,
    n272,
    n459,
    n486
  );


  xnor
  g592
  (
    n762,
    n477,
    n334,
    n332,
    n457
  );


  xor
  g593
  (
    n681,
    n302,
    n351,
    n496,
    n475
  );


  and
  g594
  (
    n779,
    n482,
    n420,
    n368,
    n293
  );


  and
  g595
  (
    n829,
    n455,
    n423,
    n337,
    n217
  );


  xor
  g596
  (
    n703,
    n187,
    n229,
    n352,
    n448
  );


  and
  g597
  (
    n733,
    n378,
    n236,
    n295,
    n491
  );


  xnor
  g598
  (
    n636,
    n275,
    n208,
    n501,
    n472
  );


  xor
  g599
  (
    n625,
    n161,
    n380,
    n409,
    n222
  );


  and
  g600
  (
    n801,
    n505,
    n451,
    n371,
    n329
  );


  or
  g601
  (
    n737,
    n444,
    n290,
    n195,
    n189
  );


  nor
  g602
  (
    n715,
    n226,
    n480,
    n443,
    n278
  );


  xnor
  g603
  (
    n691,
    n204,
    n235,
    n362,
    n477
  );


  xnor
  g604
  (
    n769,
    n486,
    n306,
    n352,
    n218
  );


  and
  g605
  (
    n672,
    n313,
    n499,
    n469,
    n430
  );


  xor
  g606
  (
    n694,
    n488,
    n224,
    n244,
    n240
  );


  nor
  g607
  (
    n675,
    n398,
    n350,
    n464,
    n357
  );


  or
  g608
  (
    n784,
    n233,
    n270,
    n164,
    n510
  );


  and
  g609
  (
    n765,
    n429,
    n314,
    n384,
    n441
  );


  xnor
  g610
  (
    n677,
    n309,
    n434,
    n257,
    n336
  );


  or
  g611
  (
    n740,
    n438,
    n221,
    n490,
    n256
  );


  nor
  g612
  (
    n771,
    n483,
    n232,
    n167,
    n425
  );


  xnor
  g613
  (
    n821,
    n431,
    n427,
    n429
  );


  or
  g614
  (
    n687,
    n500,
    n466,
    n268
  );


  and
  g615
  (
    n732,
    n382,
    n321,
    n379,
    n419
  );


  nor
  g616
  (
    n753,
    n225,
    n502,
    n309,
    n284
  );


  and
  g617
  (
    n652,
    n209,
    n231,
    n401,
    n348
  );


  xnor
  g618
  (
    n783,
    n375,
    n191,
    n172,
    n271
  );


  xor
  g619
  (
    n752,
    n397,
    n194,
    n359,
    n377
  );


  and
  g620
  (
    n676,
    n505,
    n364,
    n277,
    n356
  );


  or
  g621
  (
    n635,
    n276,
    n255,
    n180,
    n478
  );


  nor
  g622
  (
    n805,
    n189,
    n440,
    n323,
    n206
  );


  or
  g623
  (
    n734,
    n479,
    n433,
    n426,
    n467
  );


  and
  g624
  (
    n684,
    n495,
    n221,
    n478,
    n171
  );


  or
  g625
  (
    n639,
    n201,
    n296,
    n345,
    n480
  );


  nand
  g626
  (
    n710,
    n511,
    n251,
    n427,
    n510
  );


  nand
  g627
  (
    n695,
    n322,
    n353,
    n345,
    n432
  );


  and
  g628
  (
    n634,
    n497,
    n247,
    n512,
    n465
  );


  nand
  g629
  (
    n813,
    n273,
    n490,
    n365,
    n175
  );


  xnor
  g630
  (
    n623,
    n241,
    n302,
    n331,
    n494
  );


  xnor
  g631
  (
    n760,
    n476,
    n299,
    n346,
    n161
  );


  nor
  g632
  (
    n754,
    n490,
    n455,
    n475,
    n325
  );


  nor
  g633
  (
    n819,
    n260,
    n450,
    n480,
    n282
  );


  nand
  g634
  (
    n757,
    n232,
    n478,
    n485,
    n460
  );


  and
  g635
  (
    n727,
    n497,
    n230,
    n329,
    n513
  );


  nand
  g636
  (
    n828,
    n342,
    n477,
    n305,
    n396
  );


  nand
  g637
  (
    n830,
    n390,
    n205,
    n506,
    n388
  );


  and
  g638
  (
    n613,
    n453,
    n270,
    n228,
    n280
  );


  xnor
  g639
  (
    n622,
    n420,
    n238,
    n259,
    n193
  );


  or
  g640
  (
    n647,
    n165,
    n516,
    n445,
    n441
  );


  nor
  g641
  (
    n739,
    n470,
    n271,
    n205,
    n353
  );


  or
  g642
  (
    n748,
    n466,
    n421,
    n243,
    n199
  );


  nand
  g643
  (
    n797,
    n375,
    n163,
    n310,
    n444
  );


  xnor
  g644
  (
    n706,
    n404,
    n168,
    n444,
    n423
  );


  xnor
  g645
  (
    n643,
    n391,
    n303,
    n509,
    n181
  );


  nand
  g646
  (
    n713,
    n432,
    n426,
    n338,
    n340
  );


  and
  g647
  (
    n731,
    n434,
    n437,
    n248,
    n450
  );


  or
  g648
  (
    n640,
    n301,
    n492,
    n502,
    n463
  );


  or
  g649
  (
    n621,
    n452,
    n167,
    n499,
    n430
  );


  and
  g650
  (
    n673,
    n367,
    n458,
    n438,
    n428
  );


  and
  g651
  (
    n627,
    n489,
    n330,
    n445,
    n472
  );


  nand
  g652
  (
    n764,
    n516,
    n194,
    n405,
    n505
  );


  and
  g653
  (
    n607,
    n433,
    n487,
    n366,
    n214
  );


  nor
  g654
  (
    n655,
    n243,
    n237,
    n442,
    n404
  );


  xnor
  g655
  (
    n612,
    n509,
    n223,
    n166,
    n380
  );


  or
  g656
  (
    n626,
    n260,
    n394,
    n446,
    n425
  );


  xnor
  g657
  (
    n632,
    n464,
    n477,
    n453,
    n432
  );


  or
  g658
  (
    n741,
    n470,
    n355,
    n344,
    n334
  );


  xor
  g659
  (
    n756,
    n391,
    n416,
    n246,
    n227
  );


  nor
  g660
  (
    n616,
    n277,
    n495,
    n335,
    n200
  );


  nor
  g661
  (
    n660,
    n467,
    n435,
    n387,
    n230
  );


  nand
  g662
  (
    n708,
    n482,
    n204,
    n365,
    n470
  );


  nand
  g663
  (
    n716,
    n443,
    n343,
    n492,
    n308
  );


  or
  g664
  (
    n714,
    n311,
    n318,
    n458,
    n368
  );


  nand
  g665
  (
    n815,
    n206,
    n165,
    n411,
    n481
  );


  nand
  g666
  (
    n688,
    n326,
    n278,
    n236,
    n258
  );


  nor
  g667
  (
    n689,
    n422,
    n460,
    n428,
    n386
  );


  xnor
  g668
  (
    n637,
    n182,
    n359,
    n468,
    n174
  );


  xnor
  g669
  (
    n768,
    n219,
    n281,
    n430,
    n506
  );


  nor
  g670
  (
    n738,
    n446,
    n513,
    n266,
    n459
  );


  nand
  g671
  (
    n790,
    n257,
    n500,
    n515,
    n440
  );


  nor
  g672
  (
    n717,
    n181,
    n298,
    n456,
    n258
  );


  xnor
  g673
  (
    n659,
    n427,
    n200,
    n421,
    n472
  );


  nor
  g674
  (
    n642,
    n263,
    n515,
    n508,
    n512
  );


  nand
  g675
  (
    n702,
    n289,
    n216,
    n264,
    n383
  );


  and
  g676
  (
    n776,
    n435,
    n197,
    n453,
    n272
  );


  nand
  g677
  (
    n811,
    n363,
    n209,
    n249,
    n479
  );


  nand
  g678
  (
    n605,
    n254,
    n499,
    n255,
    n485
  );


  nor
  g679
  (
    n651,
    n438,
    n436,
    n212,
    n275
  );


  xor
  g680
  (
    n772,
    n176,
    n420,
    n322,
    n405
  );


  nand
  g681
  (
    n810,
    n389,
    n487,
    n201,
    n315
  );


  and
  g682
  (
    n711,
    n354,
    n274,
    n216,
    n318
  );


  xnor
  g683
  (
    n728,
    n366,
    n415,
    n417,
    n333
  );


  nand
  g684
  (
    n679,
    n388,
    n480,
    n408,
    n465
  );


  nor
  g685
  (
    n777,
    n511,
    n464,
    n177,
    n172
  );


  and
  g686
  (
    n825,
    n436,
    n482,
    n514,
    n190
  );


  nor
  g687
  (
    n709,
    n516,
    n487,
    n210,
    n517
  );


  nand
  g688
  (
    n698,
    n460,
    n483,
    n414,
    n290
  );


  xor
  g689
  (
    n742,
    n385,
    n469,
    n421,
    n418
  );


  xnor
  g690
  (
    n724,
    n498,
    n344,
    n468,
    n423
  );


  xor
  g691
  (
    n618,
    n510,
    n358,
    n268,
    n500
  );


  nand
  g692
  (
    n619,
    n374,
    n507,
    n434,
    n360
  );


  nand
  g693
  (
    n662,
    n178,
    n501,
    n491,
    n472
  );


  xor
  g694
  (
    n786,
    n516,
    n486,
    n246,
    n446
  );


  xor
  g695
  (
    n796,
    n434,
    n447,
    n325,
    n351
  );


  and
  g696
  (
    n683,
    n469,
    n349,
    n176,
    n442
  );


  nand
  g697
  (
    n668,
    n406,
    n501,
    n503,
    n245
  );


  and
  g698
  (
    n670,
    n393,
    n327,
    n187,
    n479
  );


  nand
  g699
  (
    n791,
    n331,
    n256,
    n417,
    n479
  );


  xor
  g700
  (
    n827,
    n288,
    n304,
    n504,
    n509
  );


  nand
  g701
  (
    n751,
    n287,
    n422,
    n448,
    n261
  );


  xor
  g702
  (
    n653,
    n447,
    n467,
    n396,
    n511
  );


  nand
  g703
  (
    n614,
    n174,
    n173,
    n382,
    n398
  );


  or
  g704
  (
    n658,
    n491,
    n197,
    n166,
    n319
  );


  xor
  g705
  (
    n744,
    n385,
    n317,
    n493,
    n485
  );


  xnor
  g706
  (
    n822,
    n274,
    n357,
    n441,
    n507
  );


  nor
  g707
  (
    n712,
    n412,
    n481,
    n499,
    n310
  );


  and
  g708
  (
    n816,
    n449,
    n238,
    n410,
    n300
  );


  nand
  g709
  (
    n814,
    n436,
    n492,
    n363,
    n514
  );


  nand
  g710
  (
    n818,
    n451,
    n196,
    n285,
    n316
  );


  nand
  g711
  (
    n630,
    n431,
    n376,
    n356,
    n170
  );


  xor
  g712
  (
    n770,
    n303,
    n400,
    n367,
    n376
  );


  and
  g713
  (
    n785,
    n419,
    n431,
    n286,
    n458
  );


  nor
  g714
  (
    n665,
    n293,
    n320,
    n426,
    n245
  );


  xor
  g715
  (
    n803,
    n488,
    n384,
    n207,
    n467
  );


  xnor
  g716
  (
    n656,
    n178,
    n439,
    n484,
    n423
  );


  nand
  g717
  (
    n725,
    n478,
    n320,
    n470,
    n461
  );


  nor
  g718
  (
    n792,
    n195,
    n415,
    n358,
    n259
  );


  and
  g719
  (
    n699,
    n285,
    n399,
    n437,
    n186
  );


  xor
  g720
  (
    n823,
    n503,
    n198,
    n327,
    n312
  );


  xnor
  g721
  (
    n617,
    n484,
    n450,
    n280,
    n267
  );


  nand
  g722
  (
    n800,
    n489,
    n207,
    n433,
    n507
  );


  xor
  g723
  (
    n678,
    n262,
    n324,
    n248,
    n212
  );


  nor
  g724
  (
    n826,
    n462,
    n495,
    n454,
    n349
  );


  nand
  g725
  (
    n641,
    n251,
    n433,
    n370,
    n371
  );


  and
  g726
  (
    n686,
    n229,
    n454,
    n292,
    n408
  );


  xnor
  g727
  (
    n736,
    n461,
    n426,
    n250,
    n503
  );


  nor
  g728
  (
    n664,
    n193,
    n455,
    n456,
    n319
  );


  xor
  g729
  (
    n798,
    n474,
    n462,
    n339,
    n203
  );


  xnor
  g730
  (
    n745,
    n468,
    n179,
    n224,
    n502
  );


  and
  g731
  (
    n735,
    n202,
    n364,
    n164,
    n497
  );


  nand
  g732
  (
    n750,
    n341,
    n457,
    n299,
    n465
  );


  and
  g733
  (
    n759,
    n316,
    n381,
    n493,
    n439
  );


  nor
  g734
  (
    n628,
    n413,
    n346,
    n452,
    n422
  );


  and
  g735
  (
    n761,
    n504,
    n253,
    n184,
    n330
  );


  and
  g736
  (
    n615,
    n458,
    n372,
    n354,
    n191
  );


  and
  g737
  (
    n718,
    n362,
    n341,
    n473,
    n261
  );


  nand
  g738
  (
    n806,
    n234,
    n215,
    n179,
    n185
  );


  and
  g739
  (
    n730,
    n504,
    n410,
    n279,
    n196
  );


  xnor
  g740
  (
    n690,
    n399,
    n447,
    n387,
    n381
  );


  nand
  g741
  (
    n629,
    n373,
    n188,
    n291,
    n202
  );


  and
  g742
  (
    n767,
    n184,
    n484,
    n265,
    n448
  );


  nand
  g743
  (
    n766,
    n213,
    n378,
    n315,
    n298
  );


  xnor
  g744
  (
    n778,
    n452,
    n436,
    n493,
    n483
  );


  xor
  g745
  (
    n682,
    n403,
    n214,
    n432,
    n464
  );


  or
  g746
  (
    n804,
    n474,
    n447,
    n223,
    n180
  );


  xor
  g747
  (
    n722,
    n407,
    n443,
    n300,
    n333
  );


  nand
  g748
  (
    n747,
    n513,
    n342,
    n250,
    n425
  );


  nor
  g749
  (
    n704,
    n505,
    n449,
    n471
  );


  nor
  g750
  (
    n696,
    n335,
    n235,
    n361,
    n294
  );


  xor
  g751
  (
    n749,
    n295,
    n463,
    n428,
    n488
  );


  nand
  g752
  (
    n808,
    n211,
    n323,
    n461,
    n406
  );


  xor
  g753
  (
    n820,
    n361,
    n328,
    n437,
    n489
  );


  xnor
  g754
  (
    n787,
    n459,
    n448,
    n452,
    n485
  );


  nor
  g755
  (
    n795,
    n504,
    n481,
    n515,
    n487
  );


  xnor
  g756
  (
    n782,
    n242,
    n175,
    n226,
    n494
  );


  nor
  g757
  (
    n812,
    n463,
    n446,
    n289,
    n263
  );


  xnor
  g758
  (
    n807,
    n508,
    n471,
    n169,
    n424
  );


  xor
  g759
  (
    n793,
    n401,
    n498,
    n304,
    n428
  );


  xnor
  g760
  (
    n707,
    n409,
    n339,
    n225,
    n369
  );


  nor
  g761
  (
    n663,
    n338,
    n379,
    n474,
    n513
  );


  xnor
  g762
  (
    n646,
    n228,
    n328,
    n395,
    n450
  );


  and
  g763
  (
    n620,
    n514,
    n455,
    n424,
    n475
  );


  nand
  g764
  (
    n705,
    n451,
    n213,
    n222,
    n297
  );


  xnor
  g765
  (
    n775,
    n170,
    n252,
    n459,
    n465
  );


  nor
  g766
  (
    n789,
    n449,
    n497,
    n420,
    n442
  );


  xnor
  g767
  (
    n650,
    n239,
    n162,
    n508
  );


  nand
  g768
  (
    n755,
    n383,
    n188,
    n422,
    n307
  );


  and
  g769
  (
    n609,
    n370,
    n412,
    n162,
    n475
  );


  or
  g770
  (
    n729,
    n421,
    n424,
    n454,
    n500
  );


  xor
  g771
  (
    n700,
    n473,
    n395,
    n449,
    n418
  );


  nand
  g772
  (
    n667,
    n269,
    n324,
    n296,
    n501
  );


  nor
  g773
  (
    n661,
    n314,
    n239,
    n186,
    n311
  );


  nor
  g774
  (
    n809,
    n198,
    n471,
    n220,
    n265
  );


  xnor
  g775
  (
    n721,
    n512,
    n168,
    n474,
    n337
  );


  nand
  g776
  (
    n726,
    n254,
    n392,
    n240,
    n468
  );


  and
  g777
  (
    n693,
    n411,
    n429,
    n483,
    n390
  );


  nand
  g778
  (
    n633,
    n247,
    n348,
    n297,
    n457
  );


  xnor
  g779
  (
    n624,
    n444,
    n506,
    n438,
    n445
  );


  xnor
  g780
  (
    n788,
    n305,
    n440,
    n350,
    n220
  );


  nand
  g781
  (
    n720,
    n403,
    n234,
    n374,
    n286
  );


  or
  g782
  (
    n638,
    n476,
    n498,
    n336,
    n233
  );


  nand
  g783
  (
    n611,
    n332,
    n307,
    n241,
    n203
  );


  and
  g784
  (
    n799,
    n312,
    n445,
    n266,
    n273
  );


  or
  g785
  (
    n774,
    n199,
    n457,
    n498,
    n393
  );


  and
  g786
  (
    n701,
    n215,
    n453,
    n262,
    n343
  );


  nand
  g787
  (
    n692,
    n171,
    n454,
    n451,
    n294
  );


  xnor
  g788
  (
    n763,
    n442,
    n264,
    n511,
    n488
  );


  nand
  g789
  (
    n824,
    n210,
    n496,
    n494,
    n218
  );


  nand
  g790
  (
    n610,
    n439,
    n372,
    n185,
    n440
  );


  and
  g791
  (
    n631,
    n514,
    n242,
    n276,
    n416
  );


  xnor
  g792
  (
    n780,
    n495,
    n476,
    n510,
    n267
  );


  xor
  g793
  (
    n671,
    n460,
    n284,
    n192,
    n496
  );


  or
  g794
  (
    n831,
    n279,
    n476,
    n183,
    n493
  );


  xor
  g795
  (
    n645,
    n503,
    n414,
    n217,
    n402
  );


  xnor
  g796
  (
    n685,
    n492,
    n347,
    n437,
    n507
  );


  and
  g797
  (
    n674,
    n208,
    n515,
    n347,
    n249
  );


  xnor
  g798
  (
    n666,
    n282,
    n400,
    n326,
    n430
  );


  buf
  g799
  (
    n975,
    n726
  );


  not
  g800
  (
    n951,
    n631
  );


  buf
  g801
  (
    n846,
    n618
  );


  not
  g802
  (
    n960,
    n684
  );


  buf
  g803
  (
    n832,
    n664
  );


  buf
  g804
  (
    n946,
    n722
  );


  buf
  g805
  (
    n947,
    n672
  );


  not
  g806
  (
    n838,
    n725
  );


  buf
  g807
  (
    n861,
    n698
  );


  buf
  g808
  (
    n866,
    n682
  );


  buf
  g809
  (
    n964,
    n715
  );


  buf
  g810
  (
    n987,
    n712
  );


  not
  g811
  (
    n965,
    n731
  );


  not
  g812
  (
    n952,
    n692
  );


  not
  g813
  (
    n855,
    n727
  );


  buf
  g814
  (
    n985,
    n706
  );


  not
  g815
  (
    n915,
    n693
  );


  not
  g816
  (
    n981,
    n681
  );


  not
  g817
  (
    n843,
    n757
  );


  buf
  g818
  (
    n957,
    n759
  );


  buf
  g819
  (
    n863,
    n763
  );


  buf
  g820
  (
    n848,
    n630
  );


  buf
  g821
  (
    n894,
    n653
  );


  buf
  g822
  (
    n833,
    n708
  );


  buf
  g823
  (
    n890,
    n730
  );


  buf
  g824
  (
    n953,
    n654
  );


  not
  g825
  (
    n928,
    n639
  );


  not
  g826
  (
    n884,
    n754
  );


  not
  g827
  (
    n922,
    n641
  );


  buf
  g828
  (
    n895,
    n709
  );


  buf
  g829
  (
    n902,
    n766
  );


  not
  g830
  (
    n954,
    n700
  );


  buf
  g831
  (
    n857,
    n689
  );


  buf
  g832
  (
    n977,
    n616
  );


  not
  g833
  (
    n993,
    n674
  );


  buf
  g834
  (
    n844,
    n749
  );


  buf
  g835
  (
    n925,
    n733
  );


  not
  g836
  (
    n913,
    n751
  );


  buf
  g837
  (
    n882,
    n736
  );


  buf
  g838
  (
    n865,
    n624
  );


  buf
  g839
  (
    n892,
    n694
  );


  not
  g840
  (
    n942,
    n613
  );


  not
  g841
  (
    n962,
    n655
  );


  not
  g842
  (
    n905,
    n720
  );


  buf
  g843
  (
    n917,
    n739
  );


  not
  g844
  (
    n986,
    n638
  );


  not
  g845
  (
    n883,
    n728
  );


  not
  g846
  (
    n907,
    n611
  );


  buf
  g847
  (
    n968,
    n617
  );


  not
  g848
  (
    n897,
    n647
  );


  not
  g849
  (
    n926,
    n633
  );


  buf
  g850
  (
    n851,
    n605
  );


  buf
  g851
  (
    n896,
    n711
  );


  buf
  g852
  (
    n860,
    n635
  );


  not
  g853
  (
    n856,
    n768
  );


  buf
  g854
  (
    n958,
    n666
  );


  not
  g855
  (
    n910,
    n701
  );


  not
  g856
  (
    n839,
    n756
  );


  not
  g857
  (
    n927,
    n656
  );


  buf
  g858
  (
    n978,
    n690
  );


  not
  g859
  (
    n850,
    n743
  );


  not
  g860
  (
    n867,
    n634
  );


  not
  g861
  (
    n837,
    n683
  );


  not
  g862
  (
    n912,
    n627
  );


  not
  g863
  (
    n973,
    n762
  );


  not
  g864
  (
    n885,
    n719
  );


  buf
  g865
  (
    n944,
    n608
  );


  not
  g866
  (
    n936,
    n614
  );


  buf
  g867
  (
    n983,
    n680
  );


  not
  g868
  (
    n966,
    n676
  );


  buf
  g869
  (
    n924,
    n662
  );


  buf
  g870
  (
    n916,
    n665
  );


  buf
  g871
  (
    n934,
    n644
  );


  buf
  g872
  (
    n904,
    n622
  );


  not
  g873
  (
    n845,
    n688
  );


  not
  g874
  (
    n963,
    n671
  );


  buf
  g875
  (
    n971,
    n695
  );


  buf
  g876
  (
    KeyWire_0_10,
    n612
  );


  not
  g877
  (
    n906,
    n729
  );


  not
  g878
  (
    n911,
    n747
  );


  buf
  g879
  (
    n972,
    n761
  );


  buf
  g880
  (
    n950,
    n748
  );


  buf
  g881
  (
    n872,
    n667
  );


  buf
  g882
  (
    n874,
    n691
  );


  not
  g883
  (
    n852,
    n752
  );


  buf
  g884
  (
    n938,
    n621
  );


  not
  g885
  (
    n877,
    n610
  );


  not
  g886
  (
    n976,
    n742
  );


  not
  g887
  (
    n841,
    n663
  );


  buf
  g888
  (
    n945,
    n625
  );


  not
  g889
  (
    n868,
    n760
  );


  buf
  g890
  (
    n888,
    n696
  );


  not
  g891
  (
    n920,
    n703
  );


  not
  g892
  (
    n967,
    n744
  );


  buf
  g893
  (
    n956,
    n746
  );


  buf
  g894
  (
    n876,
    n705
  );


  buf
  g895
  (
    n991,
    n737
  );


  not
  g896
  (
    n919,
    n714
  );


  not
  g897
  (
    n994,
    n649
  );


  not
  g898
  (
    n900,
    n687
  );


  not
  g899
  (
    n990,
    n673
  );


  buf
  g900
  (
    n840,
    n738
  );


  not
  g901
  (
    n870,
    n661
  );


  buf
  g902
  (
    n988,
    n628
  );


  not
  g903
  (
    n887,
    n741
  );


  buf
  g904
  (
    n881,
    n753
  );


  not
  g905
  (
    n899,
    n619
  );


  not
  g906
  (
    n889,
    n745
  );


  buf
  g907
  (
    n979,
    n629
  );


  buf
  g908
  (
    n923,
    n721
  );


  buf
  g909
  (
    n992,
    n607
  );


  not
  g910
  (
    n940,
    n697
  );


  buf
  g911
  (
    n937,
    n713
  );


  not
  g912
  (
    n969,
    n620
  );


  buf
  g913
  (
    n918,
    n660
  );


  buf
  g914
  (
    n873,
    n626
  );


  buf
  g915
  (
    n871,
    n652
  );


  buf
  g916
  (
    KeyWire_0_8,
    n686
  );


  buf
  g917
  (
    n980,
    n716
  );


  not
  g918
  (
    n995,
    n640
  );


  not
  g919
  (
    n869,
    n717
  );


  buf
  g920
  (
    n835,
    n710
  );


  buf
  g921
  (
    n974,
    n609
  );


  buf
  g922
  (
    n921,
    n637
  );


  not
  g923
  (
    n879,
    n767
  );


  buf
  g924
  (
    n903,
    n636
  );


  buf
  g925
  (
    n909,
    n732
  );


  buf
  g926
  (
    n984,
    n704
  );


  buf
  g927
  (
    n931,
    n648
  );


  not
  g928
  (
    n961,
    n678
  );


  buf
  g929
  (
    n935,
    n724
  );


  buf
  g930
  (
    n875,
    n623
  );


  buf
  g931
  (
    n949,
    n642
  );


  not
  g932
  (
    n955,
    n669
  );


  buf
  g933
  (
    n941,
    n679
  );


  buf
  g934
  (
    n948,
    n650
  );


  not
  g935
  (
    n878,
    n657
  );


  not
  g936
  (
    n854,
    n677
  );


  buf
  g937
  (
    n989,
    n615
  );


  not
  g938
  (
    n970,
    n723
  );


  buf
  g939
  (
    n836,
    n658
  );


  not
  g940
  (
    n849,
    n659
  );


  not
  g941
  (
    n842,
    n764
  );


  buf
  g942
  (
    n908,
    n668
  );


  buf
  g943
  (
    n959,
    n707
  );


  buf
  g944
  (
    n859,
    n755
  );


  not
  g945
  (
    n898,
    n702
  );


  buf
  g946
  (
    n982,
    n718
  );


  not
  g947
  (
    n891,
    n765
  );


  buf
  g948
  (
    n929,
    n734
  );


  buf
  g949
  (
    n930,
    n646
  );


  buf
  g950
  (
    n939,
    n675
  );


  buf
  g951
  (
    n901,
    n632
  );


  buf
  g952
  (
    n853,
    n740
  );


  buf
  g953
  (
    n932,
    n606
  );


  not
  g954
  (
    n858,
    n645
  );


  buf
  g955
  (
    n834,
    n758
  );


  not
  g956
  (
    n914,
    n735
  );


  not
  g957
  (
    KeyWire_0_13,
    n685
  );


  buf
  g958
  (
    n862,
    n699
  );


  buf
  g959
  (
    n886,
    n643
  );


  not
  g960
  (
    n943,
    n750
  );


  buf
  g961
  (
    n847,
    n651
  );


  buf
  g962
  (
    n864,
    n670
  );


  xnor
  g963
  (
    n998,
    n942,
    n920,
    n944,
    n872
  );


  xor
  g964
  (
    n1018,
    n876,
    n917,
    n937,
    n939
  );


  and
  g965
  (
    n1017,
    n945,
    n921,
    n836,
    n839
  );


  nor
  g966
  (
    n1006,
    n855,
    n854,
    n936,
    n911
  );


  xnor
  g967
  (
    n1020,
    n931,
    n893,
    n939,
    n849
  );


  nor
  g968
  (
    n996,
    n916,
    n934,
    n889,
    n857
  );


  and
  g969
  (
    n1014,
    n840,
    n909,
    n878,
    n846
  );


  nand
  g970
  (
    n1025,
    n924,
    n864,
    n908,
    n926
  );


  or
  g971
  (
    n1002,
    n938,
    n873,
    n928,
    n847
  );


  nor
  g972
  (
    n1015,
    n890,
    n944,
    n943,
    n912
  );


  or
  g973
  (
    n1022,
    n856,
    n841,
    n892,
    n922
  );


  nor
  g974
  (
    KeyWire_0_2,
    n930,
    n903,
    n935,
    n845
  );


  and
  g975
  (
    n1011,
    n858,
    n877,
    n844,
    n894
  );


  nor
  g976
  (
    n1003,
    n866,
    n843,
    n941,
    n923
  );


  xnor
  g977
  (
    n999,
    n902,
    n925,
    n833,
    n898
  );


  xnor
  g978
  (
    n1000,
    n883,
    n914,
    n863,
    n927
  );


  nand
  g979
  (
    n1001,
    n940,
    n901,
    n941,
    n834
  );


  nand
  g980
  (
    n1023,
    n888,
    n904,
    n870,
    n862
  );


  xnor
  g981
  (
    n997,
    n907,
    n865,
    n940,
    n837
  );


  xnor
  g982
  (
    n1010,
    n942,
    n886,
    n853,
    n881
  );


  nand
  g983
  (
    n1016,
    n842,
    n933,
    n896,
    n943
  );


  xor
  g984
  (
    n1005,
    n875,
    n860,
    n913,
    n885
  );


  xnor
  g985
  (
    n1012,
    n867,
    n906,
    n891,
    n838
  );


  xnor
  g986
  (
    n1024,
    n850,
    n887,
    n874,
    n915
  );


  nand
  g987
  (
    n1021,
    n868,
    n859,
    n897,
    n932
  );


  or
  g988
  (
    n1013,
    n879,
    n918,
    n919,
    n852
  );


  xnor
  g989
  (
    n1007,
    n832,
    n884,
    n848,
    n882
  );


  and
  g990
  (
    n1019,
    n851,
    n929,
    n861,
    n871
  );


  nand
  g991
  (
    n1004,
    n905,
    n900,
    n910,
    n899
  );


  and
  g992
  (
    n1008,
    n835,
    n895,
    n880,
    n869
  );


  not
  g993
  (
    n1026,
    n1025
  );


  buf
  g994
  (
    n1028,
    n1022
  );


  not
  g995
  (
    n1029,
    n1024
  );


  not
  g996
  (
    n1027,
    n1023
  );


  xor
  g997
  (
    n1036,
    n1027,
    n520,
    n1028,
    n521
  );


  xor
  g998
  (
    n1041,
    n525,
    n525,
    n522,
    n519
  );


  or
  g999
  (
    n1035,
    n520,
    n1027,
    n519,
    n1026
  );


  nand
  g1000
  (
    n1038,
    n521,
    n523,
    n520
  );


  xnor
  g1001
  (
    n1031,
    n1026,
    n517,
    n522,
    n524
  );


  or
  g1002
  (
    n1033,
    n1028,
    n518,
    n525
  );


  and
  g1003
  (
    n1030,
    n1027,
    n519,
    n1028
  );


  nor
  g1004
  (
    n1032,
    n524,
    n523
  );


  xnor
  g1005
  (
    n1040,
    n1026,
    n521,
    n520,
    n1027
  );


  and
  g1006
  (
    n1034,
    n517,
    n521,
    n1026,
    n519
  );


  xor
  g1007
  (
    n1039,
    n517,
    n522,
    n524
  );


  xnor
  g1008
  (
    n1037,
    n526,
    n518,
    n525
  );


  not
  g1009
  (
    n1042,
    n1031
  );


  buf
  g1010
  (
    n1046,
    n1031
  );


  not
  g1011
  (
    n1045,
    n1031
  );


  buf
  g1012
  (
    n1044,
    n1030
  );


  buf
  g1013
  (
    n1043,
    n1030
  );


  buf
  g1014
  (
    n1047,
    n1043
  );


  not
  g1015
  (
    n1049,
    n1043
  );


  not
  g1016
  (
    n1048,
    n1042
  );


  not
  g1017
  (
    n1050,
    n1042
  );


  not
  g1018
  (
    n1052,
    n527
  );


  not
  g1019
  (
    n1054,
    n1049
  );


  or
  g1020
  (
    n1055,
    n147,
    n1050
  );


  nor
  g1021
  (
    n1053,
    n1050,
    n1047,
    n148
  );


  and
  g1022
  (
    n1064,
    n147,
    n526,
    n151,
    n146
  );


  xnor
  g1023
  (
    n1059,
    n1049,
    n1048
  );


  xor
  g1024
  (
    n1061,
    n151,
    n526,
    n146,
    n149
  );


  and
  g1025
  (
    n1057,
    n144,
    n150,
    n146
  );


  and
  g1026
  (
    n1062,
    n144,
    n1049,
    n527,
    n1050
  );


  and
  g1027
  (
    n1065,
    n149,
    n145,
    n151,
    n1048
  );


  nor
  g1028
  (
    n1051,
    n147,
    n148,
    n149,
    n150
  );


  or
  g1029
  (
    n1060,
    n145,
    n147,
    n144,
    n148
  );


  xnor
  g1030
  (
    n1058,
    n144,
    n151,
    n145,
    n150
  );


  xor
  g1031
  (
    n1056,
    n1048,
    n1047,
    n149
  );


  and
  g1032
  (
    n1063,
    n150,
    n145,
    n148,
    n526
  );


  not
  g1033
  (
    n1081,
    n530
  );


  buf
  g1034
  (
    n1076,
    n1054
  );


  not
  g1035
  (
    n1071,
    n1052
  );


  not
  g1036
  (
    n1067,
    n529
  );


  not
  g1037
  (
    n1082,
    n1055
  );


  buf
  g1038
  (
    n1084,
    n532
  );


  buf
  g1039
  (
    n1066,
    n529
  );


  not
  g1040
  (
    n1078,
    n531
  );


  not
  g1041
  (
    n1074,
    n529
  );


  buf
  g1042
  (
    n1083,
    n531
  );


  not
  g1043
  (
    n1072,
    n1052
  );


  buf
  g1044
  (
    n1085,
    n1051
  );


  buf
  g1045
  (
    n1068,
    n527
  );


  or
  g1046
  (
    n1069,
    n531,
    n532,
    n530
  );


  nand
  g1047
  (
    n1070,
    n1053,
    n1054,
    n1055
  );


  nor
  g1048
  (
    n1075,
    n529,
    n1052,
    n1051,
    n530
  );


  and
  g1049
  (
    n1080,
    n528,
    n528,
    n1052,
    n1053
  );


  nor
  g1050
  (
    n1077,
    n1053,
    n1055,
    n527,
    n531
  );


  and
  g1051
  (
    n1073,
    n530,
    n528,
    n1051
  );


  nor
  g1052
  (
    n1079,
    n1053,
    n1054,
    n528,
    n1055
  );


  nor
  g1053
  (
    n1089,
    n1072,
    n798,
    n785,
    n776
  );


  nor
  g1054
  (
    n1092,
    n773,
    n787,
    n780,
    n1067
  );


  nor
  g1055
  (
    n1090,
    n788,
    n796,
    n791,
    n775
  );


  or
  g1056
  (
    n1094,
    n792,
    n774,
    n786,
    n793
  );


  xnor
  g1057
  (
    n1093,
    n784,
    n772,
    n1070,
    n790
  );


  xor
  g1058
  (
    n1095,
    n777,
    n1071,
    n783,
    n782
  );


  xor
  g1059
  (
    n1088,
    n1066,
    n778,
    n771,
    n789
  );


  nand
  g1060
  (
    n1087,
    n1069,
    n1070,
    n797,
    n781
  );


  xnor
  g1061
  (
    n1091,
    n1072,
    n770,
    n779,
    n794
  );


  xnor
  g1062
  (
    n1086,
    n1071,
    n769,
    n795,
    n1068
  );


  nand
  g1063
  (
    n1097,
    n951,
    n947,
    n948,
    n954
  );


  xor
  g1064
  (
    n1098,
    n949,
    n955,
    n1092,
    n947
  );


  xnor
  g1065
  (
    n1101,
    n952,
    n1095,
    n950,
    n948
  );


  xnor
  g1066
  (
    n1102,
    n951,
    n1094,
    n953,
    n1091
  );


  nor
  g1067
  (
    n1096,
    n945,
    n946,
    n950
  );


  xnor
  g1068
  (
    n1100,
    n954,
    n1089,
    n953,
    n1093
  );


  nor
  g1069
  (
    n1099,
    n949,
    n1090,
    n955,
    n952
  );


  xor
  g1070
  (
    n1105,
    n1101,
    n532,
    n956,
    n958
  );


  xor
  g1071
  (
    n1103,
    n533,
    n958,
    n1100,
    n532
  );


  and
  g1072
  (
    n1104,
    n1102,
    n956,
    n957
  );


  nor
  g1073
  (
    n1106,
    n960,
    n152,
    n1104
  );


  xor
  g1074
  (
    n1107,
    n960,
    n1103,
    n959
  );


  buf
  g1075
  (
    n1110,
    n1107
  );


  buf
  g1076
  (
    n1108,
    n533
  );


  nor
  g1077
  (
    n1109,
    n533,
    n533,
    n1107,
    n1106
  );


  or
  g1078
  (
    n1112,
    n1109,
    n1044,
    n534
  );


  nand
  g1079
  (
    n1111,
    n1108,
    n1110,
    n806
  );


  nor
  g1080
  (
    n1113,
    n799,
    n802,
    n804,
    n803
  );


  nor
  g1081
  (
    n1114,
    n800,
    n805,
    n801,
    n1044
  );


  and
  g1082
  (
    n1117,
    n154,
    n153,
    n1114,
    n155
  );


  nor
  g1083
  (
    n1116,
    n1112,
    n1113,
    n152,
    n153
  );


  or
  g1084
  (
    n1118,
    n154,
    n153,
    n152
  );


  nor
  g1085
  (
    n1115,
    n154,
    n154,
    n1111,
    n155
  );


  xnor
  g1086
  (
    n1130,
    n538,
    n536,
    n540
  );


  and
  g1087
  (
    n1121,
    n1117,
    n541,
    n542
  );


  or
  g1088
  (
    n1129,
    n538,
    n535,
    n539
  );


  nor
  g1089
  (
    n1120,
    n539,
    n540
  );


  xor
  g1090
  (
    n1134,
    n1115,
    n1117,
    n537
  );


  xnor
  g1091
  (
    n1119,
    n537,
    n1118,
    n541
  );


  nand
  g1092
  (
    n1122,
    n543,
    n1115
  );


  nand
  g1093
  (
    n1124,
    n542,
    n1116,
    n535
  );


  xor
  g1094
  (
    n1128,
    n537,
    n540,
    n1117
  );


  or
  g1095
  (
    n1127,
    n1118,
    n1116,
    n537
  );


  or
  g1096
  (
    KeyWire_0_9,
    n1117,
    n1115,
    n536
  );


  xor
  g1097
  (
    n1123,
    n542,
    n1116,
    n538
  );


  nor
  g1098
  (
    n1131,
    n1118,
    n534,
    n1116,
    n536
  );


  nand
  g1099
  (
    n1132,
    n535,
    n536,
    n1118,
    n539
  );


  and
  g1100
  (
    n1133,
    n539,
    n538,
    n541
  );


  xor
  g1101
  (
    n1125,
    n535,
    n542,
    n534
  );


  and
  g1102
  (
    n1194,
    n576,
    n590,
    n585,
    n1131
  );


  or
  g1103
  (
    n1171,
    n558,
    n567,
    n585,
    n584
  );


  nor
  g1104
  (
    n1160,
    n1129,
    n1120,
    n1128,
    n1130
  );


  xor
  g1105
  (
    n1142,
    n566,
    n582,
    n585,
    n571
  );


  or
  g1106
  (
    n1144,
    n589,
    n565,
    n553,
    n1121
  );


  or
  g1107
  (
    n1186,
    n548,
    n581,
    n1134,
    n574
  );


  nand
  g1108
  (
    n1197,
    n550,
    n1127,
    n1123,
    n568
  );


  xor
  g1109
  (
    n1158,
    n549,
    n557,
    n566,
    n587
  );


  xor
  g1110
  (
    n1179,
    n1123,
    n1127,
    n571,
    n546
  );


  nand
  g1111
  (
    n1147,
    n553,
    n1131,
    n548,
    n582
  );


  nand
  g1112
  (
    n1176,
    n1123,
    n558,
    n580,
    n573
  );


  and
  g1113
  (
    n1174,
    n1126,
    n589,
    n563,
    n558
  );


  nand
  g1114
  (
    n1165,
    n578,
    n1130,
    n587,
    n545
  );


  xnor
  g1115
  (
    n1190,
    n561,
    n564,
    n563,
    n554
  );


  nand
  g1116
  (
    n1149,
    n566,
    n568,
    n1122
  );


  and
  g1117
  (
    n1139,
    n1132,
    n560,
    n574,
    n1122
  );


  nand
  g1118
  (
    n1177,
    n554,
    n551,
    n570,
    n557
  );


  xor
  g1119
  (
    n1182,
    n578,
    n587,
    n586,
    n1125
  );


  nand
  g1120
  (
    n1172,
    n568,
    n569,
    n573,
    n1133
  );


  and
  g1121
  (
    n1140,
    n570,
    n569,
    n556,
    n1131
  );


  and
  g1122
  (
    n1152,
    n553,
    n578,
    n543,
    n583
  );


  and
  g1123
  (
    n1188,
    n561,
    n591,
    n586,
    n581
  );


  nor
  g1124
  (
    n1159,
    n570,
    n577,
    n550,
    n1119
  );


  and
  g1125
  (
    n1137,
    n546,
    n574,
    n572,
    n560
  );


  and
  g1126
  (
    n1196,
    n576,
    n559,
    n566,
    n1119
  );


  or
  g1127
  (
    n1183,
    n565,
    n589,
    n556,
    n588
  );


  nor
  g1128
  (
    n1175,
    n552,
    n583,
    n559,
    n551
  );


  xnor
  g1129
  (
    n1157,
    n563,
    n582,
    n560,
    n590
  );


  and
  g1130
  (
    n1169,
    n1124,
    n544,
    n569,
    n546
  );


  xor
  g1131
  (
    n1195,
    n572,
    n1134,
    n579,
    n555
  );


  xnor
  g1132
  (
    n1184,
    n549,
    n580,
    n558,
    n570
  );


  or
  g1133
  (
    n1141,
    n554,
    n581,
    n543,
    n573
  );


  or
  g1134
  (
    n1153,
    n564,
    n1125,
    n549,
    n577
  );


  nand
  g1135
  (
    n1154,
    n1130,
    n564,
    n588,
    n547
  );


  xor
  g1136
  (
    n1166,
    n567,
    n572,
    n548,
    n1120
  );


  nand
  g1137
  (
    n1164,
    n581,
    n548,
    n562,
    n567
  );


  nand
  g1138
  (
    n1170,
    n590,
    n584,
    n562,
    n549
  );


  and
  g1139
  (
    n1146,
    n576,
    n568,
    n554,
    n583
  );


  nand
  g1140
  (
    n1178,
    n1134,
    n1123,
    n574,
    n561
  );


  nor
  g1141
  (
    n1135,
    n1121,
    n1128,
    n1120,
    n555
  );


  nand
  g1142
  (
    n1193,
    n557,
    n583,
    n1121,
    n1119
  );


  and
  g1143
  (
    n1167,
    n1126,
    n586,
    n1132,
    n1121
  );


  or
  g1144
  (
    n1151,
    n1130,
    n550,
    n552,
    n556
  );


  or
  g1145
  (
    n1143,
    n567,
    n589,
    n584,
    n552
  );


  nor
  g1146
  (
    n1163,
    n555,
    n559,
    n1133,
    n576
  );


  xnor
  g1147
  (
    n1173,
    n571,
    n577,
    n1128,
    n544
  );


  or
  g1148
  (
    n1198,
    n559,
    n553,
    n1129,
    n1127
  );


  xnor
  g1149
  (
    n1191,
    n1131,
    n556,
    n563,
    n572
  );


  xor
  g1150
  (
    n1155,
    n580,
    n551,
    n545,
    n543
  );


  or
  g1151
  (
    n1138,
    n1124,
    n550,
    n579,
    n586
  );


  nor
  g1152
  (
    n1180,
    n1126,
    n544,
    n546,
    n565
  );


  or
  g1153
  (
    n1185,
    n1134,
    n575,
    n1133,
    n588
  );


  nor
  g1154
  (
    n1189,
    n1125,
    n1128,
    n590,
    n1124
  );


  nand
  g1155
  (
    n1145,
    n561,
    n575,
    n545,
    n569
  );


  or
  g1156
  (
    n1148,
    n562,
    n547,
    n544,
    n1120
  );


  nor
  g1157
  (
    n1187,
    n1122,
    n584,
    n1132,
    n580
  );


  nand
  g1158
  (
    n1192,
    n587,
    n1126,
    n557,
    n547
  );


  and
  g1159
  (
    n1168,
    n547,
    n588,
    n1132,
    n565
  );


  xnor
  g1160
  (
    n1161,
    n552,
    n1129,
    n1124,
    n573
  );


  and
  g1161
  (
    n1150,
    n1133,
    n578,
    n575,
    n571
  );


  or
  g1162
  (
    n1181,
    n564,
    n560,
    n1119,
    n1129
  );


  and
  g1163
  (
    n1162,
    n1127,
    n579,
    n545,
    n575
  );


  and
  g1164
  (
    n1136,
    n585,
    n1125,
    n555,
    n577
  );


  xor
  g1165
  (
    n1156,
    n551,
    n579,
    n562,
    n582
  );


  and
  g1166
  (
    n1199,
    n810,
    n1136,
    n811,
    n808
  );


  xor
  g1167
  (
    n1200,
    n807,
    n1135,
    n809,
    n812
  );


  not
  g1168
  (
    n1203,
    n1200
  );


  buf
  g1169
  (
    n1202,
    n1200
  );


  buf
  g1170
  (
    n1201,
    n1199
  );


  xnor
  g1171
  (
    n1206,
    n1202,
    n1074,
    n1104,
    n592
  );


  and
  g1172
  (
    n1209,
    n1075,
    n595,
    n1073,
    n1105
  );


  or
  g1173
  (
    n1204,
    n1074,
    n1201,
    n593,
    n963
  );


  xor
  g1174
  (
    n1214,
    n1105,
    n1203,
    n594,
    n591
  );


  xnor
  g1175
  (
    n1212,
    n592,
    n596,
    n1075,
    n591
  );


  xor
  g1176
  (
    n1207,
    n962,
    n961,
    n591,
    n1076
  );


  and
  g1177
  (
    n1215,
    n962,
    n594,
    n596,
    n592
  );


  and
  g1178
  (
    n1210,
    n593,
    n1203,
    n1201,
    n961
  );


  xnor
  g1179
  (
    n1205,
    n595,
    n594,
    n1201,
    n1203
  );


  nor
  g1180
  (
    n1211,
    n1202,
    n592,
    n595,
    n1201
  );


  or
  g1181
  (
    n1213,
    n595,
    n593,
    n1203,
    n594
  );


  xor
  g1182
  (
    n1208,
    n593,
    n1202,
    n1073
  );


  or
  g1183
  (
    n1234,
    n825,
    n1029,
    n1205
  );


  nor
  g1184
  (
    n1223,
    n1210,
    n1204,
    n1172,
    n1208
  );


  xnor
  g1185
  (
    n1242,
    n1208,
    n1144,
    n1207,
    n1214
  );


  xor
  g1186
  (
    n1229,
    n1175,
    n1212,
    n1147,
    n1155
  );


  and
  g1187
  (
    n1244,
    n1138,
    n157,
    n821,
    n1142
  );


  xor
  g1188
  (
    n1246,
    n1143,
    n1164,
    n1206,
    n1078
  );


  xnor
  g1189
  (
    n1236,
    n1156,
    n1045,
    n1076,
    n1171
  );


  and
  g1190
  (
    n1219,
    n1159,
    n1208,
    n1215,
    n1213
  );


  or
  g1191
  (
    n1218,
    n814,
    n1077,
    n1044,
    n1149
  );


  or
  g1192
  (
    n1226,
    n155,
    n1213,
    n1215,
    n1081
  );


  or
  g1193
  (
    n1216,
    n1081,
    n1045,
    n156,
    n1206
  );


  nor
  g1194
  (
    n1240,
    n1214,
    n1145,
    n1210,
    n1205
  );


  xor
  g1195
  (
    n1241,
    n1139,
    n1211,
    n1170,
    n1206
  );


  xnor
  g1196
  (
    n1225,
    n815,
    n1213,
    n1209,
    n1161
  );


  xnor
  g1197
  (
    n1239,
    n1214,
    n1082,
    n1158,
    n1168
  );


  and
  g1198
  (
    n1233,
    n1215,
    n1082,
    n1205,
    n1029
  );


  xor
  g1199
  (
    n1217,
    n1079,
    n155,
    n1165,
    n1212
  );


  xnor
  g1200
  (
    n1222,
    n823,
    n1148,
    n1209,
    n1151
  );


  and
  g1201
  (
    n1231,
    n1079,
    n1209,
    n1146,
    n816
  );


  nand
  g1202
  (
    n1250,
    n1204,
    n1078,
    n819,
    n1211
  );


  and
  g1203
  (
    n1221,
    n1150,
    n824,
    n964,
    n1045
  );


  or
  g1204
  (
    n1220,
    n1166,
    n1207,
    n156,
    n1169
  );


  xor
  g1205
  (
    n1224,
    n1153,
    n1141,
    n1083,
    n1080
  );


  nand
  g1206
  (
    n1232,
    n1083,
    n1174,
    n1163,
    n1080
  );


  and
  g1207
  (
    n1227,
    n156,
    n1210,
    n813,
    n1213
  );


  xnor
  g1208
  (
    n1237,
    n1056,
    n827,
    n1207
  );


  xnor
  g1209
  (
    n1228,
    n1211,
    n1209,
    n820,
    n1154
  );


  nand
  g1210
  (
    n1247,
    n822,
    n1140,
    n1208,
    n1215
  );


  and
  g1211
  (
    n1243,
    n157,
    n1214,
    n1029,
    n1173
  );


  xnor
  g1212
  (
    n1238,
    n818,
    n1212,
    n1152,
    n826
  );


  xor
  g1213
  (
    n1248,
    n1204,
    n817,
    n1167,
    n1160
  );


  nor
  g1214
  (
    n1235,
    n1045,
    n1206,
    n1211,
    n1205
  );


  nand
  g1215
  (
    n1249,
    n1210,
    n963,
    n1212,
    n1077
  );


  nor
  g1216
  (
    n1245,
    n156,
    n1162,
    n1157,
    n1204
  );


  xor
  g1217
  (
    n1230,
    n1137,
    n1174,
    n1173,
    n964
  );


  xnor
  g1218
  (
    n1285,
    n1038,
    n1179,
    n1177,
    n1040
  );


  nand
  g1219
  (
    n1279,
    n1179,
    n601,
    n1036,
    n1247
  );


  xor
  g1220
  (
    n1257,
    n1233,
    n1034,
    n603,
    n1234
  );


  or
  g1221
  (
    n1252,
    n604,
    n1046,
    n603,
    n1225
  );


  xnor
  g1222
  (
    n1278,
    n602,
    n1036,
    n597,
    n1035
  );


  nand
  g1223
  (
    n1254,
    n1246,
    n1238,
    n1034,
    n1244
  );


  nor
  g1224
  (
    n1267,
    n1032,
    n1178,
    n601,
    n599
  );


  nand
  g1225
  (
    n1263,
    n1180,
    n1178,
    n597,
    n1176
  );


  or
  g1226
  (
    n1273,
    n600,
    n158,
    n1033
  );


  or
  g1227
  (
    n1269,
    n1039,
    n1032,
    n1041,
    n597
  );


  nand
  g1228
  (
    n1258,
    n1226,
    n602,
    n1181,
    n597
  );


  nand
  g1229
  (
    n1272,
    n1041,
    n1237,
    n1175,
    n1241
  );


  nand
  g1230
  (
    n1270,
    n1032,
    n1240,
    n1216,
    n1228
  );


  xnor
  g1231
  (
    n1261,
    n159,
    n599,
    n1032,
    n1245
  );


  or
  g1232
  (
    n1283,
    n1033,
    n598,
    n601,
    n600
  );


  or
  g1233
  (
    n1266,
    n159,
    n602,
    n1218,
    n1039
  );


  nand
  g1234
  (
    n1277,
    n159,
    n1217,
    n160,
    n601
  );


  and
  g1235
  (
    n1276,
    n1038,
    n1046,
    n1036,
    n604
  );


  nand
  g1236
  (
    n1259,
    n1182,
    n158,
    n1037,
    n1232
  );


  xor
  g1237
  (
    n1256,
    n1038,
    n157,
    n1046,
    n1231
  );


  xnor
  g1238
  (
    n1284,
    n158,
    n1035,
    n1033,
    n1031
  );


  xnor
  g1239
  (
    n1260,
    n1034,
    n1222,
    n1221,
    n598
  );


  xnor
  g1240
  (
    n1281,
    n604,
    n596,
    n1229,
    n1046
  );


  xor
  g1241
  (
    n1275,
    n1219,
    n1037,
    n1035,
    n603
  );


  nand
  g1242
  (
    n1268,
    n1037,
    n1039,
    n598,
    n1034
  );


  or
  g1243
  (
    n1280,
    n1176,
    n1180,
    n1223,
    n1227
  );


  nand
  g1244
  (
    n1262,
    n1035,
    n599,
    n602,
    n1037
  );


  xnor
  g1245
  (
    n1274,
    n604,
    n1041,
    n1181,
    n1033
  );


  and
  g1246
  (
    n1255,
    n1224,
    n159,
    n1243,
    n160
  );


  or
  g1247
  (
    n1251,
    n1041,
    n1242,
    n1235,
    n596
  );


  xor
  g1248
  (
    n1265,
    n1239,
    n1040,
    n157
  );


  nor
  g1249
  (
    n1271,
    n1250,
    n1236,
    n603,
    n1248
  );


  xor
  g1250
  (
    n1264,
    n600,
    n1177,
    n1036,
    n1220
  );


  xor
  g1251
  (
    n1253,
    n1230,
    n1040,
    n599,
    n1039
  );


  xor
  g1252
  (
    n1282,
    n1249,
    n598,
    n600,
    n1038
  );


  nand
  g1253
  (
    n1298,
    n1262,
    n1275,
    n1278,
    n1263
  );


  xor
  g1254
  (
    n1310,
    n1270,
    n1277,
    n1261,
    n1273
  );


  xor
  g1255
  (
    n1309,
    n1271,
    n1272,
    n1277,
    n1261
  );


  nor
  g1256
  (
    n1293,
    n1276,
    n1282,
    n1251,
    n1263
  );


  xnor
  g1257
  (
    n1302,
    n1281,
    n1267,
    n1255,
    n1261
  );


  xnor
  g1258
  (
    KeyWire_0_14,
    n1259,
    n1274,
    n1264,
    n1273
  );


  nand
  g1259
  (
    n1303,
    n1271,
    n1274,
    n1256,
    n1268
  );


  and
  g1260
  (
    n1292,
    n1266,
    n1267,
    n1276,
    n1257
  );


  and
  g1261
  (
    n1313,
    n1269,
    n1279,
    n1254,
    n1282
  );


  nand
  g1262
  (
    n1286,
    n1283,
    n1265,
    n1270,
    n1280
  );


  nor
  g1263
  (
    n1311,
    n1267,
    n1264,
    n1255,
    n1268
  );


  or
  g1264
  (
    n1306,
    n1253,
    n1274,
    n1266,
    n1259
  );


  or
  g1265
  (
    n1289,
    n1278,
    n1271,
    n1263,
    n1275
  );


  xor
  g1266
  (
    n1305,
    n1269,
    n1272,
    n1282,
    n1262
  );


  xnor
  g1267
  (
    n1291,
    n1265,
    n1276,
    n1261,
    n1263
  );


  xnor
  g1268
  (
    n1287,
    n1277,
    n1276,
    n1273,
    n1260
  );


  nor
  g1269
  (
    n1300,
    n1264,
    n1257,
    n1253,
    n1278
  );


  nor
  g1270
  (
    n1294,
    n1268,
    n1283,
    n1252
  );


  or
  g1271
  (
    n1296,
    n1282,
    n1258,
    n1275,
    n1269
  );


  nand
  g1272
  (
    n1307,
    n1275,
    n1281,
    n1269,
    n1265
  );


  xor
  g1273
  (
    n1301,
    n1267,
    n1278,
    n1251,
    n1273
  );


  and
  g1274
  (
    n1288,
    n1279,
    n1262,
    n1270,
    n1256
  );


  nor
  g1275
  (
    n1295,
    n1254,
    n1271,
    n1252,
    n1266
  );


  or
  g1276
  (
    n1290,
    n1262,
    n1272,
    n1279
  );


  or
  g1277
  (
    n1304,
    n1280,
    n1283,
    n1281
  );


  xnor
  g1278
  (
    n1312,
    n1272,
    n1258,
    n1277,
    n1260
  );


  nor
  g1279
  (
    n1297,
    n1270,
    n1265,
    n1280,
    n1274
  );


  xor
  g1280
  (
    n1299,
    n1266,
    n1268,
    n1280,
    n1264
  );


  and
  g1281
  (
    n1336,
    n1306,
    n1062,
    n1063,
    n970
  );


  nand
  g1282
  (
    n1314,
    n994,
    n1291,
    n984,
    n1200
  );


  or
  g1283
  (
    n1325,
    n995,
    n974,
    n988,
    n1305
  );


  xnor
  g1284
  (
    KeyWire_0_1,
    n1304,
    n1059,
    n983,
    n1064
  );


  nor
  g1285
  (
    n1333,
    n989,
    n975,
    n1061,
    n992
  );


  nand
  g1286
  (
    n1326,
    n965,
    n1183,
    n1298,
    n1058
  );


  nand
  g1287
  (
    n1327,
    n985,
    n1056,
    n976,
    n1290
  );


  nor
  g1288
  (
    n1322,
    n160,
    n1058,
    n972,
    n983
  );


  xnor
  g1289
  (
    n1347,
    n1311,
    n1306,
    n981,
    n978
  );


  xor
  g1290
  (
    n1329,
    n973,
    n994,
    n1312,
    n993
  );


  and
  g1291
  (
    n1330,
    n991,
    n975,
    n1065,
    n969
  );


  or
  g1292
  (
    n1350,
    n1297,
    n1309,
    n1060,
    n1062
  );


  nor
  g1293
  (
    n1337,
    n976,
    n1183,
    n1058,
    n1313
  );


  and
  g1294
  (
    n1349,
    n1308,
    n988,
    n1284,
    n1059
  );


  or
  g1295
  (
    n1340,
    n978,
    n1293,
    n984,
    n1064
  );


  nand
  g1296
  (
    n1324,
    n991,
    n1288,
    n1058,
    n1308
  );


  and
  g1297
  (
    n1338,
    n1292,
    n831,
    n1295,
    n986
  );


  or
  g1298
  (
    n1343,
    n828,
    n1305,
    n1056,
    n160
  );


  or
  g1299
  (
    n1342,
    n1063,
    n1313,
    n968,
    n1287
  );


  and
  g1300
  (
    n1339,
    n1309,
    n1064,
    n990,
    n1303
  );


  xor
  g1301
  (
    n1317,
    n1310,
    n965,
    n970,
    n981
  );


  nand
  g1302
  (
    n1320,
    n985,
    n993,
    n1307,
    n971
  );


  or
  g1303
  (
    n1348,
    n977,
    n982,
    n1060,
    n968
  );


  and
  g1304
  (
    n1328,
    n1061,
    n1061,
    n992,
    n829
  );


  xnor
  g1305
  (
    n1319,
    n1063,
    n972,
    n979,
    n967
  );


  nor
  g1306
  (
    n1323,
    n1299,
    n1059,
    n987,
    n1310
  );


  or
  g1307
  (
    n1331,
    n830,
    n1062,
    n1289,
    n1056
  );


  xnor
  g1308
  (
    n1318,
    n1064,
    n1063,
    n1060,
    n1057
  );


  xor
  g1309
  (
    n1316,
    n1307,
    n1050,
    n973,
    n1301
  );


  nand
  g1310
  (
    n1335,
    n1057,
    n966,
    n989
  );


  or
  g1311
  (
    n1345,
    n1286,
    n990,
    n1302,
    n1182
  );


  and
  g1312
  (
    n1344,
    n986,
    n982,
    n1059,
    n1061
  );


  nor
  g1313
  (
    n1334,
    n967,
    n1300,
    n1062,
    n1065
  );


  and
  g1314
  (
    n1315,
    n1057,
    n1312,
    n995,
    n980
  );


  xor
  g1315
  (
    n1341,
    n979,
    n969,
    n1311,
    n977
  );


  xnor
  g1316
  (
    n1346,
    n980,
    n1294,
    n1057,
    n987
  );


  xnor
  g1317
  (
    n1321,
    n971,
    n1060,
    n974,
    n1296
  );


  nor
  g1318
  (
    n1361,
    n1347,
    n1189,
    n1193,
    n1331
  );


  and
  g1319
  (
    n1368,
    n1187,
    n1348,
    n1349,
    n1188
  );


  nand
  g1320
  (
    n1358,
    n1321,
    n1328,
    n1185,
    n1084
  );


  nor
  g1321
  (
    n1359,
    n1345,
    n1085,
    n1336,
    n1084
  );


  xor
  g1322
  (
    KeyWire_0_7,
    n1197,
    n1320,
    n1200,
    n1186
  );


  and
  g1323
  (
    n1355,
    n1344,
    n1191,
    n1335,
    n1192
  );


  nand
  g1324
  (
    n1357,
    n1339,
    n1315,
    n1329,
    n1333
  );


  and
  g1325
  (
    n1364,
    n1350,
    n1196,
    n1317,
    n1197
  );


  nor
  g1326
  (
    n1366,
    n1085,
    n1327,
    n1284,
    n1323
  );


  or
  g1327
  (
    n1351,
    n1186,
    n1319,
    n1322,
    n1341
  );


  xnor
  g1328
  (
    n1362,
    n1198,
    n1191,
    n1065,
    n1195
  );


  xor
  g1329
  (
    n1356,
    n1330,
    n1192,
    n1338,
    n1196
  );


  or
  g1330
  (
    n1367,
    n1190,
    n1326,
    n1340,
    n1284
  );


  xor
  g1331
  (
    n1354,
    n1318,
    n1346,
    n1184,
    n1316
  );


  xnor
  g1332
  (
    n1360,
    n1195,
    n1190,
    n1189,
    n1332
  );


  and
  g1333
  (
    n1352,
    n1337,
    n1187,
    n1325,
    n1198
  );


  xnor
  g1334
  (
    n1363,
    n1324,
    n1188,
    n1194,
    n1343
  );


  nand
  g1335
  (
    n1353,
    n1194,
    n1065,
    n1184,
    n1342
  );


  xor
  g1336
  (
    n1369,
    n1314,
    n1193,
    n1185,
    n1334
  );


  and
  g1337
  (
    n1375,
    n1355,
    n1366,
    n1367,
    n1362
  );


  nor
  g1338
  (
    n1372,
    n1285,
    n1356,
    n1369,
    n1357
  );


  or
  g1339
  (
    n1370,
    n1352,
    n1365,
    n1361,
    n1368
  );


  nand
  g1340
  (
    n1374,
    n1363,
    n1364,
    n1351,
    n1360
  );


  nand
  g1341
  (
    n1373,
    n1285,
    n1285,
    n1284,
    n1358
  );


  nor
  g1342
  (
    n1371,
    n1354,
    n1285,
    n1359,
    n1353
  );


  xor
  KeyGate_0_0
  (
    n38,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1332,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1009,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n446,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n392,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n237,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n333,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1365,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n880,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1126,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n933,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n217,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n55,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n893,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1308,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n251,
    KeyNOTWire_0_15
  );


endmodule

