

module Stat_3000_433
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1674,
  n2471,
  n2480,
  n2989,
  n2993,
  n2986,
  n2998,
  n2994,
  n2985,
  n2987,
  n2991,
  n2983,
  n3001,
  n2984,
  n2990,
  n3004,
  n2988,
  n2997,
  n2999,
  n2996,
  n3002,
  n3000,
  n3007,
  n2992,
  n2982,
  n2995,
  n3003,
  n3005,
  n3030,
  n3031,
  n3029,
  n3032
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1674;output n2471;output n2480;output n2989;output n2993;output n2986;output n2998;output n2994;output n2985;output n2987;output n2991;output n2983;output n3001;output n2984;output n2990;output n3004;output n2988;output n2997;output n2999;output n2996;output n3002;output n3000;output n3007;output n2992;output n2982;output n2995;output n3003;output n3005;output n3030;output n3031;output n3029;output n3032;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n3006;wire n3008;wire n3009;wire n3010;wire n3011;wire n3012;wire n3013;wire n3014;wire n3015;wire n3016;wire n3017;wire n3018;wire n3019;wire n3020;wire n3021;wire n3022;wire n3023;wire n3024;wire n3025;wire n3026;wire n3027;wire n3028;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n58,
    n8
  );


  not
  g1
  (
    n114,
    n16
  );


  not
  g2
  (
    n120,
    n32
  );


  not
  g3
  (
    n156,
    n9
  );


  buf
  g4
  (
    n100,
    n23
  );


  not
  g5
  (
    n133,
    n10
  );


  not
  g6
  (
    n98,
    n26
  );


  not
  g7
  (
    n153,
    n16
  );


  buf
  g8
  (
    n143,
    n28
  );


  buf
  g9
  (
    n55,
    n28
  );


  buf
  g10
  (
    n123,
    n13
  );


  buf
  g11
  (
    n61,
    n27
  );


  buf
  g12
  (
    n45,
    n20
  );


  buf
  g13
  (
    n34,
    n31
  );


  buf
  g14
  (
    n141,
    n24
  );


  buf
  g15
  (
    n44,
    n15
  );


  buf
  g16
  (
    n96,
    n6
  );


  buf
  g17
  (
    n43,
    n18
  );


  buf
  g18
  (
    n104,
    n23
  );


  buf
  g19
  (
    n99,
    n30
  );


  not
  g20
  (
    n89,
    n30
  );


  not
  g21
  (
    n145,
    n22
  );


  buf
  g22
  (
    n42,
    n25
  );


  not
  g23
  (
    n41,
    n26
  );


  buf
  g24
  (
    n50,
    n19
  );


  buf
  g25
  (
    n82,
    n1
  );


  not
  g26
  (
    n150,
    n24
  );


  not
  g27
  (
    n102,
    n31
  );


  not
  g28
  (
    n69,
    n2
  );


  not
  g29
  (
    n52,
    n27
  );


  buf
  g30
  (
    n108,
    n10
  );


  buf
  g31
  (
    n155,
    n28
  );


  buf
  g32
  (
    n74,
    n13
  );


  not
  g33
  (
    n51,
    n23
  );


  buf
  g34
  (
    n128,
    n14
  );


  buf
  g35
  (
    n140,
    n21
  );


  not
  g36
  (
    n85,
    n2
  );


  buf
  g37
  (
    n124,
    n12
  );


  not
  g38
  (
    n148,
    n3
  );


  buf
  g39
  (
    n149,
    n14
  );


  buf
  g40
  (
    n147,
    n13
  );


  buf
  g41
  (
    n75,
    n21
  );


  not
  g42
  (
    n54,
    n1
  );


  buf
  g43
  (
    n137,
    n3
  );


  buf
  g44
  (
    n121,
    n14
  );


  buf
  g45
  (
    n63,
    n20
  );


  buf
  g46
  (
    n77,
    n29
  );


  not
  g47
  (
    n97,
    n5
  );


  not
  g48
  (
    n160,
    n4
  );


  buf
  g49
  (
    n119,
    n19
  );


  buf
  g50
  (
    KeyWire_0_17,
    n9
  );


  buf
  g51
  (
    n146,
    n4
  );


  buf
  g52
  (
    n159,
    n7
  );


  not
  g53
  (
    n47,
    n17
  );


  not
  g54
  (
    n101,
    n1
  );


  not
  g55
  (
    n154,
    n11
  );


  buf
  g56
  (
    n142,
    n10
  );


  not
  g57
  (
    n127,
    n17
  );


  not
  g58
  (
    n95,
    n32
  );


  not
  g59
  (
    n135,
    n27
  );


  not
  g60
  (
    n76,
    n27
  );


  buf
  g61
  (
    n129,
    n21
  );


  not
  g62
  (
    n122,
    n16
  );


  buf
  g63
  (
    n157,
    n12
  );


  buf
  g64
  (
    n68,
    n2
  );


  not
  g65
  (
    n152,
    n26
  );


  buf
  g66
  (
    n84,
    n21
  );


  not
  g67
  (
    n139,
    n32
  );


  buf
  g68
  (
    n66,
    n4
  );


  buf
  g69
  (
    n73,
    n2
  );


  not
  g70
  (
    n136,
    n11
  );


  buf
  g71
  (
    n125,
    n20
  );


  not
  g72
  (
    n106,
    n6
  );


  buf
  g73
  (
    n94,
    n9
  );


  buf
  g74
  (
    n70,
    n26
  );


  buf
  g75
  (
    n138,
    n6
  );


  buf
  g76
  (
    n116,
    n18
  );


  not
  g77
  (
    n130,
    n25
  );


  not
  g78
  (
    n151,
    n25
  );


  buf
  g79
  (
    n109,
    n18
  );


  buf
  g80
  (
    n107,
    n28
  );


  not
  g81
  (
    n111,
    n8
  );


  buf
  g82
  (
    n110,
    n24
  );


  not
  g83
  (
    n48,
    n25
  );


  not
  g84
  (
    n126,
    n23
  );


  buf
  g85
  (
    n33,
    n29
  );


  buf
  g86
  (
    n92,
    n11
  );


  buf
  g87
  (
    n134,
    n5
  );


  buf
  g88
  (
    n78,
    n19
  );


  not
  g89
  (
    n113,
    n7
  );


  buf
  g90
  (
    n115,
    n11
  );


  buf
  g91
  (
    n93,
    n13
  );


  not
  g92
  (
    n49,
    n7
  );


  buf
  g93
  (
    n67,
    n6
  );


  not
  g94
  (
    n46,
    n22
  );


  buf
  g95
  (
    n56,
    n18
  );


  not
  g96
  (
    n118,
    n32
  );


  buf
  g97
  (
    n158,
    n22
  );


  not
  g98
  (
    n59,
    n20
  );


  not
  g99
  (
    n83,
    n5
  );


  not
  g100
  (
    n72,
    n30
  );


  not
  g101
  (
    n117,
    n29
  );


  buf
  g102
  (
    n144,
    n17
  );


  not
  g103
  (
    n57,
    n15
  );


  not
  g104
  (
    n37,
    n3
  );


  buf
  g105
  (
    n103,
    n8
  );


  not
  g106
  (
    n53,
    n16
  );


  not
  g107
  (
    n62,
    n3
  );


  not
  g108
  (
    n80,
    n7
  );


  not
  g109
  (
    n40,
    n5
  );


  not
  g110
  (
    n60,
    n17
  );


  buf
  g111
  (
    n86,
    n1
  );


  not
  g112
  (
    n132,
    n4
  );


  buf
  g113
  (
    n87,
    n22
  );


  buf
  g114
  (
    n64,
    n15
  );


  buf
  g115
  (
    n36,
    n15
  );


  buf
  g116
  (
    n65,
    n30
  );


  not
  g117
  (
    n35,
    n29
  );


  not
  g118
  (
    n131,
    n12
  );


  not
  g119
  (
    n88,
    n8
  );


  buf
  g120
  (
    n105,
    n31
  );


  buf
  g121
  (
    n71,
    n19
  );


  buf
  g122
  (
    n38,
    n10
  );


  buf
  g123
  (
    n91,
    n24
  );


  buf
  g124
  (
    n90,
    n14
  );


  not
  g125
  (
    n79,
    n31
  );


  not
  g126
  (
    n112,
    n9
  );


  not
  g127
  (
    n39,
    n12
  );


  buf
  g128
  (
    n380,
    n49
  );


  not
  g129
  (
    n283,
    n48
  );


  not
  g130
  (
    n351,
    n133
  );


  not
  g131
  (
    n332,
    n59
  );


  not
  g132
  (
    n299,
    n125
  );


  not
  g133
  (
    n447,
    n33
  );


  not
  g134
  (
    n232,
    n158
  );


  not
  g135
  (
    n313,
    n120
  );


  not
  g136
  (
    n166,
    n69
  );


  not
  g137
  (
    n344,
    n77
  );


  not
  g138
  (
    n670,
    n72
  );


  buf
  g139
  (
    n265,
    n79
  );


  buf
  g140
  (
    n656,
    n117
  );


  buf
  g141
  (
    n331,
    n103
  );


  buf
  g142
  (
    KeyWire_0_18,
    n153
  );


  buf
  g143
  (
    n168,
    n87
  );


  buf
  g144
  (
    n206,
    n132
  );


  not
  g145
  (
    n250,
    n159
  );


  not
  g146
  (
    n277,
    n115
  );


  buf
  g147
  (
    n169,
    n67
  );


  buf
  g148
  (
    n583,
    n137
  );


  not
  g149
  (
    n479,
    n38
  );


  not
  g150
  (
    n466,
    n116
  );


  not
  g151
  (
    n597,
    n71
  );


  buf
  g152
  (
    n204,
    n34
  );


  not
  g153
  (
    n573,
    n103
  );


  buf
  g154
  (
    n249,
    n85
  );


  buf
  g155
  (
    n643,
    n141
  );


  not
  g156
  (
    n360,
    n75
  );


  buf
  g157
  (
    n502,
    n57
  );


  not
  g158
  (
    n374,
    n100
  );


  buf
  g159
  (
    KeyWire_0_30,
    n65
  );


  buf
  g160
  (
    n349,
    n108
  );


  buf
  g161
  (
    n409,
    n159
  );


  not
  g162
  (
    n252,
    n139
  );


  buf
  g163
  (
    n624,
    n68
  );


  not
  g164
  (
    n602,
    n85
  );


  not
  g165
  (
    n385,
    n104
  );


  buf
  g166
  (
    n304,
    n82
  );


  buf
  g167
  (
    n207,
    n73
  );


  buf
  g168
  (
    n665,
    n147
  );


  not
  g169
  (
    n621,
    n45
  );


  buf
  g170
  (
    n419,
    n139
  );


  buf
  g171
  (
    n383,
    n141
  );


  buf
  g172
  (
    n556,
    n111
  );


  buf
  g173
  (
    n414,
    n63
  );


  buf
  g174
  (
    n375,
    n84
  );


  not
  g175
  (
    n172,
    n61
  );


  buf
  g176
  (
    n664,
    n67
  );


  buf
  g177
  (
    n623,
    n127
  );


  buf
  g178
  (
    n197,
    n37
  );


  buf
  g179
  (
    n390,
    n78
  );


  not
  g180
  (
    n552,
    n159
  );


  buf
  g181
  (
    n511,
    n40
  );


  buf
  g182
  (
    n578,
    n131
  );


  buf
  g183
  (
    n521,
    n60
  );


  not
  g184
  (
    n454,
    n48
  );


  buf
  g185
  (
    n213,
    n95
  );


  buf
  g186
  (
    n508,
    n113
  );


  not
  g187
  (
    n403,
    n110
  );


  not
  g188
  (
    n547,
    n132
  );


  not
  g189
  (
    n242,
    n155
  );


  not
  g190
  (
    n235,
    n157
  );


  buf
  g191
  (
    n572,
    n91
  );


  buf
  g192
  (
    n495,
    n75
  );


  buf
  g193
  (
    n534,
    n43
  );


  buf
  g194
  (
    n340,
    n92
  );


  buf
  g195
  (
    n259,
    n138
  );


  buf
  g196
  (
    n499,
    n66
  );


  not
  g197
  (
    n575,
    n59
  );


  not
  g198
  (
    n588,
    n43
  );


  not
  g199
  (
    n557,
    n80
  );


  buf
  g200
  (
    n494,
    n101
  );


  not
  g201
  (
    n345,
    n152
  );


  not
  g202
  (
    n367,
    n51
  );


  buf
  g203
  (
    n425,
    n54
  );


  buf
  g204
  (
    n445,
    n84
  );


  not
  g205
  (
    n382,
    n142
  );


  buf
  g206
  (
    n472,
    n143
  );


  buf
  g207
  (
    n647,
    n57
  );


  buf
  g208
  (
    n372,
    n89
  );


  not
  g209
  (
    n310,
    n139
  );


  buf
  g210
  (
    n585,
    n67
  );


  buf
  g211
  (
    n193,
    n131
  );


  not
  g212
  (
    n397,
    n152
  );


  not
  g213
  (
    n630,
    n47
  );


  buf
  g214
  (
    n203,
    n100
  );


  buf
  g215
  (
    n482,
    n59
  );


  not
  g216
  (
    n452,
    n109
  );


  not
  g217
  (
    n410,
    n144
  );


  buf
  g218
  (
    n294,
    n90
  );


  buf
  g219
  (
    n337,
    n75
  );


  not
  g220
  (
    n642,
    n88
  );


  not
  g221
  (
    n510,
    n38
  );


  not
  g222
  (
    n287,
    n93
  );


  buf
  g223
  (
    n653,
    n56
  );


  not
  g224
  (
    n526,
    n135
  );


  not
  g225
  (
    n429,
    n53
  );


  buf
  g226
  (
    n363,
    n119
  );


  not
  g227
  (
    n342,
    n121
  );


  buf
  g228
  (
    n280,
    n33
  );


  not
  g229
  (
    n481,
    n45
  );


  buf
  g230
  (
    n399,
    n71
  );


  buf
  g231
  (
    n487,
    n37
  );


  buf
  g232
  (
    n546,
    n138
  );


  buf
  g233
  (
    n171,
    n100
  );


  not
  g234
  (
    n369,
    n143
  );


  not
  g235
  (
    n335,
    n122
  );


  buf
  g236
  (
    n306,
    n151
  );


  not
  g237
  (
    n655,
    n137
  );


  buf
  g238
  (
    n343,
    n76
  );


  buf
  g239
  (
    KeyWire_0_22,
    n160
  );


  buf
  g240
  (
    n353,
    n129
  );


  buf
  g241
  (
    n542,
    n92
  );


  not
  g242
  (
    n240,
    n54
  );


  buf
  g243
  (
    KeyWire_0_28,
    n129
  );


  buf
  g244
  (
    n554,
    n91
  );


  buf
  g245
  (
    n632,
    n104
  );


  buf
  g246
  (
    n519,
    n126
  );


  buf
  g247
  (
    n317,
    n120
  );


  not
  g248
  (
    n366,
    n159
  );


  buf
  g249
  (
    n274,
    n153
  );


  buf
  g250
  (
    n210,
    n113
  );


  buf
  g251
  (
    n218,
    n60
  );


  not
  g252
  (
    n318,
    n136
  );


  not
  g253
  (
    n644,
    n116
  );


  buf
  g254
  (
    n417,
    n87
  );


  buf
  g255
  (
    n262,
    n150
  );


  buf
  g256
  (
    n569,
    n105
  );


  not
  g257
  (
    n458,
    n138
  );


  not
  g258
  (
    n501,
    n140
  );


  not
  g259
  (
    n266,
    n149
  );


  not
  g260
  (
    n229,
    n42
  );


  buf
  g261
  (
    n324,
    n140
  );


  buf
  g262
  (
    n307,
    n149
  );


  not
  g263
  (
    n416,
    n36
  );


  buf
  g264
  (
    n507,
    n34
  );


  buf
  g265
  (
    KeyWire_0_13,
    n69
  );


  not
  g266
  (
    n355,
    n119
  );


  not
  g267
  (
    n174,
    n72
  );


  buf
  g268
  (
    n222,
    n115
  );


  not
  g269
  (
    n189,
    n66
  );


  not
  g270
  (
    n500,
    n124
  );


  buf
  g271
  (
    n386,
    n114
  );


  buf
  g272
  (
    n412,
    n134
  );


  not
  g273
  (
    n347,
    n142
  );


  not
  g274
  (
    n549,
    n107
  );


  not
  g275
  (
    n650,
    n118
  );


  buf
  g276
  (
    n178,
    n56
  );


  buf
  g277
  (
    n165,
    n53
  );


  buf
  g278
  (
    n540,
    n134
  );


  buf
  g279
  (
    n606,
    n125
  );


  buf
  g280
  (
    n480,
    n111
  );


  not
  g281
  (
    n336,
    n141
  );


  buf
  g282
  (
    n405,
    n58
  );


  buf
  g283
  (
    n270,
    n141
  );


  buf
  g284
  (
    n513,
    n71
  );


  buf
  g285
  (
    n341,
    n63
  );


  not
  g286
  (
    n612,
    n87
  );


  buf
  g287
  (
    n357,
    n101
  );


  buf
  g288
  (
    n202,
    n135
  );


  buf
  g289
  (
    n555,
    n78
  );


  buf
  g290
  (
    n443,
    n125
  );


  buf
  g291
  (
    n301,
    n51
  );


  not
  g292
  (
    n492,
    n62
  );


  buf
  g293
  (
    n214,
    n112
  );


  buf
  g294
  (
    n322,
    n55
  );


  buf
  g295
  (
    n576,
    n94
  );


  buf
  g296
  (
    n600,
    n84
  );


  buf
  g297
  (
    n545,
    n56
  );


  buf
  g298
  (
    n185,
    n126
  );


  buf
  g299
  (
    n520,
    n104
  );


  buf
  g300
  (
    n544,
    n78
  );


  not
  g301
  (
    n362,
    n134
  );


  not
  g302
  (
    n496,
    n82
  );


  buf
  g303
  (
    n477,
    n39
  );


  not
  g304
  (
    n219,
    n41
  );


  buf
  g305
  (
    n231,
    n135
  );


  buf
  g306
  (
    n657,
    n128
  );


  buf
  g307
  (
    n660,
    n54
  );


  buf
  g308
  (
    n486,
    n86
  );


  buf
  g309
  (
    n463,
    n82
  );


  not
  g310
  (
    n389,
    n91
  );


  not
  g311
  (
    n626,
    n46
  );


  not
  g312
  (
    n599,
    n96
  );


  not
  g313
  (
    n581,
    n149
  );


  not
  g314
  (
    n563,
    n64
  );


  not
  g315
  (
    n288,
    n143
  );


  not
  g316
  (
    n509,
    n73
  );


  not
  g317
  (
    n640,
    n148
  );


  buf
  g318
  (
    n361,
    n116
  );


  not
  g319
  (
    n292,
    n45
  );


  not
  g320
  (
    n271,
    n112
  );


  buf
  g321
  (
    n446,
    n88
  );


  buf
  g322
  (
    n604,
    n131
  );


  not
  g323
  (
    n488,
    n61
  );


  not
  g324
  (
    n436,
    n72
  );


  not
  g325
  (
    n395,
    n108
  );


  buf
  g326
  (
    n639,
    n105
  );


  not
  g327
  (
    n170,
    n123
  );


  buf
  g328
  (
    n562,
    n89
  );


  not
  g329
  (
    n183,
    n99
  );


  not
  g330
  (
    n596,
    n130
  );


  not
  g331
  (
    n613,
    n122
  );


  not
  g332
  (
    n491,
    n65
  );


  not
  g333
  (
    n475,
    n137
  );


  buf
  g334
  (
    n348,
    n154
  );


  buf
  g335
  (
    n352,
    n41
  );


  buf
  g336
  (
    n528,
    n85
  );


  buf
  g337
  (
    n442,
    n156
  );


  not
  g338
  (
    n590,
    n153
  );


  not
  g339
  (
    n584,
    n41
  );


  not
  g340
  (
    n568,
    n52
  );


  not
  g341
  (
    n497,
    n77
  );


  not
  g342
  (
    n661,
    n156
  );


  not
  g343
  (
    n255,
    n109
  );


  not
  g344
  (
    n328,
    n38
  );


  not
  g345
  (
    n512,
    n86
  );


  buf
  g346
  (
    n393,
    n44
  );


  buf
  g347
  (
    n257,
    n145
  );


  buf
  g348
  (
    n293,
    n114
  );


  not
  g349
  (
    n560,
    n98
  );


  buf
  g350
  (
    n167,
    n82
  );


  not
  g351
  (
    n227,
    n50
  );


  buf
  g352
  (
    n236,
    n50
  );


  buf
  g353
  (
    n459,
    n48
  );


  buf
  g354
  (
    n498,
    n143
  );


  buf
  g355
  (
    n594,
    n160
  );


  not
  g356
  (
    n591,
    n117
  );


  not
  g357
  (
    n413,
    n105
  );


  not
  g358
  (
    n663,
    n73
  );


  buf
  g359
  (
    n617,
    n76
  );


  buf
  g360
  (
    KeyWire_0_26,
    n157
  );


  buf
  g361
  (
    n566,
    n146
  );


  not
  g362
  (
    n201,
    n102
  );


  buf
  g363
  (
    n634,
    n122
  );


  not
  g364
  (
    n548,
    n138
  );


  buf
  g365
  (
    n377,
    n49
  );


  buf
  g366
  (
    n421,
    n36
  );


  buf
  g367
  (
    n619,
    n130
  );


  buf
  g368
  (
    n433,
    n135
  );


  not
  g369
  (
    n457,
    n152
  );


  buf
  g370
  (
    n490,
    n63
  );


  buf
  g371
  (
    n273,
    n101
  );


  buf
  g372
  (
    n254,
    n65
  );


  not
  g373
  (
    n543,
    n78
  );


  not
  g374
  (
    n538,
    n33
  );


  buf
  g375
  (
    n672,
    n147
  );


  not
  g376
  (
    n225,
    n103
  );


  buf
  g377
  (
    n483,
    n102
  );


  not
  g378
  (
    n267,
    n123
  );


  not
  g379
  (
    n381,
    n49
  );


  not
  g380
  (
    n577,
    n62
  );


  buf
  g381
  (
    n354,
    n121
  );


  not
  g382
  (
    n633,
    n52
  );


  buf
  g383
  (
    n551,
    n100
  );


  not
  g384
  (
    n648,
    n69
  );


  buf
  g385
  (
    n531,
    n120
  );


  not
  g386
  (
    n305,
    n110
  );


  not
  g387
  (
    n541,
    n51
  );


  buf
  g388
  (
    n415,
    n48
  );


  not
  g389
  (
    n319,
    n98
  );


  buf
  g390
  (
    n320,
    n53
  );


  buf
  g391
  (
    n587,
    n98
  );


  not
  g392
  (
    n176,
    n111
  );


  buf
  g393
  (
    n586,
    n109
  );


  buf
  g394
  (
    n515,
    n92
  );


  buf
  g395
  (
    n184,
    n74
  );


  not
  g396
  (
    n198,
    n102
  );


  buf
  g397
  (
    n522,
    n94
  );


  buf
  g398
  (
    n312,
    n81
  );


  not
  g399
  (
    n455,
    n46
  );


  not
  g400
  (
    n489,
    n87
  );


  buf
  g401
  (
    n517,
    n106
  );


  not
  g402
  (
    n618,
    n62
  );


  not
  g403
  (
    n401,
    n125
  );


  not
  g404
  (
    n323,
    n65
  );


  buf
  g405
  (
    n607,
    n112
  );


  not
  g406
  (
    n408,
    n90
  );


  buf
  g407
  (
    n539,
    n45
  );


  not
  g408
  (
    n418,
    n140
  );


  buf
  g409
  (
    n286,
    n58
  );


  buf
  g410
  (
    n209,
    n150
  );


  not
  g411
  (
    n220,
    n111
  );


  not
  g412
  (
    n180,
    n97
  );


  buf
  g413
  (
    n506,
    n151
  );


  not
  g414
  (
    n290,
    n148
  );


  buf
  g415
  (
    n190,
    n103
  );


  buf
  g416
  (
    n470,
    n116
  );


  not
  g417
  (
    n298,
    n97
  );


  not
  g418
  (
    n530,
    n80
  );


  buf
  g419
  (
    n641,
    n43
  );


  buf
  g420
  (
    n253,
    n33
  );


  not
  g421
  (
    n561,
    n127
  );


  not
  g422
  (
    n609,
    n132
  );


  buf
  g423
  (
    n230,
    n102
  );


  not
  g424
  (
    n302,
    n129
  );


  not
  g425
  (
    n284,
    n150
  );


  buf
  g426
  (
    n303,
    n155
  );


  buf
  g427
  (
    n391,
    n108
  );


  not
  g428
  (
    n411,
    n81
  );


  buf
  g429
  (
    n559,
    n136
  );


  buf
  g430
  (
    n350,
    n136
  );


  buf
  g431
  (
    n478,
    n53
  );


  not
  g432
  (
    n241,
    n96
  );


  not
  g433
  (
    n666,
    n46
  );


  not
  g434
  (
    n338,
    n114
  );


  not
  g435
  (
    n620,
    n93
  );


  not
  g436
  (
    n484,
    n89
  );


  not
  g437
  (
    n662,
    n60
  );


  buf
  g438
  (
    n200,
    n158
  );


  buf
  g439
  (
    n668,
    n47
  );


  not
  g440
  (
    n321,
    n64
  );


  not
  g441
  (
    n654,
    n147
  );


  not
  g442
  (
    n394,
    n145
  );


  not
  g443
  (
    n468,
    n104
  );


  not
  g444
  (
    n275,
    n142
  );


  buf
  g445
  (
    n669,
    n47
  );


  not
  g446
  (
    n289,
    n120
  );


  buf
  g447
  (
    n423,
    n68
  );


  buf
  g448
  (
    n358,
    n153
  );


  buf
  g449
  (
    n223,
    n149
  );


  buf
  g450
  (
    n285,
    n118
  );


  not
  g451
  (
    n430,
    n86
  );


  buf
  g452
  (
    n516,
    n95
  );


  buf
  g453
  (
    n325,
    n37
  );


  not
  g454
  (
    n467,
    n81
  );


  buf
  g455
  (
    n179,
    n39
  );


  buf
  g456
  (
    n334,
    n58
  );


  buf
  g457
  (
    n282,
    n137
  );


  buf
  g458
  (
    n651,
    n44
  );


  not
  g459
  (
    n608,
    n58
  );


  buf
  g460
  (
    n364,
    n155
  );


  not
  g461
  (
    n191,
    n43
  );


  not
  g462
  (
    n631,
    n151
  );


  not
  g463
  (
    n469,
    n126
  );


  not
  g464
  (
    n432,
    n124
  );


  not
  g465
  (
    n226,
    n61
  );


  buf
  g466
  (
    n258,
    n77
  );


  not
  g467
  (
    n244,
    n64
  );


  not
  g468
  (
    n579,
    n84
  );


  buf
  g469
  (
    KeyWire_0_20,
    n35
  );


  buf
  g470
  (
    n460,
    n72
  );


  buf
  g471
  (
    n615,
    n112
  );


  not
  g472
  (
    n195,
    n110
  );


  not
  g473
  (
    n233,
    n94
  );


  buf
  g474
  (
    n625,
    n70
  );


  buf
  g475
  (
    n256,
    n93
  );


  buf
  g476
  (
    n260,
    n160
  );


  not
  g477
  (
    n427,
    n70
  );


  buf
  g478
  (
    n396,
    n134
  );


  not
  g479
  (
    n279,
    n127
  );


  not
  g480
  (
    n616,
    n47
  );


  buf
  g481
  (
    n627,
    n76
  );


  not
  g482
  (
    n309,
    n83
  );


  not
  g483
  (
    n173,
    n157
  );


  not
  g484
  (
    n217,
    n133
  );


  not
  g485
  (
    n529,
    n145
  );


  not
  g486
  (
    n314,
    n50
  );


  buf
  g487
  (
    n505,
    n79
  );


  buf
  g488
  (
    n461,
    n113
  );


  buf
  g489
  (
    n368,
    n106
  );


  buf
  g490
  (
    n246,
    n88
  );


  not
  g491
  (
    n264,
    n49
  );


  buf
  g492
  (
    n659,
    n60
  );


  buf
  g493
  (
    n658,
    n145
  );


  buf
  g494
  (
    n186,
    n52
  );


  not
  g495
  (
    n404,
    n123
  );


  buf
  g496
  (
    n444,
    n41
  );


  buf
  g497
  (
    n536,
    n83
  );


  buf
  g498
  (
    n503,
    n146
  );


  buf
  g499
  (
    n533,
    n107
  );


  buf
  g500
  (
    n645,
    n124
  );


  not
  g501
  (
    n605,
    n61
  );


  not
  g502
  (
    n504,
    n94
  );


  buf
  g503
  (
    n163,
    n114
  );


  buf
  g504
  (
    n311,
    n91
  );


  not
  g505
  (
    n199,
    n117
  );


  not
  g506
  (
    n330,
    n160
  );


  not
  g507
  (
    n300,
    n86
  );


  not
  g508
  (
    n365,
    n130
  );


  buf
  g509
  (
    n263,
    n115
  );


  not
  g510
  (
    KeyWire_0_14,
    n144
  );


  buf
  g511
  (
    n221,
    n113
  );


  not
  g512
  (
    n402,
    n154
  );


  not
  g513
  (
    n574,
    n38
  );


  buf
  g514
  (
    n346,
    n69
  );


  buf
  g515
  (
    n595,
    n34
  );


  buf
  g516
  (
    n392,
    n133
  );


  not
  g517
  (
    n182,
    n80
  );


  buf
  g518
  (
    n376,
    n77
  );


  buf
  g519
  (
    n441,
    n121
  );


  not
  g520
  (
    n378,
    n119
  );


  not
  g521
  (
    n177,
    n126
  );


  not
  g522
  (
    n181,
    n85
  );


  not
  g523
  (
    n434,
    n106
  );


  not
  g524
  (
    n564,
    n148
  );


  buf
  g525
  (
    n248,
    n39
  );


  buf
  g526
  (
    n297,
    n97
  );


  buf
  g527
  (
    n440,
    n83
  );


  buf
  g528
  (
    n224,
    n46
  );


  not
  g529
  (
    n671,
    n40
  );


  buf
  g530
  (
    n315,
    n70
  );


  not
  g531
  (
    n398,
    n155
  );


  buf
  g532
  (
    n316,
    n158
  );


  not
  g533
  (
    n439,
    n110
  );


  buf
  g534
  (
    n610,
    n42
  );


  not
  g535
  (
    n476,
    n132
  );


  buf
  g536
  (
    n228,
    n68
  );


  not
  g537
  (
    n635,
    n89
  );


  not
  g538
  (
    n356,
    n128
  );


  not
  g539
  (
    n558,
    n67
  );


  buf
  g540
  (
    n194,
    n108
  );


  buf
  g541
  (
    n636,
    n98
  );


  buf
  g542
  (
    n379,
    n118
  );


  not
  g543
  (
    n527,
    n40
  );


  buf
  g544
  (
    n388,
    n57
  );


  not
  g545
  (
    n438,
    n70
  );


  not
  g546
  (
    n339,
    n147
  );


  not
  g547
  (
    n524,
    n83
  );


  buf
  g548
  (
    n326,
    n140
  );


  not
  g549
  (
    n278,
    n115
  );


  buf
  g550
  (
    n208,
    n117
  );


  not
  g551
  (
    n550,
    n131
  );


  buf
  g552
  (
    n426,
    n156
  );


  buf
  g553
  (
    n424,
    n151
  );


  not
  g554
  (
    n518,
    n95
  );


  buf
  g555
  (
    n580,
    n92
  );


  not
  g556
  (
    n164,
    n71
  );


  buf
  g557
  (
    n603,
    n157
  );


  not
  g558
  (
    n192,
    n50
  );


  not
  g559
  (
    n308,
    n90
  );


  not
  g560
  (
    n281,
    n142
  );


  not
  g561
  (
    n514,
    n35
  );


  not
  g562
  (
    n428,
    n96
  );


  not
  g563
  (
    n451,
    n133
  );


  not
  g564
  (
    n329,
    n42
  );


  buf
  g565
  (
    n565,
    n36
  );


  not
  g566
  (
    n243,
    n74
  );


  buf
  g567
  (
    n371,
    n95
  );


  buf
  g568
  (
    n400,
    n39
  );


  not
  g569
  (
    n212,
    n144
  );


  buf
  g570
  (
    n420,
    n56
  );


  not
  g571
  (
    n359,
    n35
  );


  not
  g572
  (
    n525,
    n118
  );


  not
  g573
  (
    n589,
    n101
  );


  not
  g574
  (
    n407,
    n156
  );


  buf
  g575
  (
    n593,
    n52
  );


  not
  g576
  (
    n234,
    n107
  );


  not
  g577
  (
    n567,
    n146
  );


  not
  g578
  (
    n456,
    n76
  );


  not
  g579
  (
    n215,
    n136
  );


  not
  g580
  (
    n175,
    n119
  );


  buf
  g581
  (
    n493,
    n57
  );


  buf
  g582
  (
    n187,
    n99
  );


  buf
  g583
  (
    n239,
    n122
  );


  not
  g584
  (
    n333,
    n121
  );


  not
  g585
  (
    n272,
    n106
  );


  buf
  g586
  (
    n582,
    n35
  );


  not
  g587
  (
    n471,
    n54
  );


  not
  g588
  (
    n327,
    n150
  );


  not
  g589
  (
    n570,
    n96
  );


  not
  g590
  (
    n448,
    n37
  );


  not
  g591
  (
    n667,
    n127
  );


  not
  g592
  (
    n622,
    n128
  );


  buf
  g593
  (
    n649,
    n44
  );


  buf
  g594
  (
    n474,
    n55
  );


  not
  g595
  (
    n537,
    n51
  );


  not
  g596
  (
    n384,
    n109
  );


  buf
  g597
  (
    n449,
    n146
  );


  buf
  g598
  (
    n370,
    n124
  );


  not
  g599
  (
    n523,
    n99
  );


  not
  g600
  (
    n268,
    n139
  );


  buf
  g601
  (
    n238,
    n59
  );


  not
  g602
  (
    n437,
    n81
  );


  not
  g603
  (
    n601,
    n68
  );


  buf
  g604
  (
    n291,
    n93
  );


  not
  g605
  (
    n406,
    n80
  );


  not
  g606
  (
    n422,
    n90
  );


  buf
  g607
  (
    n473,
    n36
  );


  not
  g608
  (
    n216,
    n75
  );


  not
  g609
  (
    n276,
    n55
  );


  buf
  g610
  (
    n247,
    n66
  );


  buf
  g611
  (
    n269,
    n148
  );


  not
  g612
  (
    n462,
    n130
  );


  not
  g613
  (
    n638,
    n154
  );


  buf
  g614
  (
    n251,
    n34
  );


  not
  g615
  (
    n553,
    n74
  );


  not
  g616
  (
    n592,
    n40
  );


  not
  g617
  (
    n387,
    n154
  );


  not
  g618
  (
    n611,
    n79
  );


  buf
  g619
  (
    n646,
    n144
  );


  buf
  g620
  (
    n373,
    n99
  );


  not
  g621
  (
    n485,
    n105
  );


  not
  g622
  (
    n532,
    n158
  );


  buf
  g623
  (
    n245,
    n55
  );


  buf
  g624
  (
    n464,
    n74
  );


  not
  g625
  (
    n211,
    n63
  );


  buf
  g626
  (
    n435,
    n42
  );


  buf
  g627
  (
    n450,
    n44
  );


  buf
  g628
  (
    n453,
    n129
  );


  buf
  g629
  (
    n237,
    n79
  );


  buf
  g630
  (
    n629,
    n66
  );


  not
  g631
  (
    n465,
    n97
  );


  not
  g632
  (
    n161,
    n128
  );


  not
  g633
  (
    n628,
    n62
  );


  buf
  g634
  (
    n571,
    n152
  );


  buf
  g635
  (
    n598,
    n64
  );


  buf
  g636
  (
    n295,
    n123
  );


  buf
  g637
  (
    n296,
    n107
  );


  buf
  g638
  (
    n188,
    n73
  );


  not
  g639
  (
    n205,
    n88
  );


  not
  g640
  (
    n1448,
    n252
  );


  not
  g641
  (
    n1483,
    n554
  );


  buf
  g642
  (
    n991,
    n188
  );


  buf
  g643
  (
    n910,
    n236
  );


  not
  g644
  (
    n1533,
    n613
  );


  buf
  g645
  (
    n714,
    n266
  );


  buf
  g646
  (
    n1461,
    n316
  );


  not
  g647
  (
    n1040,
    n418
  );


  buf
  g648
  (
    n1260,
    n174
  );


  not
  g649
  (
    n726,
    n231
  );


  buf
  g650
  (
    n1098,
    n367
  );


  buf
  g651
  (
    n1010,
    n471
  );


  buf
  g652
  (
    n984,
    n574
  );


  buf
  g653
  (
    n942,
    n493
  );


  not
  g654
  (
    n948,
    n459
  );


  not
  g655
  (
    n1548,
    n239
  );


  not
  g656
  (
    n674,
    n489
  );


  not
  g657
  (
    n768,
    n171
  );


  not
  g658
  (
    n767,
    n532
  );


  not
  g659
  (
    n1068,
    n602
  );


  not
  g660
  (
    n1002,
    n207
  );


  buf
  g661
  (
    n1388,
    n468
  );


  not
  g662
  (
    n1272,
    n259
  );


  buf
  g663
  (
    n1529,
    n272
  );


  buf
  g664
  (
    n805,
    n352
  );


  not
  g665
  (
    n1380,
    n371
  );


  buf
  g666
  (
    n772,
    n322
  );


  buf
  g667
  (
    n969,
    n193
  );


  not
  g668
  (
    n1417,
    n504
  );


  buf
  g669
  (
    n1556,
    n446
  );


  buf
  g670
  (
    n1309,
    n358
  );


  buf
  g671
  (
    n797,
    n565
  );


  not
  g672
  (
    n1095,
    n340
  );


  not
  g673
  (
    n781,
    n428
  );


  not
  g674
  (
    n1487,
    n515
  );


  buf
  g675
  (
    n1603,
    n524
  );


  buf
  g676
  (
    n1201,
    n503
  );


  not
  g677
  (
    n1554,
    n446
  );


  buf
  g678
  (
    n793,
    n521
  );


  not
  g679
  (
    n1454,
    n360
  );


  not
  g680
  (
    n1072,
    n450
  );


  not
  g681
  (
    n1523,
    n294
  );


  not
  g682
  (
    n1079,
    n257
  );


  buf
  g683
  (
    n848,
    n286
  );


  not
  g684
  (
    n730,
    n241
  );


  not
  g685
  (
    n939,
    n303
  );


  not
  g686
  (
    n1270,
    n327
  );


  buf
  g687
  (
    n981,
    n557
  );


  not
  g688
  (
    n1569,
    n387
  );


  buf
  g689
  (
    n1092,
    n444
  );


  not
  g690
  (
    n1499,
    n384
  );


  not
  g691
  (
    n753,
    n425
  );


  not
  g692
  (
    n784,
    n171
  );


  not
  g693
  (
    n1504,
    n273
  );


  not
  g694
  (
    n1607,
    n488
  );


  buf
  g695
  (
    n1061,
    n221
  );


  buf
  g696
  (
    n699,
    n493
  );


  buf
  g697
  (
    n953,
    n366
  );


  buf
  g698
  (
    n1394,
    n338
  );


  not
  g699
  (
    n1050,
    n458
  );


  not
  g700
  (
    n988,
    n428
  );


  buf
  g701
  (
    n1115,
    n581
  );


  buf
  g702
  (
    n1463,
    n320
  );


  not
  g703
  (
    n1234,
    n431
  );


  not
  g704
  (
    n884,
    n482
  );


  buf
  g705
  (
    n1447,
    n513
  );


  not
  g706
  (
    n1249,
    n407
  );


  not
  g707
  (
    n945,
    n395
  );


  buf
  g708
  (
    n973,
    n440
  );


  not
  g709
  (
    n1525,
    n167
  );


  buf
  g710
  (
    n1042,
    n532
  );


  buf
  g711
  (
    n775,
    n165
  );


  not
  g712
  (
    n1467,
    n231
  );


  buf
  g713
  (
    n1178,
    n422
  );


  buf
  g714
  (
    n1303,
    n321
  );


  buf
  g715
  (
    n1426,
    n245
  );


  not
  g716
  (
    n682,
    n363
  );


  buf
  g717
  (
    n1584,
    n587
  );


  not
  g718
  (
    n1172,
    n581
  );


  buf
  g719
  (
    n1590,
    n317
  );


  not
  g720
  (
    n1104,
    n264
  );


  buf
  g721
  (
    n839,
    n550
  );


  buf
  g722
  (
    n1264,
    n326
  );


  not
  g723
  (
    n1240,
    n415
  );


  not
  g724
  (
    n961,
    n375
  );


  buf
  g725
  (
    n1100,
    n435
  );


  buf
  g726
  (
    n1204,
    n578
  );


  buf
  g727
  (
    n997,
    n442
  );


  not
  g728
  (
    n1610,
    n172
  );


  buf
  g729
  (
    n764,
    n538
  );


  not
  g730
  (
    n1220,
    n592
  );


  not
  g731
  (
    n798,
    n387
  );


  not
  g732
  (
    n941,
    n242
  );


  buf
  g733
  (
    n1352,
    n186
  );


  buf
  g734
  (
    n1030,
    n163
  );


  not
  g735
  (
    n1254,
    n178
  );


  buf
  g736
  (
    n801,
    n502
  );


  buf
  g737
  (
    n1337,
    n482
  );


  buf
  g738
  (
    n1491,
    n465
  );


  buf
  g739
  (
    n1331,
    n380
  );


  buf
  g740
  (
    n1442,
    n240
  );


  not
  g741
  (
    n1642,
    n250
  );


  not
  g742
  (
    n1216,
    n426
  );


  buf
  g743
  (
    n888,
    n549
  );


  not
  g744
  (
    n836,
    n486
  );


  buf
  g745
  (
    n1536,
    n194
  );


  buf
  g746
  (
    n1280,
    n443
  );


  not
  g747
  (
    n1415,
    n611
  );


  not
  g748
  (
    n788,
    n229
  );


  not
  g749
  (
    n1214,
    n556
  );


  not
  g750
  (
    n1118,
    n521
  );


  buf
  g751
  (
    n1592,
    n307
  );


  buf
  g752
  (
    n1205,
    n284
  );


  not
  g753
  (
    n1196,
    n421
  );


  not
  g754
  (
    n1160,
    n296
  );


  not
  g755
  (
    n677,
    n509
  );


  not
  g756
  (
    n956,
    n407
  );


  not
  g757
  (
    n883,
    n585
  );


  buf
  g758
  (
    n1009,
    n430
  );


  buf
  g759
  (
    n1387,
    n523
  );


  not
  g760
  (
    n823,
    n453
  );


  not
  g761
  (
    n739,
    n276
  );


  not
  g762
  (
    n1595,
    n169
  );


  not
  g763
  (
    n680,
    n553
  );


  buf
  g764
  (
    n1456,
    n317
  );


  buf
  g765
  (
    n1408,
    n391
  );


  not
  g766
  (
    n1063,
    n311
  );


  not
  g767
  (
    n1191,
    n170
  );


  not
  g768
  (
    KeyWire_0_31,
    n309
  );


  not
  g769
  (
    n715,
    n396
  );


  not
  g770
  (
    n1086,
    n168
  );


  buf
  g771
  (
    n1598,
    n419
  );


  buf
  g772
  (
    n874,
    n578
  );


  not
  g773
  (
    n1366,
    n466
  );


  buf
  g774
  (
    n1000,
    n479
  );


  not
  g775
  (
    n1370,
    n329
  );


  not
  g776
  (
    n1526,
    n361
  );


  not
  g777
  (
    KeyWire_0_15,
    n161
  );


  buf
  g778
  (
    n1596,
    n249
  );


  not
  g779
  (
    n1014,
    n566
  );


  buf
  g780
  (
    n935,
    n367
  );


  buf
  g781
  (
    n800,
    n363
  );


  buf
  g782
  (
    n1403,
    n588
  );


  not
  g783
  (
    n1545,
    n454
  );


  not
  g784
  (
    n806,
    n594
  );


  not
  g785
  (
    n1297,
    n378
  );


  not
  g786
  (
    n815,
    n189
  );


  buf
  g787
  (
    n887,
    n362
  );


  buf
  g788
  (
    n838,
    n353
  );


  buf
  g789
  (
    n1427,
    n422
  );


  not
  g790
  (
    n708,
    n192
  );


  buf
  g791
  (
    n1335,
    n496
  );


  not
  g792
  (
    n958,
    n545
  );


  not
  g793
  (
    n1047,
    n394
  );


  not
  g794
  (
    n1353,
    n568
  );


  not
  g795
  (
    n1345,
    n279
  );


  buf
  g796
  (
    n865,
    n345
  );


  buf
  g797
  (
    n1235,
    n363
  );


  buf
  g798
  (
    n742,
    n477
  );


  not
  g799
  (
    n1039,
    n259
  );


  buf
  g800
  (
    n1146,
    n423
  );


  not
  g801
  (
    n870,
    n422
  );


  buf
  g802
  (
    n828,
    n230
  );


  not
  g803
  (
    n1507,
    n589
  );


  buf
  g804
  (
    KeyWire_0_12,
    n414
  );


  not
  g805
  (
    n1517,
    n467
  );


  buf
  g806
  (
    n1181,
    n183
  );


  not
  g807
  (
    n1099,
    n443
  );


  buf
  g808
  (
    n1080,
    n162
  );


  not
  g809
  (
    n684,
    n216
  );


  buf
  g810
  (
    n1211,
    n442
  );


  buf
  g811
  (
    n1469,
    n608
  );


  not
  g812
  (
    n925,
    n552
  );


  buf
  g813
  (
    n1257,
    n202
  );


  buf
  g814
  (
    n1381,
    n382
  );


  not
  g815
  (
    n1488,
    n283
  );


  not
  g816
  (
    n1357,
    n216
  );


  buf
  g817
  (
    n1559,
    n559
  );


  not
  g818
  (
    n1025,
    n249
  );


  buf
  g819
  (
    n1094,
    n505
  );


  not
  g820
  (
    n922,
    n614
  );


  not
  g821
  (
    n713,
    n168
  );


  buf
  g822
  (
    n867,
    n602
  );


  not
  g823
  (
    n1489,
    n198
  );


  not
  g824
  (
    n696,
    n347
  );


  buf
  g825
  (
    n814,
    n283
  );


  not
  g826
  (
    n1550,
    n203
  );


  buf
  g827
  (
    n729,
    n370
  );


  not
  g828
  (
    n685,
    n492
  );


  not
  g829
  (
    n850,
    n603
  );


  buf
  g830
  (
    n980,
    n546
  );


  not
  g831
  (
    n1321,
    n457
  );


  not
  g832
  (
    n852,
    n564
  );


  not
  g833
  (
    n1601,
    n310
  );


  not
  g834
  (
    n1466,
    n370
  );


  buf
  g835
  (
    n1164,
    n279
  );


  not
  g836
  (
    n1162,
    n329
  );


  not
  g837
  (
    n1210,
    n595
  );


  not
  g838
  (
    n1630,
    n379
  );


  buf
  g839
  (
    n754,
    n343
  );


  buf
  g840
  (
    n1605,
    n341
  );


  buf
  g841
  (
    n782,
    n460
  );


  buf
  g842
  (
    n1011,
    n579
  );


  buf
  g843
  (
    n1486,
    n268
  );


  buf
  g844
  (
    n1473,
    n557
  );


  buf
  g845
  (
    n1393,
    n397
  );


  buf
  g846
  (
    n733,
    n559
  );


  not
  g847
  (
    n694,
    n469
  );


  not
  g848
  (
    n999,
    n480
  );


  not
  g849
  (
    n1295,
    n542
  );


  not
  g850
  (
    n1213,
    n469
  );


  not
  g851
  (
    n872,
    n178
  );


  not
  g852
  (
    n735,
    n471
  );


  buf
  g853
  (
    n1446,
    n378
  );


  buf
  g854
  (
    n1476,
    n474
  );


  buf
  g855
  (
    n1421,
    n427
  );


  buf
  g856
  (
    n902,
    n163
  );


  not
  g857
  (
    n1036,
    n534
  );


  not
  g858
  (
    n721,
    n447
  );


  buf
  g859
  (
    n1022,
    n164
  );


  not
  g860
  (
    n1278,
    n518
  );


  buf
  g861
  (
    n1096,
    n452
  );


  not
  g862
  (
    n1562,
    n227
  );


  buf
  g863
  (
    n1119,
    n487
  );


  buf
  g864
  (
    n1589,
    n361
  );


  buf
  g865
  (
    n1465,
    n166
  );


  not
  g866
  (
    n681,
    n399
  );


  not
  g867
  (
    n1378,
    n517
  );


  buf
  g868
  (
    n1224,
    n341
  );


  not
  g869
  (
    n692,
    n444
  );


  buf
  g870
  (
    n1565,
    n319
  );


  buf
  g871
  (
    n691,
    n498
  );


  not
  g872
  (
    n695,
    n535
  );


  buf
  g873
  (
    n1147,
    n249
  );


  buf
  g874
  (
    n1409,
    n455
  );


  not
  g875
  (
    n1026,
    n529
  );


  buf
  g876
  (
    n1512,
    n584
  );


  buf
  g877
  (
    n1665,
    n551
  );


  not
  g878
  (
    n1247,
    n486
  );


  not
  g879
  (
    n1308,
    n464
  );


  buf
  g880
  (
    n1246,
    n600
  );


  buf
  g881
  (
    n932,
    n212
  );


  buf
  g882
  (
    n763,
    n524
  );


  not
  g883
  (
    n1611,
    n340
  );


  buf
  g884
  (
    n987,
    n311
  );


  not
  g885
  (
    n1193,
    n573
  );


  buf
  g886
  (
    n1074,
    n348
  );


  buf
  g887
  (
    n1142,
    n456
  );


  buf
  g888
  (
    n1651,
    n214
  );


  buf
  g889
  (
    n975,
    n529
  );


  not
  g890
  (
    n1007,
    n504
  );


  not
  g891
  (
    n1399,
    n357
  );


  not
  g892
  (
    n1244,
    n501
  );


  buf
  g893
  (
    n1154,
    n450
  );


  not
  g894
  (
    n1561,
    n270
  );


  buf
  g895
  (
    n968,
    n254
  );


  buf
  g896
  (
    n1623,
    n608
  );


  buf
  g897
  (
    n1571,
    n518
  );


  buf
  g898
  (
    n1612,
    n196
  );


  buf
  g899
  (
    n1511,
    n561
  );


  buf
  g900
  (
    n847,
    n165
  );


  not
  g901
  (
    n849,
    n221
  );


  not
  g902
  (
    n1549,
    n252
  );


  not
  g903
  (
    n1481,
    n437
  );


  buf
  g904
  (
    n1645,
    n421
  );


  not
  g905
  (
    n1636,
    n313
  );


  buf
  g906
  (
    n1171,
    n335
  );


  buf
  g907
  (
    n1141,
    n165
  );


  not
  g908
  (
    n1413,
    n297
  );


  buf
  g909
  (
    n1626,
    n608
  );


  buf
  g910
  (
    n1315,
    n323
  );


  buf
  g911
  (
    n1663,
    n545
  );


  not
  g912
  (
    n1444,
    n614
  );


  not
  g913
  (
    n718,
    n196
  );


  buf
  g914
  (
    n946,
    n470
  );


  buf
  g915
  (
    n1156,
    n300
  );


  not
  g916
  (
    n740,
    n456
  );


  buf
  g917
  (
    n1459,
    n519
  );


  buf
  g918
  (
    n1312,
    n169
  );


  not
  g919
  (
    n747,
    n598
  );


  not
  g920
  (
    n936,
    n447
  );


  not
  g921
  (
    n1356,
    n507
  );


  not
  g922
  (
    n1343,
    n398
  );


  not
  g923
  (
    n1043,
    n226
  );


  buf
  g924
  (
    n1236,
    n381
  );


  not
  g925
  (
    n1208,
    n174
  );


  not
  g926
  (
    n1051,
    n308
  );


  buf
  g927
  (
    n1306,
    n614
  );


  buf
  g928
  (
    n875,
    n517
  );


  buf
  g929
  (
    n1258,
    n466
  );


  not
  g930
  (
    n1631,
    n596
  );


  buf
  g931
  (
    n1480,
    n522
  );


  buf
  g932
  (
    n1062,
    n184
  );


  buf
  g933
  (
    n1342,
    n227
  );


  not
  g934
  (
    n1494,
    n263
  );


  not
  g935
  (
    n1229,
    n523
  );


  buf
  g936
  (
    n856,
    n541
  );


  not
  g937
  (
    n1023,
    n572
  );


  buf
  g938
  (
    n1155,
    n485
  );


  buf
  g939
  (
    n1431,
    n244
  );


  buf
  g940
  (
    n1212,
    n233
  );


  not
  g941
  (
    n1652,
    n546
  );


  not
  g942
  (
    KeyWire_0_27,
    n416
  );


  not
  g943
  (
    n1033,
    n276
  );


  not
  g944
  (
    n791,
    n243
  );


  buf
  g945
  (
    n822,
    n177
  );


  not
  g946
  (
    n921,
    n209
  );


  not
  g947
  (
    n812,
    n459
  );


  buf
  g948
  (
    n1639,
    n449
  );


  not
  g949
  (
    n1316,
    n359
  );


  not
  g950
  (
    n1532,
    n302
  );


  not
  g951
  (
    n1024,
    n386
  );


  not
  g952
  (
    n900,
    n575
  );


  not
  g953
  (
    n762,
    n551
  );


  buf
  g954
  (
    n985,
    n466
  );


  buf
  g955
  (
    n982,
    n569
  );


  buf
  g956
  (
    n996,
    n431
  );


  buf
  g957
  (
    n1617,
    n331
  );


  not
  g958
  (
    n1372,
    n437
  );


  not
  g959
  (
    n1551,
    n413
  );


  not
  g960
  (
    n893,
    n469
  );


  buf
  g961
  (
    n769,
    n406
  );


  not
  g962
  (
    n1434,
    n541
  );


  buf
  g963
  (
    n1384,
    n586
  );


  not
  g964
  (
    n1328,
    n278
  );


  buf
  g965
  (
    n1097,
    n204
  );


  not
  g966
  (
    n1509,
    n179
  );


  buf
  g967
  (
    n1262,
    n217
  );


  buf
  g968
  (
    n690,
    n230
  );


  buf
  g969
  (
    n746,
    n483
  );


  buf
  g970
  (
    n1322,
    n273
  );


  not
  g971
  (
    n821,
    n429
  );


  buf
  g972
  (
    n1217,
    n183
  );


  not
  g973
  (
    n1576,
    n542
  );


  not
  g974
  (
    n977,
    n458
  );


  not
  g975
  (
    n1664,
    n397
  );


  buf
  g976
  (
    n760,
    n262
  );


  buf
  g977
  (
    n717,
    n559
  );


  not
  g978
  (
    n851,
    n534
  );


  not
  g979
  (
    n871,
    n584
  );


  buf
  g980
  (
    n860,
    n285
  );


  buf
  g981
  (
    n892,
    n395
  );


  not
  g982
  (
    n1410,
    n491
  );


  buf
  g983
  (
    n1613,
    n347
  );


  not
  g984
  (
    n1505,
    n248
  );


  not
  g985
  (
    n1064,
    n376
  );


  not
  g986
  (
    n845,
    n241
  );


  buf
  g987
  (
    n777,
    n175
  );


  buf
  g988
  (
    n1660,
    n320
  );


  not
  g989
  (
    n1304,
    n530
  );


  not
  g990
  (
    n783,
    n347
  );


  buf
  g991
  (
    n679,
    n300
  );


  buf
  g992
  (
    n1302,
    n304
  );


  buf
  g993
  (
    n1527,
    n186
  );


  not
  g994
  (
    n1256,
    n288
  );


  buf
  g995
  (
    n878,
    n577
  );


  buf
  g996
  (
    n928,
    n552
  );


  not
  g997
  (
    n700,
    n275
  );


  buf
  g998
  (
    n1150,
    n383
  );


  buf
  g999
  (
    n737,
    n193
  );


  buf
  g1000
  (
    n1075,
    n506
  );


  not
  g1001
  (
    n1519,
    n312
  );


  buf
  g1002
  (
    n1398,
    n188
  );


  not
  g1003
  (
    n1563,
    n585
  );


  buf
  g1004
  (
    n1127,
    n409
  );


  buf
  g1005
  (
    n903,
    n506
  );


  not
  g1006
  (
    n873,
    n295
  );


  not
  g1007
  (
    n1305,
    n548
  );


  buf
  g1008
  (
    n1169,
    n463
  );


  buf
  g1009
  (
    n1567,
    n174
  );


  buf
  g1010
  (
    n794,
    n538
  );


  buf
  g1011
  (
    n1558,
    n264
  );


  buf
  g1012
  (
    n869,
    n581
  );


  not
  g1013
  (
    n1177,
    n491
  );


  not
  g1014
  (
    n1471,
    n595
  );


  buf
  g1015
  (
    n1404,
    n412
  );


  not
  g1016
  (
    n1553,
    n462
  );


  buf
  g1017
  (
    n974,
    n472
  );


  buf
  g1018
  (
    n1006,
    n565
  );


  not
  g1019
  (
    n1130,
    n544
  );


  buf
  g1020
  (
    n1547,
    n535
  );


  not
  g1021
  (
    n1069,
    n420
  );


  buf
  g1022
  (
    n859,
    n457
  );


  buf
  g1023
  (
    n1005,
    n410
  );


  not
  g1024
  (
    n894,
    n375
  );


  not
  g1025
  (
    n837,
    n171
  );


  buf
  g1026
  (
    n811,
    n207
  );


  not
  g1027
  (
    n898,
    n487
  );


  buf
  g1028
  (
    n1327,
    n317
  );


  not
  g1029
  (
    n962,
    n232
  );


  not
  g1030
  (
    n1425,
    n282
  );


  buf
  g1031
  (
    n1149,
    n528
  );


  not
  g1032
  (
    n1555,
    n289
  );


  not
  g1033
  (
    n790,
    n208
  );


  buf
  g1034
  (
    n1255,
    n341
  );


  not
  g1035
  (
    n722,
    n512
  );


  not
  g1036
  (
    n1503,
    n296
  );


  not
  g1037
  (
    n1583,
    n434
  );


  not
  g1038
  (
    n1060,
    n571
  );


  not
  g1039
  (
    n1445,
    n318
  );


  not
  g1040
  (
    n1318,
    n235
  );


  buf
  g1041
  (
    n1581,
    n208
  );


  buf
  g1042
  (
    n1641,
    n401
  );


  buf
  g1043
  (
    n1239,
    n180
  );


  not
  g1044
  (
    n998,
    n202
  );


  buf
  g1045
  (
    n1338,
    n297
  );


  not
  g1046
  (
    n885,
    n555
  );


  not
  g1047
  (
    n832,
    n602
  );


  not
  g1048
  (
    n796,
    n323
  );


  buf
  g1049
  (
    n1317,
    n606
  );


  buf
  g1050
  (
    n926,
    n247
  );


  not
  g1051
  (
    n705,
    n420
  );


  buf
  g1052
  (
    n1105,
    n246
  );


  not
  g1053
  (
    n1385,
    n419
  );


  buf
  g1054
  (
    n1449,
    n427
  );


  not
  g1055
  (
    n1046,
    n200
  );


  buf
  g1056
  (
    n944,
    n433
  );


  buf
  g1057
  (
    n864,
    n316
  );


  not
  g1058
  (
    n1055,
    n464
  );


  buf
  g1059
  (
    n846,
    n221
  );


  buf
  g1060
  (
    n786,
    n554
  );


  not
  g1061
  (
    n1112,
    n612
  );


  not
  g1062
  (
    n830,
    n440
  );


  buf
  g1063
  (
    n1090,
    n338
  );


  not
  g1064
  (
    n1339,
    n432
  );


  buf
  g1065
  (
    n770,
    n440
  );


  buf
  g1066
  (
    n857,
    n335
  );


  buf
  g1067
  (
    n1197,
    n307
  );


  buf
  g1068
  (
    n1114,
    n542
  );


  buf
  g1069
  (
    n1450,
    n484
  );


  buf
  g1070
  (
    n1542,
    n607
  );


  not
  g1071
  (
    n914,
    n351
  );


  buf
  g1072
  (
    KeyWire_0_5,
    n260
  );


  buf
  g1073
  (
    n1518,
    n593
  );


  buf
  g1074
  (
    n1238,
    n571
  );


  not
  g1075
  (
    n1326,
    n556
  );


  not
  g1076
  (
    n675,
    n426
  );


  buf
  g1077
  (
    n923,
    n390
  );


  buf
  g1078
  (
    n1110,
    n203
  );


  buf
  g1079
  (
    n994,
    n562
  );


  not
  g1080
  (
    n1233,
    n604
  );


  buf
  g1081
  (
    n1502,
    n327
  );


  buf
  g1082
  (
    n1606,
    n348
  );


  not
  g1083
  (
    n1076,
    n214
  );


  buf
  g1084
  (
    n1520,
    n293
  );


  not
  g1085
  (
    n787,
    n276
  );


  buf
  g1086
  (
    n954,
    n238
  );


  buf
  g1087
  (
    n1492,
    n521
  );


  not
  g1088
  (
    n707,
    n229
  );


  buf
  g1089
  (
    n917,
    n475
  );


  buf
  g1090
  (
    n1027,
    n315
  );


  not
  g1091
  (
    n1460,
    n377
  );


  not
  g1092
  (
    n1510,
    n393
  );


  not
  g1093
  (
    n1170,
    n445
  );


  buf
  g1094
  (
    n1593,
    n214
  );


  buf
  g1095
  (
    n938,
    n483
  );


  not
  g1096
  (
    n1194,
    n471
  );


  buf
  g1097
  (
    n1325,
    n311
  );


  not
  g1098
  (
    n1673,
    n480
  );


  not
  g1099
  (
    n1332,
    n180
  );


  buf
  g1100
  (
    n1521,
    n331
  );


  not
  g1101
  (
    n731,
    n268
  );


  not
  g1102
  (
    n1279,
    n293
  );


  buf
  g1103
  (
    n1107,
    n371
  );


  not
  g1104
  (
    n1624,
    n166
  );


  not
  g1105
  (
    n1412,
    n250
  );


  buf
  g1106
  (
    n1018,
    n299
  );


  buf
  g1107
  (
    n1291,
    n307
  );


  buf
  g1108
  (
    n1324,
    n488
  );


  not
  g1109
  (
    n686,
    n452
  );


  not
  g1110
  (
    n1157,
    n355
  );


  buf
  g1111
  (
    n1198,
    n309
  );


  buf
  g1112
  (
    n756,
    n440
  );


  buf
  g1113
  (
    n1057,
    n163
  );


  not
  g1114
  (
    n1109,
    n439
  );


  not
  g1115
  (
    n1031,
    n609
  );


  not
  g1116
  (
    n1591,
    n333
  );


  buf
  g1117
  (
    n1666,
    n436
  );


  buf
  g1118
  (
    n1085,
    n354
  );


  not
  g1119
  (
    n930,
    n377
  );


  buf
  g1120
  (
    n1437,
    n373
  );


  not
  g1121
  (
    n780,
    n306
  );


  not
  g1122
  (
    n1129,
    n613
  );


  buf
  g1123
  (
    n929,
    n361
  );


  buf
  g1124
  (
    n843,
    n222
  );


  not
  g1125
  (
    n698,
    n224
  );


  buf
  g1126
  (
    n1367,
    n314
  );


  buf
  g1127
  (
    n1541,
    n258
  );


  not
  g1128
  (
    n1566,
    n609
  );


  buf
  g1129
  (
    n913,
    n289
  );


  buf
  g1130
  (
    n947,
    n600
  );


  buf
  g1131
  (
    n895,
    n210
  );


  not
  g1132
  (
    n952,
    n430
  );


  not
  g1133
  (
    n906,
    n389
  );


  buf
  g1134
  (
    n1379,
    n477
  );


  buf
  g1135
  (
    n1377,
    n444
  );


  buf
  g1136
  (
    n1106,
    n414
  );


  buf
  g1137
  (
    n1165,
    n303
  );


  not
  g1138
  (
    n1362,
    n288
  );


  not
  g1139
  (
    n841,
    n597
  );


  buf
  g1140
  (
    n1081,
    n540
  );


  not
  g1141
  (
    n1029,
    n201
  );


  not
  g1142
  (
    n1470,
    n364
  );


  not
  g1143
  (
    n1614,
    n514
  );


  not
  g1144
  (
    n1134,
    n343
  );


  buf
  g1145
  (
    n1102,
    n534
  );


  not
  g1146
  (
    n1311,
    n257
  );


  buf
  g1147
  (
    n1273,
    n590
  );


  not
  g1148
  (
    n1669,
    n590
  );


  buf
  g1149
  (
    n978,
    n590
  );


  not
  g1150
  (
    n1364,
    n478
  );


  buf
  g1151
  (
    n758,
    n244
  );


  buf
  g1152
  (
    n810,
    n436
  );


  not
  g1153
  (
    n1292,
    n300
  );


  buf
  g1154
  (
    n1203,
    n297
  );


  not
  g1155
  (
    n1375,
    n225
  );


  buf
  g1156
  (
    n1199,
    n310
  );


  not
  g1157
  (
    n972,
    n391
  );


  not
  g1158
  (
    n1135,
    n607
  );


  buf
  g1159
  (
    n889,
    n237
  );


  buf
  g1160
  (
    n1646,
    n421
  );


  buf
  g1161
  (
    n1406,
    n319
  );


  buf
  g1162
  (
    n1032,
    n315
  );


  not
  g1163
  (
    n1088,
    n588
  );


  buf
  g1164
  (
    n1493,
    n549
  );


  not
  g1165
  (
    n1649,
    n355
  );


  buf
  g1166
  (
    n1298,
    n277
  );


  not
  g1167
  (
    n1355,
    n330
  );


  not
  g1168
  (
    n711,
    n373
  );


  not
  g1169
  (
    n1158,
    n369
  );


  not
  g1170
  (
    n795,
    n224
  );


  buf
  g1171
  (
    n1552,
    n202
  );


  buf
  g1172
  (
    n789,
    n228
  );


  not
  g1173
  (
    n1346,
    n563
  );


  buf
  g1174
  (
    n840,
    n298
  );


  not
  g1175
  (
    n1560,
    n414
  );


  not
  g1176
  (
    n1168,
    n278
  );


  buf
  g1177
  (
    n1139,
    n462
  );


  not
  g1178
  (
    n1522,
    n281
  );


  buf
  g1179
  (
    n743,
    n334
  );


  buf
  g1180
  (
    n1052,
    n450
  );


  buf
  g1181
  (
    n1478,
    n220
  );


  buf
  g1182
  (
    n1428,
    n573
  );


  buf
  g1183
  (
    n1263,
    n334
  );


  not
  g1184
  (
    n1245,
    n281
  );


  buf
  g1185
  (
    n1637,
    n511
  );


  buf
  g1186
  (
    n809,
    n170
  );


  buf
  g1187
  (
    n1251,
    n567
  );


  not
  g1188
  (
    n899,
    n402
  );


  buf
  g1189
  (
    n879,
    n509
  );


  buf
  g1190
  (
    n1633,
    n164
  );


  not
  g1191
  (
    n725,
    n357
  );


  buf
  g1192
  (
    n1294,
    n500
  );


  not
  g1193
  (
    n1574,
    n580
  );


  not
  g1194
  (
    n757,
    n515
  );


  buf
  g1195
  (
    n1293,
    n548
  );


  buf
  g1196
  (
    n1041,
    n500
  );


  buf
  g1197
  (
    n1058,
    n161
  );


  buf
  g1198
  (
    n826,
    n222
  );


  not
  g1199
  (
    n891,
    n315
  );


  not
  g1200
  (
    n1622,
    n507
  );


  buf
  g1201
  (
    n955,
    n243
  );


  buf
  g1202
  (
    n1128,
    n482
  );


  not
  g1203
  (
    n1200,
    n390
  );


  not
  g1204
  (
    n1453,
    n238
  );


  not
  g1205
  (
    n1126,
    n383
  );


  not
  g1206
  (
    n728,
    n342
  );


  buf
  g1207
  (
    n723,
    n442
  );


  buf
  g1208
  (
    n741,
    n354
  );


  not
  g1209
  (
    n890,
    n605
  );


  not
  g1210
  (
    n755,
    n368
  );


  not
  g1211
  (
    n1422,
    n521
  );


  buf
  g1212
  (
    n1537,
    n401
  );


  not
  g1213
  (
    n1621,
    n574
  );


  not
  g1214
  (
    n877,
    n199
  );


  buf
  g1215
  (
    n1620,
    n589
  );


  buf
  g1216
  (
    n1336,
    n547
  );


  not
  g1217
  (
    n1084,
    n372
  );


  not
  g1218
  (
    n927,
    n246
  );


  buf
  g1219
  (
    n710,
    n480
  );


  buf
  g1220
  (
    n1455,
    n197
  );


  not
  g1221
  (
    n1059,
    n604
  );


  not
  g1222
  (
    n1661,
    n284
  );


  not
  g1223
  (
    n1373,
    n368
  );


  buf
  g1224
  (
    n862,
    n599
  );


  buf
  g1225
  (
    n1440,
    n336
  );


  buf
  g1226
  (
    n1501,
    n218
  );


  not
  g1227
  (
    n1125,
    n360
  );


  not
  g1228
  (
    n1137,
    n526
  );


  not
  g1229
  (
    n986,
    n290
  );


  not
  g1230
  (
    n829,
    n191
  );


  buf
  g1231
  (
    n886,
    n554
  );


  buf
  g1232
  (
    n1320,
    n563
  );


  buf
  g1233
  (
    n949,
    n573
  );


  not
  g1234
  (
    n1121,
    n527
  );


  buf
  g1235
  (
    n963,
    n529
  );


  not
  g1236
  (
    n1190,
    n331
  );


  buf
  g1237
  (
    n1658,
    n439
  );


  not
  g1238
  (
    n1390,
    n384
  );


  buf
  g1239
  (
    n1111,
    n403
  );


  buf
  g1240
  (
    n1082,
    n269
  );


  buf
  g1241
  (
    n1540,
    n530
  );


  buf
  g1242
  (
    n727,
    n444
  );


  not
  g1243
  (
    n1508,
    n372
  );


  buf
  g1244
  (
    n785,
    n487
  );


  buf
  g1245
  (
    n1056,
    n292
  );


  buf
  g1246
  (
    n1116,
    n348
  );


  not
  g1247
  (
    n1180,
    n270
  );


  buf
  g1248
  (
    n1575,
    n339
  );


  not
  g1249
  (
    n761,
    n525
  );


  not
  g1250
  (
    n1516,
    n221
  );


  not
  g1251
  (
    n950,
    n324
  );


  not
  g1252
  (
    n817,
    n450
  );


  buf
  g1253
  (
    n1451,
    n347
  );


  not
  g1254
  (
    n1414,
    n226
  );


  not
  g1255
  (
    n1189,
    n316
  );


  buf
  g1256
  (
    n776,
    n472
  );


  buf
  g1257
  (
    n1365,
    n229
  );


  not
  g1258
  (
    n1012,
    n518
  );


  not
  g1259
  (
    n964,
    n161
  );


  buf
  g1260
  (
    n1640,
    n383
  );


  not
  g1261
  (
    n1654,
    n520
  );


  buf
  g1262
  (
    n683,
    n382
  );


  not
  g1263
  (
    n1475,
    n386
  );


  buf
  g1264
  (
    n1392,
    n199
  );


  not
  g1265
  (
    n1672,
    n553
  );


  buf
  g1266
  (
    n1275,
    n470
  );


  buf
  g1267
  (
    n1383,
    n345
  );


  not
  g1268
  (
    n1344,
    n226
  );


  buf
  g1269
  (
    n1635,
    n201
  );


  buf
  g1270
  (
    n1604,
    n298
  );


  not
  g1271
  (
    n855,
    n424
  );


  not
  g1272
  (
    n1267,
    n596
  );


  not
  g1273
  (
    n918,
    n228
  );


  buf
  g1274
  (
    n1073,
    n423
  );


  buf
  g1275
  (
    n1250,
    n472
  );


  buf
  g1276
  (
    n792,
    n591
  );


  not
  g1277
  (
    n1230,
    n205
  );


  not
  g1278
  (
    n1215,
    n419
  );


  not
  g1279
  (
    n676,
    n555
  );


  not
  g1280
  (
    n1144,
    n403
  );


  not
  g1281
  (
    n1391,
    n290
  );


  buf
  g1282
  (
    n1538,
    n433
  );


  buf
  g1283
  (
    n701,
    n427
  );


  not
  g1284
  (
    n803,
    n219
  );


  not
  g1285
  (
    n807,
    n583
  );


  buf
  g1286
  (
    n1578,
    n456
  );


  not
  g1287
  (
    n1066,
    n251
  );


  buf
  g1288
  (
    n1227,
    n319
  );


  buf
  g1289
  (
    n702,
    n184
  );


  buf
  g1290
  (
    n1382,
    n531
  );


  not
  g1291
  (
    n1019,
    n415
  );


  not
  g1292
  (
    n1496,
    n540
  );


  buf
  g1293
  (
    n1531,
    n358
  );


  not
  g1294
  (
    n1071,
    n575
  );


  not
  g1295
  (
    n706,
    n547
  );


  not
  g1296
  (
    n1580,
    n497
  );


  buf
  g1297
  (
    n1218,
    n567
  );


  not
  g1298
  (
    n989,
    n606
  );


  not
  g1299
  (
    n1585,
    n484
  );


  buf
  g1300
  (
    n678,
    n262
  );


  buf
  g1301
  (
    n1586,
    n361
  );


  not
  g1302
  (
    n749,
    n568
  );


  not
  g1303
  (
    n1432,
    n234
  );


  buf
  g1304
  (
    n1490,
    n187
  );


  buf
  g1305
  (
    n1396,
    n344
  );


  not
  g1306
  (
    n1016,
    n531
  );


  not
  g1307
  (
    n736,
    n349
  );


  not
  g1308
  (
    n1535,
    n295
  );


  buf
  g1309
  (
    n1323,
    n299
  );


  not
  g1310
  (
    n959,
    n494
  );


  buf
  g1311
  (
    n1588,
    n457
  );


  not
  g1312
  (
    n1619,
    n301
  );


  buf
  g1313
  (
    n1120,
    n234
  );


  not
  g1314
  (
    n1655,
    n516
  );


  buf
  g1315
  (
    n1138,
    n252
  );


  buf
  g1316
  (
    n1310,
    n579
  );


  not
  g1317
  (
    n1600,
    n260
  );


  not
  g1318
  (
    n1221,
    n407
  );


  buf
  g1319
  (
    n1484,
    n499
  );


  buf
  g1320
  (
    n1330,
    n176
  );


  not
  g1321
  (
    n1259,
    n430
  );


  not
  g1322
  (
    n1159,
    n271
  );


  not
  g1323
  (
    n751,
    n537
  );


  not
  g1324
  (
    n1667,
    n441
  );


  not
  g1325
  (
    n990,
    n455
  );


  not
  g1326
  (
    n1288,
    n449
  );


  not
  g1327
  (
    n1418,
    n585
  );


  not
  g1328
  (
    n882,
    n559
  );


  not
  g1329
  (
    n738,
    n507
  );


  buf
  g1330
  (
    n1132,
    n304
  );


  buf
  g1331
  (
    n858,
    n167
  );


  buf
  g1332
  (
    n734,
    n301
  );


  buf
  g1333
  (
    n1618,
    n325
  );


  not
  g1334
  (
    n1638,
    n412
  );


  not
  g1335
  (
    n1354,
    n251
  );


  not
  g1336
  (
    KeyWire_0_1,
    n215
  );


  not
  g1337
  (
    n1017,
    n182
  );


  buf
  g1338
  (
    n1103,
    n400
  );


  not
  g1339
  (
    n1281,
    n490
  );


  not
  g1340
  (
    n1188,
    n490
  );


  buf
  g1341
  (
    n1539,
    n528
  );


  buf
  g1342
  (
    n1004,
    n226
  );


  not
  g1343
  (
    n1307,
    n190
  );


  not
  g1344
  (
    n1438,
    n268
  );


  not
  g1345
  (
    n909,
    n367
  );


  buf
  g1346
  (
    n1087,
    n593
  );


  not
  g1347
  (
    n1472,
    n546
  );


  not
  g1348
  (
    n966,
    n552
  );


  not
  g1349
  (
    n965,
    n486
  );


  not
  g1350
  (
    n802,
    n219
  );


  buf
  g1351
  (
    n1405,
    n341
  );


  not
  g1352
  (
    n1319,
    n181
  );


  not
  g1353
  (
    n1008,
    n253
  );


  buf
  g1354
  (
    n960,
    n338
  );


  buf
  g1355
  (
    n861,
    n432
  );


  not
  g1356
  (
    n1241,
    n255
  );


  not
  g1357
  (
    n1287,
    n239
  );


  not
  g1358
  (
    n1044,
    n381
  );


  not
  g1359
  (
    n940,
    n360
  );


  not
  g1360
  (
    n1300,
    n592
  );


  not
  g1361
  (
    n844,
    n560
  );


  not
  g1362
  (
    n1163,
    n594
  );


  buf
  g1363
  (
    n1500,
    n284
  );


  buf
  g1364
  (
    n1368,
    n538
  );


  buf
  g1365
  (
    n1219,
    n220
  );


  not
  g1366
  (
    n1334,
    n425
  );


  not
  g1367
  (
    n1482,
    n558
  );


  buf
  g1368
  (
    n1513,
    n265
  );


  nor
  g1369
  (
    n1648,
    n536,
    n234,
    n275,
    n597
  );


  nand
  g1370
  (
    n804,
    n424,
    n469,
    n218,
    n529
  );


  xor
  g1371
  (
    n1433,
    n277,
    n267,
    n296,
    n550
  );


  and
  g1372
  (
    n1237,
    n410,
    n267,
    n583,
    n335
  );


  nor
  g1373
  (
    n1093,
    n233,
    n253,
    n438,
    n566
  );


  and
  g1374
  (
    n881,
    n582,
    n452,
    n416,
    n577
  );


  or
  g1375
  (
    n1021,
    n401,
    n210,
    n567,
    n402
  );


  and
  g1376
  (
    n1643,
    n261,
    n222,
    n313,
    n560
  );


  nand
  g1377
  (
    n773,
    n439,
    n293,
    n526,
    n206
  );


  nand
  g1378
  (
    n1173,
    n342,
    n482,
    n385,
    n387
  );


  and
  g1379
  (
    n1632,
    n471,
    n459,
    n238,
    n568
  );


  xor
  g1380
  (
    n1458,
    n405,
    n612,
    n483,
    n169
  );


  xor
  g1381
  (
    n1101,
    n270,
    n498,
    n527,
    n530
  );


  xnor
  g1382
  (
    n1145,
    n412,
    n611,
    n245,
    n569
  );


  nand
  g1383
  (
    n1644,
    n397,
    n324,
    n387,
    n512
  );


  xor
  g1384
  (
    n1285,
    n373,
    n403,
    n582,
    n481
  );


  nor
  g1385
  (
    n1131,
    n588,
    n231,
    n364,
    n327
  );


  and
  g1386
  (
    n1546,
    n264,
    n506,
    n428,
    n610
  );


  or
  g1387
  (
    n1282,
    n558,
    n280,
    n173,
    n376
  );


  or
  g1388
  (
    n1261,
    n583,
    n498,
    n494,
    n176
  );


  xor
  g1389
  (
    n911,
    n326,
    n598,
    n544,
    n537
  );


  or
  g1390
  (
    n1077,
    n280,
    n437,
    n584,
    n374
  );


  xnor
  g1391
  (
    n759,
    n372,
    n249,
    n301,
    n185
  );


  xnor
  g1392
  (
    n1477,
    n464,
    n575,
    n603,
    n474
  );


  xor
  g1393
  (
    n1564,
    n369,
    n304,
    n481,
    n261
  );


  nand
  g1394
  (
    n1597,
    n287,
    n350,
    n265,
    n526
  );


  and
  g1395
  (
    n732,
    n500,
    n351,
    n547,
    n555
  );


  xor
  g1396
  (
    n1340,
    n368,
    n558,
    n378,
    n458
  );


  or
  g1397
  (
    n750,
    n356,
    n490,
    n298,
    n320
  );


  and
  g1398
  (
    n1514,
    n195,
    n217,
    n454,
    n514
  );


  xor
  g1399
  (
    n1123,
    n260,
    n313,
    n461,
    n417
  );


  xor
  g1400
  (
    n1045,
    n355,
    n253,
    n548,
    n272
  );


  and
  g1401
  (
    n1329,
    n411,
    n385,
    n369,
    n212
  );


  or
  g1402
  (
    n689,
    n494,
    n275,
    n549,
    n445
  );


  nand
  g1403
  (
    n745,
    n532,
    n180,
    n202,
    n173
  );


  or
  g1404
  (
    n1151,
    n478,
    n478,
    n308,
    n408
  );


  nand
  g1405
  (
    n752,
    n204,
    n517,
    n533,
    n223
  );


  nor
  g1406
  (
    n1226,
    n196,
    n435,
    n603,
    n236
  );


  or
  g1407
  (
    n748,
    n199,
    n348,
    n511,
    n175
  );


  nand
  g1408
  (
    n1192,
    n337,
    n459,
    n604,
    n198
  );


  nand
  g1409
  (
    n1117,
    n418,
    n197,
    n203,
    n445
  );


  or
  g1410
  (
    n1035,
    n468,
    n475,
    n460,
    n353
  );


  xnor
  g1411
  (
    n1557,
    n243,
    n225,
    n533,
    n195
  );


  or
  g1412
  (
    n868,
    n447,
    n291,
    n294,
    n234
  );


  xnor
  g1413
  (
    n1175,
    n350,
    n325,
    n606,
    n454
  );


  and
  g1414
  (
    n1468,
    n461,
    n204,
    n605,
    n374
  );


  xor
  g1415
  (
    n819,
    n488,
    n565,
    n512,
    n476
  );


  xor
  g1416
  (
    n1609,
    n572,
    n263,
    n589,
    n510
  );


  and
  g1417
  (
    n1314,
    n228,
    n501,
    n578,
    n262
  );


  xor
  g1418
  (
    n1416,
    n285,
    n568,
    n269,
    n256
  );


  nor
  g1419
  (
    n724,
    n343,
    n207,
    n405,
    n611
  );


  or
  g1420
  (
    n799,
    n281,
    n346,
    n501,
    n503
  );


  or
  g1421
  (
    n1602,
    n468,
    n302,
    n197,
    n510
  );


  nor
  g1422
  (
    n1299,
    n365,
    n354,
    n247,
    n371
  );


  or
  g1423
  (
    n1424,
    n242,
    n390,
    n208,
    n537
  );


  nand
  g1424
  (
    n1436,
    n603,
    n611,
    n269,
    n597
  );


  nand
  g1425
  (
    n687,
    n489,
    n495,
    n610,
    n329
  );


  nor
  g1426
  (
    n1423,
    n164,
    n318,
    n485,
    n211
  );


  and
  g1427
  (
    n863,
    n344,
    n220,
    n251,
    n189
  );


  xnor
  g1428
  (
    n896,
    n525,
    n352,
    n563,
    n595
  );


  nand
  g1429
  (
    n904,
    n336,
    n533,
    n527,
    n445
  );


  and
  g1430
  (
    n1407,
    n179,
    n588,
    n256,
    n292
  );


  xnor
  g1431
  (
    n1222,
    n201,
    n163,
    n522,
    n463
  );


  and
  g1432
  (
    n1528,
    n206,
    n453,
    n434,
    n191
  );


  nor
  g1433
  (
    n1161,
    n585,
    n580,
    n241,
    n491
  );


  xnor
  g1434
  (
    n779,
    n232,
    n366,
    n591,
    n175
  );


  nor
  g1435
  (
    n1049,
    n589,
    n188,
    n295,
    n259
  );


  and
  g1436
  (
    n1411,
    n509,
    n467,
    n161
  );


  or
  g1437
  (
    n1608,
    n321,
    n601,
    n613,
    n216
  );


  xnor
  g1438
  (
    n709,
    n606,
    n423,
    n458,
    n201
  );


  or
  g1439
  (
    n1464,
    n328,
    n587,
    n438,
    n326
  );


  xor
  g1440
  (
    n1497,
    n229,
    n278,
    n299,
    n591
  );


  xor
  g1441
  (
    n1474,
    n496,
    n185,
    n399,
    n543
  );


  nand
  g1442
  (
    n688,
    n185,
    n366,
    n284,
    n203
  );


  nor
  g1443
  (
    n1627,
    n593,
    n473,
    n230,
    n543
  );


  or
  g1444
  (
    n1248,
    n486,
    n576,
    n305,
    n222
  );


  nand
  g1445
  (
    n1020,
    n305,
    n177,
    n432,
    n263
  );


  and
  g1446
  (
    n1349,
    n312,
    n248,
    n381,
    n197
  );


  and
  g1447
  (
    n1587,
    n181,
    n451,
    n349,
    n409
  );


  or
  g1448
  (
    n693,
    n389,
    n513,
    n502,
    n476
  );


  or
  g1449
  (
    n897,
    n166,
    n605,
    n508,
    n283
  );


  nor
  g1450
  (
    n1209,
    n219,
    n301,
    n169,
    n572
  );


  nor
  g1451
  (
    n992,
    n375,
    n289,
    n228,
    n404
  );


  and
  g1452
  (
    n1053,
    n536,
    n595,
    n287,
    n491
  );


  nand
  g1453
  (
    n1048,
    n219,
    n224,
    n293,
    n596
  );


  nand
  g1454
  (
    n1485,
    n318,
    n292,
    n563,
    n591
  );


  and
  g1455
  (
    n1625,
    n384,
    n549,
    n436,
    n248
  );


  or
  g1456
  (
    n1242,
    n356,
    n447,
    n479,
    n523
  );


  or
  g1457
  (
    n719,
    n519,
    n350,
    n582,
    n179
  );


  and
  g1458
  (
    n1495,
    n231,
    n393,
    n600,
    n481
  );


  nor
  g1459
  (
    n825,
    n207,
    n504,
    n186,
    n193
  );


  nand
  g1460
  (
    n1568,
    n541,
    n238,
    n370,
    n535
  );


  xor
  g1461
  (
    n1534,
    n272,
    n411,
    n358,
    n395
  );


  xnor
  g1462
  (
    n1271,
    n282,
    n412,
    n235,
    n578
  );


  nor
  g1463
  (
    n1183,
    n364,
    n269,
    n451,
    n415
  );


  nor
  g1464
  (
    n1202,
    n466,
    n182,
    n586,
    n551
  );


  nor
  g1465
  (
    n934,
    n391,
    n287,
    n490,
    n607
  );


  xnor
  g1466
  (
    n1166,
    n455,
    n282,
    n346,
    n527
  );


  nand
  g1467
  (
    n1498,
    n291,
    n399,
    n300,
    n524
  );


  xnor
  g1468
  (
    n1195,
    n172,
    n562,
    n508,
    n236
  );


  nor
  g1469
  (
    n1582,
    n322,
    n175,
    n330,
    n377
  );


  or
  g1470
  (
    n1671,
    n213,
    n192,
    n405,
    n461
  );


  nand
  g1471
  (
    n1348,
    n601,
    n212,
    n264,
    n291
  );


  nor
  g1472
  (
    n831,
    n324,
    n297,
    n209,
    n256
  );


  nor
  g1473
  (
    n1252,
    n540,
    n405,
    n179,
    n528
  );


  nor
  g1474
  (
    n1662,
    n325,
    n205,
    n399,
    n613
  );


  or
  g1475
  (
    n1670,
    n476,
    n210,
    n308,
    n362
  );


  nor
  g1476
  (
    n901,
    n209,
    n298,
    n583,
    n389
  );


  nand
  g1477
  (
    n1653,
    n535,
    n505,
    n334,
    n376
  );


  and
  g1478
  (
    n1452,
    n503,
    n273,
    n182,
    n424
  );


  nand
  g1479
  (
    n1397,
    n165,
    n274,
    n192,
    n435
  );


  xor
  g1480
  (
    n771,
    n470,
    n258,
    n532,
    n561
  );


  nand
  g1481
  (
    n1430,
    n302,
    n420,
    n379,
    n191
  );


  xnor
  g1482
  (
    n1269,
    n313,
    n178,
    n324,
    n322
  );


  and
  g1483
  (
    n1034,
    n519,
    n367,
    n586,
    n413
  );


  nand
  g1484
  (
    n673,
    n267,
    n539,
    n174,
    n610
  );


  xor
  g1485
  (
    n1462,
    n561,
    n408,
    n530,
    n194
  );


  or
  g1486
  (
    n1286,
    n592,
    n208,
    n545,
    n544
  );


  nor
  g1487
  (
    n1228,
    n539,
    n534,
    n285,
    n414
  );


  xnor
  g1488
  (
    n1015,
    n346,
    n333,
    n502,
    n602
  );


  xor
  g1489
  (
    n971,
    n410,
    n505,
    n426
  );


  or
  g1490
  (
    n1078,
    n510,
    n514,
    n493,
    n209
  );


  nand
  g1491
  (
    n1363,
    n336,
    n476,
    n306,
    n322
  );


  xnor
  g1492
  (
    n1133,
    n237,
    n396,
    n612,
    n253
  );


  nand
  g1493
  (
    n813,
    n494,
    n261,
    n232,
    n538
  );


  nand
  g1494
  (
    n1232,
    n500,
    n572,
    n409,
    n515
  );


  xnor
  g1495
  (
    n704,
    n342,
    n306,
    n564,
    n499
  );


  xnor
  g1496
  (
    n1376,
    n416,
    n396,
    n404,
    n268
  );


  nand
  g1497
  (
    KeyWire_0_7,
    n609,
    n320,
    n434,
    n410
  );


  xor
  g1498
  (
    n995,
    n362,
    n380,
    n250,
    n511
  );


  nand
  g1499
  (
    n1647,
    n533,
    n261,
    n172,
    n237
  );


  or
  g1500
  (
    n1083,
    n319,
    n484,
    n390,
    n425
  );


  or
  g1501
  (
    n976,
    n386,
    n357,
    n242,
    n198
  );


  or
  g1502
  (
    n765,
    n495,
    n536,
    n407,
    n516
  );


  and
  g1503
  (
    n1479,
    n333,
    n162,
    n224,
    n182
  );


  xor
  g1504
  (
    n937,
    n246,
    n520,
    n498
  );


  xnor
  g1505
  (
    n1659,
    n237,
    n215,
    n569,
    n378
  );


  nor
  g1506
  (
    n1386,
    n543,
    n295,
    n386,
    n328
  );


  nand
  g1507
  (
    n834,
    n216,
    n329,
    n250,
    n230
  );


  nand
  g1508
  (
    n720,
    n305,
    n383,
    n481,
    n205
  );


  or
  g1509
  (
    n1347,
    n511,
    n392,
    n577,
    n240
  );


  or
  g1510
  (
    n1253,
    n433,
    n401,
    n492,
    n413
  );


  nand
  g1511
  (
    n1067,
    n351,
    n303,
    n183,
    n518
  );


  nand
  g1512
  (
    n1182,
    n314,
    n574,
    n338,
    n570
  );


  xnor
  g1513
  (
    n778,
    n499,
    n213,
    n579,
    n594
  );


  or
  g1514
  (
    n924,
    n513,
    n536,
    n598,
    n205
  );


  or
  g1515
  (
    n835,
    n392,
    n218,
    n266,
    n171
  );


  xor
  g1516
  (
    n1296,
    n233,
    n547,
    n187,
    n455
  );


  nor
  g1517
  (
    n1231,
    n330,
    n240,
    n448,
    n314
  );


  nor
  g1518
  (
    n1301,
    n287,
    n247,
    n283,
    n551
  );


  nand
  g1519
  (
    n774,
    n474,
    n385,
    n265,
    n252
  );


  nor
  g1520
  (
    n1179,
    n391,
    n258,
    n504,
    n266
  );


  xor
  g1521
  (
    n703,
    n428,
    n350,
    n365,
    n492
  );


  nor
  g1522
  (
    n1124,
    n488,
    n592,
    n612,
    n317
  );


  nand
  g1523
  (
    n1401,
    n420,
    n266,
    n462,
    n531
  );


  or
  g1524
  (
    n1515,
    n247,
    n235,
    n438,
    n608
  );


  xnor
  g1525
  (
    n919,
    n241,
    n487,
    n520,
    n340
  );


  nand
  g1526
  (
    n842,
    n168,
    n239,
    n178,
    n478
  );


  xnor
  g1527
  (
    n1152,
    n332,
    n497,
    n374,
    n248
  );


  nand
  g1528
  (
    n820,
    n206,
    n417,
    n508,
    n185
  );


  nor
  g1529
  (
    n1243,
    n326,
    n418,
    n384,
    n309
  );


  xor
  g1530
  (
    n697,
    n418,
    n505,
    n543,
    n342
  );


  or
  g1531
  (
    n931,
    n406,
    n463,
    n311,
    n184
  );


  nor
  g1532
  (
    n766,
    n590,
    n271,
    n423,
    n172
  );


  xor
  g1533
  (
    n1186,
    n309,
    n339,
    n232,
    n242
  );


  xor
  g1534
  (
    n905,
    n600,
    n368,
    n394,
    n516
  );


  nand
  g1535
  (
    n1657,
    n516,
    n274,
    n380,
    n392
  );


  nor
  g1536
  (
    n1374,
    n239,
    n562,
    n352,
    n499
  );


  and
  g1537
  (
    n1108,
    n307,
    n294,
    n365,
    n436
  );


  nor
  g1538
  (
    n1420,
    n610,
    n366,
    n312,
    n276
  );


  nor
  g1539
  (
    n912,
    n453,
    n180,
    n325,
    n344
  );


  xnor
  g1540
  (
    n1668,
    n263,
    n489,
    n187,
    n286
  );


  nand
  g1541
  (
    n1634,
    n273,
    n306,
    n198,
    n195
  );


  xnor
  g1542
  (
    n1333,
    n214,
    n570,
    n576,
    n286
  );


  nand
  g1543
  (
    n979,
    n290,
    n294,
    n279,
    n244
  );


  nor
  g1544
  (
    n866,
    n190,
    n408,
    n524,
    n243
  );


  and
  g1545
  (
    n1419,
    n540,
    n404,
    n485,
    n571
  );


  xnor
  g1546
  (
    n915,
    n277,
    n497,
    n554,
    n213
  );


  or
  g1547
  (
    n1350,
    n442,
    n389,
    n398,
    n379
  );


  xnor
  g1548
  (
    n907,
    n388,
    n195,
    n302,
    n599
  );


  nor
  g1549
  (
    n1389,
    n417,
    n460,
    n343,
    n200
  );


  nand
  g1550
  (
    n827,
    n566,
    n541,
    n470,
    n164
  );


  or
  g1551
  (
    n880,
    n275,
    n337,
    n431,
    n548
  );


  and
  g1552
  (
    n1594,
    n255,
    n381,
    n349,
    n177
  );


  xnor
  g1553
  (
    n1037,
    n502,
    n176,
    n374,
    n580
  );


  or
  g1554
  (
    n1570,
    n256,
    n473,
    n415,
    n270
  );


  xnor
  g1555
  (
    n818,
    n218,
    n574,
    n580,
    n184
  );


  xnor
  g1556
  (
    n1003,
    n240,
    n340,
    n577,
    n438
  );


  or
  g1557
  (
    n1206,
    n274,
    n318,
    n457,
    n211
  );


  and
  g1558
  (
    n1650,
    n213,
    n443,
    n596,
    n254
  );


  nor
  g1559
  (
    n1572,
    n173,
    n492,
    n346,
    n601
  );


  xor
  g1560
  (
    n957,
    n593,
    n542,
    n370,
    n587
  );


  nor
  g1561
  (
    n1443,
    n451,
    n419,
    n271,
    n188
  );


  xor
  g1562
  (
    n1544,
    n359,
    n392,
    n550,
    n215
  );


  or
  g1563
  (
    n1429,
    n173,
    n429,
    n191,
    n454
  );


  and
  g1564
  (
    n1174,
    n576,
    n334,
    n556,
    n523
  );


  and
  g1565
  (
    n1579,
    n475,
    n461,
    n416,
    n402
  );


  nor
  g1566
  (
    n1524,
    n167,
    n594,
    n545,
    n429
  );


  nor
  g1567
  (
    n824,
    n385,
    n220,
    n289,
    n501
  );


  nor
  g1568
  (
    n1167,
    n496,
    n291,
    n446,
    n246
  );


  or
  g1569
  (
    n1341,
    n245,
    n435,
    n513,
    n497
  );


  or
  g1570
  (
    n1054,
    n449,
    n196,
    n323,
    n489
  );


  nor
  g1571
  (
    n1187,
    n254,
    n260,
    n162,
    n217
  );


  and
  g1572
  (
    n951,
    n429,
    n363,
    n575,
    n475
  );


  and
  g1573
  (
    n1274,
    n217,
    n296,
    n177,
    n599
  );


  or
  g1574
  (
    n853,
    n604,
    n335,
    n223,
    n417
  );


  and
  g1575
  (
    n1268,
    n267,
    n432,
    n393,
    n468
  );


  xor
  g1576
  (
    n993,
    n537,
    n539,
    n288,
    n310
  );


  or
  g1577
  (
    n1089,
    n206,
    n288,
    n430,
    n355
  );


  nor
  g1578
  (
    n1153,
    n190,
    n411,
    n449,
    n210
  );


  nand
  g1579
  (
    KeyWire_0_19,
    n375,
    n365,
    n479,
    n465
  );


  xnor
  g1580
  (
    n1506,
    n290,
    n227,
    n413,
    n570
  );


  nor
  g1581
  (
    n1013,
    n400,
    n605,
    n473,
    n576
  );


  nand
  g1582
  (
    n1065,
    n254,
    n280,
    n356,
    n421
  );


  and
  g1583
  (
    n808,
    n372,
    n331,
    n369,
    n183
  );


  xnor
  g1584
  (
    n1369,
    n257,
    n552,
    n607,
    n485
  );


  xor
  g1585
  (
    n1371,
    n394,
    n274,
    n168,
    n400
  );


  and
  g1586
  (
    n1543,
    n598,
    n233,
    n332,
    n339
  );


  and
  g1587
  (
    n1266,
    n562,
    n262,
    n483,
    n553
  );


  xnor
  g1588
  (
    n1207,
    n553,
    n411,
    n388,
    n359
  );


  or
  g1589
  (
    n1351,
    n227,
    n282,
    n614,
    n522
  );


  and
  g1590
  (
    n1277,
    n215,
    n495,
    n433,
    n473
  );


  or
  g1591
  (
    n1185,
    n465,
    n400,
    n555,
    n515
  );


  xnor
  g1592
  (
    n1148,
    n285,
    n167,
    n571,
    n299
  );


  xor
  g1593
  (
    n744,
    n225,
    n353,
    n187,
    n328
  );


  xnor
  g1594
  (
    n1358,
    n564,
    n479,
    n357,
    n472
  );


  nor
  g1595
  (
    n1001,
    n354,
    n422,
    n235,
    n564
  );


  nor
  g1596
  (
    n1140,
    n582,
    n480,
    n452,
    n560
  );


  and
  g1597
  (
    n816,
    n394,
    n506,
    n388,
    n362
  );


  xor
  g1598
  (
    n1577,
    n510,
    n223,
    n465,
    n556
  );


  or
  g1599
  (
    n1359,
    n277,
    n517,
    n166,
    n379
  );


  xnor
  g1600
  (
    n1599,
    n257,
    n569,
    n425,
    n615
  );


  nand
  g1601
  (
    n1289,
    n345,
    n601,
    n199,
    n397
  );


  and
  g1602
  (
    n1628,
    n255,
    n508,
    n225,
    n474
  );


  and
  g1603
  (
    n1629,
    n336,
    n460,
    n402,
    n223
  );


  and
  g1604
  (
    n1038,
    n200,
    n443,
    n565,
    n396
  );


  or
  g1605
  (
    n1573,
    n373,
    n170,
    n496,
    n189
  );


  and
  g1606
  (
    n1091,
    n170,
    n409,
    n351,
    n484
  );


  xor
  g1607
  (
    n1361,
    n176,
    n382,
    n314,
    n557
  );


  and
  g1608
  (
    n1143,
    n212,
    n337,
    n332,
    n599
  );


  or
  g1609
  (
    n1122,
    n558,
    n581,
    n526,
    n344
  );


  xor
  g1610
  (
    n1070,
    n312,
    n358,
    n522,
    n477
  );


  nor
  g1611
  (
    n1656,
    n584,
    n380,
    n408,
    n321
  );


  nor
  g1612
  (
    n854,
    n398,
    n451,
    n359,
    n525
  );


  nor
  g1613
  (
    n1283,
    n431,
    n467,
    n192,
    n356
  );


  or
  g1614
  (
    n1530,
    n189,
    n393,
    n560,
    n453
  );


  nor
  g1615
  (
    n1313,
    n194,
    n330,
    n509,
    n539
  );


  and
  g1616
  (
    n983,
    n446,
    n398,
    n303,
    n310
  );


  nand
  g1617
  (
    n1616,
    n477,
    n609,
    n437,
    n546
  );


  nor
  g1618
  (
    n1615,
    n507,
    n194,
    n315,
    n377
  );


  nand
  g1619
  (
    n1435,
    n200,
    n339,
    n382,
    n456
  );


  and
  g1620
  (
    n1176,
    n550,
    n323,
    n514,
    n236
  );


  xor
  g1621
  (
    n970,
    n305,
    n337,
    n493,
    n395
  );


  xnor
  g1622
  (
    KeyWire_0_29,
    n245,
    n424,
    n360,
    n441
  );


  xnor
  g1623
  (
    n1265,
    n186,
    n352,
    n259,
    n345
  );


  xor
  g1624
  (
    n916,
    n441,
    n211,
    n495,
    n333
  );


  xnor
  g1625
  (
    n1136,
    n327,
    n280,
    n404,
    n265
  );


  xor
  g1626
  (
    n1402,
    n434,
    n349,
    n462,
    n279
  );


  nor
  g1627
  (
    n1457,
    n406,
    n204,
    n162,
    n388
  );


  or
  g1628
  (
    n1276,
    n364,
    n567,
    n258,
    n292
  );


  or
  g1629
  (
    n1223,
    n190,
    n463,
    n353,
    n286
  );


  xor
  g1630
  (
    n716,
    n528,
    n512,
    n376,
    n579
  );


  xnor
  g1631
  (
    n1284,
    n181,
    n272,
    n557,
    n251
  );


  xor
  g1632
  (
    n1113,
    n278,
    n587,
    n316,
    n566
  );


  or
  g1633
  (
    n920,
    n211,
    n328,
    n308,
    n519
  );


  nor
  g1634
  (
    n908,
    n332,
    n255,
    n570,
    n427
  );


  or
  g1635
  (
    n1400,
    n193,
    n271,
    n464,
    n573
  );


  and
  g1636
  (
    n1184,
    n439,
    n304,
    n531,
    n281
  );


  and
  g1637
  (
    n876,
    n448,
    n321,
    n525,
    n406
  );


  xnor
  g1638
  (
    n1441,
    n441,
    n597,
    n561,
    n448
  );


  or
  g1639
  (
    n943,
    n403,
    n586,
    n371,
    n244
  );


  nand
  g1640
  (
    n712,
    n503,
    n448,
    n544,
    n181
  );


  nor
  g1641
  (
    n1675,
    n673,
    n678,
    n676,
    n674
  );


  or
  g1642
  (
    n1674,
    n677,
    n680,
    n679,
    n675
  );


  nor
  g1643
  (
    n1676,
    n682,
    n1675,
    n683,
    n681
  );


  xor
  g1644
  (
    n1680,
    n616,
    n617
  );


  nor
  g1645
  (
    n1678,
    n615,
    n617,
    n1676
  );


  nor
  g1646
  (
    n1679,
    n1676,
    n616
  );


  and
  g1647
  (
    n1677,
    n616,
    n615,
    n618
  );


  xor
  g1648
  (
    n1686,
    n1677,
    n1679,
    n1680,
    n707
  );


  or
  g1649
  (
    n1681,
    n695,
    n704,
    n689,
    n685
  );


  and
  g1650
  (
    n1688,
    n703,
    n1679,
    n710,
    n684
  );


  nor
  g1651
  (
    n1683,
    n700,
    n705,
    n702,
    n693
  );


  or
  g1652
  (
    n1690,
    n1679,
    n1679,
    n699,
    n708
  );


  nor
  g1653
  (
    n1685,
    n692,
    n688,
    n706,
    n713
  );


  xor
  g1654
  (
    n1682,
    n709,
    n694,
    n1678,
    n712
  );


  xor
  g1655
  (
    n1687,
    n687,
    n696,
    n1680,
    n701
  );


  xnor
  g1656
  (
    n1684,
    n691,
    n711,
    n697,
    n1680
  );


  xnor
  g1657
  (
    n1689,
    n686,
    n690,
    n1680,
    n698
  );


  buf
  g1658
  (
    n1701,
    n1686
  );


  not
  g1659
  (
    n1694,
    n723
  );


  not
  g1660
  (
    n1692,
    n1686
  );


  buf
  g1661
  (
    n1693,
    n729
  );


  not
  g1662
  (
    n1703,
    n1685
  );


  buf
  g1663
  (
    n1705,
    n720
  );


  buf
  g1664
  (
    n1706,
    n722
  );


  not
  g1665
  (
    n1704,
    n730
  );


  not
  g1666
  (
    n1696,
    n1684
  );


  xor
  g1667
  (
    n1695,
    n1686,
    n1685,
    n1683,
    n726
  );


  or
  g1668
  (
    n1698,
    n1685,
    n719,
    n1687,
    n716
  );


  or
  g1669
  (
    n1700,
    n717,
    n1684,
    n1687,
    n1681
  );


  xor
  g1670
  (
    n1697,
    n1682,
    n718,
    n1686,
    n1684
  );


  and
  g1671
  (
    n1699,
    n725,
    n733,
    n727,
    n732
  );


  xor
  g1672
  (
    n1702,
    n1684,
    n715,
    n731,
    n728
  );


  xnor
  g1673
  (
    n1691,
    n714,
    n721,
    n724,
    n1685
  );


  not
  g1674
  (
    n1719,
    n1706
  );


  buf
  g1675
  (
    n1710,
    n1700
  );


  buf
  g1676
  (
    n1720,
    n1692
  );


  not
  g1677
  (
    n1718,
    n1697
  );


  not
  g1678
  (
    n1709,
    n1701
  );


  buf
  g1679
  (
    n1722,
    n1695
  );


  not
  g1680
  (
    n1707,
    n1691
  );


  buf
  g1681
  (
    n1712,
    n1693
  );


  buf
  g1682
  (
    n1717,
    n1704
  );


  not
  g1683
  (
    n1716,
    n1694
  );


  not
  g1684
  (
    n1711,
    n1698
  );


  buf
  g1685
  (
    n1714,
    n1705
  );


  buf
  g1686
  (
    n1721,
    n1703
  );


  not
  g1687
  (
    n1715,
    n1699
  );


  not
  g1688
  (
    n1713,
    n1702
  );


  buf
  g1689
  (
    n1708,
    n1696
  );


  not
  g1690
  (
    n1723,
    n1709
  );


  nor
  g1691
  (
    n1724,
    n1707,
    n1708,
    n1710
  );


  and
  g1692
  (
    n1726,
    n1711,
    n1723,
    n1724,
    n1714
  );


  or
  g1693
  (
    n1725,
    n1716,
    n1712,
    n1713,
    n1715
  );


  not
  g1694
  (
    n1727,
    n1725
  );


  xor
  g1695
  (
    n1729,
    n1727,
    n1720
  );


  buf
  g1696
  (
    KeyWire_0_11,
    n1727
  );


  nor
  g1697
  (
    n1728,
    n1727,
    n1717
  );


  and
  g1698
  (
    n1731,
    n1719,
    n1718
  );


  not
  g1699
  (
    n1733,
    n1728
  );


  buf
  g1700
  (
    n1743,
    n1731
  );


  buf
  g1701
  (
    n1746,
    n1729
  );


  buf
  g1702
  (
    n1739,
    n1731
  );


  buf
  g1703
  (
    n1734,
    n1731
  );


  buf
  g1704
  (
    n1742,
    n1730
  );


  buf
  g1705
  (
    n1738,
    n1728
  );


  not
  g1706
  (
    n1737,
    n1729
  );


  buf
  g1707
  (
    n1741,
    n1728
  );


  buf
  g1708
  (
    n1744,
    n1730
  );


  buf
  g1709
  (
    n1736,
    n1729
  );


  buf
  g1710
  (
    n1740,
    n1729
  );


  not
  g1711
  (
    n1732,
    n1730
  );


  buf
  g1712
  (
    n1745,
    n1730
  );


  not
  g1713
  (
    n1747,
    n1728
  );


  buf
  g1714
  (
    n1735,
    n1731
  );


  buf
  g1715
  (
    n1748,
    n1732
  );


  not
  g1716
  (
    n1750,
    n1732
  );


  not
  g1717
  (
    n1749,
    n1732
  );


  not
  g1718
  (
    n1751,
    n1732
  );


  nor
  g1719
  (
    n1764,
    n1744,
    n1736,
    n1734,
    n1749
  );


  nor
  g1720
  (
    n1761,
    n1749,
    n1750,
    n1751
  );


  and
  g1721
  (
    n1760,
    n1738,
    n1736,
    n1751,
    n1735
  );


  or
  g1722
  (
    n1757,
    n1751,
    n1741,
    n1748,
    n1740
  );


  and
  g1723
  (
    n1752,
    n1741,
    n1735,
    n1736,
    n1748
  );


  or
  g1724
  (
    n1766,
    n1743,
    n1743,
    n1744,
    n1742
  );


  nor
  g1725
  (
    n1753,
    n1735,
    n1748,
    n1734,
    n1738
  );


  xor
  g1726
  (
    n1758,
    n1739,
    n1744,
    n1734,
    n1733
  );


  nand
  g1727
  (
    n1755,
    n1742,
    n1733,
    n1740,
    n1743
  );


  or
  g1728
  (
    n1763,
    n1737,
    n734,
    n1742,
    n1739
  );


  nor
  g1729
  (
    n1756,
    n1738,
    n1737,
    n1740,
    n1741
  );


  nand
  g1730
  (
    n1762,
    n1733,
    n1749,
    n1737,
    n1741
  );


  or
  g1731
  (
    n1754,
    n1748,
    n1740,
    n1739,
    n1751
  );


  or
  g1732
  (
    n1759,
    n1737,
    n1749,
    n1736,
    n1743
  );


  xor
  g1733
  (
    n1765,
    n1734,
    n1742,
    n1738,
    n1739
  );


  nor
  g1734
  (
    n1767,
    n1735,
    n1733,
    n1750
  );


  nor
  g1735
  (
    n1795,
    n1758,
    n1756,
    n618,
    n636
  );


  or
  g1736
  (
    n1827,
    n650,
    n650,
    n1765,
    n644
  );


  nand
  g1737
  (
    n1803,
    n637,
    n652,
    n631,
    n662
  );


  xor
  g1738
  (
    n1773,
    n618,
    n1762,
    n658,
    n630
  );


  nand
  g1739
  (
    n1810,
    n1760,
    n1753,
    n621,
    n618
  );


  xor
  g1740
  (
    n1813,
    n648,
    n633,
    n1761,
    n653
  );


  nor
  g1741
  (
    n1788,
    n627,
    n627,
    n623,
    n620
  );


  xor
  g1742
  (
    n1789,
    n660,
    n1757,
    n635,
    n656
  );


  and
  g1743
  (
    n1826,
    n1757,
    n633,
    n1758,
    n624
  );


  xnor
  g1744
  (
    n1818,
    n642,
    n646,
    n1753,
    n619
  );


  nor
  g1745
  (
    n1786,
    n1752,
    n628,
    n653,
    n621
  );


  xor
  g1746
  (
    n1784,
    n659,
    n645,
    n636,
    n1755
  );


  and
  g1747
  (
    n1801,
    n1755,
    n620,
    n1764,
    n663
  );


  or
  g1748
  (
    n1800,
    n631,
    n665,
    n659,
    n646
  );


  nor
  g1749
  (
    n1825,
    n648,
    n631,
    n627,
    n655
  );


  and
  g1750
  (
    n1807,
    n652,
    n1759,
    n643,
    n1755
  );


  and
  g1751
  (
    n1828,
    n647,
    n658,
    n1760,
    n619
  );


  nor
  g1752
  (
    n1792,
    n662,
    n651,
    n1755,
    n642
  );


  xnor
  g1753
  (
    n1783,
    n650,
    n659,
    n640,
    n645
  );


  xnor
  g1754
  (
    n1808,
    n641,
    n646,
    n630,
    n625
  );


  nor
  g1755
  (
    n1796,
    n634,
    n1766,
    n633,
    n624
  );


  or
  g1756
  (
    n1823,
    n653,
    n629,
    n1764,
    n643
  );


  xor
  g1757
  (
    n1830,
    n663,
    n656,
    n640
  );


  or
  g1758
  (
    n1780,
    n638,
    n650,
    n644,
    n630
  );


  xor
  g1759
  (
    n1812,
    n634,
    n1762,
    n642,
    n657
  );


  or
  g1760
  (
    n1809,
    n637,
    n664,
    n644
  );


  nor
  g1761
  (
    n1779,
    n1765,
    n640,
    n1767,
    n632
  );


  or
  g1762
  (
    n1774,
    n639,
    n626,
    n1760,
    n1752
  );


  nand
  g1763
  (
    n1802,
    n626,
    n619,
    n1760,
    n1756
  );


  or
  g1764
  (
    n1798,
    n627,
    n634,
    n1761,
    n1762
  );


  nand
  g1765
  (
    n1829,
    n620,
    n1765,
    n658,
    n1754
  );


  xor
  g1766
  (
    n1794,
    n655,
    n642,
    n638,
    n644
  );


  nand
  g1767
  (
    n1787,
    n654,
    n1752,
    n661,
    n1764
  );


  xor
  g1768
  (
    n1814,
    n630,
    n640,
    n1764,
    n648
  );


  xnor
  g1769
  (
    n1811,
    n622,
    n1752,
    n639
  );


  or
  g1770
  (
    n1777,
    n1758,
    n625,
    n659,
    n636
  );


  nor
  g1771
  (
    n1804,
    n645,
    n635,
    n1767,
    n655
  );


  xnor
  g1772
  (
    n1778,
    n631,
    n1761,
    n664,
    n633
  );


  or
  g1773
  (
    n1771,
    n1754,
    n632,
    n663,
    n664
  );


  nor
  g1774
  (
    n1824,
    n632,
    n634,
    n662,
    n1763
  );


  nand
  g1775
  (
    n1797,
    n623,
    n657,
    n649
  );


  nand
  g1776
  (
    n1785,
    n657,
    n1759,
    n635,
    n625
  );


  or
  g1777
  (
    n1769,
    n1761,
    n629,
    n660,
    n647
  );


  nand
  g1778
  (
    n1791,
    n619,
    n636,
    n628,
    n1765
  );


  nand
  g1779
  (
    n1817,
    n1754,
    n638,
    n654,
    n661
  );


  nand
  g1780
  (
    n1805,
    n641,
    n641,
    n629,
    n628
  );


  xor
  g1781
  (
    n1770,
    n665,
    n1753,
    n660,
    n654
  );


  nand
  g1782
  (
    n1799,
    n625,
    n663,
    n1763,
    n629
  );


  nor
  g1783
  (
    n1820,
    n648,
    n637,
    n628,
    n1767
  );


  xor
  g1784
  (
    KeyWire_0_21,
    n657,
    n1767,
    n637,
    n651
  );


  or
  g1785
  (
    n1790,
    n632,
    n647,
    n635,
    n643
  );


  nand
  g1786
  (
    n1768,
    n647,
    n1759,
    n621,
    n1758
  );


  xnor
  g1787
  (
    n1772,
    n622,
    n653,
    n1757,
    n1766
  );


  and
  g1788
  (
    n1806,
    n622,
    n622,
    n1763,
    n658
  );


  nand
  g1789
  (
    n1822,
    n1762,
    n639,
    n643,
    n660
  );


  or
  g1790
  (
    n1815,
    n1766,
    n651,
    n641,
    n1756
  );


  xor
  g1791
  (
    n1821,
    n645,
    n661,
    n1753,
    n1756
  );


  xnor
  g1792
  (
    n1831,
    n1754,
    n661,
    n626,
    n646
  );


  nand
  g1793
  (
    n1781,
    n638,
    n654,
    n665,
    n623
  );


  nor
  g1794
  (
    n1782,
    n624,
    n649,
    n1759,
    n662
  );


  nand
  g1795
  (
    n1816,
    n656,
    n1763,
    n666,
    n620
  );


  or
  g1796
  (
    n1793,
    n652,
    n652,
    n624,
    n623
  );


  nand
  g1797
  (
    KeyWire_0_16,
    n649,
    n651,
    n1766,
    n1757
  );


  xor
  g1798
  (
    n1819,
    n665,
    n621,
    n655,
    n626
  );


  xnor
  g1799
  (
    n2071,
    n1817,
    n1345,
    n1780,
    n1407
  );


  and
  g1800
  (
    n1903,
    n882,
    n1018,
    n954,
    n1368
  );


  and
  g1801
  (
    n2027,
    n1799,
    n1802,
    n1825,
    n1809
  );


  and
  g1802
  (
    n1962,
    n1031,
    n1011,
    n1439,
    n1777
  );


  or
  g1803
  (
    n1858,
    n1773,
    n1114,
    n1161,
    n1068
  );


  xor
  g1804
  (
    n2031,
    n1473,
    n756,
    n1824,
    n1338
  );


  xor
  g1805
  (
    n1983,
    n1027,
    n1392,
    n1453,
    n777
  );


  nor
  g1806
  (
    n1868,
    n1003,
    n881,
    n1222,
    n1361
  );


  xnor
  g1807
  (
    n1979,
    n1804,
    n1053,
    n1461,
    n1022
  );


  xnor
  g1808
  (
    n1939,
    n1041,
    n1800,
    n1768,
    n752
  );


  nand
  g1809
  (
    n2050,
    n1810,
    n1502,
    n1127,
    n774
  );


  nand
  g1810
  (
    n1975,
    n1796,
    n984,
    n1108,
    n1168
  );


  xnor
  g1811
  (
    n2022,
    n873,
    n1772,
    n741,
    n840
  );


  xor
  g1812
  (
    n2019,
    n1016,
    n1248,
    n1424,
    n1088
  );


  nor
  g1813
  (
    n2012,
    n876,
    n1177,
    n1794,
    n1025
  );


  and
  g1814
  (
    n1866,
    n850,
    n1188,
    n745,
    n1769
  );


  or
  g1815
  (
    n2074,
    n771,
    n1382,
    n1814,
    n1045
  );


  xnor
  g1816
  (
    n1885,
    n833,
    n1380,
    n1265,
    n1237
  );


  and
  g1817
  (
    n1905,
    n1054,
    n1819,
    n1286,
    n883
  );


  xor
  g1818
  (
    n1911,
    n1823,
    n1397,
    n831,
    n1807
  );


  nor
  g1819
  (
    n1856,
    n1210,
    n1431,
    n1793,
    n1420
  );


  or
  g1820
  (
    n2032,
    n880,
    n1788,
    n953,
    n1831
  );


  or
  g1821
  (
    n2045,
    n1303,
    n1773,
    n1274,
    n1249
  );


  nor
  g1822
  (
    n1898,
    n1772,
    n901,
    n817,
    n804
  );


  nor
  g1823
  (
    n1849,
    n879,
    n1201,
    n1781,
    n1282
  );


  xor
  g1824
  (
    n2065,
    n1242,
    n1779,
    n1351,
    n1205
  );


  nand
  g1825
  (
    n2056,
    n1775,
    n948,
    n1228,
    n1771
  );


  and
  g1826
  (
    n2081,
    n1153,
    n938,
    n1293,
    n1098
  );


  or
  g1827
  (
    n1922,
    n1489,
    n810,
    n1203,
    n1435
  );


  and
  g1828
  (
    n1994,
    n1781,
    n928,
    n985,
    n1220
  );


  and
  g1829
  (
    n1854,
    n1813,
    n1446,
    n1809,
    n764
  );


  xnor
  g1830
  (
    n2020,
    n816,
    n761,
    n803,
    n1825
  );


  nor
  g1831
  (
    n1916,
    n784,
    n1789,
    n1415,
    n1147
  );


  nor
  g1832
  (
    n2038,
    n1307,
    n1805,
    n933,
    n1339
  );


  and
  g1833
  (
    n2064,
    n1096,
    n1279,
    n1227,
    n1250
  );


  and
  g1834
  (
    n1935,
    n1367,
    n1821,
    n1378,
    n1308
  );


  nor
  g1835
  (
    n1840,
    n1158,
    n751,
    n1384,
    n1779
  );


  nor
  g1836
  (
    n1890,
    n930,
    n1786,
    n1106,
    n1312
  );


  xnor
  g1837
  (
    n1997,
    n986,
    n1783,
    n955,
    n1829
  );


  xor
  g1838
  (
    n1883,
    n811,
    n1072,
    n1786,
    n1369
  );


  and
  g1839
  (
    n2070,
    n1807,
    n1786,
    n1046,
    n1352
  );


  nand
  g1840
  (
    n1963,
    n1207,
    n1005,
    n1191,
    n1070
  );


  nor
  g1841
  (
    n1904,
    n1778,
    n1820,
    n1814,
    n1826
  );


  nor
  g1842
  (
    n1884,
    n1329,
    n847,
    n782,
    n1261
  );


  nor
  g1843
  (
    n1954,
    n1770,
    n1049,
    n1343,
    n1787
  );


  nand
  g1844
  (
    n2021,
    n1831,
    n864,
    n799,
    n1405
  );


  xnor
  g1845
  (
    n1876,
    n1822,
    n1497,
    n1251,
    n1799
  );


  or
  g1846
  (
    n1928,
    n1831,
    n1498,
    n894,
    n746
  );


  xnor
  g1847
  (
    KeyWire_0_23,
    n1451,
    n1830,
    n1300,
    n1110
  );


  xnor
  g1848
  (
    n1842,
    n1810,
    n1146,
    n1134,
    n1014
  );


  nand
  g1849
  (
    n1908,
    n1818,
    n1442,
    n1238,
    n1193
  );


  and
  g1850
  (
    n2036,
    n1827,
    n1776,
    n1822,
    n1463
  );


  nand
  g1851
  (
    n2014,
    n1481,
    n980,
    n1798,
    n1808
  );


  xor
  g1852
  (
    n2062,
    n1795,
    n1808,
    n1777,
    n983
  );


  xor
  g1853
  (
    n2055,
    n819,
    n1162,
    n1793,
    n1104
  );


  nand
  g1854
  (
    n2048,
    n1071,
    n1801,
    n796,
    n1260
  );


  xor
  g1855
  (
    n1948,
    n895,
    n838,
    n1002,
    n1464
  );


  and
  g1856
  (
    n1834,
    n1172,
    n1362,
    n1807,
    n1321
  );


  xor
  g1857
  (
    n1932,
    n1311,
    n769,
    n970,
    n1289
  );


  or
  g1858
  (
    n2068,
    n1332,
    n1806,
    n1831,
    n1102
  );


  xnor
  g1859
  (
    n1865,
    n1257,
    n1800,
    n1215,
    n1288
  );


  nand
  g1860
  (
    n2011,
    n1319,
    n1778,
    n1008,
    n1232
  );


  or
  g1861
  (
    n1844,
    n1077,
    n910,
    n1782,
    n1820
  );


  and
  g1862
  (
    n1936,
    n1302,
    n1056,
    n1808,
    n878
  );


  nand
  g1863
  (
    n1910,
    n1240,
    n929,
    n1823,
    n808
  );


  xor
  g1864
  (
    n1847,
    n935,
    n1350,
    n1294,
    n1107
  );


  xor
  g1865
  (
    n1837,
    n1768,
    n1787,
    n832,
    n1204
  );


  and
  g1866
  (
    n1906,
    n1364,
    n1824,
    n1813,
    n792
  );


  xor
  g1867
  (
    n1949,
    n1328,
    n1811,
    n863,
    n896
  );


  nand
  g1868
  (
    n2047,
    n987,
    n1792,
    n1769,
    n849
  );


  and
  g1869
  (
    n1996,
    n1830,
    n1775,
    n740,
    n923
  );


  or
  g1870
  (
    n1832,
    n1013,
    n755,
    n1090,
    n1794
  );


  or
  g1871
  (
    n1907,
    n1044,
    n1402,
    n1322,
    n853
  );


  or
  g1872
  (
    n1917,
    n1811,
    n1797,
    n1428,
    n1801
  );


  xor
  g1873
  (
    n1895,
    n1062,
    n1069,
    n1791,
    n1433
  );


  nor
  g1874
  (
    n2061,
    n1822,
    n1495,
    n995,
    n1330
  );


  nand
  g1875
  (
    n2026,
    n1373,
    n1033,
    n1359,
    n1383
  );


  nor
  g1876
  (
    n2035,
    n1216,
    n1169,
    n1035,
    n1050
  );


  or
  g1877
  (
    n1836,
    n944,
    n1052,
    n1131,
    n1803
  );


  nand
  g1878
  (
    n2003,
    n1376,
    n1824,
    n1770,
    n1231
  );


  nand
  g1879
  (
    n1920,
    n1275,
    n800,
    n1159,
    n1082
  );


  xor
  g1880
  (
    n2028,
    n1140,
    n1366,
    n904,
    n1317
  );


  nor
  g1881
  (
    n1952,
    n1771,
    n1125,
    n1189,
    n1487
  );


  xor
  g1882
  (
    n2072,
    n1434,
    n1141,
    n1775,
    n1183
  );


  nand
  g1883
  (
    n2075,
    n775,
    n1167,
    n776,
    n1278
  );


  or
  g1884
  (
    n2073,
    n1802,
    n1026,
    n1354,
    n1135
  );


  and
  g1885
  (
    n2041,
    n1255,
    n1830,
    n1034,
    n770
  );


  or
  g1886
  (
    n1914,
    n932,
    n886,
    n835,
    n1798
  );


  and
  g1887
  (
    n2057,
    n1066,
    n860,
    n1055,
    n1449
  );


  and
  g1888
  (
    n1965,
    n1030,
    n1791,
    n1078,
    n1492
  );


  xnor
  g1889
  (
    n1915,
    n1486,
    n1186,
    n959,
    n1195
  );


  xnor
  g1890
  (
    n1871,
    n1223,
    n974,
    n972,
    n1268
  );


  nor
  g1891
  (
    n1899,
    n1809,
    n906,
    n1822,
    n1818
  );


  and
  g1892
  (
    n2025,
    n1166,
    n1400,
    n1780,
    n1097
  );


  or
  g1893
  (
    n1846,
    n1233,
    n1160,
    n783,
    n936
  );


  xnor
  g1894
  (
    n1839,
    n1173,
    n1395,
    n1824,
    n1787
  );


  xor
  g1895
  (
    n2015,
    n1040,
    n1493,
    n1187,
    n1297
  );


  nand
  g1896
  (
    n1998,
    n1085,
    n780,
    n1815,
    n1181
  );


  nand
  g1897
  (
    n1891,
    n812,
    n834,
    n1830,
    n1816
  );


  nor
  g1898
  (
    n1878,
    n1815,
    n797,
    n1170,
    n779
  );


  xor
  g1899
  (
    n1950,
    n1142,
    n1458,
    n1794,
    n975
  );


  or
  g1900
  (
    n2060,
    n1798,
    n1023,
    n1283,
    n1423
  );


  and
  g1901
  (
    n2034,
    n1047,
    n1466,
    n1820,
    n1149
  );


  xnor
  g1902
  (
    n1984,
    n1342,
    n1773,
    n1826,
    n947
  );


  nor
  g1903
  (
    n1896,
    n1176,
    n1827,
    n1007,
    n762
  );


  nand
  g1904
  (
    n2066,
    n1491,
    n1772,
    n848,
    n945
  );


  and
  g1905
  (
    n1859,
    n1800,
    n1252,
    n1246,
    n1010
  );


  or
  g1906
  (
    n2086,
    n787,
    n914,
    n1059,
    n960
  );


  nor
  g1907
  (
    n2040,
    n824,
    n1259,
    n1143,
    n924
  );


  nor
  g1908
  (
    n1925,
    n1801,
    n1484,
    n1292,
    n912
  );


  and
  g1909
  (
    n1977,
    n1112,
    n1469,
    n814,
    n1353
  );


  and
  g1910
  (
    n1900,
    n1266,
    n1409,
    n1803,
    n1129
  );


  or
  g1911
  (
    n1843,
    n1365,
    n1000,
    n1388,
    n1774
  );


  or
  g1912
  (
    n2018,
    n854,
    n1426,
    n1393,
    n1394
  );


  or
  g1913
  (
    n1959,
    n1412,
    n1811,
    n1084,
    n1828
  );


  nand
  g1914
  (
    n1845,
    n1280,
    n994,
    n1163,
    n1200
  );


  and
  g1915
  (
    n1886,
    n858,
    n1229,
    n1202,
    n1820
  );


  nand
  g1916
  (
    n1992,
    n1417,
    n1784,
    n1782,
    n1785
  );


  or
  g1917
  (
    n1995,
    n963,
    n801,
    n1042,
    n788
  );


  nand
  g1918
  (
    n1877,
    n1809,
    n1019,
    n1403,
    n1323
  );


  and
  g1919
  (
    n1833,
    n827,
    n1788,
    n1036,
    n1826
  );


  nor
  g1920
  (
    n1951,
    n1379,
    n1450,
    n1081,
    n1805
  );


  xor
  g1921
  (
    n1852,
    n1296,
    n821,
    n1819,
    n1776
  );


  xnor
  g1922
  (
    n2085,
    n1425,
    n1239,
    n1083,
    n1285
  );


  xnor
  g1923
  (
    n2084,
    n781,
    n1390,
    n1151,
    n942
  );


  nor
  g1924
  (
    n2009,
    n1812,
    n822,
    n1769,
    n1821
  );


  and
  g1925
  (
    n2013,
    n917,
    n1370,
    n964,
    n1037
  );


  nand
  g1926
  (
    n1985,
    n744,
    n891,
    n1823,
    n1375
  );


  xnor
  g1927
  (
    n1882,
    n1374,
    n1793,
    n1770,
    n861
  );


  nor
  g1928
  (
    n1881,
    n991,
    n865,
    n1782,
    n1039
  );


  xnor
  g1929
  (
    n1841,
    n967,
    n908,
    n1821,
    n1829
  );


  nor
  g1930
  (
    n1937,
    n866,
    n1101,
    n1067,
    n1117
  );


  nor
  g1931
  (
    n2079,
    n1253,
    n739,
    n749,
    n1414
  );


  and
  g1932
  (
    n1875,
    n867,
    n851,
    n1299,
    n1281
  );


  xor
  g1933
  (
    n1938,
    n1148,
    n1448,
    n1796,
    n1224
  );


  xnor
  g1934
  (
    n1919,
    n951,
    n899,
    n1803,
    n1113
  );


  nor
  g1935
  (
    n2069,
    n1263,
    n1795,
    n1816,
    n1087
  );


  and
  g1936
  (
    n1986,
    n1783,
    n1441,
    n852,
    n1236
  );


  or
  g1937
  (
    n1924,
    n748,
    n1474,
    n997,
    n1406
  );


  nand
  g1938
  (
    n2052,
    n1411,
    n1199,
    n1196,
    n1795
  );


  nor
  g1939
  (
    n2010,
    n1337,
    n1298,
    n1336,
    n1213
  );


  nor
  g1940
  (
    n1923,
    n790,
    n1119,
    n1778,
    n795
  );


  and
  g1941
  (
    n1940,
    n1109,
    n1419,
    n1138,
    n845
  );


  xor
  g1942
  (
    n2000,
    n1333,
    n1389,
    n1444,
    n856
  );


  xor
  g1943
  (
    n1870,
    n892,
    n992,
    n977,
    n1156
  );


  xnor
  g1944
  (
    n1989,
    n1128,
    n1819,
    n1465,
    n1774
  );


  nor
  g1945
  (
    n1973,
    n1796,
    n1818,
    n1398,
    n1074
  );


  and
  g1946
  (
    n1926,
    n1806,
    n943,
    n1782,
    n1269
  );


  or
  g1947
  (
    n2016,
    n1799,
    n1273,
    n1313,
    n1009
  );


  xnor
  g1948
  (
    n2033,
    n889,
    n1806,
    n1401,
    n1499
  );


  nor
  g1949
  (
    n1971,
    n1080,
    n759,
    n957,
    n1454
  );


  and
  g1950
  (
    n1943,
    n837,
    n789,
    n949,
    n1310
  );


  nand
  g1951
  (
    n1961,
    n1797,
    n1057,
    n855,
    n1496
  );


  nand
  g1952
  (
    n1946,
    n1004,
    n1422,
    n1813,
    n786
  );


  nand
  g1953
  (
    n2029,
    n898,
    n1826,
    n1346,
    n1245
  );


  xor
  g1954
  (
    n1864,
    n1784,
    n1485,
    n1827,
    n1410
  );


  and
  g1955
  (
    n1969,
    n1221,
    n1287,
    n1335,
    n1028
  );


  nor
  g1956
  (
    n2049,
    n1015,
    n1192,
    n939,
    n1116
  );


  and
  g1957
  (
    n1894,
    n1290,
    n1786,
    n807,
    n1791
  );


  and
  g1958
  (
    n2006,
    n1103,
    n907,
    n1812,
    n1121
  );


  xnor
  g1959
  (
    n2008,
    n1778,
    n1791,
    n785,
    n1301
  );


  and
  g1960
  (
    n1967,
    n1817,
    n1828,
    n1784,
    n1488
  );


  nand
  g1961
  (
    n2017,
    n1798,
    n874,
    n1235,
    n1770
  );


  or
  g1962
  (
    n1993,
    n830,
    n1413,
    n1001,
    n1154
  );


  xnor
  g1963
  (
    n1941,
    n1774,
    n1295,
    n750,
    n913
  );


  or
  g1964
  (
    n1860,
    n760,
    n1182,
    n1457,
    n1089
  );


  nor
  g1965
  (
    n1945,
    n1813,
    n1768,
    n999,
    n1219
  );


  nand
  g1966
  (
    n1851,
    n1452,
    n1243,
    n1445,
    n1387
  );


  xor
  g1967
  (
    n2053,
    n1091,
    n1371,
    n1060,
    n870
  );


  nor
  g1968
  (
    n1862,
    n1471,
    n1212,
    n809,
    n836
  );


  or
  g1969
  (
    n1991,
    n1500,
    n1075,
    n747,
    n1783
  );


  xnor
  g1970
  (
    n1850,
    n825,
    n909,
    n1785,
    n1093
  );


  and
  g1971
  (
    n1957,
    n1455,
    n981,
    n976,
    n978
  );


  xor
  g1972
  (
    n2063,
    n1797,
    n988,
    n1051,
    n1086
  );


  xor
  g1973
  (
    n1874,
    n982,
    n1811,
    n1797,
    n1122
  );


  and
  g1974
  (
    n1987,
    n1775,
    n1494,
    n869,
    n1218
  );


  xor
  g1975
  (
    n1970,
    n1475,
    n767,
    n926,
    n1360
  );


  nor
  g1976
  (
    n1909,
    n1136,
    n1774,
    n1184,
    n1157
  );


  or
  g1977
  (
    n2083,
    n1808,
    n1315,
    n1061,
    n1247
  );


  xor
  g1978
  (
    n2004,
    n962,
    n1174,
    n915,
    n829
  );


  xnor
  g1979
  (
    n1892,
    n911,
    n768,
    n952,
    n1076
  );


  nand
  g1980
  (
    n2046,
    n1171,
    n1043,
    n1421,
    n1130
  );


  nor
  g1981
  (
    n2042,
    n753,
    n1155,
    n1772,
    n1206
  );


  xor
  g1982
  (
    n2054,
    n1256,
    n862,
    n971,
    n1118
  );


  xnor
  g1983
  (
    n1912,
    n887,
    n1436,
    n1817,
    n1438
  );


  and
  g1984
  (
    n1931,
    n1271,
    n1483,
    n1825,
    n843
  );


  or
  g1985
  (
    n2080,
    n918,
    n900,
    n1447,
    n1185
  );


  xor
  g1986
  (
    n2002,
    n1175,
    n1799,
    n1144,
    n1456
  );


  xnor
  g1987
  (
    n1921,
    n1816,
    n989,
    n1792,
    n1803
  );


  xnor
  g1988
  (
    n1942,
    n763,
    n1443,
    n1126,
    n1270
  );


  nor
  g1989
  (
    n2051,
    n1779,
    n1780,
    n1178,
    n1790
  );


  and
  g1990
  (
    n1861,
    n1347,
    n743,
    n961,
    n1164
  );


  xnor
  g1991
  (
    n1955,
    n927,
    n1812,
    n1789,
    n1179
  );


  xor
  g1992
  (
    n2078,
    n1372,
    n1785,
    n1006,
    n1092
  );


  nor
  g1993
  (
    n1972,
    n805,
    n757,
    n1385,
    n1779
  );


  xor
  g1994
  (
    n2001,
    n937,
    n1111,
    n1357,
    n1768
  );


  xnor
  g1995
  (
    n1835,
    n1344,
    n1810,
    n956,
    n1099
  );


  or
  g1996
  (
    KeyWire_0_0,
    n828,
    n1795,
    n1048,
    n1467
  );


  and
  g1997
  (
    n1960,
    n1358,
    n1244,
    n1476,
    n1150
  );


  nand
  g1998
  (
    n1933,
    n1490,
    n1788,
    n1814,
    n1133
  );


  nor
  g1999
  (
    n2039,
    n1800,
    n925,
    n1197,
    n798
  );


  nor
  g2000
  (
    n1934,
    n1815,
    n1440,
    n998,
    n1829
  );


  nand
  g2001
  (
    n1976,
    n1427,
    n765,
    n844,
    n872
  );


  or
  g2002
  (
    n1974,
    n1459,
    n1038,
    n1805,
    n1792
  );


  xnor
  g2003
  (
    n1838,
    n1479,
    n1123,
    n1784,
    n754
  );


  xnor
  g2004
  (
    n1981,
    n1012,
    n1468,
    n1823,
    n1462
  );


  or
  g2005
  (
    n1913,
    n965,
    n1816,
    n1105,
    n1429
  );


  nand
  g2006
  (
    n2024,
    n1815,
    n1790,
    n1827,
    n1226
  );


  xor
  g2007
  (
    n2043,
    n1291,
    n1230,
    n950,
    n737
  );


  nor
  g2008
  (
    n1848,
    n1790,
    n773,
    n778,
    n996
  );


  nand
  g2009
  (
    n1873,
    n1773,
    n1396,
    n1145,
    n1124
  );


  nor
  g2010
  (
    n1879,
    n890,
    n1807,
    n1416,
    n1064
  );


  nor
  g2011
  (
    n1901,
    n1480,
    n1781,
    n1341,
    n1825
  );


  xor
  g2012
  (
    n1853,
    n1802,
    n736,
    n875,
    n1363
  );


  nor
  g2013
  (
    n1887,
    n1804,
    n818,
    n735,
    n1790
  );


  and
  g2014
  (
    n1902,
    n1817,
    n802,
    n1804,
    n1314
  );


  xor
  g2015
  (
    n1889,
    n1120,
    n1021,
    n1771,
    n1399
  );


  xnor
  g2016
  (
    n1982,
    n1209,
    n1482,
    n893,
    n1020
  );


  and
  g2017
  (
    n2076,
    n1132,
    n1781,
    n1829,
    n839
  );


  nand
  g2018
  (
    n2005,
    n1783,
    n1355,
    n1017,
    n888
  );


  nand
  g2019
  (
    n2023,
    n1802,
    n1277,
    n1805,
    n1139
  );


  and
  g2020
  (
    n2067,
    n941,
    n1258,
    n1214,
    n1437
  );


  xnor
  g2021
  (
    n2007,
    n1356,
    n1349,
    n794,
    n772
  );


  xor
  g2022
  (
    n2087,
    n1137,
    n1309,
    n1792,
    n1381
  );


  xnor
  g2023
  (
    n2044,
    n1814,
    n1780,
    n931,
    n823
  );


  and
  g2024
  (
    n1930,
    n868,
    n1241,
    n1100,
    n1404
  );


  xnor
  g2025
  (
    n1888,
    n1208,
    n993,
    n1032,
    n1460
  );


  nor
  g2026
  (
    n1880,
    n1198,
    n1079,
    n1165,
    n877
  );


  xor
  g2027
  (
    n1893,
    n940,
    n903,
    n990,
    n1470
  );


  or
  g2028
  (
    n1947,
    n1418,
    n871,
    n1029,
    n1306
  );


  or
  g2029
  (
    n1958,
    n1828,
    n1115,
    n1095,
    n766
  );


  xor
  g2030
  (
    n2037,
    n1194,
    n1793,
    n1276,
    n973
  );


  xor
  g2031
  (
    n1857,
    n1430,
    n1316,
    n1065,
    n793
  );


  or
  g2032
  (
    n1918,
    n791,
    n966,
    n1267,
    n902
  );


  and
  g2033
  (
    n2030,
    n1211,
    n1180,
    n1477,
    n1810
  );


  and
  g2034
  (
    n1966,
    n1320,
    n1063,
    n934,
    n841
  );


  nor
  g2035
  (
    n1897,
    n1318,
    n1094,
    n1272,
    n1348
  );


  nand
  g2036
  (
    n2082,
    n1828,
    n1777,
    n1024,
    n1327
  );


  nor
  g2037
  (
    n1964,
    n916,
    n1769,
    n1334,
    n1771
  );


  and
  g2038
  (
    n2058,
    n1262,
    n1777,
    n738,
    n1305
  );


  nand
  g2039
  (
    KeyWire_0_25,
    n1234,
    n1801,
    n1304,
    n1806
  );


  nand
  g2040
  (
    n1944,
    n813,
    n1796,
    n922,
    n1324
  );


  or
  g2041
  (
    n1869,
    n1340,
    n758,
    n1225,
    n1821
  );


  xnor
  g2042
  (
    n1978,
    n1190,
    n1326,
    n905,
    n885
  );


  nand
  g2043
  (
    n2059,
    n1391,
    n826,
    n1073,
    n1284
  );


  or
  g2044
  (
    n2077,
    n1377,
    n897,
    n1812,
    n1789
  );


  or
  g2045
  (
    n1855,
    n820,
    n1472,
    n1776,
    n1501
  );


  xor
  g2046
  (
    n1867,
    n946,
    n1776,
    n920,
    n1331
  );


  and
  g2047
  (
    n1956,
    n1386,
    n1264,
    n846,
    n919
  );


  or
  g2048
  (
    n1863,
    n1804,
    n969,
    n1787,
    n884
  );


  nand
  g2049
  (
    n1968,
    n1432,
    n806,
    n1254,
    n1819
  );


  nor
  g2050
  (
    n1999,
    n1408,
    n742,
    n842,
    n1058
  );


  and
  g2051
  (
    n1980,
    n815,
    n1794,
    n859,
    n1788
  );


  or
  g2052
  (
    n1990,
    n979,
    n1217,
    n1152,
    n857
  );


  xor
  g2053
  (
    n1872,
    n1818,
    n921,
    n1789,
    n1325
  );


  or
  g2054
  (
    n1927,
    n958,
    n1478,
    n1785,
    n968
  );


  buf
  g2055
  (
    n2088,
    n1839
  );


  not
  g2056
  (
    n2100,
    n1843
  );


  not
  g2057
  (
    n2101,
    n1841
  );


  buf
  g2058
  (
    n2093,
    n1842
  );


  not
  g2059
  (
    n2094,
    n1834
  );


  not
  g2060
  (
    n2095,
    n1838
  );


  buf
  g2061
  (
    n2091,
    n1835
  );


  not
  g2062
  (
    n2102,
    n1846
  );


  buf
  g2063
  (
    n2096,
    n1832
  );


  not
  g2064
  (
    n2090,
    n1845
  );


  buf
  g2065
  (
    n2098,
    n1847
  );


  buf
  g2066
  (
    n2092,
    n1840
  );


  buf
  g2067
  (
    n2099,
    n1836
  );


  not
  g2068
  (
    n2103,
    n1833
  );


  buf
  g2069
  (
    n2089,
    n1844
  );


  not
  g2070
  (
    n2097,
    n1837
  );


  and
  g2071
  (
    n2115,
    n2002,
    n2089,
    n1860,
    n1952
  );


  nor
  g2072
  (
    n2119,
    n2103,
    n1929,
    n1962,
    n1852
  );


  xnor
  g2073
  (
    n2128,
    n1933,
    n2001,
    n1986,
    n1956
  );


  or
  g2074
  (
    n2149,
    n1963,
    n1850,
    n2004,
    n1953
  );


  xnor
  g2075
  (
    n2106,
    n1907,
    n1999,
    n1973,
    n1989
  );


  and
  g2076
  (
    n2134,
    n2098,
    n2098,
    n2008,
    n2095
  );


  nor
  g2077
  (
    n2155,
    n2102,
    n1976,
    n1949,
    n2088
  );


  or
  g2078
  (
    n2156,
    n2028,
    n2038,
    n1982,
    n2089
  );


  nor
  g2079
  (
    n2112,
    n1984,
    n2094,
    n2005,
    n1987
  );


  or
  g2080
  (
    n2126,
    n1859,
    n2099,
    n1883,
    n1926
  );


  and
  g2081
  (
    n2138,
    n1862,
    n1931,
    n2096,
    n2021
  );


  nand
  g2082
  (
    n2153,
    n1851,
    n2094,
    n2006,
    n1897
  );


  nor
  g2083
  (
    n2167,
    n1911,
    n1889,
    n1906,
    n1886
  );


  xnor
  g2084
  (
    n2150,
    n2090,
    n1868,
    n1940,
    n1975
  );


  and
  g2085
  (
    n2116,
    n1932,
    n2017,
    n1864,
    n2089
  );


  and
  g2086
  (
    n2122,
    n2096,
    n2031,
    n1858,
    n1879
  );


  and
  g2087
  (
    n2124,
    n1854,
    n1904,
    n1944,
    n2093
  );


  xnor
  g2088
  (
    n2165,
    n1873,
    n1988,
    n2011,
    n2093
  );


  or
  g2089
  (
    n2154,
    n1857,
    n1939,
    n1855,
    n2100
  );


  or
  g2090
  (
    n2140,
    n2091,
    n2026,
    n2094,
    n2009
  );


  xor
  g2091
  (
    n2120,
    n1994,
    n2102,
    n2095,
    n2016
  );


  or
  g2092
  (
    n2158,
    n2027,
    n1894,
    n1921,
    n1892
  );


  and
  g2093
  (
    n2148,
    n1955,
    n2101,
    n1902,
    n2014
  );


  nand
  g2094
  (
    n2143,
    n2092,
    n2093,
    n1922,
    n1909
  );


  nand
  g2095
  (
    n2139,
    n1877,
    n1856,
    n1848,
    n2088
  );


  nor
  g2096
  (
    n2130,
    n1934,
    n2029,
    n1853,
    n2019
  );


  nor
  g2097
  (
    n2161,
    n1885,
    n1927,
    n2097,
    n1891
  );


  and
  g2098
  (
    n2123,
    n2024,
    n2102,
    n1971,
    n1947
  );


  nand
  g2099
  (
    n2114,
    n2094,
    n2092,
    n2100,
    n1871
  );


  and
  g2100
  (
    n2125,
    n1992,
    n2097,
    n1863,
    n1888
  );


  or
  g2101
  (
    n2141,
    n2102,
    n1887,
    n1866,
    n2032
  );


  xnor
  g2102
  (
    n2109,
    n1959,
    n1914,
    n1919,
    n2091
  );


  and
  g2103
  (
    n2118,
    n1972,
    n2090,
    n1917,
    n1995
  );


  xnor
  g2104
  (
    n2151,
    n1946,
    n2099,
    n1890,
    n1861
  );


  or
  g2105
  (
    n2144,
    n1920,
    n2093,
    n1991,
    n2097
  );


  xnor
  g2106
  (
    n2107,
    n2035,
    n1928,
    n1865,
    n1996
  );


  or
  g2107
  (
    n2146,
    n2095,
    n1980,
    n2088,
    n1936
  );


  and
  g2108
  (
    n2159,
    n1979,
    n1964,
    n1900,
    n1849
  );


  xor
  g2109
  (
    n2137,
    n1908,
    n2022,
    n2095,
    n2000
  );


  nor
  g2110
  (
    n2145,
    n1893,
    n2034,
    n1981,
    n1941
  );


  xor
  g2111
  (
    n2160,
    n2088,
    n2090,
    n1948,
    n1925
  );


  xor
  g2112
  (
    n2162,
    n1872,
    n1896,
    n1874,
    n1951
  );


  xor
  g2113
  (
    n2142,
    n2103,
    n1967,
    n1905,
    n1945
  );


  or
  g2114
  (
    n2117,
    n1942,
    n2037,
    n1913,
    n2096
  );


  xnor
  g2115
  (
    n2129,
    n1918,
    n2103,
    n1977,
    n2091
  );


  nor
  g2116
  (
    n2166,
    n1961,
    n1875,
    n1867,
    n1912
  );


  or
  g2117
  (
    n2127,
    n1960,
    n1882,
    n2089,
    n1878
  );


  xor
  g2118
  (
    n2105,
    n2098,
    n2098,
    n1970,
    n2036
  );


  and
  g2119
  (
    n2163,
    n2099,
    n2092,
    n1916,
    n1899
  );


  xnor
  g2120
  (
    n2135,
    n2018,
    n1876,
    n2097,
    n1998
  );


  nand
  g2121
  (
    n2164,
    n2003,
    n2100,
    n1923,
    n1950
  );


  nor
  g2122
  (
    n2108,
    n1966,
    n1997,
    n1903,
    n1974
  );


  or
  g2123
  (
    n2113,
    n2023,
    n1990,
    n1924,
    n1943
  );


  nand
  g2124
  (
    n2147,
    n2096,
    n1895,
    n1969,
    n1930
  );


  and
  g2125
  (
    n2104,
    n1884,
    n2101,
    n1898,
    n1968
  );


  xor
  g2126
  (
    n2157,
    n1954,
    n2010,
    n1985,
    n2101
  );


  xor
  g2127
  (
    n2132,
    n2091,
    n2092,
    n1938,
    n1993
  );


  nor
  g2128
  (
    n2136,
    n1881,
    n2012,
    n1910,
    n1901
  );


  xor
  g2129
  (
    n2110,
    n2101,
    n2020,
    n2103,
    n2015
  );


  nor
  g2130
  (
    n2133,
    n2100,
    n1935,
    n2099,
    n1957
  );


  xnor
  g2131
  (
    n2152,
    n1937,
    n2090,
    n1965,
    n2033
  );


  nor
  g2132
  (
    n2131,
    n1983,
    n2039,
    n1958,
    n2025
  );


  nor
  g2133
  (
    n2111,
    n1915,
    n2030,
    n1869,
    n1880
  );


  nor
  g2134
  (
    n2121,
    n2013,
    n1978,
    n2007,
    n1870
  );


  not
  g2135
  (
    n2359,
    n2157
  );


  not
  g2136
  (
    n2188,
    n2158
  );


  not
  g2137
  (
    n2262,
    n2156
  );


  not
  g2138
  (
    n2297,
    n2142
  );


  buf
  g2139
  (
    n2391,
    n2114
  );


  not
  g2140
  (
    n2375,
    n2117
  );


  not
  g2141
  (
    n2384,
    n2161
  );


  not
  g2142
  (
    n2405,
    n2122
  );


  not
  g2143
  (
    n2390,
    n2115
  );


  not
  g2144
  (
    n2292,
    n2137
  );


  buf
  g2145
  (
    n2382,
    n2114
  );


  not
  g2146
  (
    n2303,
    n2127
  );


  buf
  g2147
  (
    n2175,
    n2120
  );


  not
  g2148
  (
    n2234,
    n2141
  );


  buf
  g2149
  (
    n2257,
    n2110
  );


  buf
  g2150
  (
    n2369,
    n2158
  );


  buf
  g2151
  (
    n2399,
    n2120
  );


  not
  g2152
  (
    n2207,
    n2160
  );


  not
  g2153
  (
    n2247,
    n2111
  );


  not
  g2154
  (
    n2228,
    n2153
  );


  not
  g2155
  (
    n2316,
    n2149
  );


  buf
  g2156
  (
    n2256,
    n2142
  );


  buf
  g2157
  (
    n2306,
    n2042
  );


  not
  g2158
  (
    n2187,
    n2125
  );


  buf
  g2159
  (
    n2356,
    n2047
  );


  not
  g2160
  (
    n2261,
    n2130
  );


  buf
  g2161
  (
    KeyWire_0_2,
    n2148
  );


  not
  g2162
  (
    n2218,
    n2124
  );


  not
  g2163
  (
    n2330,
    n2128
  );


  not
  g2164
  (
    n2268,
    n2109
  );


  buf
  g2165
  (
    n2420,
    n2136
  );


  buf
  g2166
  (
    n2289,
    n2118
  );


  not
  g2167
  (
    n2346,
    n2129
  );


  not
  g2168
  (
    n2329,
    n2134
  );


  buf
  g2169
  (
    n2393,
    n2162
  );


  buf
  g2170
  (
    n2348,
    n2117
  );


  buf
  g2171
  (
    n2418,
    n2142
  );


  not
  g2172
  (
    n2362,
    n2144
  );


  buf
  g2173
  (
    n2370,
    n2166
  );


  buf
  g2174
  (
    n2395,
    n2044
  );


  buf
  g2175
  (
    n2322,
    n2119
  );


  buf
  g2176
  (
    n2296,
    n2162
  );


  not
  g2177
  (
    n2217,
    n2160
  );


  not
  g2178
  (
    n2194,
    n2154
  );


  buf
  g2179
  (
    n2233,
    n2110
  );


  buf
  g2180
  (
    n2349,
    n2147
  );


  buf
  g2181
  (
    n2170,
    n2107
  );


  buf
  g2182
  (
    n2396,
    n2112
  );


  buf
  g2183
  (
    n2332,
    n2148
  );


  buf
  g2184
  (
    n2220,
    n2137
  );


  not
  g2185
  (
    n2350,
    n2157
  );


  buf
  g2186
  (
    n2397,
    n2164
  );


  not
  g2187
  (
    n2229,
    n2129
  );


  not
  g2188
  (
    n2421,
    n2107
  );


  not
  g2189
  (
    n2224,
    n2150
  );


  buf
  g2190
  (
    n2291,
    n2048
  );


  not
  g2191
  (
    n2254,
    n2133
  );


  buf
  g2192
  (
    n2266,
    n2135
  );


  buf
  g2193
  (
    n2341,
    n2124
  );


  not
  g2194
  (
    n2342,
    n2157
  );


  not
  g2195
  (
    n2377,
    n2144
  );


  not
  g2196
  (
    n2172,
    n2162
  );


  not
  g2197
  (
    n2244,
    n2111
  );


  not
  g2198
  (
    n2290,
    n2118
  );


  buf
  g2199
  (
    n2237,
    n2115
  );


  not
  g2200
  (
    n2352,
    n2116
  );


  not
  g2201
  (
    n2400,
    n2129
  );


  not
  g2202
  (
    n2406,
    n2138
  );


  not
  g2203
  (
    n2408,
    n2110
  );


  not
  g2204
  (
    n2318,
    n2164
  );


  not
  g2205
  (
    n2223,
    n2165
  );


  not
  g2206
  (
    n2199,
    n2137
  );


  buf
  g2207
  (
    n2381,
    n2166
  );


  not
  g2208
  (
    n2295,
    n2163
  );


  not
  g2209
  (
    n2190,
    n2121
  );


  not
  g2210
  (
    n2325,
    n2127
  );


  buf
  g2211
  (
    n2221,
    n2130
  );


  buf
  g2212
  (
    n2317,
    n2045
  );


  buf
  g2213
  (
    n2312,
    n2138
  );


  not
  g2214
  (
    n2238,
    n2113
  );


  not
  g2215
  (
    KeyWire_0_6,
    n2136
  );


  not
  g2216
  (
    n2275,
    n2130
  );


  not
  g2217
  (
    n2222,
    n2147
  );


  not
  g2218
  (
    n2378,
    n2126
  );


  buf
  g2219
  (
    n2376,
    n2041
  );


  not
  g2220
  (
    n2271,
    n2105
  );


  not
  g2221
  (
    n2183,
    n2131
  );


  not
  g2222
  (
    n2281,
    n2139
  );


  buf
  g2223
  (
    n2209,
    n2163
  );


  not
  g2224
  (
    n2205,
    n2128
  );


  not
  g2225
  (
    n2307,
    n2133
  );


  not
  g2226
  (
    n2358,
    n2144
  );


  not
  g2227
  (
    n2351,
    n2167
  );


  buf
  g2228
  (
    n2213,
    n2106
  );


  not
  g2229
  (
    n2182,
    n2131
  );


  not
  g2230
  (
    n2284,
    n2155
  );


  not
  g2231
  (
    n2294,
    n2159
  );


  buf
  g2232
  (
    n2343,
    n2152
  );


  buf
  g2233
  (
    n2227,
    n2164
  );


  buf
  g2234
  (
    n2176,
    n2111
  );


  buf
  g2235
  (
    n2354,
    n2124
  );


  not
  g2236
  (
    n2301,
    n2119
  );


  not
  g2237
  (
    n2265,
    n2110
  );


  not
  g2238
  (
    n2302,
    n2140
  );


  not
  g2239
  (
    n2260,
    n2148
  );


  not
  g2240
  (
    n2267,
    n2150
  );


  not
  g2241
  (
    n2272,
    n2109
  );


  buf
  g2242
  (
    n2315,
    n2106
  );


  buf
  g2243
  (
    n2360,
    n2126
  );


  buf
  g2244
  (
    n2401,
    n2166
  );


  buf
  g2245
  (
    n2410,
    n2113
  );


  not
  g2246
  (
    n2327,
    n2136
  );


  not
  g2247
  (
    n2347,
    n2046
  );


  not
  g2248
  (
    n2423,
    n2125
  );


  buf
  g2249
  (
    n2285,
    n2164
  );


  buf
  g2250
  (
    n2345,
    n2159
  );


  not
  g2251
  (
    n2404,
    n2135
  );


  buf
  g2252
  (
    n2311,
    n2126
  );


  buf
  g2253
  (
    n2235,
    n2121
  );


  not
  g2254
  (
    n2252,
    n2143
  );


  not
  g2255
  (
    n2251,
    n2107
  );


  not
  g2256
  (
    n2365,
    n2141
  );


  not
  g2257
  (
    n2240,
    n2163
  );


  not
  g2258
  (
    n2246,
    n2160
  );


  buf
  g2259
  (
    n2208,
    n2140
  );


  not
  g2260
  (
    n2402,
    n2116
  );


  not
  g2261
  (
    n2214,
    n2121
  );


  buf
  g2262
  (
    n2189,
    n2122
  );


  buf
  g2263
  (
    n2200,
    n2114
  );


  buf
  g2264
  (
    n2243,
    n2120
  );


  not
  g2265
  (
    n2274,
    n2125
  );


  not
  g2266
  (
    n2344,
    n2155
  );


  not
  g2267
  (
    n2407,
    n2165
  );


  not
  g2268
  (
    n2270,
    n2122
  );


  buf
  g2269
  (
    n2269,
    n2125
  );


  buf
  g2270
  (
    n2336,
    n2104
  );


  not
  g2271
  (
    n2203,
    n2161
  );


  not
  g2272
  (
    n2409,
    n2108
  );


  not
  g2273
  (
    n2184,
    n2113
  );


  buf
  g2274
  (
    n2250,
    n2140
  );


  buf
  g2275
  (
    n2273,
    n2123
  );


  buf
  g2276
  (
    n2334,
    n2137
  );


  buf
  g2277
  (
    n2174,
    n2112
  );


  not
  g2278
  (
    n2193,
    n2104
  );


  not
  g2279
  (
    n2201,
    n2108
  );


  not
  g2280
  (
    n2185,
    n2154
  );


  buf
  g2281
  (
    n2278,
    n2156
  );


  not
  g2282
  (
    n2216,
    n2116
  );


  not
  g2283
  (
    n2263,
    n2156
  );


  not
  g2284
  (
    n2309,
    n2152
  );


  not
  g2285
  (
    n2198,
    n2123
  );


  not
  g2286
  (
    n2392,
    n2167
  );


  buf
  g2287
  (
    n2379,
    n2128
  );


  not
  g2288
  (
    n2171,
    n2158
  );


  buf
  g2289
  (
    n2245,
    n2117
  );


  not
  g2290
  (
    n2286,
    n2148
  );


  not
  g2291
  (
    n2355,
    n2114
  );


  not
  g2292
  (
    n2353,
    n2145
  );


  buf
  g2293
  (
    n2398,
    n2167
  );


  buf
  g2294
  (
    n2264,
    n2146
  );


  buf
  g2295
  (
    n2416,
    n2145
  );


  buf
  g2296
  (
    n2372,
    n2139
  );


  not
  g2297
  (
    n2298,
    n2119
  );


  not
  g2298
  (
    n2422,
    n2116
  );


  not
  g2299
  (
    n2259,
    n2141
  );


  not
  g2300
  (
    n2367,
    n2128
  );


  buf
  g2301
  (
    n2202,
    n2151
  );


  not
  g2302
  (
    n2196,
    n2156
  );


  not
  g2303
  (
    n2232,
    n2132
  );


  buf
  g2304
  (
    n2305,
    n2131
  );


  buf
  g2305
  (
    n2321,
    n2133
  );


  buf
  g2306
  (
    n2253,
    n2158
  );


  not
  g2307
  (
    n2191,
    n2112
  );


  buf
  g2308
  (
    n2282,
    n2149
  );


  not
  g2309
  (
    n2168,
    n2133
  );


  buf
  g2310
  (
    n2192,
    n2138
  );


  not
  g2311
  (
    n2197,
    n2120
  );


  buf
  g2312
  (
    n2323,
    n2127
  );


  buf
  g2313
  (
    n2279,
    n2165
  );


  buf
  g2314
  (
    n2419,
    n2108
  );


  not
  g2315
  (
    n2413,
    n2145
  );


  buf
  g2316
  (
    n2241,
    n2108
  );


  not
  g2317
  (
    n2283,
    n2153
  );


  not
  g2318
  (
    n2374,
    n2115
  );


  not
  g2319
  (
    KeyWire_0_24,
    n2111
  );


  buf
  g2320
  (
    KeyWire_0_8,
    n2161
  );


  buf
  g2321
  (
    n2339,
    n2104
  );


  not
  g2322
  (
    n2331,
    n2152
  );


  not
  g2323
  (
    n2366,
    n2109
  );


  not
  g2324
  (
    n2368,
    n2139
  );


  buf
  g2325
  (
    n2324,
    n2155
  );


  not
  g2326
  (
    n2337,
    n2130
  );


  buf
  g2327
  (
    n2206,
    n2115
  );


  not
  g2328
  (
    n2226,
    n2152
  );


  buf
  g2329
  (
    n2373,
    n2105
  );


  buf
  g2330
  (
    n2304,
    n2143
  );


  not
  g2331
  (
    n2338,
    n2153
  );


  not
  g2332
  (
    n2255,
    n2144
  );


  not
  g2333
  (
    n2319,
    n2132
  );


  buf
  g2334
  (
    n2415,
    n2109
  );


  not
  g2335
  (
    n2333,
    n2147
  );


  not
  g2336
  (
    n2389,
    n2132
  );


  buf
  g2337
  (
    n2371,
    n2105
  );


  not
  g2338
  (
    n2380,
    n2040
  );


  not
  g2339
  (
    n2411,
    n2105
  );


  buf
  g2340
  (
    n2287,
    n2127
  );


  not
  g2341
  (
    n2277,
    n2149
  );


  buf
  g2342
  (
    n2186,
    n2142
  );


  not
  g2343
  (
    n2231,
    n2122
  );


  not
  g2344
  (
    n2387,
    n2143
  );


  not
  g2345
  (
    n2364,
    n2150
  );


  not
  g2346
  (
    n2299,
    n2134
  );


  not
  g2347
  (
    n2328,
    n2106
  );


  not
  g2348
  (
    n2204,
    n2161
  );


  not
  g2349
  (
    n2177,
    n2118
  );


  not
  g2350
  (
    n2388,
    n2132
  );


  buf
  g2351
  (
    n2340,
    n2145
  );


  not
  g2352
  (
    n2249,
    n2131
  );


  not
  g2353
  (
    n2403,
    n2136
  );


  buf
  g2354
  (
    n2361,
    n2149
  );


  buf
  g2355
  (
    n2414,
    n2151
  );


  not
  g2356
  (
    n2417,
    n2117
  );


  not
  g2357
  (
    n2248,
    n2150
  );


  buf
  g2358
  (
    n2230,
    n2119
  );


  not
  g2359
  (
    n2313,
    n2162
  );


  not
  g2360
  (
    n2293,
    n2163
  );


  buf
  g2361
  (
    n2276,
    n2126
  );


  not
  g2362
  (
    n2320,
    n2107
  );


  not
  g2363
  (
    n2363,
    n2129
  );


  buf
  g2364
  (
    n2385,
    n2123
  );


  buf
  g2365
  (
    n2210,
    n2166
  );


  buf
  g2366
  (
    n2236,
    n2124
  );


  buf
  g2367
  (
    n2280,
    n2123
  );


  not
  g2368
  (
    n2225,
    n2146
  );


  buf
  g2369
  (
    n2211,
    n2104
  );


  not
  g2370
  (
    n2178,
    n2154
  );


  buf
  g2371
  (
    n2288,
    n2147
  );


  buf
  g2372
  (
    n2219,
    n2151
  );


  buf
  g2373
  (
    n2212,
    n2118
  );


  buf
  g2374
  (
    n2169,
    n2160
  );


  buf
  g2375
  (
    n2394,
    n2134
  );


  buf
  g2376
  (
    n2326,
    n2153
  );


  buf
  g2377
  (
    n2239,
    n2106
  );


  not
  g2378
  (
    n2335,
    n2135
  );


  not
  g2379
  (
    n2180,
    n2159
  );


  buf
  g2380
  (
    n2195,
    n2134
  );


  buf
  g2381
  (
    n2179,
    n2154
  );


  buf
  g2382
  (
    n2386,
    n2146
  );


  buf
  g2383
  (
    n2308,
    n2139
  );


  not
  g2384
  (
    n2181,
    n2140
  );


  not
  g2385
  (
    n2314,
    n2155
  );


  buf
  g2386
  (
    n2383,
    n2143
  );


  buf
  g2387
  (
    n2310,
    n2141
  );


  xnor
  g2388
  (
    n2412,
    n2167,
    n2135,
    n2146,
    n2121
  );


  nand
  g2389
  (
    n2300,
    n2159,
    n2157,
    n2113,
    n2112
  );


  or
  g2390
  (
    n2258,
    n2151,
    n2138,
    n2165,
    n2043
  );


  and
  g2391
  (
    n2424,
    n2168,
    n2049
  );


  not
  g2392
  (
    n2425,
    n2424
  );


  nor
  g2393
  (
    n2426,
    n2424,
    n2050
  );


  xor
  g2394
  (
    n2428,
    n2425,
    n2053
  );


  nand
  g2395
  (
    n2427,
    n2056,
    n2055,
    n2425
  );


  and
  g2396
  (
    n2429,
    n2057,
    n2052,
    n2054,
    n2051
  );


  or
  g2397
  (
    n2431,
    n2174,
    n2171,
    n1722,
    n2179
  );


  xnor
  g2398
  (
    n2435,
    n2429,
    n2173,
    n2183,
    n2176
  );


  or
  g2399
  (
    n2433,
    n2184,
    n2429,
    n2428,
    n2180
  );


  and
  g2400
  (
    n2437,
    n2177,
    n2169,
    n2429,
    n2427
  );


  nand
  g2401
  (
    n2430,
    n2175,
    n2429,
    n2178,
    n2182
  );


  xnor
  g2402
  (
    n2432,
    n2170,
    n2181,
    n2061,
    n1721
  );


  nor
  g2403
  (
    n2434,
    n2172,
    n1503,
    n2060,
    n2058
  );


  nand
  g2404
  (
    n2436,
    n2428,
    n2428,
    n2185,
    n2059
  );


  not
  g2405
  (
    n2438,
    n2434
  );


  not
  g2406
  (
    n2443,
    n2433
  );


  buf
  g2407
  (
    n2442,
    n2436
  );


  not
  g2408
  (
    n2445,
    n2435
  );


  and
  g2409
  (
    n2441,
    n2062,
    n2063,
    n2437
  );


  nor
  g2410
  (
    n2440,
    n2431,
    n2064,
    n2065
  );


  xor
  g2411
  (
    n2439,
    n2430,
    n2067,
    n2066
  );


  or
  g2412
  (
    n2444,
    n2068,
    n1726,
    n2432
  );


  not
  g2413
  (
    n2446,
    n1504
  );


  buf
  g2414
  (
    n2449,
    n2439
  );


  not
  g2415
  (
    n2452,
    n2439
  );


  not
  g2416
  (
    n2453,
    n2443
  );


  buf
  g2417
  (
    n2448,
    n2426
  );


  buf
  g2418
  (
    n2463,
    n2444
  );


  buf
  g2419
  (
    n2447,
    n2439
  );


  not
  g2420
  (
    n2451,
    n2442
  );


  not
  g2421
  (
    n2456,
    n2441
  );


  not
  g2422
  (
    n2450,
    n2443
  );


  not
  g2423
  (
    n2461,
    n2445
  );


  or
  g2424
  (
    n2465,
    n2186,
    n2441,
    n2438
  );


  or
  g2425
  (
    n2459,
    n2442,
    n2439,
    n2443
  );


  or
  g2426
  (
    n2462,
    n2444,
    n2438,
    n2445
  );


  nand
  g2427
  (
    n2458,
    n2438,
    n2441
  );


  and
  g2428
  (
    n2464,
    n2440,
    n2444,
    n2425
  );


  xnor
  g2429
  (
    n2457,
    n2445,
    n2440
  );


  or
  g2430
  (
    n2455,
    n2426,
    n2442,
    n2440
  );


  and
  g2431
  (
    n2460,
    n2444,
    n2438,
    n2445
  );


  xor
  g2432
  (
    n2454,
    n2443,
    n2426,
    n2442
  );


  nor
  g2433
  (
    n2468,
    n2465,
    n2464,
    n2457,
    n2456
  );


  xor
  g2434
  (
    n2467,
    n2461,
    n2458,
    n2459,
    n2453
  );


  and
  g2435
  (
    n2466,
    n2462,
    n2446,
    n2452,
    n2455
  );


  nand
  g2436
  (
    n2469,
    n2451,
    n2454,
    n2463,
    n2449
  );


  or
  g2437
  (
    n2470,
    n2460,
    n2448,
    n2447,
    n2450
  );


  and
  g2438
  (
    n2474,
    n2466,
    n1747,
    n1745
  );


  nor
  g2439
  (
    n2472,
    n2469,
    n1746,
    n1745,
    n1747
  );


  nand
  g2440
  (
    n2471,
    n1745,
    n1744,
    n1746,
    n2467
  );


  and
  g2441
  (
    n2475,
    n1745,
    n2470
  );


  nand
  g2442
  (
    n2476,
    n1747,
    n1746,
    n2465
  );


  xnor
  g2443
  (
    n2473,
    n2468,
    n2465,
    n2470
  );


  not
  g2444
  (
    n2477,
    n2473
  );


  buf
  g2445
  (
    n2478,
    n2472
  );


  not
  g2446
  (
    n2479,
    n2477
  );


  buf
  g2447
  (
    n2481,
    n2479
  );


  buf
  g2448
  (
    n2480,
    n2479
  );


  and
  g2449
  (
    n2482,
    n2481,
    n2069,
    n2070,
    n2071
  );


  nand
  g2450
  (
    n2483,
    n2082,
    n2076,
    n2074,
    n2482
  );


  and
  g2451
  (
    n2484,
    n2081,
    n2073,
    n2075,
    n2083
  );


  xnor
  g2452
  (
    n2485,
    n2482,
    n2077,
    n2078,
    n2079
  );


  xnor
  g2453
  (
    n2486,
    n2482,
    n2482,
    n2072,
    n2080
  );


  xor
  g2454
  (
    n2495,
    n2483,
    n1690,
    n1687
  );


  xnor
  g2455
  (
    n2490,
    n2476,
    n2479,
    n670,
    n667
  );


  nand
  g2456
  (
    n2489,
    n667,
    n1690,
    n2486,
    n1689
  );


  xor
  g2457
  (
    n2493,
    n669,
    n2475,
    n2478,
    n666
  );


  xor
  g2458
  (
    n2500,
    n1688,
    n2486,
    n2485,
    n668
  );


  xnor
  g2459
  (
    n2492,
    n2478,
    n667,
    n668,
    n669
  );


  xnor
  g2460
  (
    n2496,
    n2484,
    n2486,
    n669,
    n672
  );


  nand
  g2461
  (
    n2488,
    n2485,
    n2484,
    n666
  );


  nand
  g2462
  (
    n2498,
    n667,
    n671
  );


  xnor
  g2463
  (
    n2487,
    n1689,
    n1688,
    n2479,
    n670
  );


  and
  g2464
  (
    n2491,
    n1689,
    n671,
    n1688
  );


  and
  g2465
  (
    n2499,
    n668,
    n672,
    n2485
  );


  and
  g2466
  (
    n2501,
    n2474,
    n668,
    n2484,
    n2478
  );


  xnor
  g2467
  (
    n2497,
    n666,
    n669,
    n2483,
    n1687
  );


  nand
  g2468
  (
    n2494,
    n1689,
    n2486,
    n670,
    n2483
  );


  xnor
  g2469
  (
    n2502,
    n670,
    n672,
    n1690,
    n2483
  );


  or
  g2470
  (
    n2560,
    n2488,
    n1670,
    n1666,
    n1671
  );


  nand
  g2471
  (
    n2566,
    n1665,
    n1664,
    n1649,
    n1594
  );


  and
  g2472
  (
    n2555,
    n1522,
    n2492,
    n1625,
    n2489
  );


  nand
  g2473
  (
    n2552,
    n1630,
    n1667,
    n1552,
    n1521
  );


  and
  g2474
  (
    n2542,
    n1571,
    n1621,
    n1559,
    n1548
  );


  and
  g2475
  (
    n2508,
    n1590,
    n1666,
    n2495,
    n1567
  );


  nand
  g2476
  (
    n2512,
    n1624,
    n2500,
    n1514,
    n1664
  );


  and
  g2477
  (
    n2506,
    n2489,
    n1572,
    n1627,
    n1592
  );


  xnor
  g2478
  (
    n2534,
    n1553,
    n2502,
    n2496,
    n1545
  );


  xnor
  g2479
  (
    n2561,
    n1565,
    n2490,
    n1637
  );


  or
  g2480
  (
    n2524,
    n1526,
    n1668,
    n1609,
    n2487
  );


  xor
  g2481
  (
    n2537,
    n2496,
    n1511,
    n1507,
    n1603
  );


  xor
  g2482
  (
    n2526,
    n1596,
    n2491,
    n1554,
    n1651
  );


  and
  g2483
  (
    n2531,
    n1640,
    n1658,
    n1574,
    n1615
  );


  nor
  g2484
  (
    n2541,
    n1585,
    n1528,
    n1669,
    n1519
  );


  xor
  g2485
  (
    n2503,
    n1670,
    n2500,
    n1668,
    n1632
  );


  and
  g2486
  (
    n2504,
    n1599,
    n1646,
    n2499,
    n2495
  );


  or
  g2487
  (
    n2547,
    n1588,
    n1600,
    n1628,
    n2501
  );


  and
  g2488
  (
    n2551,
    n1669,
    n1558,
    n1619,
    n2492
  );


  or
  g2489
  (
    n2538,
    n1648,
    n1647,
    n1612,
    n1510
  );


  xor
  g2490
  (
    n2523,
    n1509,
    n1587,
    n1541,
    n1529
  );


  or
  g2491
  (
    n2540,
    n1569,
    n1655,
    n1543,
    n2499
  );


  xor
  g2492
  (
    n2565,
    n2487,
    n2187,
    n1616,
    n1629
  );


  xor
  g2493
  (
    n2521,
    n1527,
    n1520,
    n1668,
    n1666
  );


  nand
  g2494
  (
    n2527,
    n1670,
    n2493,
    n1557,
    n1668
  );


  xnor
  g2495
  (
    n2511,
    n1589,
    n1638,
    n1532,
    n1608
  );


  xor
  g2496
  (
    n2563,
    n1611,
    n1652,
    n2490,
    n1622
  );


  nor
  g2497
  (
    n2557,
    n2487,
    n1582,
    n2494,
    n1636
  );


  nand
  g2498
  (
    n2553,
    n1644,
    n1579,
    n1650,
    n1606
  );


  xor
  g2499
  (
    n2554,
    n2500,
    n2488,
    n1597,
    n1568
  );


  xnor
  g2500
  (
    n2515,
    n2497,
    n1665,
    n1657,
    n1563
  );


  xnor
  g2501
  (
    n2518,
    n2497,
    n2502,
    n1653,
    n1660
  );


  and
  g2502
  (
    n2507,
    n1605,
    n1670,
    n2490,
    n1620
  );


  nand
  g2503
  (
    n2539,
    n1515,
    n1523,
    n1536,
    n1566
  );


  xnor
  g2504
  (
    n2544,
    n1533,
    n1583,
    n1584,
    n2498
  );


  xnor
  g2505
  (
    n2558,
    n1535,
    n2499,
    n2491,
    n1560
  );


  nand
  g2506
  (
    n2536,
    n1549,
    n1601,
    n1561,
    n1581
  );


  or
  g2507
  (
    n2505,
    n2497,
    n1671,
    n2492,
    n1662
  );


  xor
  g2508
  (
    n2514,
    n1531,
    n1617,
    n1564,
    n1551
  );


  nand
  g2509
  (
    n2529,
    n1614,
    n1595,
    n1671,
    n1661
  );


  xnor
  g2510
  (
    n2550,
    n1576,
    n1642,
    n1659,
    n1604
  );


  nor
  g2511
  (
    n2556,
    n1556,
    n2501,
    n2493,
    n1580
  );


  xor
  g2512
  (
    n2543,
    n1534,
    n1634,
    n2499,
    n1643
  );


  xnor
  g2513
  (
    n2520,
    n2497,
    n2488,
    n1525,
    n1573
  );


  and
  g2514
  (
    n2516,
    n1663,
    n1664,
    n1610,
    n1555
  );


  nor
  g2515
  (
    n2562,
    n1665,
    n2501,
    n1669,
    n1570
  );


  or
  g2516
  (
    n2510,
    n1607,
    n1667,
    n1578,
    n1575
  );


  and
  g2517
  (
    n2548,
    n1635,
    n1645,
    n1506,
    n1665
  );


  and
  g2518
  (
    n2532,
    n2495,
    n2496,
    n1602,
    n1669
  );


  xnor
  g2519
  (
    n2546,
    n1654,
    n1626,
    n1539,
    n1513
  );


  nor
  g2520
  (
    n2517,
    n2502,
    n1623,
    n2488,
    n1671
  );


  xor
  g2521
  (
    n2535,
    n2487,
    n2492,
    n1591,
    n1544
  );


  nor
  g2522
  (
    n2530,
    n2494,
    n2495,
    n2501,
    n2491
  );


  xnor
  g2523
  (
    n2564,
    n1577,
    n2498,
    n2489,
    n2496
  );


  and
  g2524
  (
    n2519,
    n1538,
    n1516,
    n1547,
    n1631
  );


  or
  g2525
  (
    n2513,
    n1518,
    n2489,
    n1633,
    n1667
  );


  nand
  g2526
  (
    n2528,
    n2498,
    n1618,
    n1664,
    n2494
  );


  and
  g2527
  (
    n2545,
    n1542,
    n2491,
    n1666,
    n1586
  );


  xnor
  g2528
  (
    n2522,
    n2493,
    n1593,
    n1641,
    n1546
  );


  and
  g2529
  (
    n2509,
    n1512,
    n1550,
    n1517,
    n1505
  );


  nor
  g2530
  (
    n2549,
    n1613,
    n1508,
    n1562,
    n2502
  );


  nand
  g2531
  (
    n2559,
    n1524,
    n1530,
    n1656,
    n1537
  );


  xor
  g2532
  (
    n2525,
    n2493,
    n1540,
    n1667,
    n2498
  );


  nand
  g2533
  (
    n2533,
    n1639,
    n1598,
    n2500,
    n2494
  );


  nand
  g2534
  (
    n2806,
    n2251,
    n2550,
    n2357,
    n2318
  );


  nor
  g2535
  (
    n2673,
    n2528,
    n2262,
    n2404,
    n2562
  );


  xor
  g2536
  (
    n2785,
    n2314,
    n2377,
    n2541,
    n2254
  );


  xnor
  g2537
  (
    n2651,
    n2560,
    n2279,
    n2355,
    n2328
  );


  xnor
  g2538
  (
    n2778,
    n2287,
    n2508,
    n2522,
    n2364
  );


  xnor
  g2539
  (
    n2708,
    n2331,
    n2514,
    n2534,
    n2322
  );


  xor
  g2540
  (
    n2751,
    n2335,
    n2319,
    n2275,
    n2258
  );


  or
  g2541
  (
    n2764,
    n2409,
    n2547,
    n2524,
    n2269
  );


  xor
  g2542
  (
    n2781,
    n2263,
    n2566,
    n2390,
    n2514
  );


  or
  g2543
  (
    n2570,
    n2325,
    n2556,
    n2221,
    n2566
  );


  nor
  g2544
  (
    n2747,
    n2263,
    n2385,
    n2277,
    n2543
  );


  or
  g2545
  (
    n2592,
    n2287,
    n2403,
    n2209,
    n2253
  );


  xnor
  g2546
  (
    n2780,
    n2318,
    n2418,
    n2304,
    n2382
  );


  or
  g2547
  (
    n2646,
    n2535,
    n2362,
    n2415,
    n2345
  );


  or
  g2548
  (
    n2754,
    n2337,
    n2311,
    n2365,
    n2278
  );


  xnor
  g2549
  (
    n2640,
    n2556,
    n2551,
    n2405,
    n2303
  );


  xor
  g2550
  (
    n2614,
    n2368,
    n2537,
    n2319,
    n2383
  );


  and
  g2551
  (
    n2576,
    n2268,
    n2279,
    n2337,
    n2544
  );


  or
  g2552
  (
    n2740,
    n2378,
    n2413,
    n2229,
    n2311
  );


  nand
  g2553
  (
    n2627,
    n2358,
    n2523,
    n2373,
    n2310
  );


  nand
  g2554
  (
    n2571,
    n2416,
    n2365,
    n2259,
    n2418
  );


  or
  g2555
  (
    n2761,
    n2423,
    n2282,
    n2321,
    n2522
  );


  or
  g2556
  (
    n2729,
    n2309,
    n2272,
    n2190,
    n2247
  );


  xnor
  g2557
  (
    n2741,
    n2328,
    n2552,
    n2419,
    n2400
  );


  and
  g2558
  (
    n2587,
    n2359,
    n2245,
    n2372,
    n2252
  );


  nor
  g2559
  (
    n2767,
    n2319,
    n2281,
    n2530,
    n2346
  );


  nor
  g2560
  (
    n2677,
    n2529,
    n2283,
    n2294,
    n2516
  );


  xor
  g2561
  (
    n2691,
    n2192,
    n2195,
    n2520,
    n2545
  );


  xnor
  g2562
  (
    n2765,
    n2564,
    n2307,
    n2558,
    n2295
  );


  nor
  g2563
  (
    n2804,
    n2289,
    n2286,
    n2533,
    n2285
  );


  or
  g2564
  (
    n2714,
    n2313,
    n2399,
    n2260,
    n2288
  );


  or
  g2565
  (
    n2567,
    n2357,
    n2364,
    n2547,
    n2407
  );


  nand
  g2566
  (
    n2750,
    n2270,
    n2414,
    n2272,
    n2507
  );


  and
  g2567
  (
    n2688,
    n2292,
    n2352,
    n2249,
    n2416
  );


  nor
  g2568
  (
    n2628,
    n2367,
    n2553,
    n2307,
    n2532
  );


  nand
  g2569
  (
    n2649,
    n2294,
    n2305,
    n2556,
    n2255
  );


  nor
  g2570
  (
    n2744,
    n2523,
    n2519,
    n2248,
    n2266
  );


  nand
  g2571
  (
    n2577,
    n2309,
    n2352,
    n2290,
    n2303
  );


  and
  g2572
  (
    n2757,
    n2259,
    n2360,
    n2376,
    n2326
  );


  nor
  g2573
  (
    n2784,
    n2246,
    n2421,
    n2329,
    n2507
  );


  xor
  g2574
  (
    n2656,
    n2216,
    n2250,
    n2402,
    n2509
  );


  nor
  g2575
  (
    n2706,
    n2415,
    n2387,
    n2267,
    n2297
  );


  xor
  g2576
  (
    n2760,
    n2207,
    n2331,
    n2559,
    n2256
  );


  and
  g2577
  (
    n2600,
    n2369,
    n2339,
    n2261,
    n2338
  );


  and
  g2578
  (
    n2623,
    n2189,
    n2331,
    n2390,
    n2292
  );


  nand
  g2579
  (
    n2632,
    n2199,
    n2526,
    n2382,
    n2419
  );


  nor
  g2580
  (
    n2642,
    n2421,
    n2542,
    n2322,
    n2553
  );


  xor
  g2581
  (
    n2715,
    n2384,
    n2222,
    n2512,
    n2372
  );


  xnor
  g2582
  (
    n2589,
    n2294,
    n2512,
    n2380,
    n2300
  );


  xor
  g2583
  (
    n2805,
    n2410,
    n2283,
    n2316,
    n2503
  );


  xor
  g2584
  (
    n2783,
    n2342,
    n2321,
    n2196,
    n2340
  );


  or
  g2585
  (
    n2618,
    n2398,
    n2344,
    n2325,
    n2518
  );


  nor
  g2586
  (
    n2652,
    n2536,
    n2365,
    n2362,
    n2524
  );


  or
  g2587
  (
    n2680,
    n2374,
    n2220,
    n2402,
    n2521
  );


  xor
  g2588
  (
    n2599,
    n2295,
    n2266,
    n2548,
    n2505
  );


  xnor
  g2589
  (
    n2746,
    n2563,
    n2249,
    n2547,
    n2398
  );


  xor
  g2590
  (
    n2768,
    n2251,
    n2371,
    n2308,
    n2316
  );


  and
  g2591
  (
    n2631,
    n2331,
    n2290,
    n2298,
    n2347
  );


  or
  g2592
  (
    n2572,
    n2535,
    n2348,
    n2404,
    n2363
  );


  nor
  g2593
  (
    n2772,
    n2276,
    n2418,
    n2291,
    n2390
  );


  xor
  g2594
  (
    n2724,
    n2293,
    n2297,
    n2421,
    n2359
  );


  or
  g2595
  (
    n2758,
    n2296,
    n2303,
    n2420,
    n2388
  );


  xnor
  g2596
  (
    n2734,
    n2253,
    n2408,
    n2250,
    n2551
  );


  xor
  g2597
  (
    n2616,
    n2386,
    n2512,
    n2334,
    n2210
  );


  xor
  g2598
  (
    n2634,
    n2338,
    n2341,
    n2387,
    n2518
  );


  nand
  g2599
  (
    n2648,
    n2388,
    n2381,
    n2377,
    n2511
  );


  and
  g2600
  (
    n2670,
    n2408,
    n2530,
    n2542,
    n2360
  );


  nand
  g2601
  (
    n2683,
    n2288,
    n2343,
    n2518,
    n2233
  );


  xor
  g2602
  (
    n2813,
    n2548,
    n2327,
    n2336,
    n2291
  );


  nand
  g2603
  (
    n2786,
    n2298,
    n2554,
    n2566,
    n2341
  );


  nor
  g2604
  (
    n2613,
    n2266,
    n2561,
    n2278,
    n2212
  );


  xnor
  g2605
  (
    n2735,
    n2401,
    n2366,
    n2254,
    n2252
  );


  nor
  g2606
  (
    n2626,
    n2550,
    n2277,
    n2279,
    n2323
  );


  xnor
  g2607
  (
    n2591,
    n2345,
    n2340,
    n2400,
    n2298
  );


  and
  g2608
  (
    n2748,
    n2334,
    n2552,
    n2370,
    n2371
  );


  and
  g2609
  (
    n2569,
    n2397,
    n2289,
    n2240,
    n2320
  );


  or
  g2610
  (
    n2625,
    n2296,
    n2353,
    n2349,
    n2505
  );


  nand
  g2611
  (
    n2713,
    n2550,
    n2269,
    n2408,
    n2293
  );


  or
  g2612
  (
    n2581,
    n2536,
    n2266,
    n2333,
    n2273
  );


  or
  g2613
  (
    n2568,
    n2517,
    n2386,
    n2519,
    n2516
  );


  xnor
  g2614
  (
    n2803,
    n2364,
    n2524,
    n2552,
    n2543
  );


  or
  g2615
  (
    n2742,
    n2301,
    n2382,
    n2402,
    n2248
  );


  nand
  g2616
  (
    n2624,
    n2269,
    n2386,
    n2247,
    n2513
  );


  or
  g2617
  (
    n2689,
    n2312,
    n2375,
    n2350,
    n2356
  );


  nand
  g2618
  (
    n2816,
    n2347,
    n2204,
    n2194,
    n2503
  );


  xnor
  g2619
  (
    n2728,
    n2368,
    n2411,
    n2336,
    n2420
  );


  nor
  g2620
  (
    n2698,
    n2271,
    n2263,
    n2538,
    n2540
  );


  xnor
  g2621
  (
    n2654,
    n2293,
    n2255,
    n2554,
    n2307
  );


  or
  g2622
  (
    n2661,
    n2300,
    n2536,
    n2540,
    n2415
  );


  xor
  g2623
  (
    n2791,
    n2553,
    n2225,
    n2267,
    n2369
  );


  xnor
  g2624
  (
    n2702,
    n2297,
    n2563,
    n2392,
    n2205
  );


  xnor
  g2625
  (
    n2718,
    n2537,
    n2373,
    n2521,
    n2262
  );


  nor
  g2626
  (
    n2774,
    n2317,
    n2332,
    n2545,
    n2517
  );


  nor
  g2627
  (
    n2723,
    n2525,
    n2525,
    n2420,
    n2193
  );


  nor
  g2628
  (
    n2789,
    n2313,
    n2274,
    n2250,
    n2268
  );


  nor
  g2629
  (
    n2611,
    n2416,
    n2534,
    n2341,
    n2544
  );


  nand
  g2630
  (
    n2710,
    n2503,
    n2256,
    n2275,
    n2242
  );


  xor
  g2631
  (
    n2787,
    n2414,
    n2563,
    n2422,
    n2318
  );


  or
  g2632
  (
    n2704,
    n2270,
    n2380,
    n2504,
    n2330
  );


  nand
  g2633
  (
    n2641,
    n2546,
    n2084,
    n2545,
    n2344
  );


  nand
  g2634
  (
    n2779,
    n2521,
    n2555,
    n2557,
    n2537
  );


  xnor
  g2635
  (
    n2603,
    n2423,
    n2256,
    n2357,
    n2324
  );


  xnor
  g2636
  (
    n2597,
    n2197,
    n2359,
    n2261,
    n2274
  );


  xnor
  g2637
  (
    n2666,
    n2392,
    n2411,
    n2563,
    n2404
  );


  and
  g2638
  (
    n2655,
    n2535,
    n2373,
    n2267,
    n2376
  );


  xnor
  g2639
  (
    n2753,
    n2379,
    n2515,
    n2539,
    n2203
  );


  or
  g2640
  (
    n2749,
    n2422,
    n2413,
    n2276,
    n2400
  );


  nand
  g2641
  (
    n2653,
    n2334,
    n2361,
    n2389,
    n2300
  );


  or
  g2642
  (
    n2762,
    n2520,
    n2375,
    n2344,
    n2552
  );


  xnor
  g2643
  (
    n2808,
    n2508,
    n2332,
    n2252,
    n2327
  );


  nand
  g2644
  (
    n2590,
    n2329,
    n2315,
    n2423,
    n2358
  );


  xor
  g2645
  (
    n2726,
    n2330,
    n2328,
    n2297,
    n2311
  );


  and
  g2646
  (
    n2658,
    n2342,
    n2306,
    n2264,
    n2387
  );


  nand
  g2647
  (
    n2739,
    n2284,
    n2292,
    n2538,
    n2323
  );


  xnor
  g2648
  (
    n2582,
    n2557,
    n2280,
    n2314,
    n2306
  );


  nor
  g2649
  (
    n2637,
    n2330,
    n2269,
    n2543,
    n2524
  );


  and
  g2650
  (
    n2812,
    n2523,
    n2369,
    n2299,
    n2541
  );


  or
  g2651
  (
    n2583,
    n2259,
    n2386,
    n2417,
    n2378
  );


  and
  g2652
  (
    n2815,
    n2413,
    n2387,
    n2349,
    n2318
  );


  xnor
  g2653
  (
    n2707,
    n2520,
    n2405,
    n2257,
    n2409
  );


  or
  g2654
  (
    n2671,
    n2279,
    n2398,
    n2366,
    n2354
  );


  or
  g2655
  (
    n2716,
    n2509,
    n2379,
    n2284,
    n2253
  );


  or
  g2656
  (
    n2630,
    n2389,
    n2549,
    n2403,
    n2284
  );


  nor
  g2657
  (
    n2681,
    n2372,
    n2391,
    n2358,
    n2280
  );


  nor
  g2658
  (
    n2811,
    n2327,
    n2282,
    n2317,
    n2370
  );


  and
  g2659
  (
    n2604,
    n2511,
    n2265,
    n2270,
    n2349
  );


  nor
  g2660
  (
    n2766,
    n2406,
    n2353,
    n2268,
    n2380
  );


  nand
  g2661
  (
    n2644,
    n2553,
    n2549,
    n2357,
    n2363
  );


  and
  g2662
  (
    n2795,
    n2299,
    n2381,
    n2248,
    n2315
  );


  nand
  g2663
  (
    n2732,
    n2217,
    n2514,
    n2557,
    n2351
  );


  xnor
  g2664
  (
    n2737,
    n2399,
    n2370,
    n2556,
    n2407
  );


  nand
  g2665
  (
    n2731,
    n2324,
    n2358,
    n2306,
    n2251
  );


  and
  g2666
  (
    n2793,
    n2368,
    n2410,
    n2394,
    n2248
  );


  xor
  g2667
  (
    n2687,
    n2412,
    n2517,
    n2393,
    n2280
  );


  nor
  g2668
  (
    n2650,
    n2282,
    n2361,
    n2555,
    n2335
  );


  xnor
  g2669
  (
    n2776,
    n2405,
    n2368,
    n2385,
    n2319
  );


  nor
  g2670
  (
    n2579,
    n2322,
    n2191,
    n2370,
    n2367
  );


  nand
  g2671
  (
    n2711,
    n2558,
    n2271,
    n2325,
    n2234
  );


  xnor
  g2672
  (
    n2679,
    n2332,
    n2329,
    n2369,
    n2198
  );


  and
  g2673
  (
    n2700,
    n2333,
    n2378,
    n2419,
    n2376
  );


  xor
  g2674
  (
    n2612,
    n2226,
    n2270,
    n2539,
    n2342
  );


  xor
  g2675
  (
    n2788,
    n2392,
    n2551,
    n2351,
    n2534
  );


  nor
  g2676
  (
    n2660,
    n2235,
    n2516,
    n2336,
    n2273
  );


  nor
  g2677
  (
    n2598,
    n2408,
    n2423,
    n2549,
    n2555
  );


  nor
  g2678
  (
    n2730,
    n2211,
    n2527,
    n2532,
    n2529
  );


  nor
  g2679
  (
    n2807,
    n2363,
    n2508,
    n2557,
    n2506
  );


  xor
  g2680
  (
    n2782,
    n2365,
    n2285,
    n2271,
    n2320
  );


  xnor
  g2681
  (
    n2697,
    n2283,
    n2347,
    n2355,
    n2549
  );


  nor
  g2682
  (
    n2821,
    n2532,
    n2510,
    n2323,
    n2565
  );


  and
  g2683
  (
    n2763,
    n2565,
    n2414,
    n2533,
    n2337
  );


  and
  g2684
  (
    n2745,
    n2565,
    n2290,
    n2394,
    n2347
  );


  or
  g2685
  (
    n2743,
    n2283,
    n2353,
    n2562,
    n2346
  );


  nand
  g2686
  (
    n2676,
    n2201,
    n2546,
    n2326,
    n2276
  );


  and
  g2687
  (
    n2619,
    n2373,
    n2561,
    n2564,
    n2542
  );


  nor
  g2688
  (
    n2574,
    n2507,
    n2417,
    n2403,
    n2296
  );


  nor
  g2689
  (
    n2797,
    n2506,
    n2396,
    n2361,
    n2528
  );


  or
  g2690
  (
    n2622,
    n2258,
    n2547,
    n2415,
    n2252
  );


  xor
  g2691
  (
    n2722,
    n2538,
    n2420,
    n2272,
    n2515
  );


  xnor
  g2692
  (
    n2659,
    n2406,
    n2404,
    n2302,
    n2508
  );


  nor
  g2693
  (
    n2692,
    n2348,
    n2561,
    n2258,
    n2539
  );


  nand
  g2694
  (
    n2596,
    n2298,
    n2231,
    n2340,
    n2314
  );


  and
  g2695
  (
    n2798,
    n2286,
    n2529,
    n2249,
    n2352
  );


  and
  g2696
  (
    n2703,
    n2565,
    n2281,
    n2393,
    n2396
  );


  nand
  g2697
  (
    n2586,
    n2551,
    n2422,
    n2310,
    n2249
  );


  and
  g2698
  (
    n2810,
    n2258,
    n2412,
    n2379,
    n2389
  );


  and
  g2699
  (
    n2799,
    n2566,
    n2519,
    n2315,
    n2254
  );


  or
  g2700
  (
    n2809,
    n2410,
    n2505,
    n2366,
    n2416
  );


  and
  g2701
  (
    n2667,
    n2308,
    n2312,
    n2286,
    n2313
  );


  xor
  g2702
  (
    n2769,
    n2541,
    n2272,
    n2384,
    n2385
  );


  xor
  g2703
  (
    n2738,
    n2522,
    n2511,
    n2292,
    n2419
  );


  nor
  g2704
  (
    n2664,
    n2296,
    n2308,
    n2291,
    n2526
  );


  nand
  g2705
  (
    n2736,
    n2257,
    n2402,
    n2371,
    n2397
  );


  or
  g2706
  (
    n2725,
    n2377,
    n2378,
    n2285,
    n2555
  );


  xnor
  g2707
  (
    n2756,
    n2255,
    n2310,
    n2206,
    n2559
  );


  xnor
  g2708
  (
    n2588,
    n2320,
    n2324,
    n2301,
    n2259
  );


  nor
  g2709
  (
    n2759,
    n2514,
    n2401,
    n2333,
    n2284
  );


  and
  g2710
  (
    n2792,
    n2558,
    n2399,
    n2381,
    n2299
  );


  xor
  g2711
  (
    n2593,
    n2251,
    n2280,
    n2325,
    n2260
  );


  nor
  g2712
  (
    n2775,
    n2507,
    n2542,
    n2354,
    n2352
  );


  or
  g2713
  (
    n2771,
    n2398,
    n2383,
    n2418,
    n2545
  );


  xnor
  g2714
  (
    n2682,
    n2510,
    n2329,
    n2303,
    n2263
  );


  xor
  g2715
  (
    n2690,
    n2412,
    n2395,
    n2228,
    n2321
  );


  xnor
  g2716
  (
    n2721,
    n2531,
    n2267,
    n2539,
    n2320
  );


  and
  g2717
  (
    n2796,
    n2275,
    n2333,
    n2372,
    n2504
  );


  nand
  g2718
  (
    n2573,
    n2546,
    n2527,
    n2394,
    n2525
  );


  nand
  g2719
  (
    n2610,
    n2232,
    n2540,
    n2382,
    n2293
  );


  xnor
  g2720
  (
    n2607,
    n2397,
    n2560,
    n2302,
    n2346
  );


  or
  g2721
  (
    n2605,
    n2526,
    n2265,
    n2282,
    n2375
  );


  or
  g2722
  (
    n2645,
    n2299,
    n2306,
    n2515,
    n2214
  );


  xnor
  g2723
  (
    n2701,
    n2383,
    n2362,
    n2351,
    n2414
  );


  nor
  g2724
  (
    n2647,
    n2528,
    n2260,
    n2188,
    n2338
  );


  xor
  g2725
  (
    n2665,
    n2395,
    n2305,
    n2273,
    n2215
  );


  xnor
  g2726
  (
    n2672,
    n2273,
    n2208,
    n2366,
    n2544
  );


  nand
  g2727
  (
    n2636,
    n2289,
    n2388,
    n2374,
    n2559
  );


  xor
  g2728
  (
    n2584,
    n2527,
    n2288,
    n2531,
    n2411
  );


  xor
  g2729
  (
    n2615,
    n2305,
    n2537,
    n2377,
    n2395
  );


  nand
  g2730
  (
    n2585,
    n2311,
    n2523,
    n2543,
    n2302
  );


  xnor
  g2731
  (
    n2773,
    n2530,
    n2236,
    n2513,
    n2406
  );


  nor
  g2732
  (
    n2608,
    n2289,
    n2512,
    n2264,
    n2256
  );


  and
  g2733
  (
    n2601,
    n2308,
    n2312,
    n2381,
    n2290
  );


  xor
  g2734
  (
    n2777,
    n2375,
    n2274,
    n2309,
    n2349
  );


  or
  g2735
  (
    n2638,
    n2417,
    n2326,
    n2339,
    n2257
  );


  or
  g2736
  (
    n2595,
    n2243,
    n2562,
    n2309,
    n2401
  );


  and
  g2737
  (
    n2814,
    n2510,
    n2335,
    n2342,
    n2384
  );


  xor
  g2738
  (
    n2705,
    n2531,
    n2391,
    n2367,
    n2278
  );


  and
  g2739
  (
    n2643,
    n2223,
    n2516,
    n2360,
    n2362
  );


  nor
  g2740
  (
    n2800,
    n2417,
    n2371,
    n2262,
    n2527
  );


  and
  g2741
  (
    n2794,
    n2345,
    n2337,
    n2564,
    n2534
  );


  and
  g2742
  (
    n2817,
    n2301,
    n2395,
    n2339,
    n2533
  );


  nor
  g2743
  (
    n2819,
    n2513,
    n2503,
    n2247,
    n2396
  );


  nand
  g2744
  (
    n2686,
    n2295,
    n2285,
    n2393,
    n2261
  );


  or
  g2745
  (
    KeyWire_0_3,
    n2295,
    n2515,
    n2304,
    n2540
  );


  and
  g2746
  (
    n2578,
    n2541,
    n2413,
    n2519,
    n2237
  );


  or
  g2747
  (
    n2678,
    n2317,
    n2525,
    n2554,
    n2422
  );


  or
  g2748
  (
    n2717,
    n2343,
    n2324,
    n2544,
    n2250
  );


  nand
  g2749
  (
    n2755,
    n2239,
    n2562,
    n2310,
    n2510
  );


  xnor
  g2750
  (
    n2685,
    n2406,
    n2383,
    n2403,
    n2384
  );


  and
  g2751
  (
    n2617,
    n2335,
    n2509,
    n2271,
    n2389
  );


  nand
  g2752
  (
    n2602,
    n2410,
    n2548,
    n2388,
    n2287
  );


  xor
  g2753
  (
    n2580,
    n2412,
    n2559,
    n2400,
    n2317
  );


  nand
  g2754
  (
    n2674,
    n2302,
    n2536,
    n2350,
    n2409
  );


  nor
  g2755
  (
    n2594,
    n2264,
    n2261,
    n2356,
    n2230
  );


  xor
  g2756
  (
    n2635,
    n2396,
    n2346,
    n2312,
    n2528
  );


  and
  g2757
  (
    n2669,
    n2247,
    n2550,
    n2504,
    n2506
  );


  nor
  g2758
  (
    n2620,
    n2376,
    n2561,
    n2355,
    n2275
  );


  xor
  g2759
  (
    n2727,
    n2265,
    n2354,
    n2509,
    n2521
  );


  or
  g2760
  (
    n2621,
    n2307,
    n2520,
    n2361,
    n2200
  );


  and
  g2761
  (
    n2712,
    n2262,
    n2281,
    n2350
  );


  or
  g2762
  (
    n2770,
    n2530,
    n2407,
    n2379,
    n2202
  );


  xnor
  g2763
  (
    n2719,
    n2316,
    n2219,
    n2348,
    n2291
  );


  xnor
  g2764
  (
    n2733,
    n2374,
    n2526,
    n2564,
    n2344
  );


  xnor
  g2765
  (
    n2802,
    n2227,
    n2294,
    n2304,
    n2558
  );


  xnor
  g2766
  (
    n2699,
    n2394,
    n2355,
    n2286,
    n2511
  );


  nand
  g2767
  (
    n2695,
    n2257,
    n2401,
    n2407,
    n2529
  );


  and
  g2768
  (
    n2662,
    n2360,
    n2367,
    n2323,
    n2336
  );


  xor
  g2769
  (
    n2657,
    n2327,
    n2264,
    n2364,
    n2305
  );


  nor
  g2770
  (
    n2668,
    n2380,
    n2274,
    n2343,
    n2321
  );


  nand
  g2771
  (
    n2606,
    n2504,
    n2393,
    n2277,
    n2392
  );


  or
  g2772
  (
    KeyWire_0_10,
    n2560,
    n2356,
    n2359,
    n2554
  );


  nand
  g2773
  (
    n2790,
    n2316,
    n2300,
    n2301,
    n2304
  );


  and
  g2774
  (
    n2694,
    n2548,
    n2345,
    n2278,
    n2254
  );


  and
  g2775
  (
    n2818,
    n2532,
    n2322,
    n2276,
    n2535
  );


  and
  g2776
  (
    n2575,
    n2260,
    n2313,
    n2340,
    n2341
  );


  and
  g2777
  (
    n2675,
    n2253,
    n2546,
    n2391,
    n2339
  );


  and
  g2778
  (
    n2684,
    n2390,
    n2218,
    n2518,
    n2411
  );


  xor
  g2779
  (
    n2709,
    n2255,
    n2277,
    n2348,
    n2391
  );


  xor
  g2780
  (
    n2696,
    n2334,
    n2522,
    n2505,
    n2328
  );


  nor
  g2781
  (
    n2629,
    n2399,
    n2374,
    n2506,
    n2314
  );


  nand
  g2782
  (
    n2720,
    n2288,
    n2213,
    n2538,
    n2330
  );


  xnor
  g2783
  (
    n2663,
    n2287,
    n2238,
    n2350,
    n2332
  );


  nand
  g2784
  (
    n2752,
    n2265,
    n2356,
    n2351,
    n2268
  );


  xor
  g2785
  (
    n2639,
    n2533,
    n2315,
    n2531,
    n2241
  );


  and
  g2786
  (
    n2609,
    n2224,
    n2385,
    n2326,
    n2354
  );


  or
  g2787
  (
    n2820,
    n2421,
    n2397,
    n2405,
    n2513
  );


  nor
  g2788
  (
    n2693,
    n2560,
    n2338,
    n2244,
    n2517
  );


  xor
  g2789
  (
    n2633,
    n2363,
    n2409,
    n2353,
    n2343
  );


  or
  g2790
  (
    n2891,
    n2816,
    n2741,
    n2739,
    n2787
  );


  and
  g2791
  (
    n2953,
    n2758,
    n2730,
    n2763,
    n2720
  );


  xnor
  g2792
  (
    n2961,
    n2719,
    n2786,
    n2766,
    n2817
  );


  nor
  g2793
  (
    n2949,
    n2812,
    n2587,
    n2722,
    n2575
  );


  and
  g2794
  (
    n2852,
    n2739,
    n2816,
    n2737,
    n2700
  );


  or
  g2795
  (
    n2941,
    n2771,
    n2821,
    n2805,
    n2698
  );


  nor
  g2796
  (
    n2877,
    n2793,
    n2819,
    n2800,
    n2772
  );


  or
  g2797
  (
    n2978,
    n2705,
    n2772,
    n2724,
    n2764
  );


  nor
  g2798
  (
    n2972,
    n2659,
    n2693,
    n2680,
    n2725
  );


  xnor
  g2799
  (
    n2955,
    n2819,
    n2799,
    n2644,
    n2765
  );


  nor
  g2800
  (
    n2944,
    n2722,
    n2589,
    n2707,
    n2746
  );


  xnor
  g2801
  (
    n2836,
    n2802,
    n2740,
    n2818,
    n2670
  );


  nand
  g2802
  (
    n2837,
    n2816,
    n2704,
    n2602,
    n2755
  );


  nor
  g2803
  (
    n2937,
    n2797,
    n2786,
    n2764,
    n2780
  );


  nand
  g2804
  (
    n2959,
    n2697,
    n2782,
    n2637,
    n2752
  );


  xor
  g2805
  (
    n2911,
    n2716,
    n2677,
    n2625,
    n2729
  );


  xnor
  g2806
  (
    n2971,
    n2683,
    n2751,
    n2817,
    n2768
  );


  and
  g2807
  (
    n2881,
    n2818,
    n2747,
    n2740,
    n2791
  );


  nor
  g2808
  (
    n2948,
    n2819,
    n2591,
    n2743,
    n2717
  );


  nand
  g2809
  (
    n2981,
    n2657,
    n2774,
    n2700,
    n2803
  );


  nor
  g2810
  (
    n2843,
    n2692,
    n2777,
    n2733
  );


  xnor
  g2811
  (
    n2918,
    n2746,
    n2691,
    n2596,
    n2753
  );


  xor
  g2812
  (
    n2938,
    n2623,
    n2777,
    n2728,
    n2719
  );


  and
  g2813
  (
    n2897,
    n2643,
    n2821,
    n2749,
    n2763
  );


  nor
  g2814
  (
    n2925,
    n2782,
    n2737,
    n2792,
    n2761
  );


  xnor
  g2815
  (
    n2892,
    n2701,
    n2756,
    n2821,
    n2700
  );


  xnor
  g2816
  (
    n2970,
    n2799,
    n2716,
    n2717,
    n2808
  );


  or
  g2817
  (
    n2863,
    n2748,
    n2752,
    n2698,
    n2778
  );


  nor
  g2818
  (
    n2858,
    n2620,
    n2813,
    n2086
  );


  and
  g2819
  (
    n2825,
    n2085,
    n2674,
    n2702,
    n2804
  );


  and
  g2820
  (
    n2969,
    n2715,
    n2773,
    n2686,
    n2783
  );


  nand
  g2821
  (
    n2962,
    n2796,
    n2604,
    n2736,
    n2751
  );


  nor
  g2822
  (
    n2872,
    n2802,
    n2720,
    n2715,
    n2726
  );


  xnor
  g2823
  (
    n2915,
    n2603,
    n2750,
    n2761,
    n2713
  );


  or
  g2824
  (
    n2976,
    n2724,
    n2810,
    n2756,
    n2798
  );


  or
  g2825
  (
    n2920,
    n2694,
    n2738,
    n2760,
    n2687
  );


  xnor
  g2826
  (
    n2869,
    n2728,
    n2785,
    n2822,
    n2739
  );


  nor
  g2827
  (
    n2980,
    n2569,
    n2630,
    n2758,
    n2788
  );


  nand
  g2828
  (
    n2875,
    n2729,
    n2820,
    n2786,
    n2760
  );


  xor
  g2829
  (
    n2874,
    n2802,
    n2584,
    n2727,
    n2632
  );


  nand
  g2830
  (
    n2845,
    n2730,
    n2792,
    n2704,
    n2804
  );


  and
  g2831
  (
    n2979,
    n2627,
    n2780,
    n2806
  );


  nor
  g2832
  (
    n2841,
    n2735,
    n2718,
    n2628,
    n2792
  );


  nor
  g2833
  (
    n2934,
    n2808,
    n2621,
    n2655,
    n2578
  );


  or
  g2834
  (
    n2857,
    n2776,
    n2735,
    n2751,
    n2794
  );


  or
  g2835
  (
    n2943,
    n2704,
    n2732,
    n2756,
    n2727
  );


  nand
  g2836
  (
    n2859,
    n2800,
    n2771,
    n2709,
    n2725
  );


  nor
  g2837
  (
    n2936,
    n2700,
    n2706,
    n2759,
    n2774
  );


  or
  g2838
  (
    n2888,
    n2811,
    n2799,
    n2749,
    n2791
  );


  or
  g2839
  (
    n2975,
    n2711,
    n2711,
    n2619,
    n2769
  );


  nor
  g2840
  (
    n2939,
    n2695,
    n2717,
    n2705,
    n2698
  );


  xnor
  g2841
  (
    n2870,
    n2615,
    n2754,
    n2714,
    n2789
  );


  nand
  g2842
  (
    n2902,
    n2705,
    n2585,
    n2576,
    n2778
  );


  nand
  g2843
  (
    n2904,
    n2696,
    n2087,
    n2765,
    n2667
  );


  and
  g2844
  (
    n2833,
    n2732,
    n2581,
    n2629,
    n2766
  );


  xnor
  g2845
  (
    n2896,
    n2790,
    n2679,
    n2593,
    n2793
  );


  xor
  g2846
  (
    n2831,
    n2776,
    n2795,
    n2577,
    n2809
  );


  xor
  g2847
  (
    n2930,
    n2765,
    n2728,
    n2791,
    n2815
  );


  xor
  g2848
  (
    n2847,
    n2811,
    n2734,
    n2820
  );


  xnor
  g2849
  (
    n2899,
    n2731,
    n2741,
    n2706,
    n2808
  );


  and
  g2850
  (
    n2974,
    n2740,
    n2760,
    n2642,
    n2658
  );


  and
  g2851
  (
    n2910,
    n2744,
    n2711,
    n2725,
    n2583
  );


  or
  g2852
  (
    n2883,
    n2743,
    n2725,
    n2811,
    n2737
  );


  xnor
  g2853
  (
    n2885,
    n2650,
    n2769,
    n2754,
    n2802
  );


  xor
  g2854
  (
    n2827,
    n2704,
    n2586,
    n2814,
    n2816
  );


  nand
  g2855
  (
    n2823,
    n2684,
    n2744,
    n2821,
    n2612
  );


  nand
  g2856
  (
    n2924,
    n2708,
    n2662,
    n2747,
    n2803
  );


  nand
  g2857
  (
    n2846,
    n2810,
    n2721,
    n2712,
    n2710
  );


  nand
  g2858
  (
    n2878,
    n2672,
    n2712,
    n2779,
    n2814
  );


  or
  g2859
  (
    n2940,
    n2742,
    n2707,
    n2571,
    n2720
  );


  and
  g2860
  (
    n2916,
    n2710,
    n2703,
    n2773,
    n2803
  );


  or
  g2861
  (
    n2855,
    n2781,
    n2804,
    n2639,
    n2649
  );


  xor
  g2862
  (
    n2965,
    n2714,
    n2708,
    n2709,
    n2622
  );


  or
  g2863
  (
    n2849,
    n2598,
    n2771,
    n2774,
    n2708
  );


  nand
  g2864
  (
    n2942,
    n2818,
    n2788,
    n2624,
    n2763
  );


  nand
  g2865
  (
    n2868,
    n2732,
    n2782,
    n2708,
    n2772
  );


  xnor
  g2866
  (
    n2861,
    n2759,
    n2758,
    n2801,
    n2812
  );


  xor
  g2867
  (
    n2906,
    n2789,
    n2716,
    n2742,
    n2780
  );


  xor
  g2868
  (
    n2945,
    n2656,
    n2817,
    n2797,
    n2784
  );


  or
  g2869
  (
    n2935,
    n2722,
    n2815,
    n2791,
    n2790
  );


  nand
  g2870
  (
    n2917,
    n2608,
    n2736,
    n2702,
    n2734
  );


  nor
  g2871
  (
    n2828,
    n2748,
    n2779,
    n2718,
    n2727
  );


  xor
  g2872
  (
    n2856,
    n2770,
    n2744,
    n2782,
    n2767
  );


  xor
  g2873
  (
    n2829,
    n2799,
    n2777,
    n2707,
    n2616
  );


  and
  g2874
  (
    n2826,
    n2567,
    n2648,
    n2681,
    n2790
  );


  nor
  g2875
  (
    n2882,
    n2800,
    n2749,
    n2626,
    n2712
  );


  and
  g2876
  (
    n2864,
    n2701,
    n2723,
    n2706,
    n2768
  );


  xor
  g2877
  (
    n2956,
    n2638,
    n2776,
    n2617,
    n2770
  );


  nand
  g2878
  (
    n2914,
    n2783,
    n2798,
    n2580,
    n2745
  );


  and
  g2879
  (
    n2851,
    n2688,
    n2689,
    n2822,
    n2713
  );


  nor
  g2880
  (
    n2867,
    n2812,
    n2723,
    n2794,
    n2590
  );


  nand
  g2881
  (
    n2893,
    n2705,
    n2814,
    n2721,
    n2573
  );


  nor
  g2882
  (
    n2963,
    n2699,
    n2737,
    n2806,
    n2805
  );


  xnor
  g2883
  (
    n2931,
    n2781,
    n2574,
    n2794,
    n2815
  );


  xnor
  g2884
  (
    n2900,
    n2698,
    n2599,
    n2719,
    n2767
  );


  and
  g2885
  (
    n2968,
    n2720,
    n2661,
    n2728,
    n2718
  );


  or
  g2886
  (
    n2926,
    n2775,
    n2607,
    n2745,
    n2810
  );


  and
  g2887
  (
    n2865,
    n2763,
    n2772,
    n2822,
    n2755
  );


  xnor
  g2888
  (
    n2905,
    n2717,
    n2797,
    n2775,
    n2807
  );


  or
  g2889
  (
    n2922,
    n2769,
    n2818,
    n2775,
    n2614
  );


  xnor
  g2890
  (
    n2838,
    n2699,
    n2778,
    n2606,
    n2785
  );


  nor
  g2891
  (
    n2947,
    n2779,
    n2757,
    n2748,
    n2770
  );


  nor
  g2892
  (
    n2973,
    n2641,
    n2768,
    n2813,
    n2702
  );


  nand
  g2893
  (
    n2886,
    n2426,
    n2746,
    n2817,
    n2762
  );


  nor
  g2894
  (
    n2932,
    n2745,
    n2634,
    n2812,
    n2595
  );


  xor
  g2895
  (
    n2933,
    n2715,
    n2809,
    n2652,
    n2709
  );


  nand
  g2896
  (
    n2832,
    n2605,
    n2676,
    n2811,
    n2767
  );


  nor
  g2897
  (
    n2890,
    n2752,
    n2631,
    n2663,
    n2803
  );


  xor
  g2898
  (
    n2840,
    n2762,
    n2743,
    n2819,
    n2707
  );


  xor
  g2899
  (
    n2927,
    n2796,
    n2601,
    n2757,
    n2815
  );


  and
  g2900
  (
    n2950,
    n2789,
    n2609,
    n2735,
    n2703
  );


  nand
  g2901
  (
    n2895,
    n2701,
    n2572,
    n2726,
    n2801
  );


  nand
  g2902
  (
    n2880,
    n2759,
    n2758,
    n2731,
    n2699
  );


  nor
  g2903
  (
    n2887,
    n2800,
    n2734,
    n2729,
    n2653
  );


  and
  g2904
  (
    n2866,
    n2568,
    n2730,
    n2701,
    n2723
  );


  xnor
  g2905
  (
    n2928,
    n2747,
    n2796,
    n2804
  );


  nor
  g2906
  (
    n2889,
    n2807,
    n2775,
    n2784,
    n2735
  );


  and
  g2907
  (
    n2830,
    n2703,
    n2740,
    n2731,
    n2773
  );


  and
  g2908
  (
    n2860,
    n2747,
    n2646,
    n2786,
    n2766
  );


  xnor
  g2909
  (
    n2958,
    n2732,
    n2750,
    n2781,
    n2741
  );


  nor
  g2910
  (
    n2921,
    n2748,
    n2801,
    n2795,
    n2813
  );


  and
  g2911
  (
    n2967,
    n2734,
    n2754,
    n2733,
    n2738
  );


  and
  g2912
  (
    n2908,
    n2668,
    n2635,
    n2673,
    n2594
  );


  xnor
  g2913
  (
    n2884,
    n2742,
    n2778,
    n2753,
    n2733
  );


  and
  g2914
  (
    n2903,
    n2753,
    n2754,
    n2794,
    n2759
  );


  xor
  g2915
  (
    n2850,
    n2771,
    n2715,
    n2783,
    n2807
  );


  and
  g2916
  (
    n2977,
    n2675,
    n2738,
    n2810,
    n2709
  );


  and
  g2917
  (
    n2907,
    n2760,
    n2750,
    n2749,
    n2755
  );


  nor
  g2918
  (
    n2901,
    n2736,
    n2741,
    n2721,
    n2762
  );


  xnor
  g2919
  (
    n2929,
    n2739,
    n2806,
    n2793,
    n2768
  );


  xor
  g2920
  (
    n2960,
    n2722,
    n2579,
    n2710,
    n2785
  );


  xor
  g2921
  (
    n2898,
    n2787,
    n2761,
    n2597,
    n2766
  );


  or
  g2922
  (
    n2871,
    n2678,
    n2682,
    n2787,
    n2784
  );


  nand
  g2923
  (
    n2923,
    n672,
    n2795,
    n2690,
    n2785
  );


  xnor
  g2924
  (
    n2913,
    n2762,
    n2666,
    n2792,
    n2729
  );


  xor
  g2925
  (
    n2954,
    n2779,
    n2767,
    n2809,
    n2703
  );


  xor
  g2926
  (
    n2835,
    n2745,
    n2770,
    n2633,
    n2651
  );


  nand
  g2927
  (
    n2854,
    n2795,
    n2781,
    n2724,
    n2756
  );


  nor
  g2928
  (
    n2879,
    n2660,
    n2764,
    n2726,
    n2807
  );


  xor
  g2929
  (
    n2853,
    n2774,
    n2723,
    n2610,
    n2805
  );


  and
  g2930
  (
    n2842,
    n2710,
    n2699,
    n2798,
    n2712
  );


  and
  g2931
  (
    n2964,
    n2714,
    n2730,
    n2713,
    n2647
  );


  and
  g2932
  (
    n2862,
    n2592,
    n2820,
    n2743,
    n2724
  );


  nand
  g2933
  (
    n2873,
    n2769,
    n2731,
    n2822,
    n2714
  );


  nor
  g2934
  (
    n2946,
    n2685,
    n2613,
    n2738,
    n2761
  );


  or
  g2935
  (
    n2951,
    n2640,
    n2789,
    n2797,
    n2706
  );


  and
  g2936
  (
    KeyWire_0_4,
    n2793,
    n2654,
    n2726,
    n2588
  );


  and
  g2937
  (
    n2912,
    n2752,
    n2801,
    n2721,
    n2582
  );


  and
  g2938
  (
    n2966,
    n2755,
    n2611,
    n2718,
    n2808
  );


  nand
  g2939
  (
    n2844,
    n2798,
    n2773,
    n2750,
    n2713
  );


  or
  g2940
  (
    n2848,
    n2805,
    n2716,
    n2744,
    n2757
  );


  nand
  g2941
  (
    n2952,
    n2790,
    n2719,
    n2664,
    n2776
  );


  or
  g2942
  (
    n2919,
    n2736,
    n2814,
    n2727,
    n2645
  );


  nor
  g2943
  (
    n2834,
    n2753,
    n2765,
    n2764,
    n2780
  );


  or
  g2944
  (
    n2876,
    n2733,
    n2751,
    n2636,
    n2600
  );


  xor
  g2945
  (
    n2894,
    n2671,
    n2784,
    n2711,
    n2787
  );


  nor
  g2946
  (
    n2824,
    n2742,
    n2783,
    n2570,
    n2757
  );


  or
  g2947
  (
    n2909,
    n2665,
    n2809,
    n2702,
    n2788
  );


  xor
  g2948
  (
    n2957,
    n2746,
    n2618,
    n2669,
    n2788
  );


  and
  g2949
  (
    n2987,
    n2838,
    n2909,
    n2830,
    n2861
  );


  and
  g2950
  (
    n3000,
    n2839,
    n2917,
    n2864,
    n2891
  );


  xor
  g2951
  (
    n2996,
    n2855,
    n2873,
    n2849,
    n2910
  );


  and
  g2952
  (
    n2997,
    n2831,
    n2859,
    n2869,
    n2874
  );


  or
  g2953
  (
    n3002,
    n2828,
    n2883,
    n2842,
    n2878
  );


  or
  g2954
  (
    n2984,
    n2846,
    n2890,
    n2852,
    n2867
  );


  and
  g2955
  (
    n2983,
    n2834,
    n2880,
    n2871,
    n2919
  );


  xnor
  g2956
  (
    n3007,
    n2882,
    n2857,
    n2835,
    n2901
  );


  or
  g2957
  (
    n2988,
    n2920,
    n2898,
    n2826,
    n2856
  );


  xor
  g2958
  (
    n2985,
    n2833,
    n2923,
    n2851,
    n2823
  );


  xnor
  g2959
  (
    n3006,
    n2912,
    n2914,
    n2860,
    n2848
  );


  xnor
  g2960
  (
    n3003,
    n2885,
    n2926,
    n2866,
    n2900
  );


  or
  g2961
  (
    n2982,
    n2875,
    n2922,
    n2870,
    n2824
  );


  nor
  g2962
  (
    n2992,
    n2925,
    n2887,
    n2894,
    n2841
  );


  xor
  g2963
  (
    n2991,
    n2908,
    n2840,
    n2876,
    n2899
  );


  and
  g2964
  (
    n3001,
    n2906,
    n2888,
    n2921,
    n2877
  );


  and
  g2965
  (
    n2995,
    n2863,
    n2902,
    n2913,
    n2896
  );


  xor
  g2966
  (
    n2986,
    n2832,
    n2916,
    n2911,
    n2907
  );


  or
  g2967
  (
    n3004,
    n2868,
    n2827,
    n2903,
    n2904
  );


  xor
  g2968
  (
    n2999,
    n2879,
    n2884,
    n2886,
    n2844
  );


  nor
  g2969
  (
    n2990,
    n2915,
    n2845,
    n2847,
    n2897
  );


  nand
  g2970
  (
    n2989,
    n2865,
    n2836,
    n2854,
    n2858
  );


  xnor
  g2971
  (
    n2994,
    n2862,
    n2850,
    n2895,
    n2881
  );


  or
  g2972
  (
    KeyWire_0_9,
    n2905,
    n2825,
    n2837,
    n2924
  );


  and
  g2973
  (
    n2998,
    n2892,
    n2829,
    n2893,
    n2889
  );


  nand
  g2974
  (
    n2993,
    n2918,
    n2872,
    n2853,
    n2843
  );


  nor
  g2975
  (
    n3008,
    n2928,
    n2927,
    n3007,
    n2929
  );


  nand
  g2976
  (
    n3011,
    n2933,
    n3008,
    n1672
  );


  nor
  g2977
  (
    n3012,
    n3008,
    n2931,
    n1672,
    n1673
  );


  xor
  g2978
  (
    n3009,
    n1673,
    n2932,
    n1672
  );


  and
  g2979
  (
    n3010,
    n2930,
    n1673,
    n3008
  );


  or
  g2980
  (
    n3028,
    n2963,
    n2942,
    n3012,
    n3010
  );


  xor
  g2981
  (
    n3019,
    n3009,
    n2977,
    n2972,
    n2957
  );


  and
  g2982
  (
    n3026,
    n2969,
    n2939,
    n2950,
    n2949
  );


  xnor
  g2983
  (
    n3013,
    n2936,
    n2937,
    n2944,
    n2973
  );


  or
  g2984
  (
    n3014,
    n2974,
    n2961,
    n3011
  );


  xor
  g2985
  (
    n3027,
    n2964,
    n2971,
    n3010,
    n3012
  );


  or
  g2986
  (
    n3018,
    n2965,
    n2981,
    n2955,
    n2948
  );


  or
  g2987
  (
    n3023,
    n2952,
    n2968,
    n2954,
    n3009
  );


  nor
  g2988
  (
    n3015,
    n2980,
    n3011,
    n2959,
    n2970
  );


  nand
  g2989
  (
    n3021,
    n2946,
    n2934,
    n2958,
    n2941
  );


  and
  g2990
  (
    n3022,
    n2975,
    n2978,
    n2960,
    n2943
  );


  or
  g2991
  (
    n3017,
    n2966,
    n2979,
    n2935,
    n2953
  );


  xnor
  g2992
  (
    n3025,
    n2962,
    n3009,
    n3010,
    n3012
  );


  and
  g2993
  (
    n3020,
    n2951,
    n3012,
    n3010,
    n2956
  );


  xor
  g2994
  (
    n3016,
    n2938,
    n2967,
    n2947,
    n3009
  );


  and
  g2995
  (
    n3024,
    n3011,
    n2945,
    n2976,
    n2940
  );


  nand
  g2996
  (
    n3029,
    n3027,
    n3028,
    n3014,
    n3024
  );


  xnor
  g2997
  (
    n3031,
    n3022,
    n3020,
    n3023,
    n3025
  );


  nor
  g2998
  (
    n3032,
    n3013,
    n3017,
    n3021,
    n3026
  );


  or
  g2999
  (
    n3030,
    n3019,
    n3018,
    n3016,
    n3015
  );


  xor
  KeyGate_0_0
  (
    n1988,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n967,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n2242,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n2822,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n2839,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n833,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n2357,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1439,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n2215,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n3005,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n2801,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1730,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1290,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n261,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n196,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n1028,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1776,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n81,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n637,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n1225,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n652,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1775,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n535,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1929,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n2173,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1953,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n162,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n933,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n431,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1360,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n614,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1395,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


