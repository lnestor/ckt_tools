

module Stat_100_42
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n116,
  n115,
  n114,
  n107,
  n101,
  n125,
  n119,
  n103,
  n112,
  n111,
  n117,
  n129,
  n113,
  n126,
  n109,
  n110,
  n132,
  n120,
  n104,
  n102,
  n122,
  n131,
  n105,
  n128,
  n123,
  n108,
  n130,
  n124,
  n118,
  n121,
  n127,
  n106,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n116;output n115;output n114;output n107;output n101;output n125;output n119;output n103;output n112;output n111;output n117;output n129;output n113;output n126;output n109;output n110;output n132;output n120;output n104;output n102;output n122;output n131;output n105;output n128;output n123;output n108;output n130;output n124;output n118;output n121;output n127;output n106;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  not
  g0
  (
    n41,
    n8
  );


  buf
  g1
  (
    n38,
    n6
  );


  buf
  g2
  (
    n55,
    n2
  );


  not
  g3
  (
    n51,
    n11
  );


  not
  g4
  (
    n52,
    n9
  );


  buf
  g5
  (
    n56,
    n8
  );


  buf
  g6
  (
    n49,
    n9
  );


  not
  g7
  (
    n36,
    n10
  );


  buf
  g8
  (
    n42,
    n10
  );


  not
  g9
  (
    n37,
    n8
  );


  not
  g10
  (
    n60,
    n3
  );


  not
  g11
  (
    n50,
    n6
  );


  buf
  g12
  (
    n33,
    n7
  );


  buf
  g13
  (
    n58,
    n7
  );


  buf
  g14
  (
    n40,
    n10
  );


  buf
  g15
  (
    n48,
    n8
  );


  buf
  g16
  (
    n54,
    n9
  );


  buf
  g17
  (
    n46,
    n9
  );


  not
  g18
  (
    n34,
    n1
  );


  not
  g19
  (
    n59,
    n11
  );


  buf
  g20
  (
    n57,
    n7
  );


  buf
  g21
  (
    n45,
    n5
  );


  not
  g22
  (
    n39,
    n10
  );


  not
  g23
  (
    n47,
    n6
  );


  not
  g24
  (
    n35,
    n11
  );


  buf
  g25
  (
    n61,
    n4
  );


  not
  g26
  (
    n53,
    n6
  );


  not
  g27
  (
    n43,
    n7
  );


  not
  g28
  (
    n44,
    n11
  );


  buf
  g29
  (
    n68,
    n33
  );


  not
  g30
  (
    n66,
    n37
  );


  not
  g31
  (
    n69,
    n35
  );


  not
  g32
  (
    n67,
    n37
  );


  buf
  g33
  (
    n64,
    n37
  );


  not
  g34
  (
    n63,
    n36
  );


  not
  g35
  (
    n65,
    n37
  );


  not
  g36
  (
    n62,
    n34
  );


  nand
  g37
  (
    n79,
    n20,
    n29,
    n67,
    n17
  );


  or
  g38
  (
    n98,
    n21,
    n23,
    n69
  );


  and
  g39
  (
    n76,
    n30,
    n68,
    n25,
    n15
  );


  or
  g40
  (
    n87,
    n39,
    n65,
    n66,
    n14
  );


  or
  g41
  (
    n86,
    n38,
    n38,
    n23,
    n39
  );


  nor
  g42
  (
    n73,
    n68,
    n12,
    n21
  );


  xnor
  g43
  (
    n95,
    n19,
    n29,
    n28
  );


  nor
  g44
  (
    n94,
    n62,
    n25,
    n38,
    n16
  );


  and
  g45
  (
    n72,
    n26,
    n24,
    n68,
    n65
  );


  nor
  g46
  (
    n91,
    n63,
    n28,
    n40,
    n22
  );


  or
  g47
  (
    n77,
    n39,
    n30,
    n66,
    n15
  );


  nand
  g48
  (
    n96,
    n32,
    n64,
    n14,
    n63
  );


  nand
  g49
  (
    n83,
    n67,
    n62,
    n23,
    n69
  );


  nand
  g50
  (
    n70,
    n27,
    n67,
    n22
  );


  or
  g51
  (
    n97,
    n27,
    n31,
    n30,
    n17
  );


  or
  g52
  (
    n89,
    n28,
    n24,
    n12,
    n13
  );


  xnor
  g53
  (
    n82,
    n22,
    n14,
    n27,
    n68
  );


  and
  g54
  (
    n93,
    n16,
    n22,
    n31,
    n62
  );


  nor
  g55
  (
    n100,
    n64,
    n23,
    n13
  );


  nand
  g56
  (
    n88,
    n18,
    n63,
    n65
  );


  xor
  g57
  (
    n78,
    n40,
    n19,
    n64,
    n30
  );


  and
  g58
  (
    n75,
    n28,
    n40,
    n29,
    n26
  );


  and
  g59
  (
    n85,
    n19,
    n15,
    n17,
    n62
  );


  xnor
  g60
  (
    n84,
    n14,
    n19,
    n64,
    n27
  );


  or
  g61
  (
    n80,
    n66,
    n65,
    n24,
    n25
  );


  nand
  g62
  (
    n99,
    n18,
    n16,
    n31,
    n20
  );


  xnor
  g63
  (
    n74,
    n20,
    n26,
    n39,
    n21
  );


  xnor
  g64
  (
    n81,
    n25,
    n66,
    n16,
    n32
  );


  xnor
  g65
  (
    n92,
    n18,
    n38,
    n24,
    n15
  );


  xnor
  g66
  (
    n71,
    n18,
    n12,
    n13,
    n20
  );


  nor
  g67
  (
    n90,
    n21,
    n31,
    n26,
    n17
  );


  nand
  g68
  (
    n118,
    n95,
    n94,
    n57,
    n43
  );


  xnor
  g69
  (
    n126,
    n48,
    n61,
    n93,
    n59
  );


  xnor
  g70
  (
    n132,
    n47,
    n99,
    n100,
    n56
  );


  nand
  g71
  (
    n129,
    n54,
    n42,
    n71,
    n48
  );


  xnor
  g72
  (
    n110,
    n45,
    n47,
    n98,
    n44
  );


  xor
  g73
  (
    n109,
    n96,
    n85,
    n86,
    n88
  );


  and
  g74
  (
    n125,
    n55,
    n60,
    n80,
    n41
  );


  xnor
  g75
  (
    n127,
    n41,
    n44,
    n53,
    n90
  );


  nor
  g76
  (
    n114,
    n73,
    n60,
    n91,
    n54
  );


  and
  g77
  (
    n120,
    n81,
    n43,
    n48,
    n41
  );


  nand
  g78
  (
    n111,
    n99,
    n51,
    n74,
    n40
  );


  and
  g79
  (
    n113,
    n57,
    n82,
    n100,
    n41
  );


  xnor
  g80
  (
    AntiSAT_key_wire,
    n51,
    n46,
    n45,
    n56
  );


  nor
  g81
  (
    n105,
    n51,
    n99,
    n49
  );


  or
  g82
  (
    n121,
    n98,
    n54,
    n57,
    n60
  );


  nor
  g83
  (
    n103,
    n92,
    n58,
    n79,
    n76
  );


  xnor
  g84
  (
    n131,
    n54,
    n46,
    n59,
    n50
  );


  xnor
  g85
  (
    n106,
    n97,
    n56,
    n99,
    n58
  );


  nand
  g86
  (
    n116,
    n47,
    n53,
    n77,
    n46
  );


  xor
  g87
  (
    n115,
    n78,
    n44,
    n100,
    n98
  );


  and
  g88
  (
    n124,
    n98,
    n89,
    n43,
    n48
  );


  or
  g89
  (
    n104,
    n55,
    n50,
    n53,
    n61
  );


  xnor
  g90
  (
    n102,
    n42,
    n70,
    n50,
    n49
  );


  nand
  g91
  (
    n101,
    n45,
    n60,
    n59,
    n69
  );


  and
  g92
  (
    n107,
    n42,
    n44,
    n52,
    n58
  );


  xor
  g93
  (
    n122,
    n58,
    n32,
    n53,
    n59
  );


  xnor
  g94
  (
    n130,
    n83,
    n100,
    n61,
    n55
  );


  and
  g95
  (
    n123,
    n84,
    n45,
    n57,
    n51
  );


  xnor
  g96
  (
    n108,
    n87,
    n47,
    n42,
    n43
  );


  or
  g97
  (
    n117,
    n50,
    n46,
    n52,
    n61
  );


  nand
  g98
  (
    n119,
    n72,
    n49,
    n52
  );


  and
  g99
  (
    n112,
    n75,
    n55,
    n32,
    n56
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n128,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

