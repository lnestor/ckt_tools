// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_4000_363 written by SynthGen on 2021/04/05 11:24:27
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_4000_363 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1259, n1256, n1252, n1247, n1236, n1251, n1249, n1253,
 n1262, n1242, n1248, n1260, n1235, n1261, n1238, n1246,
 n1263, n1264, n1254, n1268, n1245, n1316, n1295, n1630,
 n1631, n1731, n1727, n1728, n1732, n1729, n1734, n4032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1259, n1256, n1252, n1247, n1236, n1251, n1249, n1253,
 n1262, n1242, n1248, n1260, n1235, n1261, n1238, n1246,
 n1263, n1264, n1254, n1268, n1245, n1316, n1295, n1630,
 n1631, n1731, n1727, n1728, n1732, n1729, n1734, n4032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1237, n1239, n1240, n1241, n1243, n1244,
 n1250, n1255, n1257, n1258, n1265, n1266, n1267, n1269,
 n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
 n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
 n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
 n1294, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
 n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
 n1311, n1312, n1313, n1314, n1315, n1317, n1318, n1319,
 n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
 n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
 n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
 n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
 n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
 n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
 n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
 n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
 n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
 n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
 n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
 n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
 n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
 n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
 n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
 n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
 n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
 n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
 n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
 n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
 n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
 n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
 n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
 n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
 n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
 n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
 n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
 n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
 n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
 n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
 n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
 n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
 n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
 n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
 n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
 n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
 n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
 n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
 n1624, n1625, n1626, n1627, n1628, n1629, n1632, n1633,
 n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
 n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
 n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
 n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
 n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
 n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
 n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
 n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
 n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
 n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
 n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
 n1722, n1723, n1724, n1725, n1726, n1730, n1733, n1735,
 n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
 n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
 n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
 n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
 n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
 n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
 n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
 n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
 n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
 n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
 n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
 n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
 n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
 n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
 n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
 n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
 n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
 n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
 n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
 n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
 n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
 n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
 n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
 n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
 n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
 n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
 n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
 n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
 n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
 n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
 n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
 n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
 n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
 n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
 n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
 n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
 n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
 n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
 n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
 n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
 n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
 n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
 n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
 n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
 n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
 n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
 n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
 n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
 n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
 n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
 n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
 n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
 n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
 n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
 n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
 n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
 n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
 n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
 n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
 n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
 n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
 n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
 n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
 n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
 n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
 n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
 n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
 n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
 n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
 n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
 n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
 n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
 n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
 n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
 n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
 n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
 n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
 n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
 n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
 n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
 n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
 n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
 n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
 n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
 n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
 n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
 n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
 n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
 n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
 n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
 n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
 n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
 n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
 n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
 n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495,
 n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
 n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
 n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
 n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
 n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535,
 n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
 n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
 n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
 n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
 n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
 n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
 n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
 n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
 n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
 n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615,
 n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
 n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
 n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
 n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
 n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655,
 n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
 n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
 n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
 n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
 n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695,
 n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
 n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
 n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
 n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
 n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735,
 n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
 n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
 n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
 n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
 n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775,
 n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
 n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
 n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
 n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
 n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815,
 n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
 n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
 n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
 n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
 n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855,
 n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
 n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
 n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
 n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
 n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
 n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
 n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
 n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
 n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
 n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
 n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
 n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
 n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
 n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
 n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
 n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
 n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
 n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
 n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
 n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
 n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
 n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
 n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
 n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
 n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
 n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
 n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
 n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
 n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
 n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
 n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
 n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
 n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
 n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
 n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
 n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
 n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
 n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
 n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
 n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
 n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
 n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
 n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
 n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
 n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
 n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
 n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
 n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
 n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
 n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
 n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
 n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
 n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
 n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
 n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
 n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
 n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
 n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
 n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
 n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
 n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
 n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
 n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
 n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
 n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
 n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
 n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
 n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
 n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
 n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
 n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
 n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
 n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
 n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
 n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
 n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
 n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
 n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
 n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
 n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
 n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
 n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
 n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
 n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
 n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
 n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
 n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
 n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
 n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
 n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
 n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
 n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
 n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
 n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
 n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
 n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
 n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
 n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
 n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
 n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
 n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
 n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
 n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
 n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
 n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
 n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
 n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
 n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
 n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
 n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
 n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
 n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
 n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
 n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
 n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
 n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
 n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
 n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
 n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
 n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
 n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
 n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
 n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
 n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
 n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
 n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
 n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
 n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
 n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
 n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
 n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
 n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
 n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
 n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
 n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
 n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
 n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
 n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
 n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
 n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
 n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
 n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
 n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
 n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
 n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
 n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
 n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031;

buf  g0 (n93, n7);
buf  g1 (n61, n18);
buf  g2 (n45, n31);
buf  g3 (n103, n9);
buf  g4 (n41, n8);
buf  g5 (n121, n16);
not  g6 (n84, n23);
not  g7 (n113, n19);
buf  g8 (n33, n31);
not  g9 (n155, n3);
not  g10 (n57, n17);
not  g11 (n97, n22);
not  g12 (n56, n11);
buf  g13 (n36, n15);
buf  g14 (n75, n1);
buf  g15 (n108, n21);
buf  g16 (n85, n10);
buf  g17 (n59, n17);
not  g18 (n47, n18);
not  g19 (n82, n12);
buf  g20 (n128, n11);
buf  g21 (n55, n17);
buf  g22 (n154, n32);
buf  g23 (n109, n9);
not  g24 (n115, n10);
not  g25 (n34, n13);
buf  g26 (n86, n12);
buf  g27 (n153, n14);
not  g28 (n80, n12);
buf  g29 (n149, n24);
not  g30 (n39, n1);
buf  g31 (n124, n8);
buf  g32 (n35, n8);
not  g33 (n116, n20);
not  g34 (n92, n23);
not  g35 (n105, n27);
buf  g36 (n79, n26);
not  g37 (n134, n30);
buf  g38 (n148, n15);
not  g39 (n68, n26);
not  g40 (n156, n9);
not  g41 (n157, n5);
not  g42 (n69, n4);
buf  g43 (n62, n20);
buf  g44 (n83, n28);
buf  g45 (n72, n25);
buf  g46 (n54, n5);
not  g47 (n110, n26);
buf  g48 (n64, n29);
not  g49 (n147, n4);
buf  g50 (n71, n16);
buf  g51 (n131, n2);
not  g52 (n48, n6);
not  g53 (n143, n3);
not  g54 (n133, n24);
not  g55 (n90, n6);
not  g56 (n76, n27);
not  g57 (n138, n14);
not  g58 (n150, n4);
not  g59 (n117, n15);
buf  g60 (n137, n3);
not  g61 (n63, n29);
not  g62 (n49, n12);
buf  g63 (n98, n32);
not  g64 (n42, n5);
not  g65 (n120, n21);
buf  g66 (n66, n22);
not  g67 (n58, n23);
not  g68 (n158, n13);
buf  g69 (n70, n2);
buf  g70 (n37, n6);
buf  g71 (n73, n22);
not  g72 (n159, n5);
buf  g73 (n52, n21);
buf  g74 (n146, n7);
buf  g75 (n118, n15);
not  g76 (n130, n29);
not  g77 (n102, n2);
not  g78 (n145, n10);
not  g79 (n87, n25);
buf  g80 (n114, n31);
not  g81 (n99, n2);
not  g82 (n81, n14);
not  g83 (n95, n30);
not  g84 (n125, n27);
buf  g85 (n67, n13);
not  g86 (n46, n19);
buf  g87 (n51, n7);
not  g88 (n144, n30);
buf  g89 (n142, n20);
not  g90 (n152, n16);
not  g91 (n44, n25);
buf  g92 (n135, n31);
not  g93 (n123, n11);
not  g94 (n53, n28);
not  g95 (n50, n9);
not  g96 (n40, n26);
buf  g97 (n38, n20);
buf  g98 (n160, n10);
buf  g99 (n126, n16);
buf  g100 (n107, n32);
buf  g101 (n151, n8);
buf  g102 (n140, n21);
not  g103 (n43, n1);
not  g104 (n139, n6);
not  g105 (n89, n24);
not  g106 (n127, n13);
not  g107 (n65, n22);
buf  g108 (n112, n24);
not  g109 (n94, n19);
buf  g110 (n74, n25);
not  g111 (n96, n1);
not  g112 (n129, n3);
not  g113 (n136, n4);
not  g114 (n60, n14);
buf  g115 (n122, n29);
buf  g116 (n104, n32);
not  g117 (n101, n28);
buf  g118 (n78, n30);
buf  g119 (n91, n17);
not  g120 (n106, n27);
buf  g121 (n77, n28);
not  g122 (n132, n18);
buf  g123 (n119, n7);
buf  g124 (n88, n23);
not  g125 (n111, n18);
not  g126 (n100, n11);
buf  g127 (n141, n19);
buf  g128 (n608, n143);
buf  g129 (n528, n75);
not  g130 (n482, n41);
buf  g131 (n635, n42);
not  g132 (n553, n146);
buf  g133 (n177, n124);
buf  g134 (n449, n42);
buf  g135 (n604, n140);
not  g136 (n171, n100);
not  g137 (n455, n140);
buf  g138 (n265, n50);
not  g139 (n296, n95);
buf  g140 (n316, n156);
buf  g141 (n367, n57);
not  g142 (n654, n153);
buf  g143 (n308, n128);
not  g144 (n485, n134);
buf  g145 (n162, n110);
not  g146 (n650, n86);
buf  g147 (n352, n94);
not  g148 (n343, n153);
not  g149 (n490, n80);
buf  g150 (n474, n120);
buf  g151 (n203, n109);
buf  g152 (n440, n122);
not  g153 (n665, n100);
not  g154 (n472, n109);
buf  g155 (n561, n129);
buf  g156 (n327, n39);
not  g157 (n401, n37);
not  g158 (n235, n62);
buf  g159 (n286, n136);
buf  g160 (n494, n118);
not  g161 (n576, n125);
buf  g162 (n234, n90);
not  g163 (n473, n60);
not  g164 (n639, n66);
buf  g165 (n621, n56);
not  g166 (n543, n90);
not  g167 (n463, n110);
buf  g168 (n573, n117);
not  g169 (n217, n85);
buf  g170 (n532, n145);
buf  g171 (n446, n54);
not  g172 (n627, n83);
buf  g173 (n632, n126);
buf  g174 (n272, n122);
not  g175 (n434, n57);
not  g176 (n338, n101);
not  g177 (n525, n131);
buf  g178 (n527, n40);
buf  g179 (n429, n139);
not  g180 (n205, n128);
buf  g181 (n392, n111);
buf  g182 (n218, n153);
not  g183 (n199, n84);
buf  g184 (n242, n103);
buf  g185 (n206, n48);
not  g186 (n366, n80);
buf  g187 (n521, n72);
not  g188 (n393, n76);
buf  g189 (n247, n84);
not  g190 (n230, n51);
buf  g191 (n280, n89);
buf  g192 (n559, n48);
not  g193 (n351, n119);
not  g194 (n496, n103);
buf  g195 (n166, n76);
not  g196 (n606, n68);
not  g197 (n184, n55);
buf  g198 (n661, n69);
not  g199 (n465, n108);
not  g200 (n670, n124);
not  g201 (n198, n57);
not  g202 (n303, n68);
not  g203 (n536, n107);
not  g204 (n486, n135);
buf  g205 (n666, n43);
not  g206 (n418, n114);
buf  g207 (n223, n142);
buf  g208 (n384, n116);
not  g209 (n570, n93);
buf  g210 (n477, n150);
buf  g211 (n616, n92);
not  g212 (n186, n136);
not  g213 (n513, n152);
buf  g214 (n614, n54);
not  g215 (n438, n99);
not  g216 (n520, n58);
buf  g217 (n535, n112);
not  g218 (n179, n152);
buf  g219 (n398, n73);
buf  g220 (n295, n96);
buf  g221 (n191, n106);
not  g222 (n596, n79);
not  g223 (n554, n58);
buf  g224 (n309, n110);
buf  g225 (n350, n45);
buf  g226 (n450, n125);
buf  g227 (n504, n111);
not  g228 (n181, n153);
not  g229 (n298, n71);
buf  g230 (n590, n79);
not  g231 (n574, n156);
not  g232 (n619, n102);
buf  g233 (n228, n96);
buf  g234 (n461, n64);
not  g235 (n617, n133);
buf  g236 (n363, n118);
buf  g237 (n251, n87);
buf  g238 (n588, n61);
buf  g239 (n385, n41);
buf  g240 (n211, n134);
buf  g241 (n187, n60);
buf  g242 (n625, n53);
buf  g243 (n657, n156);
buf  g244 (n537, n108);
buf  g245 (n193, n97);
buf  g246 (n297, n115);
buf  g247 (n368, n38);
buf  g248 (n376, n36);
buf  g249 (n315, n121);
buf  g250 (n618, n69);
not  g251 (n388, n122);
buf  g252 (n224, n127);
not  g253 (n329, n117);
not  g254 (n200, n94);
not  g255 (n600, n99);
not  g256 (n479, n97);
not  g257 (n499, n123);
not  g258 (n413, n47);
not  g259 (n257, n155);
not  g260 (n607, n112);
not  g261 (n353, n108);
not  g262 (n647, n63);
buf  g263 (n163, n65);
not  g264 (n495, n139);
buf  g265 (n567, n92);
buf  g266 (n545, n124);
buf  g267 (n260, n43);
buf  g268 (n514, n148);
buf  g269 (n173, n127);
buf  g270 (n386, n114);
not  g271 (n256, n98);
buf  g272 (n360, n156);
buf  g273 (n245, n60);
not  g274 (n491, n44);
not  g275 (n314, n104);
not  g276 (n506, n86);
buf  g277 (n221, n48);
buf  g278 (n213, n120);
buf  g279 (n640, n138);
not  g280 (n471, n63);
buf  g281 (n266, n144);
buf  g282 (n595, n144);
buf  g283 (n562, n72);
not  g284 (n522, n78);
not  g285 (n404, n99);
not  g286 (n175, n93);
not  g287 (n427, n46);
not  g288 (n551, n133);
not  g289 (n441, n151);
not  g290 (n507, n78);
not  g291 (n248, n79);
buf  g292 (n509, n147);
buf  g293 (n410, n151);
not  g294 (n356, n129);
buf  g295 (n344, n69);
not  g296 (n526, n140);
not  g297 (n176, n54);
not  g298 (n340, n116);
buf  g299 (n470, n86);
buf  g300 (n663, n40);
not  g301 (n273, n75);
buf  g302 (n458, n146);
not  g303 (n359, n123);
buf  g304 (n210, n146);
buf  g305 (n197, n121);
not  g306 (n655, n129);
buf  g307 (n500, n82);
not  g308 (n331, n73);
buf  g309 (n544, n84);
not  g310 (n364, n55);
not  g311 (n337, n137);
buf  g312 (n530, n101);
buf  g313 (n538, n77);
not  g314 (n291, n74);
buf  g315 (n660, n160);
not  g316 (n301, n44);
not  g317 (n498, n94);
buf  g318 (n254, n61);
buf  g319 (n444, n46);
buf  g320 (n539, n49);
not  g321 (n659, n59);
not  g322 (n671, n113);
buf  g323 (n307, n105);
buf  g324 (n326, n145);
not  g325 (n510, n70);
not  g326 (n282, n95);
buf  g327 (n375, n56);
buf  g328 (n488, n66);
buf  g329 (n423, n59);
not  g330 (n585, n106);
not  g331 (n229, n92);
buf  g332 (n231, n121);
not  g333 (n658, n60);
buf  g334 (n630, n116);
not  g335 (n335, n158);
not  g336 (n633, n120);
buf  g337 (n597, n134);
buf  g338 (n239, n39);
buf  g339 (n227, n111);
buf  g340 (n412, n51);
buf  g341 (n610, n50);
buf  g342 (n558, n47);
buf  g343 (n243, n129);
buf  g344 (n373, n116);
not  g345 (n594, n56);
buf  g346 (n267, n58);
not  g347 (n165, n65);
buf  g348 (n653, n109);
buf  g349 (n263, n158);
buf  g350 (n183, n71);
not  g351 (n249, n33);
buf  g352 (n253, n141);
not  g353 (n548, n118);
buf  g354 (n382, n120);
buf  g355 (n403, n43);
buf  g356 (n383, n107);
buf  g357 (n432, n87);
not  g358 (n428, n93);
not  g359 (n246, n118);
not  g360 (n212, n137);
buf  g361 (n613, n83);
not  g362 (n583, n57);
buf  g363 (n518, n52);
buf  g364 (n226, n96);
not  g365 (n207, n89);
buf  g366 (n405, n70);
not  g367 (n399, n88);
not  g368 (n628, n130);
not  g369 (n542, n141);
not  g370 (n365, n36);
buf  g371 (n484, n69);
buf  g372 (n264, n77);
buf  g373 (n631, n67);
not  g374 (n185, n58);
not  g375 (n419, n98);
buf  g376 (n390, n83);
buf  g377 (n642, n105);
not  g378 (n512, n74);
buf  g379 (n349, n65);
buf  g380 (n285, n77);
not  g381 (n409, n119);
buf  g382 (n531, n52);
not  g383 (n667, n81);
not  g384 (n323, n50);
buf  g385 (n577, n158);
not  g386 (n581, n135);
not  g387 (n648, n56);
buf  g388 (n189, n154);
buf  g389 (n268, n160);
not  g390 (n277, n89);
not  g391 (n330, n121);
buf  g392 (n233, n79);
buf  g393 (n371, n53);
buf  g394 (n417, n44);
not  g395 (n415, n36);
not  g396 (n250, n159);
buf  g397 (n241, n132);
buf  g398 (n565, n130);
buf  g399 (n487, n155);
not  g400 (n300, n115);
not  g401 (n319, n101);
not  g402 (n466, n142);
not  g403 (n435, n154);
buf  g404 (n283, n91);
not  g405 (n644, n66);
not  g406 (n219, n34);
not  g407 (n194, n135);
buf  g408 (n400, n130);
not  g409 (n420, n68);
not  g410 (n407, n148);
buf  g411 (n445, n149);
not  g412 (n334, n88);
not  g413 (n270, n104);
not  g414 (n476, n102);
not  g415 (n481, n126);
not  g416 (n192, n108);
not  g417 (n209, n90);
not  g418 (n555, n152);
buf  g419 (n168, n105);
buf  g420 (n261, n133);
buf  g421 (n589, n138);
buf  g422 (n238, n64);
buf  g423 (n305, n36);
not  g424 (n511, n143);
buf  g425 (n310, n82);
buf  g426 (n453, n34);
not  g427 (n582, n157);
not  g428 (n439, n150);
not  g429 (n497, n33);
not  g430 (n584, n49);
buf  g431 (n336, n63);
not  g432 (n624, n95);
not  g433 (n519, n87);
buf  g434 (n304, n80);
not  g435 (n372, n105);
buf  g436 (n232, n115);
buf  g437 (n201, n88);
not  g438 (n288, n45);
not  g439 (n467, n78);
buf  g440 (n575, n83);
not  g441 (n215, n122);
buf  g442 (n566, n90);
buf  g443 (n178, n99);
buf  g444 (n430, n96);
not  g445 (n195, n38);
not  g446 (n318, n148);
not  g447 (n225, n91);
not  g448 (n387, n149);
not  g449 (n172, n33);
buf  g450 (n169, n45);
buf  g451 (n389, n70);
not  g452 (n593, n148);
buf  g453 (n603, n141);
not  g454 (n651, n104);
buf  g455 (n456, n64);
buf  g456 (n609, n140);
buf  g457 (n317, n128);
buf  g458 (n332, n126);
not  g459 (n598, n125);
not  g460 (n402, n64);
not  g461 (n451, n35);
not  g462 (n508, n76);
buf  g463 (n208, n42);
buf  g464 (n259, n142);
buf  g465 (n550, n52);
not  g466 (n641, n67);
buf  g467 (n649, n103);
buf  g468 (n668, n84);
not  g469 (n188, n135);
buf  g470 (n347, n130);
buf  g471 (n502, n134);
not  g472 (n411, n45);
not  g473 (n174, n38);
buf  g474 (n569, n35);
buf  g475 (n443, n53);
not  g476 (n333, n81);
buf  g477 (n377, n157);
buf  g478 (n292, n117);
not  g479 (n167, n82);
not  g480 (n560, n65);
not  g481 (n447, n133);
not  g482 (n448, n127);
not  g483 (n556, n102);
buf  g484 (n611, n149);
buf  g485 (n483, n112);
not  g486 (n396, n104);
not  g487 (n541, n88);
buf  g488 (n454, n51);
buf  g489 (n517, n42);
not  g490 (n369, n41);
buf  g491 (n416, n59);
not  g492 (n284, n55);
not  g493 (n460, n50);
not  g494 (n599, n112);
buf  g495 (n634, n54);
buf  g496 (n237, n39);
buf  g497 (n252, n95);
not  g498 (n341, n113);
buf  g499 (n492, n46);
not  g500 (n564, n138);
not  g501 (n516, n40);
not  g502 (n636, n34);
buf  g503 (n302, n150);
buf  g504 (n170, n111);
not  g505 (n580, n33);
buf  g506 (n442, n63);
not  g507 (n276, n113);
buf  g508 (n294, n34);
not  g509 (n287, n123);
not  g510 (n459, n149);
buf  g511 (n493, n145);
not  g512 (n328, n146);
buf  g513 (n629, n144);
buf  g514 (n348, n44);
not  g515 (n214, n128);
buf  g516 (n626, n39);
buf  g517 (n320, n61);
not  g518 (n339, n53);
buf  g519 (n279, n52);
buf  g520 (n572, n47);
not  g521 (n397, n125);
not  g522 (n269, n114);
not  g523 (n408, n37);
buf  g524 (n258, n154);
not  g525 (n325, n85);
not  g526 (n362, n73);
buf  g527 (n503, n157);
not  g528 (n462, n106);
buf  g529 (n354, n92);
buf  g530 (n299, n86);
buf  g531 (n421, n37);
not  g532 (n244, n160);
buf  g533 (n312, n137);
not  g534 (n505, n71);
buf  g535 (n380, n94);
buf  g536 (n620, n81);
not  g537 (n216, n62);
not  g538 (n645, n147);
buf  g539 (n433, n41);
not  g540 (n646, n106);
not  g541 (n592, n113);
buf  g542 (n424, n159);
buf  g543 (n236, n89);
buf  g544 (n391, n151);
buf  g545 (n355, n71);
buf  g546 (n534, n147);
buf  g547 (n370, n77);
buf  g548 (n313, n78);
buf  g549 (n255, n67);
not  g550 (n568, n114);
not  g551 (n220, n132);
not  g552 (n605, n110);
buf  g553 (n346, n119);
not  g554 (n306, n80);
buf  g555 (n547, n67);
buf  g556 (n515, n101);
buf  g557 (n571, n144);
buf  g558 (n357, n97);
buf  g559 (n395, n158);
not  g560 (n468, n66);
not  g561 (n601, n47);
not  g562 (n281, n155);
buf  g563 (n374, n72);
buf  g564 (n656, n109);
not  g565 (n475, n37);
not  g566 (n378, n98);
not  g567 (n240, n75);
not  g568 (n190, n119);
not  g569 (n361, n35);
buf  g570 (n422, n103);
not  g571 (n480, n142);
buf  g572 (n615, n107);
not  g573 (n222, n155);
buf  g574 (n612, n48);
buf  g575 (n652, n154);
not  g576 (n602, n62);
buf  g577 (n342, n100);
buf  g578 (n489, n143);
not  g579 (n164, n102);
not  g580 (n290, n124);
not  g581 (n426, n132);
buf  g582 (n274, n51);
not  g583 (n381, n55);
not  g584 (n436, n40);
buf  g585 (n623, n117);
not  g586 (n643, n136);
buf  g587 (n271, n91);
not  g588 (n664, n62);
buf  g589 (n549, n141);
buf  g590 (n324, n159);
not  g591 (n523, n76);
buf  g592 (n275, n85);
buf  g593 (n662, n59);
buf  g594 (n202, n139);
buf  g595 (n464, n74);
buf  g596 (n196, n87);
buf  g597 (n563, n38);
not  g598 (n478, n138);
not  g599 (n579, n61);
not  g600 (n591, n136);
not  g601 (n587, n115);
not  g602 (n452, n82);
buf  g603 (n557, n137);
buf  g604 (n524, n72);
buf  g605 (n379, n49);
buf  g606 (n546, n131);
buf  g607 (n262, n150);
not  g608 (n289, n131);
buf  g609 (n469, n151);
not  g610 (n321, n159);
buf  g611 (n529, n93);
not  g612 (n414, n100);
not  g613 (n437, n147);
not  g614 (n622, n126);
not  g615 (n180, n139);
buf  g616 (n637, n85);
not  g617 (n204, n70);
not  g618 (n669, n152);
buf  g619 (n457, n132);
buf  g620 (n394, n73);
not  g621 (n293, n145);
not  g622 (n540, n143);
not  g623 (n578, n49);
not  g624 (n552, n46);
not  g625 (n345, n123);
buf  g626 (n425, n75);
buf  g627 (n322, n43);
not  g628 (n586, n157);
not  g629 (n311, n127);
buf  g630 (n278, n74);
buf  g631 (n638, n68);
not  g632 (n161, n91);
not  g633 (n533, n107);
buf  g634 (n358, n81);
not  g635 (n182, n35);
not  g636 (n501, n98);
buf  g637 (n406, n97);
buf  g638 (n431, n131);
nand g639 (n1126, n476, n579, n466, n203);
nor  g640 (n749, n529, n642, n519, n638);
nor  g641 (n935, n273, n666, n439, n573);
nand g642 (n809, n446, n388, n592, n375);
or   g643 (n855, n474, n276, n390, n632);
and  g644 (n959, n227, n198, n387, n512);
xnor g645 (n1019, n575, n246, n664, n379);
xor  g646 (n715, n279, n382, n325, n274);
xor  g647 (n687, n215, n569, n432, n632);
xor  g648 (n728, n382, n434, n659, n525);
nor  g649 (n1002, n448, n199, n652, n393);
xor  g650 (n1015, n286, n524, n431, n175);
nor  g651 (n1068, n518, n327, n427, n265);
or   g652 (n1027, n216, n307, n356, n340);
xnor g653 (n1146, n586, n473, n348, n542);
and  g654 (n859, n252, n259, n639, n274);
nor  g655 (n927, n297, n299, n596, n316);
nand g656 (n1088, n383, n474, n344, n641);
xnor g657 (n784, n255, n535, n591, n393);
and  g658 (n762, n425, n508, n477, n445);
and  g659 (n810, n523, n528, n275, n418);
nor  g660 (n1122, n480, n592, n616, n251);
xnor g661 (n999, n391, n655, n163, n525);
nor  g662 (n985, n552, n266, n570, n623);
or   g663 (n729, n404, n515, n625, n634);
and  g664 (n778, n439, n244, n521, n274);
nor  g665 (n837, n299, n370, n218, n410);
xor  g666 (n904, n511, n527, n318, n394);
nand g667 (n1058, n404, n562, n546, n257);
nor  g668 (n1040, n454, n217, n317, n354);
nand g669 (n1057, n258, n301, n263, n595);
and  g670 (n843, n346, n660, n227, n506);
nand g671 (n848, n298, n312, n550, n226);
nor  g672 (n720, n488, n654, n444, n340);
and  g673 (n709, n353, n248, n546, n552);
nand g674 (n673, n202, n389, n520, n656);
and  g675 (n681, n212, n509, n400, n353);
xnor g676 (n1152, n414, n236, n652, n284);
nand g677 (n953, n472, n399, n553, n597);
or   g678 (n968, n602, n574, n622, n219);
xor  g679 (n1093, n456, n268, n528, n515);
nor  g680 (n845, n531, n620, n501, n662);
xnor g681 (n733, n547, n332, n618, n288);
xor  g682 (n731, n417, n542, n581, n279);
nand g683 (n773, n462, n287, n343, n546);
xor  g684 (n917, n259, n197, n645, n229);
nand g685 (n834, n495, n397, n377, n615);
nor  g686 (n975, n245, n609, n544, n486);
and  g687 (n829, n620, n289, n319, n523);
xnor g688 (n746, n457, n320, n488, n622);
nand g689 (n994, n614, n469, n545, n667);
and  g690 (n833, n388, n411, n273, n578);
or   g691 (n777, n385, n329, n333, n668);
or   g692 (n692, n268, n482, n457, n637);
and  g693 (n942, n342, n451, n564, n270);
and  g694 (n915, n447, n451, n471, n630);
or   g695 (n701, n460, n416, n438, n528);
and  g696 (n782, n330, n513, n566, n209);
or   g697 (n831, n590, n584, n652, n453);
xnor g698 (n721, n482, n239, n539, n468);
and  g699 (n940, n518, n657, n457, n376);
nor  g700 (n871, n538, n579, n534, n633);
nand g701 (n865, n309, n359, n189, n278);
or   g702 (n956, n581, n519, n241, n276);
and  g703 (n813, n420, n352, n233, n493);
or   g704 (n1157, n220, n423, n485, n517);
and  g705 (n1113, n283, n386, n269, n344);
xor  g706 (n876, n440, n362, n658, n517);
xor  g707 (n839, n664, n261, n209, n303);
and  g708 (n769, n205, n405, n663, n322);
xor  g709 (n965, n364, n355, n577, n370);
nand g710 (n913, n210, n548, n656, n295);
or   g711 (n1063, n565, n374, n305, n338);
and  g712 (n901, n328, n272, n519, n464);
xor  g713 (n753, n289, n467, n418, n594);
nor  g714 (n1052, n299, n427, n193, n243);
xnor g715 (n735, n613, n605, n486, n665);
or   g716 (n847, n287, n251, n647, n537);
nand g717 (n1062, n526, n215, n297, n636);
xor  g718 (n883, n230, n302, n585, n337);
xnor g719 (n1096, n558, n557, n670, n617);
nor  g720 (n947, n560, n435, n661, n624);
nand g721 (n991, n217, n467, n308, n261);
and  g722 (n711, n578, n382, n368, n442);
and  g723 (n1082, n218, n293, n643, n598);
nand g724 (n874, n292, n210, n419, n587);
xnor g725 (n1109, n649, n179, n214, n432);
or   g726 (n805, n465, n455, n268, n317);
or   g727 (n1117, n426, n545, n522, n355);
xor  g728 (n678, n290, n459, n496, n652);
nor  g729 (n868, n362, n429, n213, n237);
xor  g730 (n811, n462, n426, n341, n200);
xnor g731 (n877, n579, n637, n235, n500);
xnor g732 (n1094, n228, n321, n628, n203);
or   g733 (n807, n219, n568, n286, n254);
nand g734 (n747, n571, n391, n498, n523);
xnor g735 (n1049, n263, n529, n501, n610);
and  g736 (n960, n533, n238, n398, n258);
xor  g737 (n911, n424, n588, n606, n510);
and  g738 (n1086, n603, n572, n366, n356);
and  g739 (n791, n419, n422, n396, n610);
and  g740 (n1147, n464, n358, n283, n561);
nand g741 (n768, n243, n548, n527, n642);
xor  g742 (n864, n285, n193, n578, n502);
nand g743 (n986, n629, n282, n265, n495);
xnor g744 (n952, n237, n556, n507, n266);
nor  g745 (n1044, n617, n469, n529, n349);
nand g746 (n841, n208, n451, n573, n635);
or   g747 (n821, n489, n367, n516, n535);
and  g748 (n995, n223, n419, n322, n387);
nor  g749 (n724, n294, n571, n643, n248);
nand g750 (n785, n445, n250, n391, n364);
or   g751 (n1038, n648, n587, n394, n272);
nor  g752 (n706, n337, n408, n395, n439);
or   g753 (n1030, n514, n544, n425, n555);
nand g754 (n1118, n240, n640, n295, n241);
nor  g755 (n825, n242, n461, n608, n354);
xnor g756 (n1016, n411, n410, n612, n424);
or   g757 (n802, n594, n265, n552, n329);
xnor g758 (n1130, n178, n354, n286, n663);
xor  g759 (n844, n644, n305, n285, n551);
and  g760 (n686, n522, n242, n281, n330);
nor  g761 (n1025, n352, n364, n529, n206);
xnor g762 (n1110, n397, n426, n367, n305);
and  g763 (n693, n228, n635, n383, n489);
xor  g764 (n861, n177, n328, n542, n379);
or   g765 (n1042, n344, n301, n559, n635);
nand g766 (n938, n287, n610, n391, n268);
xor  g767 (n967, n363, n264, n550, n303);
xnor g768 (n740, n655, n670, n493, n560);
xnor g769 (n688, n621, n576, n357, n350);
xor  g770 (n817, n479, n663, n330, n659);
or   g771 (n727, n279, n580, n539, n537);
xor  g772 (n714, n490, n284, n290, n576);
nand g773 (n774, n378, n478, n239, n509);
xor  g774 (n838, n272, n608, n327, n478);
xor  g775 (n886, n242, n223, n192, n658);
or   g776 (n1100, n366, n406, n440, n200);
or   g777 (n689, n564, n316, n477, n240);
nand g778 (n1033, n384, n412, n670, n663);
nand g779 (n808, n449, n421, n588, n204);
nand g780 (n980, n311, n277, n453, n362);
nand g781 (n897, n459, n351, n271, n597);
xor  g782 (n976, n537, n517, n598, n311);
nand g783 (n966, n336, n488, n299, n416);
nor  g784 (n1144, n275, n214, n471, n414);
xor  g785 (n931, n205, n563, n571, n405);
or   g786 (n754, n256, n420, n452, n571);
and  g787 (n744, n350, n413, n583, n487);
and  g788 (n1132, n373, n181, n448, n283);
nor  g789 (n1077, n641, n608, n588, n654);
nor  g790 (n923, n415, n558, n645, n468);
or   g791 (n1155, n253, n535, n595);
or   g792 (n770, n444, n474, n609, n536);
xnor g793 (n981, n428, n407, n204, n522);
or   g794 (n1036, n577, n465, n624, n293);
and  g795 (n766, n594, n195, n560, n221);
xnor g796 (n957, n451, n208, n375, n452);
xnor g797 (n800, n470, n506, n201, n338);
and  g798 (n779, n244, n430, n354, n551);
nand g799 (n707, n651, n490, n342, n271);
and  g800 (n1056, n194, n480, n569, n301);
nand g801 (n962, n256, n613, n656, n547);
nor  g802 (n1123, n492, n213, n503, n208);
nor  g803 (n925, n365, n605, n350, n398);
nor  g804 (n875, n332, n618, n270, n463);
nor  g805 (n1031, n166, n650, n408, n195);
and  g806 (n900, n416, n646, n282, n434);
xnor g807 (n892, n476, n654, n635, n477);
or   g808 (n713, n568, n260, n566, n582);
or   g809 (n708, n648, n201, n359, n280);
xor  g810 (n984, n446, n371, n366, n452);
xnor g811 (n1151, n228, n584, n375, n638);
xor  g812 (n699, n526, n559, n276, n585);
and  g813 (n930, n349, n653, n604, n281);
xor  g814 (n819, n436, n606, n238, n356);
xor  g815 (n939, n280, n340, n489, n339);
nand g816 (n842, n250, n401, n664, n356);
xnor g817 (n878, n436, n433, n279, n483);
xor  g818 (n826, n550, n338, n374, n211);
nor  g819 (n910, n367, n585, n225, n328);
and  g820 (n1134, n324, n504, n619, n371);
and  g821 (n1081, n404, n540, n332, n536);
nand g822 (n1129, n641, n502, n260, n226);
xnor g823 (n1020, n576, n557, n521, n206);
nand g824 (n973, n236, n380, n193, n614);
nor  g825 (n691, n617, n517, n374, n233);
nor  g826 (n790, n222, n570, n370, n492);
or   g827 (n716, n450, n469, n540, n197);
xor  g828 (n792, n382, n252, n234, n491);
or   g829 (n1143, n310, n341, n562, n620);
or   g830 (n1000, n224, n369, n314, n627);
nor  g831 (n1097, n370, n583, n291, n458);
nand g832 (n884, n561, n524, n303, n657);
nand g833 (n788, n222, n310, n412, n567);
nor  g834 (n972, n267, n544, n583, n231);
or   g835 (n964, n460, n258, n584, n473);
and  g836 (n1128, n347, n538, n249, n398);
xor  g837 (n1125, n472, n478, n200, n586);
and  g838 (n1099, n445, n603, n499, n249);
or   g839 (n739, n294, n548, n330, n555);
xnor g840 (n1069, n230, n305, n357, n626);
nor  g841 (n989, n390, n463, n409, n312);
and  g842 (n1131, n420, n576, n442, n358);
nor  g843 (n899, n515, n229, n296, n492);
xnor g844 (n906, n218, n336, n654, n660);
nor  g845 (n896, n339, n220, n434, n314);
or   g846 (n830, n237, n498, n432, n569);
nand g847 (n869, n486, n414, n403, n669);
or   g848 (n1017, n199, n196, n668, n376);
nand g849 (n1046, n547, n262, n371, n483);
nor  g850 (n801, n361, n252, n650, n479);
nand g851 (n1035, n446, n358, n459, n246);
and  g852 (n870, n533, n565, n337, n628);
xor  g853 (n717, n543, n235, n615, n462);
xor  g854 (n1053, n631, n326, n449, n570);
and  g855 (n1139, n213, n172, n622, n581);
and  g856 (n786, n437, n325, n617, n504);
xnor g857 (n993, n353, n461, n618, n502);
xor  g858 (n974, n573, n402, n334, n545);
nand g859 (n889, n361, n577, n320, n619);
xor  g860 (n863, n533, n666, n450, n422);
nand g861 (n794, n516, n463, n502, n387);
nand g862 (n887, n497, n473, n188, n232);
and  g863 (n951, n436, n401, n368, n240);
and  g864 (n853, n509, n369, n417, n207);
nor  g865 (n902, n209, n486, n211, n510);
and  g866 (n705, n381, n167, n559, n285);
and  g867 (n955, n384, n420, n532, n496);
xnor g868 (n695, n217, n468, n292, n479);
and  g869 (n682, n444, n236, n437, n380);
nor  g870 (n684, n426, n435, n363, n582);
xor  g871 (n1090, n331, n484, n229, n365);
and  g872 (n704, n300, n161, n644, n513);
nand g873 (n1029, n428, n534, n632, n449);
nor  g874 (n1003, n409, n222, n421, n627);
and  g875 (n1119, n512, n392, n417, n522);
xor  g876 (n1066, n372, n649, n360, n415);
xor  g877 (n1012, n650, n405, n423, n562);
nand g878 (n836, n613, n590, n347, n484);
nand g879 (n1112, n619, n653, n514, n633);
nand g880 (n885, n287, n607, n423, n282);
or   g881 (n905, n389, n496, n376, n668);
xnor g882 (n1149, n456, n405, n466, n607);
xnor g883 (n763, n303, n216, n265, n554);
nand g884 (n916, n343, n271, n563, n328);
and  g885 (n932, n362, n457, n418, n599);
xor  g886 (n926, n400, n278, n384, n660);
xnor g887 (n949, n631, n348, n491, n372);
nand g888 (n1045, n224, n647, n601, n360);
and  g889 (n1032, n511, n291, n377, n623);
nor  g890 (n1138, n335, n538, n527, n183);
nand g891 (n755, n225, n615, n465, n204);
and  g892 (n1091, n207, n307, n645, n438);
xor  g893 (n1013, n295, n277, n290, n607);
or   g894 (n1084, n346, n667, n358, n243);
nand g895 (n954, n381, n440, n619, n168);
nor  g896 (n1095, n469, n390, n602, n388);
xor  g897 (n872, n227, n593, n386, n625);
nand g898 (n1010, n302, n253, n638, n226);
nand g899 (n1106, n556, n385, n452, n424);
nor  g900 (n856, n563, n430, n435, n575);
xnor g901 (n1048, n403, n507, n262, n234);
nor  g902 (n685, n417, n491, n562, n345);
nor  g903 (n798, n579, n374, n171, n233);
nor  g904 (n990, n460, n325, n630, n443);
nand g905 (n726, n441, n357, n514, n256);
xor  g906 (n1098, n394, n251, n532, n642);
nor  g907 (n780, n314, n255, n640, n306);
xnor g908 (n849, n267, n366, n564, n234);
xor  g909 (n946, n257, n485, n352, n412);
or   g910 (n674, n463, n349, n643, n500);
xor  g911 (n759, n304, n455, n197, n516);
and  g912 (n795, n329, n647, n547, n304);
and  g913 (n1028, n478, n302, n347, n633);
nand g914 (n852, n359, n397, n281, n596);
xnor g915 (n1055, n345, n400, n296, n393);
nor  g916 (n862, n378, n208, n274, n202);
xnor g917 (n987, n232, n264, n225, n331);
xnor g918 (n1023, n248, n526, n476, n254);
or   g919 (n867, n587, n657, n367, n464);
xor  g920 (n761, n636, n378, n428, n215);
xor  g921 (n1070, n211, n306, n205, n667);
nand g922 (n977, n472, n525, n176, n590);
nand g923 (n732, n611, n238, n549, n225);
nand g924 (n846, n531, n498, n523, n342);
xor  g925 (n982, n247, n316, n582, n249);
xnor g926 (n1089, n649, n246, n591, n631);
xnor g927 (n922, n372, n603, n308, n551);
xor  g928 (n950, n553, n580, n399, n505);
nand g929 (n971, n474, n380, n492, n428);
nor  g930 (n1136, n515, n611, n373, n454);
and  g931 (n1124, n292, n436, n437, n343);
or   g932 (n1103, n239, n621, n499, n269);
nand g933 (n745, n395, n186, n170, n219);
or   g934 (n696, n557, n651, n311, n653);
nand g935 (n969, n508, n574, n468, n213);
or   g936 (n1142, n180, n419, n289, n645);
and  g937 (n803, n422, n633, n310, n216);
nand g938 (n1073, n524, n568, n311, n321);
nor  g939 (n827, n625, n164, n441, n604);
nand g940 (n775, n383, n616, n651, n658);
nand g941 (n734, n266, n614, n324, n626);
xnor g942 (n992, n456, n232, n313, n326);
nor  g943 (n700, n503, n261, n470, n605);
nand g944 (n928, n235, n326, n317, n343);
xnor g945 (n1115, n516, n493, n668, n199);
and  g946 (n858, n404, n276, n410, n494);
nor  g947 (n880, n612, n600, n558);
or   g948 (n1101, n462, n498, n341, n563);
or   g949 (n933, n304, n254, n622, n513);
nor  g950 (n676, n269, n409, n371, n350);
xnor g951 (n1153, n281, n427, n572, n618);
nor  g952 (n1026, n580, n278, n442, n665);
xor  g953 (n757, n203, n307, n406, n408);
nand g954 (n1051, n485, n210, n256, n454);
xor  g955 (n924, n433, n490, n539, n248);
xnor g956 (n797, n666, n253, n588, n497);
nand g957 (n748, n558, n278, n379, n346);
xnor g958 (n944, n361, n396, n560, n650);
and  g959 (n814, n365, n308, n506, n241);
or   g960 (n1145, n583, n338, n526, n387);
and  g961 (n1054, n480, n629, n567, n506);
xor  g962 (n672, n264, n669, n612, n329);
or   g963 (n679, n334, n572, n270, n377);
or   g964 (n937, n433, n220, n304, n199);
nand g965 (n1047, n269, n368, n608, n628);
or   g966 (n822, n418, n471, n589, n255);
nand g967 (n703, n507, n298, n206, n584);
xnor g968 (n816, n283, n593, n230, n567);
and  g969 (n1011, n500, n378, n389, n224);
and  g970 (n997, n388, n482, n296, n315);
xnor g971 (n1050, n202, n323, n621, n312);
xor  g972 (n888, n471, n270, n553, n664);
nor  g973 (n963, n534, n505, n297, n295);
nor  g974 (n948, n363, n429, n323, n425);
xor  g975 (n1137, n195, n435, n628, n259);
nor  g976 (n1102, n196, n389, n221, n335);
nor  g977 (n898, n282, n626, n401, n284);
nor  g978 (n1135, n430, n606, n595, n267);
xnor g979 (n767, n531, n360, n317, n630);
nand g980 (n1114, n597, n629, n589, n313);
or   g981 (n882, n455, n661, n448, n198);
or   g982 (n1121, n277, n290, n217, n597);
or   g983 (n783, n549, n554, n565, n392);
xor  g984 (n860, n302, n660, n607, n294);
nor  g985 (n1083, n551, n424, n626, n640);
nand g986 (n771, n540, n537, n432, n252);
or   g987 (n789, n438, n394, n327, n613);
and  g988 (n907, n288, n477, n349, n251);
nand g989 (n1156, n434, n291, n413, n411);
xnor g990 (n1018, n657, n641, n399, n308);
and  g991 (n894, n173, n545, n518, n490);
nor  g992 (n694, n541, n347, n629, n355);
xor  g993 (n893, n401, n623, n300, n211);
nor  g994 (n718, n570, n390, n294, n438);
and  g995 (n970, n162, n580, n554, n266);
nand g996 (n1061, n566, n344, n634, n495);
and  g997 (n820, n514, n510, n651, n549);
nor  g998 (n675, n423, n476, n400, n369);
nor  g999 (n1150, n313, n507, n206, n264);
xnor g1000 (n1072, n322, n273, n223, n320);
and  g1001 (n680, n623, n443, n325, n288);
xor  g1002 (n854, n611, n479, n585, n503);
xor  g1003 (n764, n449, n194, n255, n616);
nor  g1004 (n1021, n262, n319, n599, n345);
nor  g1005 (n912, n565, n625, n624, n599);
nand g1006 (n765, n554, n203, n530, n196);
or   g1007 (n1127, n307, n272, n319, n586);
xnor g1008 (n804, n620, n267, n543, n481);
xnor g1009 (n1133, n231, n245, n443);
or   g1010 (n1001, n331, n646, n598, n323);
nand g1011 (n1022, n413, n226, n415, n646);
nand g1012 (n1108, n327, n429, n241, n497);
xor  g1013 (n903, n601, n323, n501, n541);
xor  g1014 (n857, n310, n348, n489, n353);
and  g1015 (n812, n601, n300, n609, n335);
and  g1016 (n793, n503, n662, n339, n383);
or   g1017 (n772, n306, n293, n351, n301);
and  g1018 (n702, n351, n644, n561, n495);
nand g1019 (n698, n643, n357, n174, n263);
and  g1020 (n1037, n467, n373, n525, n512);
xor  g1021 (n919, n250, n321, n348, n249);
xor  g1022 (n758, n574, n421, n244, n408);
xor  g1023 (n1075, n397, n667, n589, n361);
nor  g1024 (n909, n413, n437, n292, n508);
xnor g1025 (n1074, n395, n409, n555, n485);
nand g1026 (n806, n662, n591, n480, n454);
and  g1027 (n988, n271, n298, n316, n572);
nor  g1028 (n1116, n494, n656, n639, n665);
nand g1029 (n998, n614, n273, n355, n319);
and  g1030 (n1005, n368, n442, n466, n655);
nand g1031 (n737, n415, n447, n466, n602);
xor  g1032 (n799, n602, n600, n376, n214);
xor  g1033 (n850, n606, n333, n483, n286);
or   g1034 (n941, n306, n557, n385, n318);
nand g1035 (n983, n336, n592, n288, n235);
xor  g1036 (n1078, n505, n483, n518, n548);
or   g1037 (n929, n254, n402, n193, n441);
or   g1038 (n866, n333, n484, n459, n535);
nor  g1039 (n891, n487, n277, n453, n212);
xnor g1040 (n914, n291, n407, n577, n497);
or   g1041 (n1104, n567, n508, n530, n453);
xor  g1042 (n934, n410, n470, n369, n194);
or   g1043 (n881, n247, n488, n232, n359);
xor  g1044 (n1024, n345, n636, n574, n360);
nor  g1045 (n835, n482, n315, n324, n219);
or   g1046 (n1004, n406, n247, n511, n464);
nor  g1047 (n840, n309, n627, n377, n407);
nand g1048 (n879, n300, n594, n341, n403);
or   g1049 (n828, n534, n637, n592, n520);
or   g1050 (n1107, n575, n566, n448, n624);
or   g1051 (n1085, n631, n586, n421, n399);
and  g1052 (n1071, n223, n411, n458, n596);
xor  g1053 (n908, n194, n533, n207, n621);
nor  g1054 (n1141, n260, n245, n528, n364);
xnor g1055 (n1006, n634, n504, n380, n556);
xor  g1056 (n751, n505, n246, n322, n450);
xor  g1057 (n1064, n564, n412, n250, n334);
xor  g1058 (n945, n342, n589, n393, n289);
nor  g1059 (n743, n649, n467, n165, n637);
nor  g1060 (n996, n659, n481, n416, n541);
xnor g1061 (n730, n598, n262, n429, n431);
xnor g1062 (n873, n293, n540, n207, n509);
xnor g1063 (n722, n609, n240, n541, n242);
xnor g1064 (n1140, n539, n313, n231, n200);
nand g1065 (n920, n494, n326, n559, n195);
and  g1066 (n1076, n536, n275, n169, n340);
xor  g1067 (n738, n520, n662, n632, n210);
or   g1068 (n1154, n318, n375, n324, n481);
nand g1069 (n1079, n441, n636, n427, n640);
and  g1070 (n958, n501, n315, n532, n587);
nor  g1071 (n1092, n484, n599, n475, n431);
nand g1072 (n725, n458, n385, n334, n569);
xor  g1073 (n750, n553, n321, n542, n499);
xor  g1074 (n736, n446, n475, n309, n653);
xnor g1075 (n1039, n601, n461, n475, n639);
xnor g1076 (n741, n536, n227, n336, n634);
or   g1077 (n677, n275, n239, n512, n472);
or   g1078 (n1043, n261, n552, n611, n214);
and  g1079 (n895, n351, n259, n381, n615);
nand g1080 (n742, n422, n561, n531, n431);
and  g1081 (n710, n312, n524, n447, n257);
nor  g1082 (n760, n285, n543, n465, n284);
nand g1083 (n781, n659, n549, n519, n603);
and  g1084 (n978, n231, n555, n456, n333);
nand g1085 (n1059, n204, n392, n297, n538);
or   g1086 (n918, n581, n544, n236, n494);
xnor g1087 (n1120, n578, n510, n646, n473);
nor  g1088 (n832, n314, n201, n527, n243);
or   g1089 (n1041, n215, n221, n298, n445);
xnor g1090 (n1148, n414, n395, n430, n372);
and  g1091 (n1087, n280, n648, n201, n309);
nand g1092 (n690, n331, n185, n669, n244);
and  g1093 (n723, n425, n184, n593, n600);
xnor g1094 (n1060, n191, n630, n229, n443);
nand g1095 (n936, n363, n318, n499, n237);
or   g1096 (n796, n639, n258, n669, n280);
xnor g1097 (n1009, n220, n543, n253, n247);
xnor g1098 (n1111, n337, n320, n238, n440);
or   g1099 (n890, n209, n521, n504, n610);
and  g1100 (n752, n205, n493, n666, n379);
or   g1101 (n815, n260, n648, n612, n257);
xor  g1102 (n1067, n198, n365, n568, n582);
and  g1103 (n1105, n591, n593, n573, n665);
and  g1104 (n1007, n496, n604, n373, n661);
nor  g1105 (n697, n605, n638, n458, n216);
xnor g1106 (n921, n475, n521, n511, n661);
and  g1107 (n818, n487, n296, n386, n513);
and  g1108 (n979, n187, n604, n234, n658);
and  g1109 (n823, n616, n550, n196, n197);
and  g1110 (n719, n396, n433, n444, n202);
or   g1111 (n961, n406, n386, n352, n439);
or   g1112 (n824, n530, n556, n520, n575);
nand g1113 (n943, n402, n530, n346, n481);
xor  g1114 (n1034, n500, n447, n222, n218);
or   g1115 (n1080, n335, n221, n315, n491);
nor  g1116 (n1014, n596, n460, n228, n487);
or   g1117 (n712, n339, n212, n642, n407);
xor  g1118 (n776, n670, n546, n450, n461);
xnor g1119 (n1008, n403, n263, n182, n532);
xor  g1120 (n1065, n384, n332, n190, n396);
or   g1121 (n683, n655, n233, n627, n644);
xnor g1122 (n851, n470, n398, n198, n381);
and  g1123 (n787, n455, n647, n402, n230);
or   g1124 (n756, n224, n212, n590, n392);
buf  g1125 (n1168, n684);
buf  g1126 (n1161, n688);
not  g1127 (n1180, n693);
buf  g1128 (n1172, n679);
not  g1129 (n1185, n689);
buf  g1130 (n1181, n699);
buf  g1131 (n1176, n690);
buf  g1132 (n1174, n692);
not  g1133 (n1167, n673);
buf  g1134 (n1173, n696);
buf  g1135 (n1163, n691);
not  g1136 (n1175, n694);
not  g1137 (n1183, n678);
not  g1138 (n1160, n682);
buf  g1139 (n1179, n677);
buf  g1140 (n1164, n681);
not  g1141 (n1166, n697);
buf  g1142 (n1162, n685);
buf  g1143 (n1178, n676);
not  g1144 (n1169, n683);
not  g1145 (n1159, n675);
not  g1146 (n1184, n672);
not  g1147 (n1182, n698);
buf  g1148 (n1171, n674);
not  g1149 (n1177, n687);
not  g1150 (n1158, n680);
not  g1151 (n1165, n695);
buf  g1152 (n1170, n686);
buf  g1153 (n1191, n1159);
buf  g1154 (n1188, n700);
nand g1155 (n1192, n1158, n1160);
nand g1156 (n1187, n1159, n1159, n706, n701);
nand g1157 (n1189, n707, n1158, n710, n703);
and  g1158 (n1186, n705, n712, n709, n704);
xor  g1159 (n1190, n1158, n708, n711, n702);
buf  g1160 (n1207, n1187);
not  g1161 (n1199, n1187);
buf  g1162 (n1201, n1187);
not  g1163 (n1193, n713);
buf  g1164 (n1204, n1189);
buf  g1165 (n1208, n1186);
buf  g1166 (n1194, n1188);
not  g1167 (n1197, n1188);
not  g1168 (n1205, n716);
not  g1169 (n1202, n1186);
buf  g1170 (n1198, n714);
buf  g1171 (n1203, n1187);
not  g1172 (n1196, n717);
buf  g1173 (n1195, n1188);
nand g1174 (n1206, n1189, n718, n715, n1186);
xor  g1175 (n1200, n1186, n1189, n1188);
buf  g1176 (n1214, n1196);
buf  g1177 (n1222, n719);
buf  g1178 (n1211, n1194);
buf  g1179 (n1216, n1193);
not  g1180 (n1220, n1195);
not  g1181 (n1215, n1195);
buf  g1182 (n1217, n1196);
not  g1183 (n1210, n1193);
not  g1184 (n1219, n1195);
not  g1185 (n1224, n1195);
buf  g1186 (n1218, n1194);
not  g1187 (n1212, n721);
not  g1188 (n1213, n1193);
not  g1189 (n1209, n1194);
and  g1190 (n1223, n720, n1194);
xnor g1191 (n1221, n1193, n722, n1196);
buf  g1192 (n1225, n1215);
buf  g1193 (n1233, n1212);
buf  g1194 (n1230, n1213);
buf  g1195 (n1231, n1214);
not  g1196 (n1229, n1211);
not  g1197 (n1227, n1209);
not  g1198 (n1226, n1215);
not  g1199 (n1228, n1215);
not  g1200 (n1234, n1215);
not  g1201 (n1232, n1210);
nor  g1202 (n1235, n828, n804, n1226, n727);
nor  g1203 (n1258, n748, n776, n812, n1233);
xor  g1204 (n1265, n780, n829, n1228, n741);
and  g1205 (n1239, n738, n1226, n824, n1233);
nor  g1206 (n1270, n797, n775, n781, n757);
or   g1207 (n1263, n742, n765, n782, n736);
or   g1208 (n1248, n818, n799, n770, n1225);
xor  g1209 (n1261, n806, n1231, n801, n752);
xnor g1210 (n1246, n729, n723, n1229, n756);
nor  g1211 (n1241, n761, n779, n1227, n732);
xnor g1212 (n1259, n789, n1231, n815, n726);
xor  g1213 (n1262, n784, n800, n814, n1232);
xor  g1214 (n1264, n737, n745, n1229, n787);
nand g1215 (n1267, n743, n731, n766, n777);
nor  g1216 (n1243, n1227, n791, n817, n755);
xor  g1217 (n1238, n767, n763, n1234, n1231);
and  g1218 (n1242, n802, n747, n751, n810);
xor  g1219 (n1255, n730, n768, n754, n769);
nor  g1220 (n1251, n809, n813, n807, n808);
or   g1221 (n1249, n1233, n1230, n1226, n1227);
nor  g1222 (n1247, n739, n825, n1226, n803);
nand g1223 (n1253, n1228, n771, n728, n774);
or   g1224 (n1244, n798, n733, n821, n740);
and  g1225 (n1236, n785, n735, n744, n811);
nand g1226 (n1257, n773, n1225, n1233, n772);
xor  g1227 (n1268, n1229, n823, n792, n1232);
or   g1228 (n1250, n764, n750, n746, n1228);
nor  g1229 (n1254, n793, n816, n1230, n724);
nand g1230 (n1266, n749, n1230, n1231);
or   g1231 (n1269, n796, n833, n758, n832);
nand g1232 (n1252, n1225, n725, n1228, n778);
xor  g1233 (n1271, n831, n805, n790, n786);
xor  g1234 (n1240, n1229, n795, n822, n1225);
xnor g1235 (n1237, n794, n1227, n762, n759);
xor  g1236 (n1256, n760, n1232, n753, n820);
and  g1237 (n1260, n1232, n788, n830, n827);
xor  g1238 (n1245, n826, n819, n783, n734);
buf  g1239 (n1276, n1256);
not  g1240 (n1280, n1258);
buf  g1241 (n1273, n839);
not  g1242 (n1277, n1261);
not  g1243 (n1278, n1263);
buf  g1244 (n1279, n1257);
not  g1245 (n1274, n1262);
buf  g1246 (n1275, n835);
nand g1247 (n1281, n834, n837, n1265, n1264);
nand g1248 (n1272, n836, n1260, n1259, n838);
nand g1249 (n1312, n1181, n1162, n847, n1278);
or   g1250 (n1299, n1183, n1177, n845, n1172);
and  g1251 (n1307, n1274, n1171, n851, n1163);
xor  g1252 (n1304, n1171, n1278, n1281, n1168);
xnor g1253 (n1315, n1171, n1163, n1185, n1280);
nor  g1254 (n1285, n1169, n1179, n1275, n1161);
xor  g1255 (n1310, n1173, n1162, n1174, n1170);
xor  g1256 (n1297, n1275, n1162, n1273, n1185);
xor  g1257 (n1314, n1279, n1167, n1177, n1170);
and  g1258 (n1318, n1168, n1274, n1185, n1183);
xor  g1259 (n1282, n1279, n1181, n1175);
xnor g1260 (n1302, n1276, n1280, n1182, n1172);
xnor g1261 (n1298, n1164, n848, n1165, n1176);
xor  g1262 (n1316, n1273, n1167, n841, n1173);
nand g1263 (n1294, n840, n1172, n1175, n1275);
nor  g1264 (n1306, n1277, n1277, n1174, n1181);
xor  g1265 (n1308, n1166, n1168, n1161, n1276);
or   g1266 (n1288, n1280, n1165, n1176, n1181);
nand g1267 (n1309, n1167, n849, n1180, n1277);
and  g1268 (n1286, n1278, n1177, n1272);
or   g1269 (n1290, n843, n850, n1171, n1179);
xnor g1270 (n1313, n1182, n1166, n1277);
xnor g1271 (n1301, n1182, n1178, n1276, n1160);
and  g1272 (n1311, n1169, n1279, n1176, n1164);
nand g1273 (n1305, n844, n1274, n1184, n1167);
or   g1274 (n1293, n1183, n1184, n1165, n1272);
xor  g1275 (n1303, n1274, n1160, n1179, n1174);
xor  g1276 (n1291, n846, n1178, n1184, n1180);
and  g1277 (n1283, n1165, n1272, n1180, n1183);
nor  g1278 (n1317, n1169, n1161, n1273, n1278);
xnor g1279 (n1292, n1176, n1184, n1169, n1164);
nand g1280 (n1289, n1185, n852, n1273, n1275);
and  g1281 (n1284, n1276, n1175, n1173, n1182);
nand g1282 (n1287, n1174, n1180, n1279, n1178);
nand g1283 (n1295, n1173, n1179, n1163, n1168);
xnor g1284 (n1296, n1166, n1170, n1172, n1280);
nand g1285 (n1300, n1178, n1170, n1177, n842);
not  g1286 (n1326, n1220);
not  g1287 (n1345, n864);
buf  g1288 (n1331, n1219);
not  g1289 (n1322, n857);
not  g1290 (n1330, n1224);
not  g1291 (n1343, n859);
buf  g1292 (n1319, n1297);
not  g1293 (n1352, n1191);
not  g1294 (n1341, n858);
buf  g1295 (n1338, n862);
xor  g1296 (n1350, n869, n1218, n1190, n1295);
xor  g1297 (n1332, n1216, n1316, n1318, n1223);
xor  g1298 (n1353, n1216, n1317, n861, n867);
nand g1299 (n1348, n856, n1305, n1292, n1306);
or   g1300 (n1337, n1289, n1217, n1293, n1298);
nand g1301 (n1328, n1284, n1301, n1224, n1223);
or   g1302 (n1324, n1222, n1310, n872, n1217);
nand g1303 (n1329, n1198, n1290, n1197, n1216);
and  g1304 (n1320, n1221, n1303, n865, n1288);
nand g1305 (n1347, n1198, n1221, n1286, n1287);
nor  g1306 (n1321, n1291, n1220, n1314, n1223);
nand g1307 (n1351, n1221, n1218, n1192, n1191);
or   g1308 (n1327, n1224, n1191, n1217, n854);
xor  g1309 (n1325, n853, n1219, n1220, n871);
nand g1310 (n1349, n1307, n1309, n1192, n1294);
or   g1311 (n1339, n1222, n1308, n1313, n1198);
or   g1312 (n1334, n1311, n1190, n1192, n1222);
xnor g1313 (n1335, n1219, n1285, n1197, n1218);
nand g1314 (n1340, n1197, n1220, n1219, n1223);
and  g1315 (n1336, n1315, n1191, n870, n1217);
xnor g1316 (n1346, n1296, n1300, n1197, n1222);
and  g1317 (n1323, n1304, n1190, n1312, n1221);
xnor g1318 (n1344, n1198, n855, n868, n1190);
and  g1319 (n1342, n1302, n860, n1299, n866);
nor  g1320 (n1333, n1216, n1192, n863, n1218);
not  g1321 (n1369, n1342);
buf  g1322 (n1478, n1319);
buf  g1323 (n1396, n1329);
buf  g1324 (n1454, n1349);
buf  g1325 (n1481, n1202);
not  g1326 (n1488, n1332);
buf  g1327 (n1443, n1335);
not  g1328 (n1381, n1333);
not  g1329 (n1492, n1322);
buf  g1330 (n1378, n1350);
not  g1331 (n1382, n1203);
buf  g1332 (n1441, n1348);
buf  g1333 (n1384, n1325);
not  g1334 (n1458, n1204);
buf  g1335 (n1417, n1337);
not  g1336 (n1426, n1352);
not  g1337 (n1372, n879);
not  g1338 (n1422, n1343);
not  g1339 (n1468, n1341);
not  g1340 (n1392, n1200);
buf  g1341 (n1432, n1326);
not  g1342 (n1462, n1208);
not  g1343 (n1425, n1334);
not  g1344 (n1364, n1343);
not  g1345 (n1387, n1326);
buf  g1346 (n1354, n1234);
not  g1347 (n1389, n1348);
buf  g1348 (n1436, n874);
not  g1349 (n1459, n1202);
buf  g1350 (n1471, n1334);
not  g1351 (n1457, n1205);
not  g1352 (n1404, n1346);
not  g1353 (n1439, n1328);
buf  g1354 (n1398, n1332);
not  g1355 (n1376, n1320);
buf  g1356 (n1446, n877);
buf  g1357 (n1435, n1234);
not  g1358 (n1405, n1333);
not  g1359 (n1409, n1204);
not  g1360 (n1423, n1327);
not  g1361 (n1402, n1203);
not  g1362 (n1361, n1340);
not  g1363 (n1368, n1328);
buf  g1364 (n1480, n1323);
buf  g1365 (n1415, n1328);
buf  g1366 (n1479, n1207);
not  g1367 (n1356, n1339);
buf  g1368 (n1453, n1335);
not  g1369 (n1367, n1350);
buf  g1370 (n1430, n1329);
not  g1371 (n1391, n873);
buf  g1372 (n1449, n1342);
not  g1373 (n1493, n1203);
buf  g1374 (n1442, n1325);
not  g1375 (n1450, n1320);
not  g1376 (n1377, n1337);
buf  g1377 (n1489, n1199);
buf  g1378 (n1447, n1326);
not  g1379 (n1456, n1200);
buf  g1380 (n1464, n1338);
buf  g1381 (n1421, n1342);
not  g1382 (n1485, n1330);
not  g1383 (n1401, n1207);
not  g1384 (n1461, n1329);
not  g1385 (n1483, n1349);
buf  g1386 (n1419, n1351);
buf  g1387 (n1357, n1333);
not  g1388 (n1466, n1339);
buf  g1389 (n1487, n1208);
not  g1390 (n1473, n1348);
buf  g1391 (n1491, n1351);
not  g1392 (n1411, n1331);
not  g1393 (n1395, n1322);
buf  g1394 (n1451, n1344);
not  g1395 (n1444, n1343);
buf  g1396 (n1388, n1319);
buf  g1397 (n1375, n1319);
not  g1398 (n1403, n1319);
not  g1399 (n1490, n1341);
buf  g1400 (n1358, n1347);
buf  g1401 (n1379, n1204);
buf  g1402 (n1374, n1206);
buf  g1403 (n1365, n1324);
buf  g1404 (n1460, n1344);
not  g1405 (n1427, n1199);
buf  g1406 (n1418, n1327);
buf  g1407 (n1472, n1207);
not  g1408 (n1400, n1346);
buf  g1409 (n1474, n1328);
not  g1410 (n1465, n1206);
buf  g1411 (n1420, n1199);
buf  g1412 (n1407, n1208);
not  g1413 (n1394, n1323);
buf  g1414 (n1383, n1342);
not  g1415 (n1467, n1331);
buf  g1416 (n1406, n1348);
buf  g1417 (n1385, n1345);
not  g1418 (n1363, n880);
buf  g1419 (n1477, n1321);
buf  g1420 (n1428, n1340);
not  g1421 (n1373, n1343);
not  g1422 (n1455, n1331);
not  g1423 (n1362, n1351);
buf  g1424 (n1360, n1334);
not  g1425 (n1412, n1321);
not  g1426 (n1482, n1345);
buf  g1427 (n1366, n1320);
not  g1428 (n1359, n875);
not  g1429 (n1429, n1321);
buf  g1430 (n1397, n1340);
buf  g1431 (n1414, n1208);
buf  g1432 (n1433, n1335);
buf  g1433 (n1438, n1353);
buf  g1434 (n1486, n1347);
buf  g1435 (n1390, n1201);
buf  g1436 (n1440, n1323);
buf  g1437 (n1476, n1330);
not  g1438 (n1475, n876);
buf  g1439 (n1393, n1346);
buf  g1440 (n1355, n1325);
not  g1441 (n1413, n1331);
buf  g1442 (n1484, n1324);
not  g1443 (n1445, n1350);
xnor g1444 (n1408, n1203, n1353, n1352, n1336);
and  g1445 (n1424, n1349, n1346, n1350, n1207);
or   g1446 (n1410, n1205, n878, n1341, n1333);
nor  g1447 (n1452, n1337, n1201, n1330, n1329);
nand g1448 (n1463, n1327, n1338, n1206, n1325);
or   g1449 (n1416, n1205, n1199, n1339, n1344);
xnor g1450 (n1380, n1347, n1326, n1349, n1200);
nor  g1451 (n1370, n1347, n1324, n1322, n1345);
nand g1452 (n1399, n1336, n1323, n1352);
nand g1453 (n1469, n1335, n1324, n1205, n1353);
nor  g1454 (n1470, n1201, n1336, n1234, n1337);
or   g1455 (n1434, n1327, n1345, n1200, n1338);
xnor g1456 (n1431, n1334, n1202, n1321, n1201);
or   g1457 (n1437, n1332, n1339, n1351, n1330);
and  g1458 (n1371, n1340, n1206, n1332, n1202);
and  g1459 (n1448, n1344, n1204, n1322, n1338);
or   g1460 (n1386, n1320, n1353, n1341, n1336);
nor  g1461 (n1507, n1477, n1471, n1356, n1457);
xor  g1462 (n1542, n1485, n1420, n1465, n1417);
and  g1463 (n1531, n1382, n1408, n1428, n1437);
xor  g1464 (n1509, n1475, n1467, n1483, n1381);
and  g1465 (n1503, n1482, n1479, n1471);
and  g1466 (n1528, n1454, n1471, n1387, n1477);
nor  g1467 (n1512, n1482, n1400, n1446, n1481);
and  g1468 (n1500, n1455, n1479, n1365, n1474);
xnor g1469 (n1549, n1461, n1473, n1484, n1463);
xnor g1470 (n1543, n1467, n1481, n1393, n1465);
nor  g1471 (n1530, n1369, n1454, n1476, n1482);
nand g1472 (n1535, n1481, n1448, n1378, n1380);
nor  g1473 (n1518, n1484, n1360, n1433, n1460);
xnor g1474 (n1495, n1383, n1462, n1469, n1441);
nor  g1475 (n1519, n1456, n1462, n1464, n1454);
nand g1476 (n1504, n1462, n1459, n1480, n1391);
xor  g1477 (n1501, n1478, n1466, n1421, n1480);
xor  g1478 (n1541, n1439, n1458, n1447, n1457);
xor  g1479 (n1553, n1410, n1452, n1416, n1389);
and  g1480 (n1521, n1469, n1398, n1463, n1375);
nor  g1481 (n1525, n1458, n1481, n1396, n1355);
xnor g1482 (n1497, n1468, n1411, n1451, n1404);
and  g1483 (n1502, n1440, n1461, n1443, n1464);
xor  g1484 (n1533, n1419, n1476, n1403, n1453);
nor  g1485 (n1547, n1478, n1465, n1413, n1429);
xnor g1486 (n1494, n1395, n1459, n1461, n1474);
nor  g1487 (n1498, n1422, n1485, n1470, n1388);
xor  g1488 (n1550, n1483, n1452, n1470, n1468);
and  g1489 (n1536, n1392, n1485, n1480, n1478);
xnor g1490 (n1524, n1480, n1465, n1450, n1386);
or   g1491 (n1505, n1409, n1401, n1357, n1371);
xnor g1492 (n1508, n1370, n1462, n1423, n1459);
nor  g1493 (n1551, n1384, n1427, n1374, n1377);
nor  g1494 (n1522, n1469, n1354, n1451, n1459);
and  g1495 (n1539, n1476, n1484, n1367, n1466);
nand g1496 (n1496, n1451, n1452, n1412, n1463);
or   g1497 (n1516, n1452, n1442, n1464, n1456);
xnor g1498 (n1548, n1364, n1456, n1372, n1397);
xnor g1499 (n1529, n1362, n1468, n1373, n1406);
xnor g1500 (n1520, n1478, n883, n881, n1477);
and  g1501 (n1540, n1455, n1475, n1483, n1471);
and  g1502 (n1511, n1477, n1385, n1468, n1460);
and  g1503 (n1526, n1472, n1424, n1361, n1425);
and  g1504 (n1515, n1405, n1484, n1457, n1464);
nand g1505 (n1513, n882, n1358, n1458, n1407);
xor  g1506 (n1510, n1466, n1472, n1457, n1453);
nor  g1507 (n1517, n1432, n1479, n1418, n1473);
and  g1508 (n1499, n1467, n1444, n1454, n1430);
nand g1509 (n1527, n1460, n1473, n1470, n1366);
and  g1510 (n1537, n884, n1453, n1475, n1460);
and  g1511 (n1534, n1456, n1453, n1445, n1467);
nor  g1512 (n1545, n1472, n1402, n1455, n1390);
nand g1513 (n1523, n1476, n1414, n1475, n1359);
or   g1514 (n1544, n1451, n1394, n1431, n1469);
or   g1515 (n1546, n1473, n1438, n1483, n1472);
xor  g1516 (n1514, n1435, n1470, n1426, n1379);
and  g1517 (n1506, n1363, n1482, n1463, n1399);
or   g1518 (n1538, n1368, n1415, n1376, n1449);
xnor g1519 (n1552, n1458, n1466, n1434, n1474);
xor  g1520 (n1532, n1455, n1461, n1436, n1474);
nor  g1521 (n1570, n936, n1514, n1498, n961);
nor  g1522 (n1564, n1003, n1043, n1053, n1540);
and  g1523 (n1590, n1007, n891, n972, n1529);
nand g1524 (n1565, n963, n1523, n1046, n986);
nor  g1525 (n1578, n1517, n1526, n956, n1009);
and  g1526 (n1585, n1035, n994, n1503, n920);
or   g1527 (n1609, n895, n924, n1023, n1056);
nand g1528 (n1596, n1064, n1020, n903, n1021);
and  g1529 (n1602, n1025, n1525, n1028, n966);
xor  g1530 (n1586, n915, n942, n1551, n983);
or   g1531 (n1581, n1001, n887, n989, n1022);
or   g1532 (n1613, n997, n1041, n974, n907);
xnor g1533 (n1580, n968, n999, n967, n1058);
and  g1534 (n1587, n978, n950, n925, n1524);
or   g1535 (n1600, n1061, n933, n1005, n1018);
or   g1536 (n1577, n944, n943, n976, n1539);
and  g1537 (n1604, n1063, n1004, n977, n1033);
nand g1538 (n1594, n1553, n1049, n1530, n1037);
or   g1539 (n1569, n1002, n906, n1510, n1507);
nor  g1540 (n1589, n1537, n905, n938, n1062);
xor  g1541 (n1601, n1031, n1532, n888, n1533);
nor  g1542 (n1595, n1014, n1511, n991, n995);
xor  g1543 (n1608, n953, n1057, n1546, n975);
and  g1544 (n1572, n945, n1547, n921, n929);
and  g1545 (n1582, n984, n1522, n1505, n1029);
xnor g1546 (n1605, n1535, n1036, n982, n939);
nand g1547 (n1611, n960, n912, n1052, n1051);
and  g1548 (n1566, n1059, n1518, n987, n970);
xnor g1549 (n1562, n1030, n914, n934, n940);
xnor g1550 (n1554, n1048, n1015, n1013, n898);
nor  g1551 (n1558, n901, n1548, n1543, n1000);
xor  g1552 (n1559, n1550, n1012, n958, n904);
nor  g1553 (n1603, n1509, n1545, n969, n1496);
xnor g1554 (n1591, n957, n1516, n1027, n1527);
xor  g1555 (n1557, n1008, n955, n896, n998);
nor  g1556 (n1599, n910, n949, n892, n1050);
or   g1557 (n1598, n885, n911, n980, n1011);
or   g1558 (n1593, n1513, n1047, n981, n1506);
nand g1559 (n1556, n922, n1040, n1017, n897);
and  g1560 (n1588, n935, n1552, n1042, n923);
and  g1561 (n1575, n952, n959, n1494, n941);
nor  g1562 (n1561, n894, n899, n1054, n1034);
or   g1563 (n1560, n1536, n919, n909, n926);
and  g1564 (n1584, n979, n1541, n930, n985);
and  g1565 (n1563, n947, n954, n916, n908);
nand g1566 (n1573, n946, n951, n900, n1010);
nand g1567 (n1597, n993, n992, n917, n1534);
or   g1568 (n1610, n893, n1519, n1060, n1499);
nor  g1569 (n1571, n1500, n1026, n1495, n1508);
or   g1570 (n1606, n971, n902, n1512, n918);
nand g1571 (n1607, n1039, n937, n1504, n965);
xor  g1572 (n1576, n988, n1549, n962, n1016);
and  g1573 (n1612, n1024, n1045, n948, n1528);
nor  g1574 (n1592, n964, n890, n996, n931);
nand g1575 (n1583, n913, n889, n1542, n1544);
and  g1576 (n1579, n932, n1038, n1006, n928);
xnor g1577 (n1574, n1501, n927, n1538, n1055);
nand g1578 (n1568, n886, n1520, n1515, n1032);
or   g1579 (n1555, n990, n1497, n1521, n1531);
nand g1580 (n1567, n973, n1044, n1502, n1019);
not  g1581 (n1614, n1554);
not  g1582 (n1615, n1554);
not  g1583 (n1618, n1555);
buf  g1584 (n1616, n1555);
not  g1585 (n1617, n1554);
not  g1586 (n1619, n1555);
nand g1587 (n1621, n1615, n1614);
nand g1588 (n1620, n1068, n1067, n1065, n1066);
xor  g1589 (n1624, n1487, n1488, n1621);
and  g1590 (n1622, n1486, n1069, n1488, n1070);
nor  g1591 (n1623, n1071, n1486, n1621);
nand g1592 (n1626, n1485, n1620, n1487);
or   g1593 (n1625, n1487, n1486, n1621);
and  g1594 (n1628, n1488, n1489, n1625);
xor  g1595 (n1629, n1557, n1556, n1622, n1625);
xnor g1596 (n1631, n1559, n1489, n1072);
and  g1597 (n1632, n1558, n1490, n1557);
nand g1598 (n1630, n1556, n1624, n1558, n1559);
xnor g1599 (n1627, n1558, n1623, n1556, n1489);
not  g1600 (n1636, n1629);
buf  g1601 (n1635, n1630);
not  g1602 (n1633, n1631);
not  g1603 (n1634, n1632);
not  g1604 (n1644, n1562);
not  g1605 (n1649, n1565);
xnor g1606 (n1648, n1633, n1635, n1636);
xnor g1607 (n1641, n1636, n1564);
xor  g1608 (n1652, n1559, n1635, n1561);
or   g1609 (n1639, n1635, n1636, n1634);
and  g1610 (n1651, n1563, n1079, n1633);
nor  g1611 (n1650, n1074, n1636, n1633);
xnor g1612 (n1640, n1565, n1633, n1563);
xor  g1613 (n1646, n1561, n1560, n1073);
xor  g1614 (n1643, n1565, n1563, n1566);
nor  g1615 (n1642, n1561, n1566, n1635);
xor  g1616 (n1647, n1075, n1564, n1634);
and  g1617 (n1645, n1562, n1078, n1560);
xnor g1618 (n1638, n1077, n1076, n1634);
and  g1619 (n1637, n1634, n1560, n1562);
or   g1620 (n1679, n1083, n1589, n1601, n1580);
and  g1621 (n1673, n1596, n1649, n1092, n1094);
or   g1622 (n1664, n1603, n1573, n1604, n1585);
nand g1623 (n1714, n1648, n1586, n1651, n1570);
or   g1624 (n1666, n1640, n1082, n1597, n1603);
or   g1625 (n1700, n1099, n1640, n1107, n1573);
nand g1626 (n1676, n1603, n1592, n1602, n1589);
or   g1627 (n1702, n1578, n1593, n1091, n1597);
and  g1628 (n1672, n1603, n1606, n1576, n1588);
xor  g1629 (n1705, n1651, n1588, n1568, n1605);
nand g1630 (n1697, n1594, n1590, n1575, n1647);
and  g1631 (n1683, n1641, n1577, n1637, n1604);
xnor g1632 (n1707, n1602, n1644, n1638, n1597);
xnor g1633 (n1656, n1574, n1584, n1582, n1093);
nor  g1634 (n1665, n1652, n1578, n1596, n1575);
or   g1635 (n1694, n1106, n1583, n1080);
or   g1636 (n1709, n1581, n1582, n1602, n1650);
nand g1637 (n1701, n1637, n1648, n1575, n1573);
and  g1638 (n1660, n1651, n1111, n1604, n1590);
or   g1639 (n1692, n1595, n1085, n1590, n1638);
nor  g1640 (n1661, n1642, n1644, n1605, n1084);
nor  g1641 (n1653, n1569, n1645, n1646, n1591);
nor  g1642 (n1713, n1607, n1589, n1643, n1582);
and  g1643 (n1657, n1586, n1579, n1602, n1641);
nand g1644 (n1659, n1576, n1607, n1572, n1645);
and  g1645 (n1698, n1647, n1647, n1640, n1593);
xor  g1646 (n1655, n1587, n1648, n1577, n1567);
xor  g1647 (n1685, n1637, n1579, n1598, n1597);
and  g1648 (n1677, n1606, n1585, n1646, n1095);
xor  g1649 (n1704, n1638, n1594, n1096, n1604);
or   g1650 (n1708, n1574, n1605, n1579, n1583);
nor  g1651 (n1671, n1581, n1650, n1593, n1585);
or   g1652 (n1690, n1648, n1571, n1570, n1105);
or   g1653 (n1706, n1588, n1599, n1586, n1598);
nand g1654 (n1662, n1598, n1600, n1109, n1086);
nand g1655 (n1658, n1600, n1581, n1641, n1587);
xnor g1656 (n1682, n1592, n1576, n1601, n1586);
xor  g1657 (n1691, n1577, n1577, n1608, n1580);
nand g1658 (n1696, n1584, n1583, n1573, n1643);
xnor g1659 (n1675, n1569, n1642, n1578, n1566);
xor  g1660 (n1670, n1580, n1088, n1102, n1637);
xnor g1661 (n1716, n1576, n1579, n1596, n1584);
or   g1662 (n1703, n1645, n1600, n1601, n1640);
xor  g1663 (n1681, n1568, n1599, n1638, n1607);
or   g1664 (n1654, n1108, n1584, n1639, n1101);
and  g1665 (n1678, n1081, n1642, n1649, n1646);
and  g1666 (n1688, n1595, n1568, n1574, n1592);
xor  g1667 (n1684, n1601, n1599, n1587, n1591);
nand g1668 (n1687, n1591, n1581, n1585, n1652);
xnor g1669 (n1667, n1651, n1639, n1649, n1643);
or   g1670 (n1686, n1650, n1595, n1592, n1090);
nor  g1671 (n1693, n1571, n1575, n1605, n1607);
nor  g1672 (n1695, n1087, n1098, n1650, n1110);
and  g1673 (n1663, n1646, n1644, n1594, n1580);
or   g1674 (n1715, n1643, n1606, n1572, n1644);
xor  g1675 (n1689, n1594, n1591, n1578, n1649);
xor  g1676 (n1699, n1582, n1089, n1103, n1645);
xnor g1677 (n1674, n1642, n1639, n1567, n1593);
xor  g1678 (n1668, n1590, n1639, n1567, n1606);
and  g1679 (n1711, n1588, n1599, n1647, n1652);
and  g1680 (n1712, n1569, n1652, n1587, n1574);
xor  g1681 (n1680, n1598, n1641, n1600, n1097);
xor  g1682 (n1669, n1100, n1104, n1572, n1596);
xor  g1683 (n1710, n1571, n1589, n1595, n1570);
nor  g1684 (n1719, n1117, n1112, n1116, n1119);
nor  g1685 (n1720, n671, n1115, n1653, n1118);
nand g1686 (n1717, n671, n671, n1653, n1113);
and  g1687 (n1718, n1653, n1653, n671, n1114);
not  g1688 (n1725, n1120);
buf  g1689 (n1721, n1719);
not  g1690 (n1723, n1719);
not  g1691 (n1724, n1122);
nor  g1692 (n1722, n1717, n1718, n1719, n1121);
xor  g1693 (n1734, n1129, n1132, n1130, n1491);
xor  g1694 (n1730, n1127, n1138, n1133, n1721);
nor  g1695 (n1733, n1721, n1721, n1722, n1128);
and  g1696 (n1729, n1136, n1125, n1491, n1137);
xor  g1697 (n1726, n1722, n1140, n1723, n1131);
or   g1698 (n1727, n1722, n1141, n1723, n1491);
or   g1699 (n1731, n1123, n1135, n1491, n1134);
xnor g1700 (n1732, n1723, n1490, n1139);
or   g1701 (n1728, n1126, n1124, n1490, n1142);
not  g1702 (n1737, n1734);
buf  g1703 (n1735, n1733);
buf  g1704 (n1736, n1732);
not  g1705 (n1744, n1609);
buf  g1706 (n1740, n1609);
buf  g1707 (n1748, n1737);
not  g1708 (n1746, n1608);
buf  g1709 (n1743, n1735);
not  g1710 (n1739, n1736);
buf  g1711 (n1741, n1737);
not  g1712 (n1747, n1737);
or   g1713 (n1738, n1737, n1736);
xnor g1714 (n1745, n1609, n1735, n1736);
xnor g1715 (n1742, n1735, n1608, n1609);
buf  g1716 (n1752, n1738);
not  g1717 (n1782, n1745);
not  g1718 (n1788, n1740);
not  g1719 (n1762, n1741);
not  g1720 (n1777, n1747);
buf  g1721 (n1787, n1611);
not  g1722 (n1757, n1748);
buf  g1723 (n1756, n1741);
not  g1724 (n1761, n1739);
not  g1725 (n1790, n1742);
buf  g1726 (n1759, n1743);
not  g1727 (n1792, n1619);
not  g1728 (n1755, n1744);
buf  g1729 (n1763, n1720);
not  g1730 (n1766, n1746);
buf  g1731 (n1758, n1147);
buf  g1732 (n1778, n1618);
not  g1733 (n1754, n1740);
buf  g1734 (n1750, n1739);
buf  g1735 (n1783, n1740);
buf  g1736 (n1780, n1611);
not  g1737 (n1770, n1748);
buf  g1738 (n1776, n1720);
buf  g1739 (n1753, n1617);
not  g1740 (n1779, n1618);
not  g1741 (n1785, n1719);
not  g1742 (n1784, n1745);
not  g1743 (n1769, n1617);
buf  g1744 (n1771, n1742);
buf  g1745 (n1767, n1224);
not  g1746 (n1774, n1746);
buf  g1747 (n1760, n1617);
buf  g1748 (n1764, n1145);
nand g1749 (n1775, n1619, n1611, n1740, n1744);
or   g1750 (n1791, n1738, n1748, n1619, n1745);
or   g1751 (n1781, n1747, n1616, n1742);
nor  g1752 (n1786, n1748, n1741, n1738);
and  g1753 (n1772, n1610, n1144, n1720);
and  g1754 (n1789, n1146, n1747, n1739);
and  g1755 (n1749, n1617, n1618, n1610, n1612);
or   g1756 (n1765, n1744, n1610, n1618);
nor  g1757 (n1768, n1741, n1743, n1747, n1143);
nand g1758 (n1751, n1745, n1611, n1743, n1746);
xnor g1759 (n1773, n1743, n1619, n1746, n1744);
buf  g1760 (n1931, n1667);
buf  g1761 (n1810, n1789);
buf  g1762 (n1862, n1713);
not  g1763 (n1905, n1681);
buf  g1764 (n1849, n1711);
buf  g1765 (n1897, n1755);
buf  g1766 (n1963, n1697);
not  g1767 (n1929, n1707);
not  g1768 (n1887, n1708);
buf  g1769 (n1815, n1763);
not  g1770 (n1816, n1751);
not  g1771 (n1855, n1771);
not  g1772 (n1911, n1659);
not  g1773 (n1818, n1685);
not  g1774 (n1966, n1692);
not  g1775 (n1962, n1783);
not  g1776 (n1960, n1671);
not  g1777 (n1872, n1768);
not  g1778 (n1885, n1772);
not  g1779 (n1893, n1782);
not  g1780 (n1842, n1715);
buf  g1781 (n1965, n1707);
buf  g1782 (n1813, n1699);
not  g1783 (n1941, n1788);
buf  g1784 (n1899, n1672);
not  g1785 (n1914, n1678);
buf  g1786 (n1826, n1693);
buf  g1787 (n1809, n1705);
not  g1788 (n1841, n1779);
buf  g1789 (n1950, n1664);
buf  g1790 (n1793, n1666);
not  g1791 (n1945, n1791);
buf  g1792 (n1891, n1664);
not  g1793 (n1860, n1758);
not  g1794 (n1829, n1787);
buf  g1795 (n1835, n1704);
not  g1796 (n1875, n1687);
buf  g1797 (n1877, n1699);
not  g1798 (n1811, n1750);
not  g1799 (n1854, n1688);
buf  g1800 (n1820, n1686);
not  g1801 (n1902, n1709);
not  g1802 (n1932, n1691);
buf  g1803 (n1967, n1701);
and  g1804 (n1853, n1762, n1710, n1770);
and  g1805 (n1928, n1762, n1781, n1773);
and  g1806 (n1817, n1692, n1662, n1788);
nand g1807 (n1839, n1787, n1683, n1781);
nor  g1808 (n1830, n1688, n1772, n1686);
and  g1809 (n1852, n1782, n1664, n1694);
or   g1810 (n1868, n1704, n1684, n1698);
and  g1811 (n1884, n1707, n1776, n1706);
xor  g1812 (n1900, n1754, n1760, n1680);
xor  g1813 (n1947, n1783, n1689, n1765);
xor  g1814 (n1863, n1666, n1764, n1781);
xor  g1815 (n1892, n1701, n1791, n1694);
xor  g1816 (n1903, n1659, n1675, n1750);
xor  g1817 (n1861, n1779, n1682, n1690);
and  g1818 (n1926, n1752, n1708, n1785);
and  g1819 (n1883, n1760, n1675, n1702);
xnor g1820 (n1959, n1674, n1774, n1758);
xor  g1821 (n1922, n1688, n1710, n1775);
and  g1822 (n1869, n1711, n1792, n1702);
xnor g1823 (n1857, n1788, n1753, n1700);
xnor g1824 (n1888, n1753, n1780, n1673);
xnor g1825 (n1848, n1683, n1763, n1660);
xor  g1826 (n1951, n1668, n1655, n1787);
nor  g1827 (n1890, n1781, n1712, n1703);
nand g1828 (n1954, n1661, n1752, n1712);
nand g1829 (n1867, n1666, n1701, n1613);
xnor g1830 (n1808, n1783, n1669, n1788);
xor  g1831 (n1968, n1612, n1792, n1148);
nand g1832 (n1904, n1766, n1775, n1703);
nor  g1833 (n1834, n1670, n1752, n1656);
nand g1834 (n1805, n1762, n1772, n1716);
or   g1835 (n1844, n1701, n1724, n1751);
xor  g1836 (n1946, n1776, n1714, n1778);
and  g1837 (n1843, n1686, n1663, n1786);
nor  g1838 (n1798, n1765, n1761, n1776);
and  g1839 (n1851, n1690, n1784, n1791);
and  g1840 (n1803, n1764, n1714, n1660);
nor  g1841 (n1889, n1612, n1679, n1697);
xnor g1842 (n1952, n1689, n1671, n1774);
xnor g1843 (n1832, n1785, n1777, n1656);
xor  g1844 (n1801, n1666, n1712, n1658);
xnor g1845 (n1920, n1790, n1673, n1677);
and  g1846 (n1964, n1749, n1757, n1695);
and  g1847 (n1870, n1670, n1749, n1716);
xor  g1848 (n1955, n1749, n1770, n1774);
nand g1849 (n1910, n1775, n1773, n1768);
and  g1850 (n1824, n1715, n1789, n1655);
xnor g1851 (n1876, n1708, n1784, n1673);
or   g1852 (n1953, n1770, n1703, n1672);
xor  g1853 (n1925, n1754, n1668, n1792);
nand g1854 (n1794, n1790, n1756, n1706);
xor  g1855 (n1819, n1673, n1782, n1674);
xor  g1856 (n1938, n1674, n1682, n1709);
nor  g1857 (n1838, n1683, n1755, n1657);
or   g1858 (n1865, n1676, n1675, n1757);
and  g1859 (n1896, n1678, n1716, n1657);
xnor g1860 (n1812, n1697, n1689, n1657);
nand g1861 (n1907, n1769, n1713, n1693);
or   g1862 (n1921, n1703, n1660, n1612);
xor  g1863 (n1912, n1663, n1761, n1709);
xnor g1864 (n1961, n1789, n1659, n1755);
xnor g1865 (n1934, n1658, n1696, n1665);
nand g1866 (n1800, n1695, n1674, n1764);
xor  g1867 (n1933, n1711, n1762, n1778);
xor  g1868 (n1825, n1780, n1710, n1685);
nand g1869 (n1847, n1702, n1773, n1686);
xnor g1870 (n1942, n1769, n1713, n1613);
nand g1871 (n1856, n1661, n1699, n1668);
or   g1872 (n1827, n1785, n1661, n1696);
or   g1873 (n1886, n1695, n1765, n1769);
nor  g1874 (n1799, n1777, n1694, n1778);
xor  g1875 (n1878, n1668, n1676, n1671);
xor  g1876 (n1837, n1663, n1770, n1658);
xor  g1877 (n1958, n1667, n1789, n1763);
nand g1878 (n1822, n1684, n1680, n1786);
nor  g1879 (n1831, n1723, n1714, n1774);
and  g1880 (n1802, n1754, n1709, n1759);
nand g1881 (n1845, n1669, n1694, n1711);
xor  g1882 (n1919, n1681, n1779, n1698);
xor  g1883 (n1898, n1784, n1654, n1669);
nor  g1884 (n1858, n1769, n1777, n1677);
nand g1885 (n1930, n1695, n1767, n1751);
xnor g1886 (n1956, n1780, n1613, n1680);
xnor g1887 (n1821, n1782, n1792, n1707);
nand g1888 (n1901, n1713, n1767, n1784);
nand g1889 (n1871, n1676, n1786, n1679);
nand g1890 (n1939, n1693, n1771, n1678);
xor  g1891 (n1949, n1724, n1698, n1760);
and  g1892 (n1795, n1702, n1654, n1750);
xnor g1893 (n1948, n1776, n1691, n1700);
and  g1894 (n1906, n1700, n1661, n1766);
xnor g1895 (n1895, n1751, n1753, n1691);
nor  g1896 (n1796, n1706, n1791, n1665);
xnor g1897 (n1807, n1787, n1750, n1670);
nand g1898 (n1944, n1757, n1691, n1786);
and  g1899 (n1916, n1760, n1671, n1756);
or   g1900 (n1806, n1757, n1783, n1761);
nor  g1901 (n1927, n1714, n1659, n1654);
nand g1902 (n1866, n1687, n1705, n1716);
or   g1903 (n1859, n1696, n1692, n1685);
nand g1904 (n1850, n1665, n1753, n1756);
xnor g1905 (n1874, n1715, n1758, n1712);
nand g1906 (n1909, n1778, n1682, n1658);
and  g1907 (n1836, n1676, n1660, n1677);
and  g1908 (n1882, n1785, n1767, n1681);
xor  g1909 (n1957, n1662, n1667);
or   g1910 (n1833, n1767, n1690, n1699);
xor  g1911 (n1924, n1715, n1775, n1662);
xor  g1912 (n1894, n1749, n1790);
xnor g1913 (n1915, n1679, n1759, n1780);
or   g1914 (n1923, n1685, n1779, n1687);
nand g1915 (n1828, n1698, n1677, n1655);
nor  g1916 (n1913, n1706, n1613, n1678);
nor  g1917 (n1797, n1773, n1768, n1697);
xnor g1918 (n1940, n1708, n1684, n1766);
nand g1919 (n1823, n1656, n1681, n1696);
xor  g1920 (n1814, n1690, n1704, n1777);
nor  g1921 (n1846, n1756, n1755, n1692);
or   g1922 (n1873, n1705, n1670, n1672);
and  g1923 (n1943, n1663, n1705, n1758);
and  g1924 (n1936, n1662, n1669, n1656);
and  g1925 (n1917, n1684, n1700, n1664);
and  g1926 (n1864, n1752, n1693, n1704);
xnor g1927 (n1937, n1680, n1771, n1724);
xor  g1928 (n1918, n1710, n1761, n1768);
xor  g1929 (n1880, n1689, n1759, n1672);
and  g1930 (n1935, n1771, n1763, n1765);
and  g1931 (n1804, n1654, n1683, n1766);
xor  g1932 (n1881, n1682, n1688, n1679);
and  g1933 (n1908, n1687, n1764, n1759);
nand g1934 (n1840, n1754, n1655, n1657);
and  g1935 (n1879, n1665, n1772, n1675);
buf  g1936 (n2392, n1917);
not  g1937 (n2365, n1852);
not  g1938 (n2252, n1957);
not  g1939 (n2481, n1913);
buf  g1940 (n2218, n1866);
not  g1941 (n2595, n1827);
not  g1942 (n1994, n1890);
buf  g1943 (n2107, n1865);
not  g1944 (n2568, n1919);
not  g1945 (n2228, n1836);
buf  g1946 (n2339, n1909);
not  g1947 (n2317, n1888);
not  g1948 (n2634, n1899);
buf  g1949 (n2198, n1811);
not  g1950 (n2533, n1955);
buf  g1951 (n2180, n1914);
buf  g1952 (n2214, n1901);
buf  g1953 (n2665, n1861);
not  g1954 (n2263, n1824);
buf  g1955 (n2261, n1885);
buf  g1956 (n2462, n1916);
buf  g1957 (n2189, n1921);
buf  g1958 (n2213, n1892);
buf  g1959 (n2201, n1830);
not  g1960 (n2331, n1898);
not  g1961 (n2642, n1809);
buf  g1962 (n2325, n1887);
buf  g1963 (n2227, n1943);
buf  g1964 (n2540, n1796);
not  g1965 (n2357, n1949);
buf  g1966 (n2610, n1845);
buf  g1967 (n2211, n1838);
not  g1968 (n2465, n1870);
not  g1969 (n2097, n1894);
not  g1970 (n1975, n1893);
not  g1971 (n2284, n1948);
not  g1972 (n2262, n1937);
buf  g1973 (n2271, n1834);
not  g1974 (n2329, n1842);
buf  g1975 (n2453, n1887);
buf  g1976 (n2618, n1968);
buf  g1977 (n2447, n1880);
not  g1978 (n2008, n1834);
buf  g1979 (n2327, n1919);
not  g1980 (n2583, n1926);
buf  g1981 (n2323, n1821);
not  g1982 (n2353, n1871);
not  g1983 (n2613, n1872);
buf  g1984 (n2435, n1855);
not  g1985 (n1971, n1859);
buf  g1986 (n2506, n1827);
buf  g1987 (n2174, n1874);
buf  g1988 (n2575, n1840);
buf  g1989 (n2140, n1949);
not  g1990 (n2059, n1885);
buf  g1991 (n2159, n1918);
not  g1992 (n2643, n1844);
buf  g1993 (n2494, n1831);
not  g1994 (n2298, n1903);
buf  g1995 (n2579, n1869);
not  g1996 (n2199, n1821);
not  g1997 (n1997, n1799);
not  g1998 (n2443, n1905);
not  g1999 (n1989, n1844);
buf  g2000 (n2585, n1808);
buf  g2001 (n2376, n1893);
buf  g2002 (n2032, n1927);
buf  g2003 (n2235, n1958);
buf  g2004 (n2286, n1942);
not  g2005 (n2086, n1923);
not  g2006 (n2369, n1873);
not  g2007 (n2248, n1941);
not  g2008 (n2429, n1838);
not  g2009 (n2398, n1833);
buf  g2010 (n2547, n1962);
buf  g2011 (n2525, n1833);
not  g2012 (n2310, n1950);
not  g2013 (n2204, n1797);
buf  g2014 (n2270, n1947);
not  g2015 (n2153, n1940);
not  g2016 (n2608, n1799);
not  g2017 (n2596, n1801);
not  g2018 (n2394, n1828);
not  g2019 (n2428, n1825);
buf  g2020 (n2015, n1810);
not  g2021 (n2431, n1807);
buf  g2022 (n2217, n1875);
buf  g2023 (n2469, n1945);
buf  g2024 (n2129, n1806);
not  g2025 (n2282, n1872);
not  g2026 (n2010, n1799);
not  g2027 (n2170, n1919);
not  g2028 (n2126, n1859);
buf  g2029 (n2434, n1911);
buf  g2030 (n2114, n1918);
not  g2031 (n2108, n1857);
not  g2032 (n2389, n1868);
not  g2033 (n2444, n1919);
buf  g2034 (n2076, n1866);
buf  g2035 (n2621, n1954);
not  g2036 (n2121, n1909);
not  g2037 (n1974, n1938);
buf  g2038 (n2515, n1853);
not  g2039 (n2315, n1946);
buf  g2040 (n2073, n1895);
buf  g2041 (n2337, n1881);
buf  g2042 (n2000, n1817);
not  g2043 (n2512, n1815);
not  g2044 (n2498, n1917);
not  g2045 (n2130, n1891);
not  g2046 (n2401, n1801);
buf  g2047 (n2638, n1798);
buf  g2048 (n2106, n1856);
buf  g2049 (n2313, n1945);
buf  g2050 (n2532, n1937);
buf  g2051 (n2002, n1915);
buf  g2052 (n2251, n1899);
buf  g2053 (n2667, n1841);
buf  g2054 (n2306, n1800);
buf  g2055 (n2240, n1909);
not  g2056 (n2562, n1877);
not  g2057 (n2203, n1888);
not  g2058 (n2524, n1830);
buf  g2059 (n2105, n1802);
buf  g2060 (n2028, n1802);
buf  g2061 (n2060, n1965);
not  g2062 (n2499, n1797);
buf  g2063 (n2332, n1928);
buf  g2064 (n2517, n1884);
buf  g2065 (n2082, n1921);
not  g2066 (n2290, n1966);
not  g2067 (n2619, n1800);
buf  g2068 (n1991, n1888);
buf  g2069 (n2661, n1839);
buf  g2070 (n2034, n1808);
buf  g2071 (n2652, n1929);
not  g2072 (n2529, n1957);
buf  g2073 (n2183, n1914);
buf  g2074 (n2446, n1941);
not  g2075 (n2190, n1899);
not  g2076 (n2078, n1796);
not  g2077 (n2171, n1924);
buf  g2078 (n2182, n1880);
buf  g2079 (n2336, n1895);
not  g2080 (n2662, n1825);
buf  g2081 (n2287, n1885);
not  g2082 (n2479, n1942);
not  g2083 (n2194, n1837);
buf  g2084 (n2269, n1841);
not  g2085 (n2496, n1920);
not  g2086 (n2119, n1266);
buf  g2087 (n2388, n1842);
buf  g2088 (n2425, n1950);
not  g2089 (n2344, n1820);
buf  g2090 (n2226, n1856);
buf  g2091 (n2048, n1946);
not  g2092 (n2186, n1826);
not  g2093 (n2391, n1943);
buf  g2094 (n2403, n1936);
not  g2095 (n2314, n1906);
not  g2096 (n2449, n1913);
not  g2097 (n1992, n1878);
not  g2098 (n1990, n1815);
buf  g2099 (n2501, n1889);
not  g2100 (n2188, n1860);
not  g2101 (n2589, n1831);
not  g2102 (n2197, n1946);
not  g2103 (n2224, n1879);
buf  g2104 (n2022, n1874);
buf  g2105 (n2592, n1951);
not  g2106 (n2253, n1804);
not  g2107 (n2648, n1814);
not  g2108 (n2301, n1818);
not  g2109 (n1996, n1884);
not  g2110 (n2626, n1960);
buf  g2111 (n2143, n1925);
buf  g2112 (n2483, n1795);
buf  g2113 (n2548, n1886);
not  g2114 (n2320, n1848);
buf  g2115 (n2658, n1915);
not  g2116 (n2164, n1886);
buf  g2117 (n2138, n1865);
not  g2118 (n2461, n1891);
buf  g2119 (n2635, n1806);
not  g2120 (n2509, n1822);
not  g2121 (n2244, n1820);
not  g2122 (n2422, n1805);
buf  g2123 (n2536, n1795);
not  g2124 (n2233, n1877);
buf  g2125 (n2399, n1843);
buf  g2126 (n2531, n1798);
buf  g2127 (n2307, n1877);
not  g2128 (n1982, n1937);
not  g2129 (n2590, n1823);
not  g2130 (n2013, n1794);
buf  g2131 (n2406, n1915);
not  g2132 (n2081, n1847);
buf  g2133 (n2045, n1854);
not  g2134 (n2036, n1818);
buf  g2135 (n2205, n1848);
not  g2136 (n2497, n1947);
buf  g2137 (n2463, n1796);
not  g2138 (n2448, n1905);
not  g2139 (n2510, n1967);
not  g2140 (n2354, n1840);
not  g2141 (n2003, n1492);
not  g2142 (n2131, n1955);
buf  g2143 (n2351, n1918);
buf  g2144 (n2322, n1886);
not  g2145 (n2393, n1842);
buf  g2146 (n2451, n1957);
buf  g2147 (n2311, n1911);
not  g2148 (n2571, n1894);
not  g2149 (n2220, n1962);
buf  g2150 (n2330, n1848);
not  g2151 (n2324, n1493);
buf  g2152 (n2419, n1810);
buf  g2153 (n2192, n1964);
not  g2154 (n2124, n1819);
not  g2155 (n2424, n1959);
buf  g2156 (n2272, n1817);
not  g2157 (n2390, n1827);
not  g2158 (n2578, n1813);
not  g2159 (n2472, n1965);
not  g2160 (n2454, n1897);
buf  g2161 (n2297, n1862);
buf  g2162 (n2241, n1871);
not  g2163 (n2305, n1149);
buf  g2164 (n2614, n1836);
not  g2165 (n2110, n1837);
buf  g2166 (n2551, n1860);
buf  g2167 (n2576, n1832);
buf  g2168 (n2360, n1940);
buf  g2169 (n2041, n1859);
not  g2170 (n2407, n1831);
not  g2171 (n2413, n1942);
buf  g2172 (n2522, n1887);
buf  g2173 (n2649, n1626);
not  g2174 (n2377, n1860);
buf  g2175 (n1972, n1912);
not  g2176 (n2574, n1855);
buf  g2177 (n2066, n1816);
not  g2178 (n2542, n1920);
buf  g2179 (n2484, n1902);
buf  g2180 (n2582, n1961);
not  g2181 (n1999, n1869);
not  g2182 (n2474, n1881);
not  g2183 (n2264, n1904);
not  g2184 (n2061, n1906);
buf  g2185 (n2385, n1806);
not  g2186 (n2116, n1807);
buf  g2187 (n2599, n1872);
buf  g2188 (n2437, n1879);
buf  g2189 (n2663, n1928);
buf  g2190 (n2641, n1915);
buf  g2191 (n2176, n1893);
not  g2192 (n2538, n1807);
not  g2193 (n2489, n1829);
buf  g2194 (n2096, n1799);
not  g2195 (n1979, n1819);
buf  g2196 (n2230, n1922);
not  g2197 (n2523, n1934);
buf  g2198 (n2260, n1821);
not  g2199 (n2257, n1800);
not  g2200 (n2659, n1883);
not  g2201 (n2294, n1871);
buf  g2202 (n2504, n1893);
buf  g2203 (n2633, n1929);
not  g2204 (n2379, n1880);
buf  g2205 (n1986, n1831);
not  g2206 (n2612, n1876);
not  g2207 (n2668, n1923);
buf  g2208 (n2242, n1910);
buf  g2209 (n2346, n1825);
not  g2210 (n2070, n1843);
buf  g2211 (n1988, n1938);
not  g2212 (n2067, n1931);
buf  g2213 (n2442, n1961);
buf  g2214 (n2586, n1819);
not  g2215 (n2025, n1853);
not  g2216 (n2291, n1833);
not  g2217 (n2040, n1822);
not  g2218 (n2647, n1925);
not  g2219 (n2450, n1829);
not  g2220 (n2094, n1844);
buf  g2221 (n2200, n1492);
buf  g2222 (n2602, n1797);
not  g2223 (n2366, n1922);
not  g2224 (n2486, n1849);
not  g2225 (n2128, n1834);
not  g2226 (n2057, n1820);
buf  g2227 (n2095, n1964);
buf  g2228 (n2557, n1855);
not  g2229 (n2539, n1928);
not  g2230 (n2009, n1958);
buf  g2231 (n2611, n1912);
buf  g2232 (n2615, n1938);
buf  g2233 (n2175, n1843);
buf  g2234 (n2012, n1798);
not  g2235 (n2495, n1959);
buf  g2236 (n2292, n1824);
buf  g2237 (n2671, n1869);
buf  g2238 (n2445, n1907);
buf  g2239 (n2459, n1839);
buf  g2240 (n2372, n1804);
not  g2241 (n2342, n1493);
not  g2242 (n2587, n1812);
not  g2243 (n2091, n1807);
buf  g2244 (n2187, n1803);
buf  g2245 (n2072, n1804);
not  g2246 (n2223, n1850);
buf  g2247 (n2243, n1932);
not  g2248 (n2145, n1939);
buf  g2249 (n2139, n1929);
buf  g2250 (n2238, n1870);
not  g2251 (n2427, n1911);
not  g2252 (n2083, n1949);
not  g2253 (n2518, n1812);
not  g2254 (n2505, n1876);
buf  g2255 (n2056, n1936);
buf  g2256 (n2559, n1493);
buf  g2257 (n2544, n1873);
not  g2258 (n2480, n1841);
buf  g2259 (n2556, n1810);
buf  g2260 (n2285, n1851);
not  g2261 (n2033, n1962);
buf  g2262 (n2185, n1935);
buf  g2263 (n2299, n1837);
buf  g2264 (n2184, n1932);
not  g2265 (n2426, n1867);
not  g2266 (n2573, n1812);
buf  g2267 (n2640, n1848);
buf  g2268 (n2092, n1933);
buf  g2269 (n2239, n1907);
not  g2270 (n2349, n1890);
buf  g2271 (n2380, n1879);
not  g2272 (n2309, n1865);
buf  g2273 (n2087, n1968);
not  g2274 (n1981, n1968);
buf  g2275 (n2566, n1923);
buf  g2276 (n2383, n1951);
buf  g2277 (n2440, n1845);
not  g2278 (n2038, n1887);
buf  g2279 (n2229, n1850);
not  g2280 (n2490, n1821);
buf  g2281 (n1998, n1880);
not  g2282 (n2347, n1948);
buf  g2283 (n1970, n1853);
buf  g2284 (n2416, n1811);
buf  g2285 (n2333, n1830);
buf  g2286 (n2630, n1835);
buf  g2287 (n2043, n1906);
not  g2288 (n2520, n1900);
not  g2289 (n2606, n1943);
not  g2290 (n2172, n1911);
buf  g2291 (n2456, n1916);
buf  g2292 (n2374, n1965);
not  g2293 (n2004, n1859);
buf  g2294 (n2420, n1861);
buf  g2295 (n2069, n1903);
not  g2296 (n2439, n1889);
buf  g2297 (n2122, n1924);
buf  g2298 (n2558, n1878);
buf  g2299 (n2312, n1839);
buf  g2300 (n2020, n1815);
buf  g2301 (n2234, n1892);
not  g2302 (n2415, n1794);
buf  g2303 (n2651, n1968);
not  g2304 (n2650, n1841);
not  g2305 (n2473, n1852);
not  g2306 (n2166, n1882);
buf  g2307 (n2279, n1954);
not  g2308 (n2316, n1884);
buf  g2309 (n2546, n1855);
buf  g2310 (n2588, n1803);
not  g2311 (n2155, n1846);
not  g2312 (n2103, n1928);
buf  g2313 (n2055, n1898);
buf  g2314 (n2476, n1849);
not  g2315 (n2267, n1874);
buf  g2316 (n2047, n1809);
buf  g2317 (n2364, n1904);
not  g2318 (n2245, n1894);
buf  g2319 (n2207, n1922);
not  g2320 (n2039, n1867);
buf  g2321 (n2053, n1844);
not  g2322 (n2629, n1851);
not  g2323 (n2597, n1861);
not  g2324 (n2084, n1917);
not  g2325 (n2146, n1857);
buf  g2326 (n2196, n1906);
buf  g2327 (n2514, n1957);
not  g2328 (n2137, n1941);
buf  g2329 (n2386, n1813);
not  g2330 (n2016, n1875);
not  g2331 (n2466, n1891);
buf  g2332 (n2405, n1909);
not  g2333 (n2414, n1945);
not  g2334 (n2127, n1956);
not  g2335 (n2165, n1931);
buf  g2336 (n2280, n1896);
buf  g2337 (n2623, n1930);
not  g2338 (n2584, n1944);
not  g2339 (n1976, n1953);
buf  g2340 (n2570, n1925);
not  g2341 (n2338, n1826);
not  g2342 (n2646, n1912);
not  g2343 (n2616, n1858);
buf  g2344 (n2293, n1903);
not  g2345 (n2156, n1913);
buf  g2346 (n2268, n1829);
buf  g2347 (n2378, n1918);
not  g2348 (n2464, n1832);
buf  g2349 (n2163, n1936);
not  g2350 (n2516, n1941);
not  g2351 (n2017, n1867);
not  g2352 (n2370, n1802);
buf  g2353 (n2117, n1930);
not  g2354 (n2421, n1881);
buf  g2355 (n2179, n1835);
buf  g2356 (n1987, n1850);
buf  g2357 (n2281, n1932);
buf  g2358 (n2064, n1815);
buf  g2359 (n2526, n1924);
not  g2360 (n2565, n1816);
buf  g2361 (n2289, n1950);
buf  g2362 (n2631, n1958);
buf  g2363 (n2071, n1949);
not  g2364 (n2527, n1810);
buf  g2365 (n2049, n1914);
not  g2366 (n2550, n1270);
not  g2367 (n2343, n1897);
not  g2368 (n2035, n1908);
not  g2369 (n2162, n1956);
buf  g2370 (n2144, n1814);
buf  g2371 (n1969, n1882);
buf  g2372 (n2617, n1822);
buf  g2373 (n2381, n1951);
not  g2374 (n2100, n1901);
buf  g2375 (n2237, n1806);
buf  g2376 (n2161, n1823);
buf  g2377 (n2113, n1836);
buf  g2378 (n2249, n1905);
buf  g2379 (n2193, n1958);
buf  g2380 (n2598, n1904);
not  g2381 (n2259, n1922);
buf  g2382 (n2181, n1849);
not  g2383 (n2236, n1878);
buf  g2384 (n2632, n1856);
buf  g2385 (n1973, n1889);
buf  g2386 (n2304, n1867);
buf  g2387 (n2037, n1897);
buf  g2388 (n2555, n1795);
buf  g2389 (n2063, n1492);
buf  g2390 (n2455, n1932);
buf  g2391 (n2118, n1948);
not  g2392 (n2031, n1894);
not  g2393 (n2488, n1846);
buf  g2394 (n2604, n1914);
not  g2395 (n2079, n1870);
buf  g2396 (n2191, n1895);
not  g2397 (n2508, n1905);
buf  g2398 (n2098, n1843);
buf  g2399 (n2537, n1896);
not  g2400 (n2624, n1829);
not  g2401 (n2026, n1835);
not  g2402 (n2356, n1862);
not  g2403 (n2177, n1851);
buf  g2404 (n2511, n1948);
buf  g2405 (n2382, n1847);
buf  g2406 (n2296, n1840);
not  g2407 (n2561, n1896);
not  g2408 (n2099, n1935);
not  g2409 (n2209, n1944);
buf  g2410 (n2141, n1846);
not  g2411 (n2023, n1935);
not  g2412 (n2136, n1876);
not  g2413 (n2250, n1901);
not  g2414 (n2402, n1801);
not  g2415 (n2580, n1900);
not  g2416 (n2132, n1952);
buf  g2417 (n2085, n1900);
buf  g2418 (n2014, n1939);
buf  g2419 (n2355, n1804);
not  g2420 (n2352, n1953);
buf  g2421 (n2068, n1947);
not  g2422 (n2655, n1892);
buf  g2423 (n2627, n1943);
buf  g2424 (n1980, n1965);
not  g2425 (n2150, n1837);
not  g2426 (n2335, n1492);
buf  g2427 (n2657, n1940);
buf  g2428 (n2300, n1890);
not  g2429 (n2265, n1802);
not  g2430 (n2154, n1864);
buf  g2431 (n2090, n1827);
not  g2432 (n2669, n1866);
buf  g2433 (n2395, n1931);
buf  g2434 (n2371, n1898);
not  g2435 (n2168, n1938);
buf  g2436 (n2521, n1861);
not  g2437 (n2042, n1963);
not  g2438 (n1993, n1795);
buf  g2439 (n2654, n1493);
not  g2440 (n2549, n1826);
buf  g2441 (n2423, n1626);
not  g2442 (n2216, n1828);
not  g2443 (n2011, n1913);
buf  g2444 (n2030, n1945);
not  g2445 (n2088, n1936);
not  g2446 (n2644, n1886);
buf  g2447 (n2288, n1896);
not  g2448 (n2148, n1835);
not  g2449 (n2475, n1271);
not  g2450 (n2543, n1793);
buf  g2451 (n1995, n1818);
buf  g2452 (n2433, n1902);
buf  g2453 (n2362, n1853);
not  g2454 (n2027, n1950);
buf  g2455 (n2275, n1824);
not  g2456 (n2477, n1877);
buf  g2457 (n2115, n1803);
not  g2458 (n2065, n1870);
buf  g2459 (n2373, n1956);
not  g2460 (n2276, n1931);
buf  g2461 (n2564, n1863);
buf  g2462 (n2178, n1900);
not  g2463 (n2410, n1817);
not  g2464 (n2277, n1963);
buf  g2465 (n2303, n1864);
not  g2466 (n2258, n1814);
buf  g2467 (n2554, n1907);
buf  g2468 (n2572, n1818);
buf  g2469 (n2636, n1864);
buf  g2470 (n2302, n1899);
buf  g2471 (n2221, n1868);
buf  g2472 (n2387, n1267);
not  g2473 (n2493, n1961);
not  g2474 (n2215, n1954);
buf  g2475 (n2195, n1952);
buf  g2476 (n2120, n1858);
not  g2477 (n2452, n1963);
not  g2478 (n2397, n1923);
not  g2479 (n2104, n1927);
not  g2480 (n2620, n1903);
buf  g2481 (n2513, n1820);
not  g2482 (n2334, n1910);
not  g2483 (n2222, n1930);
not  g2484 (n2058, n1934);
buf  g2485 (n2664, n1891);
buf  g2486 (n2125, n1916);
buf  g2487 (n2052, n1872);
buf  g2488 (n2247, n1955);
not  g2489 (n2173, n1888);
not  g2490 (n2123, n1912);
buf  g2491 (n2255, n1884);
buf  g2492 (n2492, n1885);
buf  g2493 (n1985, n1882);
not  g2494 (n2458, n1967);
not  g2495 (n2021, n1939);
buf  g2496 (n2308, n1926);
buf  g2497 (n2560, n1809);
not  g2498 (n2169, n1823);
not  g2499 (n2001, n1889);
not  g2500 (n2563, n1934);
not  g2501 (n2545, n1925);
buf  g2502 (n2231, n1934);
not  g2503 (n2018, n1840);
buf  g2504 (n2457, n1865);
buf  g2505 (n2274, n1879);
buf  g2506 (n2005, n1904);
not  g2507 (n2503, n1794);
not  g2508 (n2147, n1883);
not  g2509 (n2502, n1863);
buf  g2510 (n2409, n1816);
buf  g2511 (n2266, n1873);
not  g2512 (n2607, n1954);
buf  g2513 (n2670, n1878);
not  g2514 (n2232, n1268);
not  g2515 (n2432, n1892);
buf  g2516 (n2417, n1910);
buf  g2517 (n2135, n1805);
not  g2518 (n2341, n1793);
not  g2519 (n2054, n1838);
buf  g2520 (n2321, n1847);
buf  g2521 (n2007, n1897);
not  g2522 (n2051, n1953);
not  g2523 (n2044, n1857);
not  g2524 (n2637, n1845);
not  g2525 (n2318, n1868);
not  g2526 (n2569, n1863);
not  g2527 (n2202, n1842);
not  g2528 (n2430, n1805);
buf  g2529 (n2603, n1956);
buf  g2530 (n2363, n1803);
buf  g2531 (n2567, n1933);
not  g2532 (n2672, n1883);
not  g2533 (n2609, n1882);
buf  g2534 (n1977, n1793);
buf  g2535 (n2350, n1868);
buf  g2536 (n2077, n1951);
not  g2537 (n2530, n1813);
buf  g2538 (n2438, n1796);
not  g2539 (n2278, n1946);
not  g2540 (n2470, n1858);
buf  g2541 (n2319, n1952);
not  g2542 (n2412, n1857);
not  g2543 (n2006, n1866);
buf  g2544 (n2046, n1967);
not  g2545 (n2460, n1908);
not  g2546 (n2593, n1854);
not  g2547 (n2500, n1801);
buf  g2548 (n2348, n1962);
not  g2549 (n2152, n1963);
buf  g2550 (n2328, n1910);
not  g2551 (n2111, n1824);
buf  g2552 (n2605, n1916);
not  g2553 (n2581, n1847);
not  g2554 (n2660, n1952);
buf  g2555 (n2436, n1929);
not  g2556 (n2418, n1875);
buf  g2557 (n2552, n1937);
not  g2558 (n2206, n1800);
buf  g2559 (n2133, n1935);
buf  g2560 (n2485, n1626);
buf  g2561 (n2367, n1961);
buf  g2562 (n2361, n1832);
not  g2563 (n2019, n1920);
buf  g2564 (n2408, n1874);
buf  g2565 (n2591, n1926);
not  g2566 (n2600, n1812);
not  g2567 (n2639, n1826);
not  g2568 (n2246, n1940);
not  g2569 (n2102, n1881);
buf  g2570 (n2478, n1830);
buf  g2571 (n2283, n1852);
buf  g2572 (n2468, n1908);
buf  g2573 (n2149, n1933);
not  g2574 (n2340, n1959);
not  g2575 (n2273, n1814);
buf  g2576 (n2295, n1953);
buf  g2577 (n2404, n1838);
buf  g2578 (n2384, n1939);
not  g2579 (n2225, n1898);
not  g2580 (n2368, n1927);
buf  g2581 (n2628, n1902);
buf  g2582 (n2254, n1794);
buf  g2583 (n1978, n1825);
buf  g2584 (n2208, n1828);
buf  g2585 (n2358, n1873);
not  g2586 (n2622, n1921);
buf  g2587 (n2375, n1808);
not  g2588 (n2507, n1836);
buf  g2589 (n2471, n1839);
buf  g2590 (n2029, n1964);
buf  g2591 (n2093, n1832);
buf  g2592 (n2359, n1862);
buf  g2593 (n2553, n1960);
not  g2594 (n2112, n1816);
not  g2595 (n2109, n1959);
not  g2596 (n2666, n1817);
buf  g2597 (n2653, n1822);
buf  g2598 (n2528, n1852);
not  g2599 (n2411, n1834);
buf  g2600 (n1984, n1966);
not  g2601 (n2519, n1933);
not  g2602 (n2541, n1863);
not  g2603 (n1983, n1930);
not  g2604 (n2210, n1811);
not  g2605 (n2594, n1858);
not  g2606 (n2024, n1883);
buf  g2607 (n2645, n1828);
not  g2608 (n2491, n1964);
not  g2609 (n2212, n1851);
not  g2610 (n2345, n1833);
buf  g2611 (n2535, n1967);
not  g2612 (n2219, n1797);
buf  g2613 (n2151, n1907);
buf  g2614 (n2656, n1864);
not  g2615 (n2400, n1871);
not  g2616 (n2089, n1808);
not  g2617 (n2080, n1966);
not  g2618 (n2157, n1876);
buf  g2619 (n2577, n1811);
buf  g2620 (n2062, n1860);
buf  g2621 (n2075, n1890);
buf  g2622 (n2487, n1819);
not  g2623 (n2050, n1862);
buf  g2624 (n2134, n1850);
buf  g2625 (n2074, n1926);
buf  g2626 (n2256, n1960);
not  g2627 (n2101, n1944);
not  g2628 (n2142, n1269);
not  g2629 (n2441, n1854);
not  g2630 (n2158, n1869);
buf  g2631 (n2167, n1908);
not  g2632 (n2396, n1845);
buf  g2633 (n2326, n1793);
nand g2634 (n2482, n1849, n1813, n1944, n1902);
or   g2635 (n2534, n1924, n1947, n1805, n1856);
or   g2636 (n2160, n1921, n1854, n1927, n1846);
nor  g2637 (n2467, n1901, n1823, n1955, n1960);
and  g2638 (n2601, n1917, n1920, n1966, n1895);
or   g2639 (n2625, n1942, n1875, n1798, n1809);
not  g2640 (n2728, n2519);
buf  g2641 (n3136, n2571);
not  g2642 (n3571, n2217);
not  g2643 (n3401, n2433);
not  g2644 (n3004, n2261);
not  g2645 (n2990, n2035);
buf  g2646 (n2963, n2408);
not  g2647 (n3414, n2107);
not  g2648 (n2937, n2367);
not  g2649 (n3518, n2485);
not  g2650 (n2770, n2652);
not  g2651 (n3357, n2398);
buf  g2652 (n3513, n2601);
buf  g2653 (n3652, n2638);
buf  g2654 (n2707, n2036);
not  g2655 (n2698, n2223);
buf  g2656 (n3593, n2645);
buf  g2657 (n2799, n2223);
buf  g2658 (n3020, n2536);
buf  g2659 (n2734, n1997);
buf  g2660 (n2959, n2101);
buf  g2661 (n2817, n2592);
not  g2662 (n3084, n2565);
buf  g2663 (n2995, n2022);
not  g2664 (n3028, n2236);
not  g2665 (n3076, n2486);
not  g2666 (n3460, n2095);
not  g2667 (n3480, n2481);
buf  g2668 (n3651, n2397);
not  g2669 (n3496, n2529);
not  g2670 (n2700, n2409);
buf  g2671 (n2679, n2106);
not  g2672 (n2845, n2426);
buf  g2673 (n3201, n2423);
buf  g2674 (n2816, n2391);
buf  g2675 (n3233, n2405);
buf  g2676 (n2885, n2263);
not  g2677 (n2904, n2014);
not  g2678 (n3333, n2000);
not  g2679 (n3386, n2001);
buf  g2680 (n3575, n2578);
not  g2681 (n2871, n2401);
buf  g2682 (n2964, n2049);
not  g2683 (n2810, n2460);
not  g2684 (n3286, n2479);
buf  g2685 (n3230, n2212);
buf  g2686 (n3300, n2543);
buf  g2687 (n3596, n2604);
buf  g2688 (n3334, n2094);
not  g2689 (n3183, n2605);
not  g2690 (n3462, n2260);
not  g2691 (n2865, n2429);
not  g2692 (n2684, n2470);
not  g2693 (n2968, n2258);
not  g2694 (n2717, n2563);
not  g2695 (n3110, n2129);
buf  g2696 (n3628, n2432);
buf  g2697 (n2892, n2630);
not  g2698 (n2715, n2009);
buf  g2699 (n2880, n2129);
buf  g2700 (n3093, n2539);
not  g2701 (n2912, n2372);
buf  g2702 (n3337, n2257);
not  g2703 (n3471, n2268);
not  g2704 (n2784, n2093);
not  g2705 (n2697, n2617);
not  g2706 (n3425, n2182);
buf  g2707 (n2926, n1995);
buf  g2708 (n3244, n2479);
not  g2709 (n3162, n2577);
buf  g2710 (n2850, n2459);
not  g2711 (n3666, n2353);
buf  g2712 (n2730, n1976);
not  g2713 (n3132, n1996);
buf  g2714 (n3205, n2306);
buf  g2715 (n3235, n2371);
not  g2716 (n3590, n2635);
not  g2717 (n3431, n2568);
not  g2718 (n2778, n2652);
not  g2719 (n3182, n2087);
buf  g2720 (n3508, n1996);
buf  g2721 (n3646, n2222);
not  g2722 (n3295, n2032);
not  g2723 (n2745, n2245);
not  g2724 (n2765, n2338);
not  g2725 (n3068, n2578);
not  g2726 (n2686, n2198);
not  g2727 (n2681, n2331);
not  g2728 (n3341, n2629);
not  g2729 (n2879, n2272);
buf  g2730 (n3040, n2468);
buf  g2731 (n2861, n2433);
buf  g2732 (n2965, n1969);
not  g2733 (n3143, n2533);
buf  g2734 (n2801, n2539);
not  g2735 (n3660, n2641);
not  g2736 (n3152, n2113);
buf  g2737 (n3291, n1998);
buf  g2738 (n3215, n2629);
not  g2739 (n3070, n2154);
buf  g2740 (n3461, n2632);
buf  g2741 (n2984, n2091);
not  g2742 (n3053, n2453);
buf  g2743 (n3606, n2218);
buf  g2744 (n3000, n2449);
buf  g2745 (n3487, n2174);
buf  g2746 (n2824, n2194);
buf  g2747 (n3256, n2067);
buf  g2748 (n2873, n2362);
not  g2749 (n3622, n2428);
buf  g2750 (n2827, n2584);
buf  g2751 (n2790, n2371);
not  g2752 (n3335, n2370);
not  g2753 (n3641, n2451);
not  g2754 (n2867, n2320);
buf  g2755 (n3557, n2363);
not  g2756 (n2915, n2360);
buf  g2757 (n3186, n2498);
buf  g2758 (n3368, n2254);
buf  g2759 (n2872, n2664);
buf  g2760 (n3503, n2046);
buf  g2761 (n2989, n2070);
buf  g2762 (n2754, n2305);
buf  g2763 (n3281, n2271);
buf  g2764 (n3079, n2152);
buf  g2765 (n3495, n2395);
buf  g2766 (n2907, n2418);
buf  g2767 (n3451, n2280);
buf  g2768 (n3077, n2196);
not  g2769 (n2676, n2227);
buf  g2770 (n3612, n2131);
buf  g2771 (n3473, n2242);
buf  g2772 (n3686, n2469);
not  g2773 (n3365, n2381);
not  g2774 (n3608, n2046);
not  g2775 (n3366, n2238);
buf  g2776 (n3305, n2347);
not  g2777 (n3217, n2326);
buf  g2778 (n2929, n2281);
buf  g2779 (n3320, n2200);
buf  g2780 (n2952, n2110);
buf  g2781 (n3679, n2318);
buf  g2782 (n2882, n2042);
buf  g2783 (n2977, n2526);
not  g2784 (n3313, n2533);
buf  g2785 (n3009, n2411);
not  g2786 (n3214, n2074);
not  g2787 (n3511, n2091);
buf  g2788 (n2894, n2289);
buf  g2789 (n3675, n2491);
not  g2790 (n3400, n2454);
buf  g2791 (n2962, n2394);
buf  g2792 (n3550, n2464);
not  g2793 (n3393, n2517);
not  g2794 (n3052, n2456);
not  g2795 (n3038, n1981);
not  g2796 (n3617, n2350);
buf  g2797 (n3275, n2212);
not  g2798 (n2769, n2330);
not  g2799 (n2789, n2273);
buf  g2800 (n3671, n2005);
buf  g2801 (n3510, n2579);
not  g2802 (n3683, n2477);
buf  g2803 (n3031, n2497);
not  g2804 (n3553, n2242);
buf  g2805 (n3445, n2307);
not  g2806 (n3197, n2051);
buf  g2807 (n2750, n1980);
buf  g2808 (n3198, n2523);
buf  g2809 (n3269, n2578);
not  g2810 (n3263, n2381);
not  g2811 (n3155, n2238);
buf  g2812 (n3193, n2099);
buf  g2813 (n3620, n2453);
buf  g2814 (n2840, n2465);
not  g2815 (n3072, n2100);
not  g2816 (n3689, n2602);
buf  g2817 (n3229, n2266);
not  g2818 (n3113, n2230);
not  g2819 (n2719, n2274);
not  g2820 (n3432, n2523);
buf  g2821 (n2890, n2248);
not  g2822 (n3655, n2199);
buf  g2823 (n3149, n2536);
buf  g2824 (n3434, n2667);
not  g2825 (n2759, n2007);
not  g2826 (n3219, n2653);
buf  g2827 (n2802, n2577);
buf  g2828 (n2924, n2602);
buf  g2829 (n3658, n2064);
not  g2830 (n3424, n2440);
buf  g2831 (n2819, n2603);
not  g2832 (n3029, n2409);
not  g2833 (n2691, n2036);
not  g2834 (n3456, n2563);
buf  g2835 (n2888, n2250);
not  g2836 (n2785, n2071);
buf  g2837 (n2991, n2179);
not  g2838 (n3100, n2239);
not  g2839 (n3248, n2190);
not  g2840 (n3170, n2609);
buf  g2841 (n3164, n2432);
buf  g2842 (n3342, n2149);
not  g2843 (n3437, n2096);
not  g2844 (n2948, n2408);
not  g2845 (n2976, n2206);
buf  g2846 (n3045, n2208);
buf  g2847 (n3454, n2514);
not  g2848 (n3018, n2518);
buf  g2849 (n3607, n2082);
not  g2850 (n2967, n2516);
buf  g2851 (n3088, n2022);
buf  g2852 (n3290, n2281);
buf  g2853 (n3345, n2169);
buf  g2854 (n3125, n2070);
not  g2855 (n3667, n2427);
not  g2856 (n3016, n2672);
not  g2857 (n3243, n2225);
buf  g2858 (n3552, n2065);
not  g2859 (n2726, n1975);
buf  g2860 (n3479, n2086);
not  g2861 (n3207, n2079);
buf  g2862 (n2881, n2588);
buf  g2863 (n3528, n2251);
buf  g2864 (n3145, n2266);
buf  g2865 (n2951, n2374);
buf  g2866 (n3589, n2643);
buf  g2867 (n3124, n2537);
not  g2868 (n3429, n2577);
buf  g2869 (n3287, n2388);
not  g2870 (n2826, n2107);
buf  g2871 (n3331, n2385);
buf  g2872 (n2988, n2526);
buf  g2873 (n2744, n2073);
buf  g2874 (n3411, n2312);
buf  g2875 (n2866, n2524);
buf  g2876 (n3481, n2012);
buf  g2877 (n2766, n2137);
not  g2878 (n2847, n2245);
not  g2879 (n2943, n2642);
not  g2880 (n3024, n2630);
buf  g2881 (n3301, n2484);
not  g2882 (n3466, n2474);
not  g2883 (n2993, n2663);
buf  g2884 (n3267, n2624);
buf  g2885 (n3316, n2099);
buf  g2886 (n3150, n2275);
buf  g2887 (n3184, n2166);
buf  g2888 (n3399, n2256);
not  g2889 (n3035, n2092);
buf  g2890 (n2944, n2262);
buf  g2891 (n3647, n2019);
not  g2892 (n3138, n2302);
not  g2893 (n3396, n2276);
buf  g2894 (n3063, n2214);
buf  g2895 (n3225, n2167);
not  g2896 (n3584, n2313);
buf  g2897 (n2955, n2378);
buf  g2898 (n3604, n2317);
buf  g2899 (n3529, n2190);
buf  g2900 (n3677, n2034);
not  g2901 (n3385, n2118);
buf  g2902 (n3379, n2568);
not  g2903 (n2994, n2418);
buf  g2904 (n3500, n2615);
not  g2905 (n3436, n2368);
buf  g2906 (n3003, n2412);
not  g2907 (n3586, n2585);
not  g2908 (n3468, n2295);
buf  g2909 (n3426, n2616);
buf  g2910 (n3327, n2080);
not  g2911 (n3177, n2637);
not  g2912 (n3315, n2421);
buf  g2913 (n2986, n2644);
buf  g2914 (n3339, n2021);
buf  g2915 (n3619, n2253);
buf  g2916 (n2807, n2490);
not  g2917 (n2982, n2399);
not  g2918 (n3567, n2627);
buf  g2919 (n3044, n2138);
not  g2920 (n3092, n2201);
not  g2921 (n2763, n2109);
buf  g2922 (n3506, n2403);
not  g2923 (n3592, n2098);
buf  g2924 (n2875, n2429);
not  g2925 (n2891, n2269);
buf  g2926 (n2786, n1993);
not  g2927 (n2673, n2003);
not  g2928 (n3352, n2444);
not  g2929 (n3600, n2244);
not  g2930 (n3283, n2196);
buf  g2931 (n2781, n2216);
buf  g2932 (n3369, n2157);
buf  g2933 (n3277, n2407);
buf  g2934 (n3325, n2122);
not  g2935 (n2808, n2316);
buf  g2936 (n3657, n2336);
buf  g2937 (n3416, n2110);
not  g2938 (n3624, n2625);
buf  g2939 (n3037, n2493);
not  g2940 (n3493, n2143);
not  g2941 (n3535, n2340);
buf  g2942 (n2958, n2572);
buf  g2943 (n3169, n2349);
not  g2944 (n3080, n2062);
buf  g2945 (n2946, n2180);
buf  g2946 (n3408, n2316);
not  g2947 (n3157, n2567);
not  g2948 (n2695, n2365);
not  g2949 (n2849, n2209);
not  g2950 (n3098, n2394);
not  g2951 (n3580, n2580);
buf  g2952 (n3258, n2463);
not  g2953 (n2748, n2559);
buf  g2954 (n3603, n2117);
not  g2955 (n2812, n2131);
not  g2956 (n3474, n2327);
buf  g2957 (n2868, n2243);
buf  g2958 (n3464, n2266);
buf  g2959 (n2978, n2128);
buf  g2960 (n3087, n1982);
buf  g2961 (n3662, n2423);
buf  g2962 (n3034, n2373);
not  g2963 (n2806, n2069);
buf  g2964 (n2788, n2585);
buf  g2965 (n3563, n2209);
not  g2966 (n3234, n1987);
not  g2967 (n2947, n1972);
buf  g2968 (n3463, n2552);
not  g2969 (n2838, n2078);
not  g2970 (n3616, n2457);
not  g2971 (n3459, n2584);
buf  g2972 (n3645, n2305);
buf  g2973 (n3351, n2054);
buf  g2974 (n3273, n2291);
buf  g2975 (n3171, n2287);
buf  g2976 (n3525, n1725);
buf  g2977 (n3423, n2439);
buf  g2978 (n3579, n2450);
not  g2979 (n3112, n2543);
not  g2980 (n2889, n2504);
buf  g2981 (n3505, n2298);
not  g2982 (n2960, n2092);
buf  g2983 (n3635, n2304);
buf  g2984 (n3326, n2204);
not  g2985 (n3490, n2558);
buf  g2986 (n2966, n2498);
buf  g2987 (n2914, n2146);
not  g2988 (n3472, n2124);
not  g2989 (n2804, n2648);
buf  g2990 (n3404, n2233);
buf  g2991 (n3324, n2614);
not  g2992 (n3439, n2109);
not  g2993 (n3610, n2471);
not  g2994 (n3644, n2653);
buf  g2995 (n3440, n2528);
buf  g2996 (n2877, n2515);
buf  g2997 (n3328, n2012);
not  g2998 (n2767, n2052);
buf  g2999 (n3661, n2067);
buf  g3000 (n3421, n2634);
buf  g3001 (n3498, n2541);
buf  g3002 (n3049, n2580);
not  g3003 (n3378, n2027);
not  g3004 (n2740, n2549);
not  g3005 (n2841, n2173);
buf  g3006 (n2999, n2318);
buf  g3007 (n3344, n2501);
not  g3008 (n2851, n2145);
not  g3009 (n2809, n2105);
not  g3010 (n2800, n2285);
not  g3011 (n3137, n2101);
not  g3012 (n3522, n2299);
not  g3013 (n3173, n2579);
not  g3014 (n2737, n2310);
buf  g3015 (n3241, n2477);
not  g3016 (n3254, n2101);
not  g3017 (n3135, n2635);
buf  g3018 (n3298, n2604);
not  g3019 (n3191, n2347);
not  g3020 (n2940, n2044);
buf  g3021 (n3422, n2063);
buf  g3022 (n3541, n2278);
buf  g3023 (n3476, n2126);
not  g3024 (n2859, n2135);
not  g3025 (n3467, n2308);
buf  g3026 (n2874, n2426);
not  g3027 (n3682, n2512);
buf  g3028 (n3103, n2427);
not  g3029 (n2961, n2519);
buf  g3030 (n3159, n2542);
not  g3031 (n2900, n2191);
not  g3032 (n3515, n2112);
buf  g3033 (n2975, n2644);
buf  g3034 (n3289, n2469);
not  g3035 (n2677, n2392);
not  g3036 (n2870, n2516);
buf  g3037 (n3653, n2569);
buf  g3038 (n3636, n2535);
buf  g3039 (n2839, n2219);
buf  g3040 (n3502, n2533);
not  g3041 (n2795, n2383);
not  g3042 (n3014, n2466);
not  g3043 (n2797, n2072);
not  g3044 (n3625, n1976);
not  g3045 (n3073, n2217);
not  g3046 (n3066, n2482);
not  g3047 (n3388, n2051);
not  g3048 (n3309, n2374);
not  g3049 (n2909, n2600);
not  g3050 (n3687, n1725);
not  g3051 (n3151, n2087);
not  g3052 (n3226, n2409);
not  g3053 (n3587, n2528);
not  g3054 (n2934, n2103);
not  g3055 (n2729, n2052);
and  g3056 (n2743, n2448, n2033, n2672, n2427);
nor  g3057 (n2886, n2017, n2527, n2611, n1983);
and  g3058 (n3486, n2307, n2588, n2056, n2160);
nand g3059 (n3268, n2081, n2488, n2228, n2406);
nand g3060 (n3544, n1978, n2021, n2443, n2286);
nand g3061 (n3370, n2475, n2327, n2290, n2502);
nand g3062 (n3321, n2166, n2648, n2150, n2128);
nor  g3063 (n3444, n2443, n2406, n1979, n2300);
nand g3064 (n3623, n2006, n2660, n2610, n2393);
nand g3065 (n3123, n2494, n2245, n2445, n2085);
or   g3066 (n3250, n2175, n2544, n2520, n2476);
nand g3067 (n3175, n2522, n2055, n2589, n2322);
xor  g3068 (n3097, n2534, n2336, n2593, n2109);
xor  g3069 (n2974, n2481, n2459, n2615, n2132);
nand g3070 (n3008, n2608, n2569, n2543, n2288);
or   g3071 (n3349, n2518, n2077, n2297, n2419);
xnor g3072 (n3433, n2450, n2184, n2015, n2437);
nand g3073 (n3394, n2366, n2424, n2100, n2206);
nor  g3074 (n2722, n2376, n2345, n2468, n1985);
xor  g3075 (n3047, n2461, n2659, n2534, n2441);
nor  g3076 (n3621, n2662, n2594, n2119, n2670);
xor  g3077 (n2830, n2315, n2134, n2312, n2116);
or   g3078 (n3140, n2027, n2180, n2331, n2134);
and  g3079 (n3308, n2448, n2013, n2621, n2043);
nor  g3080 (n3189, n2380, n2082, n2520, n2094);
xor  g3081 (n3237, n2246, n2523, n2168, n2362);
or   g3082 (n2818, n2447, n2369, n2360, n2306);
xor  g3083 (n3144, n2538, n2228, n2018, n2004);
nand g3084 (n3684, n2458, n2367, n2625, n2021);
nand g3085 (n2735, n2562, n2532, n2360, n2520);
nand g3086 (n3240, n2110, n2284, n1991, n2669);
or   g3087 (n3319, n2446, n2298, n2177, n2389);
nor  g3088 (n2761, n2483, n2016, n2597, n1150);
nand g3089 (n3158, n2657, n2461, n2122, n2168);
nand g3090 (n2935, n2278, n2584, n2048, n2579);
nand g3091 (n2749, n2137, n2444, n2275, n2531);
and  g3092 (n2774, n2669, n2309, n2400, n2570);
nand g3093 (n3074, n2278, n2091, n2093, n2657);
xor  g3094 (n3364, n2518, n2440, n2130, n2011);
or   g3095 (n3247, n2495, n2097, n2319, n2435);
xnor g3096 (n3601, n2332, n2014, n2120, n2351);
xnor g3097 (n2724, n2261, n2167, n2671, n2127);
xnor g3098 (n3353, n2629, n2075, n1990, n2529);
xor  g3099 (n2688, n2415, n2121, n2463, n2220);
nand g3100 (n3134, n2286, n1977, n2407, n2576);
nand g3101 (n3649, n2250, n2646, n2425, n2566);
nand g3102 (n3668, n2509, n2472, n2296, n2373);
and  g3103 (n3071, n2581, n2364, n2237, n2436);
and  g3104 (n2689, n2009, n2120, n2159, n2276);
or   g3105 (n3489, n2142, n2251, n2543, n2364);
or   g3106 (n3428, n2312, n2321, n2358, n2092);
or   g3107 (n2713, n2564, n2173, n2029, n2318);
or   g3108 (n2752, n2386, n2529, n2498, n2243);
xnor g3109 (n2683, n2082, n2225, n2189, n2066);
and  g3110 (n3259, n2183, n2408, n2316, n2401);
xnor g3111 (n3648, n2535, n2521, n2303, n2069);
xnor g3112 (n2949, n2409, n2289, n2451, n2260);
nand g3113 (n3499, n2525, n2510, n2620, n2249);
or   g3114 (n2864, n2460, n2395, n2358, n2172);
xnor g3115 (n3279, n2610, n2473, n2037, n2307);
or   g3116 (n3245, n1969, n1987, n2339, n1986);
and  g3117 (n3665, n2235, n2516, n2211, n2425);
and  g3118 (n3311, n2458, n2541, n1997, n2385);
or   g3119 (n2848, n2593, n2147, n2366, n2464);
and  g3120 (n2853, n2091, n2207, n2152, n2171);
xor  g3121 (n2723, n2267, n2300, n2179, n2403);
xor  g3122 (n3566, n2263, n2043, n2317, n2195);
or   g3123 (n3221, n2591, n2563, n1992, n2355);
xor  g3124 (n3120, n1995, n2483, n2507, n2453);
or   g3125 (n2702, n2390, n2525, n2449, n2033);
and  g3126 (n3163, n2398, n2469, n2174, n1972);
nand g3127 (n3101, n2452, n2661, n2294, n2374);
nor  g3128 (n3545, n2117, n2486, n2296, n2410);
nand g3129 (n3395, n2449, n2233, n2557, n2591);
or   g3130 (n3517, n2231, n2084, n2281, n2205);
xor  g3131 (n3293, n2666, n2183, n2415, n2552);
and  g3132 (n2998, n2301, n2191, n2223, n2603);
xnor g3133 (n2736, n2656, n2496, n2012, n2597);
xnor g3134 (n3390, n2202, n2143, n2133, n2097);
nand g3135 (n3211, n2595, n2560, n2325, n2571);
or   g3136 (n2869, n2148, n2288, n2047, n2545);
or   g3137 (n3167, n2077, n2159, n2189, n2103);
nand g3138 (n3094, n2343, n2650, n2483, n2363);
xnor g3139 (n3354, n2083, n2258, n1988, n2032);
and  g3140 (n3470, n2275, n2623, n2010, n2218);
nand g3141 (n3059, n2598, n2672, n2331, n2399);
xnor g3142 (n3494, n2170, n2352, n2287, n2432);
xor  g3143 (n3501, n2299, n2545, n2100, n2633);
nor  g3144 (n3389, n2377, n2584, n2162, n2030);
and  g3145 (n3266, n2644, n2527, n2197, n2238);
and  g3146 (n2931, n2538, n2176, n2182, n2013);
nor  g3147 (n3469, n2384, n2079, n2428, n2051);
nand g3148 (n2985, n2586, n2167, n1985, n2127);
nand g3149 (n2741, n2018, n2609, n2037, n2515);
and  g3150 (n2843, n2083, n2476, n2052, n2592);
or   g3151 (n3203, n2342, n2360, n2639, n2064);
and  g3152 (n3520, n2170, n2211, n2645, n2596);
xnor g3153 (n3484, n2108, n2086, n2301, n2491);
xor  g3154 (n3446, n2090, n2224, n2421, n2024);
xnor g3155 (n3294, n2454, n2124, n2247, n2607);
nor  g3156 (n2798, n2078, n2495, n2170, n2664);
nor  g3157 (n3096, n2650, n2227, n1281, n2122);
xnor g3158 (n3210, n2397, n2377, n2424, n2540);
or   g3159 (n3148, n2367, n2467, n2478, n2658);
xor  g3160 (n3449, n2646, n2224, n2264, n2462);
xnor g3161 (n2918, n2596, n2325, n2039, n2037);
nor  g3162 (n2979, n2181, n2136, n2088, n2254);
nor  g3163 (n2887, n2148, n1971, n2159, n2548);
or   g3164 (n2858, n2503, n2348, n2071, n2632);
nor  g3165 (n3042, n2435, n2230, n2527, n2188);
nor  g3166 (n3156, n2185, n2407, n2564, n2422);
and  g3167 (n2762, n1988, n2265, n2290, n2643);
or   g3168 (n2708, n2511, n2055, n2581, n2598);
nand g3169 (n3027, n2291, n2042, n2253, n2570);
xor  g3170 (n3430, n1975, n2054, n2205, n2537);
nand g3171 (n3373, n2192, n2067, n2554, n2242);
or   g3172 (n2954, n2619, n1984, n2641, n2249);
xnor g3173 (n3450, n2354, n2648, n2431, n2293);
xor  g3174 (n3418, n2422, n1984, n2509, n2199);
and  g3175 (n2941, n2346, n2020, n2550, n2103);
xor  g3176 (n2895, n2499, n2513, n2641, n2535);
and  g3177 (n3630, n2321, n2490, n2229, n2305);
nor  g3178 (n3435, n2280, n2410, n2492, n2050);
and  g3179 (n3627, n1983, n2231, n2370, n2019);
nand g3180 (n3391, n2029, n2040, n2663, n2566);
xnor g3181 (n2682, n2520, n2330, n2487, n2504);
xnor g3182 (n3139, n2525, n2413, n2487, n2344);
nor  g3183 (n3192, n2389, n2574, n2058, n2611);
nand g3184 (n2680, n2556, n2424, n2380, n2207);
nor  g3185 (n3676, n2338, n2358, n2295, n2503);
and  g3186 (n3067, n1986, n2114, n2158, n2473);
xor  g3187 (n2813, n2618, n2497, n2640, n2164);
nor  g3188 (n2690, n2442, n2018, n2163, n2650);
and  g3189 (n3504, n2436, n2631, n2158, n2632);
or   g3190 (n3054, n2065, n2147, n2124, n2504);
nand g3191 (n2842, n2183, n1970, n2562, n2341);
xnor g3192 (n3565, n2262, n2313, n2551, n2349);
xor  g3193 (n3208, n2576, n2315, n2586, n2231);
nand g3194 (n3046, n2165, n2108, n2203, n2301);
xor  g3195 (n2772, n1991, n2507, n2134, n2418);
xor  g3196 (n3121, n2239, n2284, n2149, n2022);
and  g3197 (n2701, n2353, n2587, n2515, n2456);
xnor g3198 (n2791, n2642, n2597, n2165, n2359);
nand g3199 (n3099, n2445, n2207, n2513, n2405);
xor  g3200 (n3497, n2237, n2499, n2161, n2460);
xor  g3201 (n3249, n2352, n2467, n2586, n2018);
or   g3202 (n2738, n2196, n2273, n2171, n2132);
nor  g3203 (n2936, n2350, n2420, n2378, n2376);
xnor g3204 (n3239, n1998, n2017, n2038, n2020);
xor  g3205 (n3222, n2488, n2182, n2115, n2292);
or   g3206 (n3637, n2049, n2243, n2148, n2176);
xor  g3207 (n2899, n2528, n2398, n2436, n2107);
xnor g3208 (n3447, n2649, n2522, n2028, n2144);
xor  g3209 (n3115, n2635, n2336, n2338, n2270);
nand g3210 (n2751, n2341, n2572, n2357, n2002);
or   g3211 (n3402, n2614, n2532, n2517, n2274);
xor  g3212 (n3599, n2211, n2152, n2633, n2216);
nand g3213 (n3160, n2029, n2404, n2270, n2647);
or   g3214 (n2732, n2422, n2172, n2229, n2205);
nor  g3215 (n3632, n2570, n2358, n2606, n2387);
and  g3216 (n2862, n2181, n2624, n2026, n2060);
and  g3217 (n3374, n2012, n2112, n2114, n2041);
xor  g3218 (n2893, n2613, n2273, n2314, n2017);
xnor g3219 (n2860, n2591, n2590, n2292, n2468);
or   g3220 (n3188, n2221, n2158, n2596, n2041);
and  g3221 (n2897, n2519, n2665, n2576, n2160);
nand g3222 (n3129, n2234, n1991, n2075, n2061);
nor  g3223 (n3336, n2419, n2249, n2011, n2089);
nand g3224 (n2919, n2261, n2354, n2260, n2605);
nor  g3225 (n2720, n2531, n2310, n1970, n2031);
nand g3226 (n2925, n2430, n2041, n2061, n2311);
xnor g3227 (n2777, n2466, n2257, n2244, n2514);
xor  g3228 (n3538, n2404, n2510, n2302, n2142);
xor  g3229 (n3306, n2432, n2345, n2169, n2052);
or   g3230 (n3602, n2580, n2558, n2352, n2095);
and  g3231 (n3001, n2075, n2440, n1982, n2114);
xor  g3232 (n3105, n2669, n2201, n2583, n2213);
nand g3233 (n2796, n2664, n2116, n2448, n2222);
nand g3234 (n3307, n2611, n2032, n2375, n2076);
and  g3235 (n3238, n2028, n2206, n1969, n2099);
xnor g3236 (n3507, n2205, n2630, n2502, n2670);
and  g3237 (n3270, n2225, n2130, n2451, n1978);
nand g3238 (n2828, n2428, n2073, n2160, n2150);
nor  g3239 (n3438, n2439, n2300, n2153, n2608);
xor  g3240 (n3174, n1989, n2472, n2383, n2512);
nand g3241 (n3537, n2057, n2615, n1993, n2006);
or   g3242 (n3427, n1984, n2240, n2281, n2188);
and  g3243 (n3585, n2570, n2472, n2430, n2025);
nand g3244 (n2922, n1984, n2671, n1995, n2140);
nor  g3245 (n2727, n2050, n2290, n2023);
nand g3246 (n3010, n2203, n2590, n2186, n2338);
nor  g3247 (n2983, n2031, n1990, n2340, n2416);
xor  g3248 (n2820, n2599, n2626, n2314, n2140);
nor  g3249 (n3312, n2064, n2670, n2509, n2480);
xnor g3250 (n2794, n2282, n2038, n2257, n1994);
and  g3251 (n2910, n2437, n2034, n1986, n2187);
xnor g3252 (n2823, n2573, n2482, n2618, n2393);
and  g3253 (n3292, n2094, n2465, n2458, n1999);
nand g3254 (n3262, n2046, n2090, n2623, n2308);
and  g3255 (n3033, n2036, n2010, n1975, n2125);
xnor g3256 (n3371, n2617, n2541, n2035, n2636);
or   g3257 (n3021, n2651, n2159, n2335, n2494);
or   g3258 (n3492, n2384, n2607, n2470, n2314);
xor  g3259 (n3179, n2264, n2045, n2495, n2662);
xor  g3260 (n3332, n2366, n2193, n2368, n2485);
and  g3261 (n3108, n2285, n2083, n2218, n2455);
xor  g3262 (n2831, n2454, n2241, n2128, n2319);
and  g3263 (n2792, n2522, n2185, n2139, n2345);
xor  g3264 (n3442, n2429, n2274, n2592, n2390);
and  g3265 (n3534, n2183, n2235, n2239, n2119);
or   g3266 (n2706, n2392, n2000, n2102, n2166);
or   g3267 (n3271, n2187, n2006, n1988, n2128);
xnor g3268 (n3236, n2456, n2289, n2101, n2387);
xnor g3269 (n2992, n2198, n2148, n2038, n2362);
or   g3270 (n3681, n1724, n1992, n2212, n2210);
xor  g3271 (n3588, n2634, n2057, n2534, n2144);
xor  g3272 (n3670, n2104, n2268, n2557, n2539);
or   g3273 (n3128, n2601, n2249, n2433, n2126);
xnor g3274 (n3547, n1981, n2654, n2202, n2283);
or   g3275 (n2956, n2209, n2154, n2640, n1994);
xor  g3276 (n3296, n2530, n2070, n2228, n2127);
xor  g3277 (n3420, n2302, n2600, n2090, n2279);
xor  g3278 (n2718, n2550, n2668, n2175, n2121);
or   g3279 (n2923, n2318, n2574, n2568, n2660);
xnor g3280 (n3019, n2178, n2535, n2186, n2076);
and  g3281 (n3025, n2484, n2453, n2447, n2482);
nor  g3282 (n3085, n2527, n2490, n2279, n2554);
nor  g3283 (n3591, n2573, n2512, n2227, n2312);
or   g3284 (n3410, n2648, n2463, n2378, n2043);
xnor g3285 (n2908, n2008, n2481, n2621, n2431);
xor  g3286 (n3199, n2560, n2619, n2304, n2079);
xor  g3287 (n3011, n2118, n2151, n2630, n2620);
xor  g3288 (n3548, n2122, n2442, n2405, n2219);
nand g3289 (n3405, n1980, n2457, n2555, n2123);
or   g3290 (n3477, n2206, n2599, n1996, n1979);
xnor g3291 (n3482, n2324, n2252, n2203, n2389);
xnor g3292 (n3465, n2660, n2395, n2476, n2105);
xor  g3293 (n3611, n2464, n2369, n2413, n2577);
nor  g3294 (n3075, n2209, n1281, n2575, n2384);
xor  g3295 (n3669, n2085, n2595, n2009, n2339);
and  g3296 (n3272, n2553, n2295, n2554, n2669);
nand g3297 (n3255, n2119, n2567, n2365, n2073);
nand g3298 (n3104, n2027, n2246, n2390, n2665);
nand g3299 (n3091, n2066, n2461, n2447, n2420);
nand g3300 (n3064, n2342, n2532, n2246, n2306);
nor  g3301 (n3176, n2142, n2659, n2105, n2414);
nor  g3302 (n2753, n2220, n2631, n2425, n2585);
nor  g3303 (n3614, n2186, n2412, n2402, n2328);
xor  g3304 (n3419, n2266, n2337, n2410, n2039);
nor  g3305 (n3251, n2553, n2372, n1993, n2116);
xnor g3306 (n3549, n2567, n2443, n2069, n1977);
and  g3307 (n3348, n2073, n2176, n2228, n2553);
xnor g3308 (n3261, n2244, n2024, n2198, n2191);
xnor g3309 (n3690, n2059, n2368, n2098, n2446);
xnor g3310 (n2938, n2588, n2633, n2355, n2501);
xor  g3311 (n2855, n2003, n2113, n2450, n2220);
nor  g3312 (n3346, n2382, n2455, n2065, n2332);
nor  g3313 (n2675, n2333, n2220, n2262, n2440);
and  g3314 (n3232, n2322, n2270, n2037, n2296);
and  g3315 (n2814, n2048, n2311, n2441, n2485);
or   g3316 (n3343, n2364, n2030, n2447, n2214);
or   g3317 (n3013, n2104, n2533, n2106, n2057);
and  g3318 (n2833, n2478, n2256, n2115, n2282);
nor  g3319 (n2933, n2315, n2505, n2334, n2581);
nor  g3320 (n2716, n2549, n2627, n2028, n2141);
nand g3321 (n3597, n2247, n2276, n2548, n2564);
xnor g3322 (n3483, n2559, n2264, n2574, n2641);
and  g3323 (n3392, n1995, n2084, n2292);
or   g3324 (n3441, n2240, n2058, n1999, n2064);
nand g3325 (n2911, n2201, n2412, n2376, n2636);
xnor g3326 (n2878, n2291, n2471, n2000, n2622);
or   g3327 (n3127, n2323, n2592, n2216, n2339);
and  g3328 (n2710, n2002, n2572, n2420, n2272);
nand g3329 (n3181, n2619, n2332, n2590, n2658);
xnor g3330 (n3133, n2375, n2357, n1281, n2045);
or   g3331 (n2939, n2333, n2345, n2446, n2426);
xnor g3332 (n2950, n2391, n2158, n2173, n2487);
or   g3333 (n3457, n2613, n2561, n2119, n2661);
and  g3334 (n3223, n2272, n2127, n2293, n2600);
nor  g3335 (n3015, n2255, n2189, n2460, n2024);
xor  g3336 (n3323, n2387, n2302, n2429, n2337);
xor  g3337 (n3274, n2637, n2606, n2499, n2561);
xnor g3338 (n2757, n2646, n2479, n2059, n2271);
xnor g3339 (n3384, n2497, n2063, n2549, n2089);
xnor g3340 (n2776, n2374, n2132, n2068, n2298);
and  g3341 (n2846, n2187, n2156, n2352, n2449);
or   g3342 (n3224, n2200, n2136, n2620, n2224);
and  g3343 (n2721, n2664, n2264, n2510, n2317);
nand g3344 (n3194, n2547, n2661, n2214, n2106);
nand g3345 (n2930, n2645, n2178, n2593, n2088);
xor  g3346 (n3242, n2034, n2369, n2136, n2588);
xnor g3347 (n3165, n2045, n2192, n2177, n2373);
nor  g3348 (n2793, n2326, n2267, n2472, n2276);
and  g3349 (n3317, n2081, n2118, n2403, n2598);
xor  g3350 (n3202, n2356, n2141, n2248, n2161);
or   g3351 (n2815, n2417, n2314, n2188, n2466);
nor  g3352 (n2782, n2524, n2020, n2006, n1988);
xor  g3353 (n2711, n2373, n2389, n2617, n2189);
or   g3354 (n2945, n2045, n2537, n2299, n2420);
xnor g3355 (n3412, n2506, n2546, n1980, n1999);
or   g3356 (n3551, n2139, n2438, n2108);
nand g3357 (n2739, n2613, n2503, n2335, n2467);
nand g3358 (n2883, n2670, n2048, n2564, n2359);
nand g3359 (n3299, n2371, n2671, n2247, n2089);
nand g3360 (n2771, n2399, n2353, n2168, n2528);
and  g3361 (n3131, n2125, n2023, n2226, n2241);
nand g3362 (n2696, n2628, n2591, n2157, n2040);
and  g3363 (n3536, n2278, n2482, n2546, n1999);
nand g3364 (n3282, n2184, n2511, n2289, n2372);
xor  g3365 (n3055, n2551, n1976, n2261, n2117);
nand g3366 (n3265, n2230, n2448, n2471, n2135);
or   g3367 (n3329, n2143, n2001, n2563, n1151);
or   g3368 (n3111, n2421, n2333, n2370, n2025);
xnor g3369 (n2775, n2379, n2020, n2505, n2425);
nand g3370 (n2709, n2502, n2344, n2053, n2507);
and  g3371 (n3453, n2202, n2368, n2149, n2293);
and  g3372 (n3556, n2229, n2161, n2477, n2255);
nor  g3373 (n2768, n2537, n2552, n2286, n2493);
nor  g3374 (n3168, n2530, n2462, n2582, n2212);
nor  g3375 (n3577, n2436, n2589, n2607, n2546);
and  g3376 (n3288, n2339, n2137, n1998, n2480);
xor  g3377 (n3178, n2335, n2296, n2393, n2651);
nor  g3378 (n2832, n2151, n2007, n2230, n2439);
or   g3379 (n3172, n2388, n2130, n2254, n2143);
and  g3380 (n2901, n2156, n2363, n2236, n2499);
or   g3381 (n3304, n2252, n2478, n2434, n2647);
nor  g3382 (n2687, n2328, n2169, n2565, n2111);
and  g3383 (n3640, n2219, n2084, n2351, n2199);
xor  g3384 (n3057, n2659, n2146, n2643, n2197);
nand g3385 (n3069, n2150, n2506, n2117, n2233);
or   g3386 (n3253, n2326, n2098, n2423, n2615);
or   g3387 (n3039, n2629, n2524, n2277, n2153);
nand g3388 (n2905, n2334, n2022, n2309, n2115);
nor  g3389 (n2969, n2394, n2356, n2489, n2610);
and  g3390 (n3458, n2351, n2381, n2256, n2551);
nand g3391 (n3114, n2234, n2237, n2106, n2210);
xor  g3392 (n3407, n2011, n2265, n2310, n2033);
or   g3393 (n3509, n2607, n2030, n2016, n2337);
xor  g3394 (n3117, n2540, n2330, n2606, n2636);
nand g3395 (n3650, n1993, n2626, n2337, n2372);
xor  g3396 (n2854, n2309, n2435, n2098, n2624);
xor  g3397 (n2953, n2195, n2199, n2634, n2488);
xor  g3398 (n3142, n2556, n2571, n2093, n2263);
and  g3399 (n3519, n2594, n2634, n2016, n2378);
and  g3400 (n3231, n2505, n2622, n1978, n2273);
and  g3401 (n3488, n2200, n2547, n2462, n2178);
or   g3402 (n3206, n2416, n2216, n2089, n2452);
and  g3403 (n3081, n2536, n2221, n1981, n2214);
and  g3404 (n2942, n2229, n2053, n2161, n2521);
or   g3405 (n3539, n2149, n1973, n2382, n2210);
nor  g3406 (n2758, n2654, n2379, n2465, n2193);
xor  g3407 (n3598, n2491, n2365, n2349, n2062);
xor  g3408 (n2857, n2125, n2044, n2461, n2019);
xnor g3409 (n3375, n2172, n2283, n2135, n2181);
and  g3410 (n2779, n2344, n2003, n2654, n1983);
nand g3411 (n3322, n2666, n2396, n2054, n1979);
and  g3412 (n3659, n2023, n2002, n2538, n2328);
nand g3413 (n3691, n2316, n2604, n2599, n2190);
nor  g3414 (n3026, n2074, n2568, n2324, n2411);
nand g3415 (n3634, n2557, n2333, n2479, n2139);
nand g3416 (n3533, n2113, n2068, n2546, n2558);
nand g3417 (n3212, n2610, n2396, n2086, n2375);
nand g3418 (n3146, n2177, n2053, n2295, n2300);
and  g3419 (n2731, n2121, n2665, n2059, n2541);
or   g3420 (n3362, n2123, n2297, n1985, n1974);
nor  g3421 (n3526, n2565, n2071, n2208, n2580);
xnor g3422 (n3367, n2162, n2155, n2414, n2138);
nor  g3423 (n3338, n2323, n1994, n2049, n2009);
or   g3424 (n2970, n2594, n2474, n1974, n2431);
xnor g3425 (n3516, n2309, n2284, n2642, n2290);
nor  g3426 (n3455, n2210, n2457, n2621, n2491);
xor  g3427 (n3062, n2259, n1983, n2340, n2619);
nand g3428 (n2997, n2624, n2523, n2181, n2190);
and  g3429 (n3578, n2062, n2076, n2617, n2026);
and  g3430 (n3560, n2036, n2075, n2511, n2509);
nand g3431 (n3562, n2346, n2566, n2649, n2653);
nand g3432 (n3555, n2234, n2506, n2356, n2439);
or   g3433 (n3082, n2301, n2055, n2513, n1973);
xor  g3434 (n3443, n2658, n2489, n2008, n2043);
xor  g3435 (n3372, n2157, n2516, n2417, n2097);
or   g3436 (n3356, n2061, n2154, n2457, n2025);
nand g3437 (n3017, n2575, n2243, n1996, n2478);
nor  g3438 (n2746, n2090, n2123, n2194, n2473);
xnor g3439 (n3195, n2513, n2639, n2385, n2221);
nand g3440 (n3264, n2434, n2222, n2555, n1152);
or   g3441 (n3654, n2095, n2626, n2258, n2470);
and  g3442 (n3564, n2001, n2651, n2413, n2595);
xor  g3443 (n3166, n2576, n2129, n2663, n2060);
or   g3444 (n3633, n2662, n2285, n2640, n2434);
or   g3445 (n3090, n2060, n2361, n2320, n2113);
nand g3446 (n3036, n2492, n2397, n2331, n2058);
xor  g3447 (n3576, n2192, n2480, n2336, n2517);
or   g3448 (n3276, n2521, n2130, n2085, n2269);
xor  g3449 (n3478, n2559, n2184, n1997, n2526);
nand g3450 (n3559, n2514, n2386, n2063, n2010);
nand g3451 (n3050, n2174, n2361, n2367, n2279);
xor  g3452 (n3629, n2040, n2349, n2400, n2366);
nand g3453 (n3012, n2265, n2421, n2497, n2468);
nor  g3454 (n3355, n2047, n2391, n2442, n2096);
and  g3455 (n3398, n2232, n2365, n2217, n2417);
xnor g3456 (n3376, n2194, n2063, n2268, n2473);
nand g3457 (n3116, n2111, n2213, n2401, n2604);
nor  g3458 (n3452, n2519, n2175, n2529, n2116);
nor  g3459 (n3685, n1986, n2463, n2392, n2608);
or   g3460 (n3106, n2455, n2267, n2030, n2530);
or   g3461 (n3196, n2242, n1974, n2514, n2085);
xor  g3462 (n2692, n2626, n2196, n1980, n2108);
nand g3463 (n3491, n2324, n2144, n2341, n2450);
xnor g3464 (n3638, n2310, n2581, n2343, n2355);
xor  g3465 (n2896, n2469, n2672, n2141, n2321);
xor  g3466 (n3297, n2153, n2094, n2445, n2097);
xnor g3467 (n2898, n2067, n2215, n2164, n2384);
nand g3468 (n2903, n2351, n2203, n2668, n2647);
nand g3469 (n3618, n2442, n2620, n2292, n2405);
and  g3470 (n3688, n2438, n2056, n2265, n2028);
nand g3471 (n2852, n2233, n2572, n2363, n2280);
and  g3472 (n2884, n2361, n2315, n1973, n2377);
xor  g3473 (n3673, n2170, n2244, n2561, n2656);
nand g3474 (n3257, n2029, n2277, n2068, n2197);
and  g3475 (n2980, n2095, n2139, n2322, n2652);
or   g3476 (n2981, n2627, n2559, n2644, n2655);
and  g3477 (n3595, n2444, n2162, n2065, n2464);
xor  g3478 (n3531, n2419, n1970, n2599, n2298);
nand g3479 (n3403, n2160, n1997, n2253, n2490);
and  g3480 (n2733, n2656, n2612, n2552, n2193);
and  g3481 (n3086, n2153, n2251, n2042, n2489);
or   g3482 (n3568, n2112, n2268, n2133, n2044);
xor  g3483 (n3582, n2193, n2144, n2667, n2376);
xor  g3484 (n3130, n2424, n2154, n2245, n2456);
or   g3485 (n3102, n2639, n2493, n2566, n2475);
nor  g3486 (n3006, n2138, n2671, n2201, n1725);
or   g3487 (n3350, n2465, n2194, n2510, n2147);
and  g3488 (n2957, n2307, n2579, n2215, n2279);
xnor g3489 (n3285, n2126, n2280, n2600, n2259);
xnor g3490 (n3406, n2485, n2259, n2107, n2083);
xnor g3491 (n3302, n2642, n2240, n2005, n2415);
nand g3492 (n2703, n2486, n2665, n2004, n2657);
nor  g3493 (n3475, n2501, n2000, n2329, n2163);
xor  g3494 (n3089, n2346, n2184, n1994, n2500);
and  g3495 (n3023, n2105, n2589, n2657, n2353);
or   g3496 (n3561, n2656, n1992, n2359, n1990);
and  g3497 (n3005, n2483, n1973, n2152, n1974);
nand g3498 (n3361, n2132, n2500, n2622, n2236);
or   g3499 (n3615, n2346, n2087, n2380, n2040);
or   g3500 (n3122, n2381, n2299, n2467, n1976);
and  g3501 (n3347, n2459, n2532, n2386, n2606);
xor  g3502 (n3656, n2124, n2393, n2311, n2452);
or   g3503 (n3161, n2286, n2035, n2291, n2317);
xor  g3504 (n2783, n1985, n2522, n2145, n2357);
and  g3505 (n2837, n2308, n2182, n1979, n2334);
nand g3506 (n2920, n2308, n2262, n2508, n2470);
nand g3507 (n3642, n2547, n2272, n2391, n2362);
or   g3508 (n3051, n2305, n2388, n2608, n2248);
nand g3509 (n3583, n2294, n2445, n2126, n2613);
xnor g3510 (n3417, n2044, n2416, n2259, n2275);
xor  g3511 (n3359, n2235, n2271, n2155, n1972);
or   g3512 (n3674, n2344, n2628, n2269, n2662);
and  g3513 (n2876, n2542, n2419, n2555, n2057);
xnor g3514 (n3514, n160, n2080, n2614, n2147);
and  g3515 (n3260, n2285, n2260, n2102, n2287);
or   g3516 (n2825, n2416, n2146, n2145, n2628);
and  g3517 (n3118, n2631, n2329, n2636, n2141);
nor  g3518 (n3680, n2348, n2165, n2074, n2390);
or   g3519 (n3415, n2103, n2484, n2451, n2225);
xor  g3520 (n3065, n2004, n2176, n2011, n2379);
xor  g3521 (n3056, n1982, n2426, n2583, n2334);
xnor g3522 (n2704, n2088, n2232, n2321, n2586);
or   g3523 (n3220, n2645, n2666, n2477, n2558);
xnor g3524 (n3278, n2404, n2014, n2140, n2164);
or   g3525 (n2725, n2342, n2480, n2263, n2088);
nand g3526 (n3190, n2521, n2382, n2204, n2150);
xnor g3527 (n2836, n2080, n2667, n2618, n2508);
xor  g3528 (n3310, n2444, n2013, n2437, n2256);
or   g3529 (n3377, n2079, n2252, n2544, n2383);
nor  g3530 (n2747, n2297, n2587, n2219, n2517);
xnor g3531 (n2972, n2590, n2077, n2508, n2668);
and  g3532 (n3246, n2112, n2551, n2282, n2319);
xor  g3533 (n3340, n2504, n2655, n2226, n2163);
or   g3534 (n3532, n2056, n2427, n2015, n2202);
and  g3535 (n3485, n2347, n2016, n2553, n2361);
and  g3536 (n3303, n2179, n2414, n2413, n2109);
xor  g3537 (n3570, n2031, n2489, n1989, n2582);
or   g3538 (n2921, n2180, n2343, n2246, n2415);
xor  g3539 (n3204, n2198, n2015, n2602, n2236);
xnor g3540 (n3672, n2585, n2492, n2542, n2638);
nor  g3541 (n3043, n2129, n1971, n2133, n2046);
nor  g3542 (n2760, n2653, n1975, n2635, n2303);
or   g3543 (n3387, n2100, n2019, n1971, n2131);
and  g3544 (n2674, n2471, n1981, n2303, n2120);
or   g3545 (n3639, n2026, n2121, n2068, n2562);
xor  g3546 (n2780, n2327, n2151, n1991, n2093);
xor  g3547 (n3609, n2195, n2102, n2371, n2348);
nand g3548 (n3678, n2639, n2131, n2544, n2164);
xnor g3549 (n3530, n2603, n2179, n2500, n2380);
or   g3550 (n2803, n2169, n2637, n2511, n2609);
and  g3551 (n3330, n2408, n2078, n2587, n2282);
nand g3552 (n3213, n2204, n2013, n2594, n2227);
or   g3553 (n3058, n2582, n2155, n2621, n2239);
nor  g3554 (n3147, n2185, n2293, n2254, n2104);
xnor g3555 (n3383, n2494, n2180, n2134, n2173);
or   g3556 (n2685, n2402, n2498, n2213, n2383);
nand g3557 (n3209, n2241, n2540, n2247, n2571);
xnor g3558 (n2971, n2441, n2222, n2459, n2008);
nor  g3559 (n3227, n2069, n2503, n2474, n2306);
xor  g3560 (n3512, n2668, n2578, n2569, n2051);
or   g3561 (n2834, n2399, n2232, n2655, n2171);
or   g3562 (n3061, n2066, n2649, n2652, n2375);
xor  g3563 (n2805, n2406, n2573, n2643, n2623);
xor  g3564 (n3360, n2597, n2359, n2550, n2618);
nand g3565 (n3109, n2496, n2506, n2082, n2557);
or   g3566 (n3524, n2138, n2507, n2428, n2120);
and  g3567 (n3187, n2387, n2589, n2377, n2430);
nor  g3568 (n2773, n2096, n2325, n2433, n2574);
xor  g3569 (n3542, n2595, n2070, n2001, n2593);
xnor g3570 (n2787, n2605, n2177, n2524, n2253);
and  g3571 (n3626, n2625, n2417, n2534, n2403);
nor  g3572 (n3523, n1977, n2086, n2072, n2575);
xnor g3573 (n2902, n2569, n2175, n2223, n2647);
nor  g3574 (n3041, n2157, n2601, n2496, n2369);
or   g3575 (n2932, n2207, n2323, n2335, n2174);
xor  g3576 (n2856, n2515, n2661, n2114, n2235);
nand g3577 (n3032, n2251, n2502, n2562, n2200);
nand g3578 (n3141, n2099, n2640, n2466, n2658);
and  g3579 (n3664, n2133, n2545, n2061, n2320);
or   g3580 (n2699, n2274, n2462, n2320, n2171);
xor  g3581 (n3218, n2370, n2294, n2601, n2538);
and  g3582 (n3358, n2087, n2271, n2252, n2525);
xnor g3583 (n3119, n2208, n2355, n2602, n2151);
and  g3584 (n3381, n2208, n2215, n2406, n2311);
xor  g3585 (n3554, n2269, n2072, n2486, n2654);
or   g3586 (n2705, n2437, n2007, n2026, n2596);
nand g3587 (n3185, n2288, n1971, n1982, n2651);
nor  g3588 (n3048, n2487, n2166, n2218, n2454);
or   g3589 (n2742, n2115, n2168, n1998, n2401);
nor  g3590 (n3280, n2062, n2396, n2111, n1969);
nand g3591 (n3382, n2042, n2667, n2545, n2049);
nor  g3592 (n3581, n2402, n2025, n2004, n2250);
and  g3593 (n3318, n2501, n2027, n2430, n2248);
xnor g3594 (n3594, n2053, n2155, n2304, n2008);
nand g3595 (n3613, n2332, n2422, n2074, n2612);
or   g3596 (n2678, n2526, n2005, n2297, n2221);
nand g3597 (n3200, n2392, n2192, n2329, n2047);
or   g3598 (n3107, n2165, n2616, n2328, n2500);
xnor g3599 (n3083, n2123, n2050, n2540, n2548);
xnor g3600 (n2822, n2411, n2573, n2021, n2560);
or   g3601 (n3228, n2476, n2303, n2211, n2556);
xnor g3602 (n3413, n2078, n2475, n2410, n1970);
and  g3603 (n3573, n2234, n2024, n2270, n2250);
nor  g3604 (n3095, n2003, n2455, n2452, n2622);
or   g3605 (n2928, n2056, n2032, n2226, n1972);
and  g3606 (n2996, n2313, n2102, n2238, n2446);
nand g3607 (n3216, n2412, n2435, n2080, n1989);
and  g3608 (n2917, n2118, n2443, n2655, n2382);
nand g3609 (n3284, n2605, n2356, n2110, n2204);
nand g3610 (n3558, n2549, n2322, n2031, n2542);
xnor g3611 (n2906, n2224, n2232, n2625, n2495);
nand g3612 (n3643, n2458, n2197, n2484, n2277);
or   g3613 (n3397, n2633, n2226, n1987, n2047);
and  g3614 (n2844, n2398, n1977, n2156, n2505);
or   g3615 (n2712, n2343, n2609, n2137, n2237);
and  g3616 (n3631, n2163, n2488, n2077, n2474);
nor  g3617 (n3078, n2326, n2217, n2072, n2423);
or   g3618 (n2927, n2402, n2560, n2111, n2054);
xor  g3619 (n3543, n2347, n2554, n2284, n2142);
or   g3620 (n3574, n2010, n2041, n2172, n2404);
nor  g3621 (n2764, n2583, n2258, n2255, n2567);
and  g3622 (n3540, n2050, n1987, n2492, n2434);
nand g3623 (n2987, n2357, n2364, n2125, n2213);
and  g3624 (n3572, n2096, n2475, n2548, n2354);
xor  g3625 (n2913, n2395, n2039, n2575, n2496);
and  g3626 (n2693, n2530, n2587, n2319, n2544);
nand g3627 (n3363, n2015, n2162, n2081, n2058);
xnor g3628 (n2755, n2583, n2324, n2638, n2017);
nor  g3629 (n3314, n2539, n1725, n2060, n2611);
xnor g3630 (n3448, n2418, n2034, n2145, n2007);
xnor g3631 (n2714, n2294, n2660, n2494, n2650);
xnor g3632 (n2694, n2627, n2350, n2136, n2414);
xnor g3633 (n3569, n2555, n2048, n2195, n2002);
or   g3634 (n3007, n2431, n2400, n2646, n2140);
nor  g3635 (n3252, n2561, n2081, n2277, n2582);
or   g3636 (n3521, n2059, n2330, n2649, n2354);
or   g3637 (n2863, n2385, n2076, n2092, n2407);
or   g3638 (n3154, n1992, n2156, n2379, n2623);
nor  g3639 (n2821, n2616, n2663, n2531, n2267);
xor  g3640 (n3060, n2547, n2394, n2035, n2342);
xnor g3641 (n2756, n2288, n2493, n2257, n2556);
xnor g3642 (n3153, n2215, n2187, n2186, n2146);
nor  g3643 (n3126, n2614, n1978, n2441, n2313);
nor  g3644 (n3663, n2666, n2341, n2033, n2005);
nor  g3645 (n2835, n2135, n2531, n2536, n2565);
xnor g3646 (n3527, n2188, n2283, n2612, n2327);
or   g3647 (n3002, n1990, n2283, n2241, n2323);
xnor g3648 (n2829, n2055, n2071, n2518, n2255);
or   g3649 (n3030, n2400, n2396, n2104, n2612);
and  g3650 (n3546, n2659, n2598, n2066, n2397);
or   g3651 (n2811, n2329, n2287, n2191, n2637);
and  g3652 (n2916, n2240, n2178, n2350, n2304);
nand g3653 (n3409, n2348, n2631, n2185, n2438);
xnor g3654 (n3180, n2014, n2231, n2388, n2325);
or   g3655 (n3380, n2340, n2632, n2039, n2638);
or   g3656 (n3605, n2167, n1989, n2386, n2411);
nand g3657 (n2973, n2616, n2038, n2603, n2550);
xnor g3658 (n3022, n2508, n2512, n2481, n2628);
nor  g3659 (n3846, n3157, n3579, n2919, n3653);
xor  g3660 (n3826, n3041, n3318, n3283, n2941);
or   g3661 (n3921, n2835, n3369, n2925, n3547);
nor  g3662 (n3861, n3396, n2871, n3247, n2860);
xnor g3663 (n3791, n3432, n3486, n2734, n3112);
xnor g3664 (n3831, n3201, n3429, n3515, n2795);
and  g3665 (n3919, n3505, n2720, n3365, n3359);
and  g3666 (n3825, n3550, n3402, n3648, n3049);
xnor g3667 (n3705, n3634, n3578, n3100, n3356);
and  g3668 (n3816, n3458, n3424, n3035, n1156);
nor  g3669 (n3761, n3339, n2740, n3358, n2881);
and  g3670 (n3813, n2966, n3683, n3421, n3021);
xnor g3671 (n3827, n3073, n3517, n3186, n3127);
nand g3672 (n3901, n3573, n3625, n3665, n3563);
and  g3673 (n3867, n3596, n3109, n3604, n2764);
xor  g3674 (n3693, n3471, n3128, n3328, n2710);
and  g3675 (n3805, n3137, n3162, n3158, n2991);
and  g3676 (n3737, n2873, n3262, n3067, n2988);
and  g3677 (n3771, n2984, n2797, n3628, n2981);
or   g3678 (n3824, n2895, n3131, n2975, n3587);
nor  g3679 (n3923, n2690, n3263, n2911, n2728);
xnor g3680 (n3702, n3541, n3534, n3110, n3267);
xor  g3681 (n3763, n3626, n2769, n3388, n3172);
nand g3682 (n3893, n3450, n3274, n2800, n3592);
nor  g3683 (n3830, n3609, n3643, n2942, n3619);
nor  g3684 (n3767, n3005, n3046, n3491, n3030);
xor  g3685 (n3730, n2774, n3667, n3446, n3302);
xor  g3686 (n3868, n3558, n2808, n3122, n3232);
and  g3687 (n3853, n3497, n2688, n3160, n3449);
nand g3688 (n3741, n3464, n2711, n2922, n3200);
and  g3689 (n3880, n2807, n3617, n2707, n2876);
or   g3690 (n3806, n3395, n3567, n3312, n3176);
xnor g3691 (n3896, n3593, n2824, n3639, n2888);
nor  g3692 (n3872, n2719, n2915, n3011, n3144);
nand g3693 (n3745, n3173, n2683, n3528, n3164);
xnor g3694 (n3715, n2940, n3299, n3152, n2947);
nor  g3695 (n3821, n3509, n3616, n3083, n3612);
xor  g3696 (n3822, n3280, n2977, n3048, n1155);
xor  g3697 (n3938, n2801, n2994, n3469, n3300);
xnor g3698 (n3696, n3437, n3430, n2892, n3641);
xor  g3699 (n3749, n2777, n3384, n3661, n2717);
nand g3700 (n3738, n3598, n2883, n3036, n3649);
or   g3701 (n3905, n2681, n3080, n2877, n3107);
nand g3702 (n3692, n3051, n3602, n3198, n2902);
xor  g3703 (n3753, n3346, n3583, n3423, n2741);
nand g3704 (n3908, n2843, n3669, n2833, n2898);
xor  g3705 (n3823, n3405, n3595, n2909, n3624);
nor  g3706 (n3764, n2766, n3495, n2920, n3039);
xor  g3707 (n3852, n2682, n3079, n2775, n3679);
nand g3708 (n3718, n2901, n3009, n3268, n3484);
nand g3709 (n3708, n2897, n2936, n3307, n2948);
nand g3710 (n3719, n3234, n3203, n2862, n2803);
nor  g3711 (n3910, n2692, n3310, n3655, n3088);
nand g3712 (n3784, n3305, n3472, n2964, n3143);
xor  g3713 (n3781, n3062, n3650, n3306, n3297);
xnor g3714 (n3931, n3214, n2930, n3440, n2983);
nand g3715 (n3788, n2864, n3136, n3527, n3332);
nor  g3716 (n3935, n3488, n3452, n3493, n2673);
nor  g3717 (n3726, n2913, n2768, n2950, n2841);
nor  g3718 (n3770, n3411, n3197, n3687, n2910);
xnor g3719 (n3913, n3383, n3293, n2962, n3278);
and  g3720 (n3841, n2933, n3363, n2890, n3185);
nand g3721 (n3717, n3545, n3013, n3644, n3415);
nor  g3722 (n3716, n2736, n3585, n3081, n2802);
xor  g3723 (n3774, n2928, n3148, n3058, n2995);
nand g3724 (n3725, n3668, n3174, n2997, n3499);
or   g3725 (n3890, n3569, n3347, n3000, n3442);
nor  g3726 (n3766, n2973, n2904, n3032, n2754);
xnor g3727 (n3851, n2842, n3673, n3038, n3555);
nor  g3728 (n3734, n3364, n2989, n3019, n3508);
or   g3729 (n3817, n3553, n3150, n2786, n3237);
or   g3730 (n3814, n2693, n2951, n3231, n3163);
or   g3731 (n3721, n3489, n3529, n2675, n3003);
xor  g3732 (n3916, n3542, n3235, n2771, n3105);
nor  g3733 (n3808, n2882, n3253, n2755, n3375);
or   g3734 (n3795, n2894, n2870, n3037, n3590);
xnor g3735 (n3724, n3536, n3001, n3108, n3243);
xnor g3736 (n3947, n2861, n3685, n2838, n3480);
nor  g3737 (n3906, n3129, n3091, n2739, n2779);
xnor g3738 (n3862, n3465, n3582, n3256, n2935);
xnor g3739 (n3800, n2931, n2684, n3304, n3457);
or   g3740 (n3902, n3010, n3360, n2691, n3290);
xor  g3741 (n3865, n3059, n3504, n2980, n3398);
or   g3742 (n3903, n2794, n3654, n3317, n3345);
nor  g3743 (n3731, n3277, n3689, n2853, n2694);
xor  g3744 (n3869, n3169, n2970, n3324, n2831);
and  g3745 (n3836, n2763, n2799, n3171, n3140);
nand g3746 (n3927, n2677, n3281, n3540, n3351);
xnor g3747 (n3765, n2954, n3225, n2722, n2963);
nor  g3748 (n3915, n3621, n2697, n2784, n3184);
xor  g3749 (n3797, n3258, n3089, n3434, n3546);
xor  g3750 (n3735, n3187, n2958, n3390, n3223);
and  g3751 (n3727, n3586, n2818, n3327, n2780);
xnor g3752 (n3899, n2965, n3314, n3287, n2709);
xnor g3753 (n3736, n3024, n3463, n2804, n3221);
nor  g3754 (n3850, n3334, n3647, n3678, n3603);
or   g3755 (n3842, n3142, n3126, n3266, n1153);
xnor g3756 (n3875, n3132, n2701, n3113, n2715);
or   g3757 (n3942, n2772, n2891, n3551, n3584);
nand g3758 (n3818, n3072, n3608, n2937, n2686);
nor  g3759 (n3754, n3566, n2678, n3543, n3260);
or   g3760 (n3946, n3660, n3286, n3279, n3168);
nand g3761 (n3828, n3194, n3211, n3349, n3412);
and  g3762 (n3874, n3404, n3382, n2744, n3094);
and  g3763 (n3837, n3613, n3228, n2749, n3439);
and  g3764 (n3709, n3510, n3216, n3156, n3213);
and  g3765 (n3720, n2730, n3677, n3554, n3418);
and  g3766 (n3897, n3076, n3385, n3012, n2817);
or   g3767 (n3739, n3645, n2943, n2745, n3063);
nand g3768 (n3887, n2836, n3664, n2858, n2792);
and  g3769 (n3809, n3294, n3022, n3193, n3614);
nand g3770 (n3891, n3303, n3248, n2905, n3180);
and  g3771 (n3934, n3372, n2986, n2923, n3652);
xnor g3772 (n3710, n2826, n3047, n2696, n2885);
and  g3773 (n3787, n2731, n3182, n3015, n3682);
nand g3774 (n3752, n3065, n2849, n3496, n3154);
nor  g3775 (n3914, n3366, n2729, n3270, n2960);
nor  g3776 (n3932, n3333, n3477, n3672, n2751);
and  g3777 (n3870, n2899, n3224, n2706, n3061);
xnor g3778 (n3885, n2813, n3064, n3670, n2687);
xor  g3779 (n3697, n3289, n3084, n3060, n3101);
xnor g3780 (n3740, n3313, n3007, n3663, n3111);
or   g3781 (n3900, n3120, n3686, n2815, n2753);
xnor g3782 (n3775, n3362, n3427, n3478, n3335);
xnor g3783 (n3712, n3556, n2814, n3570, n3045);
xnor g3784 (n3786, n3519, n3642, n2781, n3078);
nor  g3785 (n3760, n2727, n3119, n3521, n2793);
or   g3786 (n3911, n2934, n3259, n3229, n3539);
nand g3787 (n3698, n2713, n3151, n3097, n3291);
and  g3788 (n3783, n3462, n3227, n3331, n3330);
nand g3789 (n3815, n3134, n3040, n3588, n2773);
xor  g3790 (n3807, n2912, n2982, n3114, n3605);
xnor g3791 (n3796, n2839, n3622, n3371, n3391);
and  g3792 (n3922, n3085, n3295, n3298, n3145);
xnor g3793 (n3839, n3407, n3531, n3657, n3118);
nand g3794 (n3832, n3601, n3638, n3461, n2956);
or   g3795 (n3884, n3524, n2829, n3288, n3627);
xor  g3796 (n3892, n3386, n2938, n2880, n3594);
xor  g3797 (n3776, n3031, n3138, n3336, n2855);
nor  g3798 (n3804, n3219, n3181, n2993, n3431);
nand g3799 (n3819, n2893, n3568, n3075, n2822);
xnor g3800 (n3773, n3629, n2712, n3125, n3139);
nand g3801 (n3713, n1154, n3240, n3376, n3092);
or   g3802 (n3912, n3506, n3296, n2906, n2783);
nor  g3803 (n3943, n3500, n3141, n2828, n3341);
nand g3804 (n3793, n2702, n3204, n2680, n2949);
nand g3805 (n3909, n3321, n2998, n3352, n3435);
or   g3806 (n3742, n3130, n2733, n2825, n3178);
xnor g3807 (n3920, n3257, n3264, n3285, n3238);
nand g3808 (n3729, n3308, n3445, n2752, n2821);
and  g3809 (n3746, n3323, n3271, n2872, n3470);
xnor g3810 (n3873, n3350, n3265, n2689, n3466);
or   g3811 (n3835, n3205, n3244, n3675, n2850);
xor  g3812 (n3700, n2830, n2924, n3018, n2747);
nor  g3813 (n3703, n3436, n3473, n2921, n2874);
nor  g3814 (n3847, n3218, n3475, n3438, n3460);
xnor g3815 (n3706, n2896, n3190, n3241, n2700);
xor  g3816 (n3769, n3146, n3017, n3389, n2714);
xor  g3817 (n3858, n3513, n3183, n2926, n3456);
xor  g3818 (n3782, n2990, n3272, n3153, n3444);
nor  g3819 (n3778, n3410, n3252, n3284, n3206);
xnor g3820 (n3886, n3576, n3514, n3104, n2770);
and  g3821 (n3732, n2889, n2790, n3482, n3215);
xnor g3822 (n3755, n3406, n2732, n2757, n3454);
and  g3823 (n3768, n2699, n3188, n3357, n3467);
xor  g3824 (n3723, n2854, n3526, n3530, n2916);
xor  g3825 (n3871, n3564, n3671, n3618, n2743);
or   g3826 (n3744, n3419, n3319, n3557, n3034);
and  g3827 (n3779, n3422, n3161, n3525, n2834);
xor  g3828 (n3711, n3249, n2791, n3548, n3116);
or   g3829 (n3801, n3106, n3518, n3633, n2978);
nor  g3830 (n3695, n3147, n2999, n3053, n2987);
nor  g3831 (n3803, n3503, n3367, n2789, n3552);
and  g3832 (n3904, n3082, n3490, n3124, n3662);
nor  g3833 (n3895, n3052, n3507, n2868, n3275);
and  g3834 (n3859, n3635, n3315, n3378, n3561);
xnor g3835 (n3882, n3043, n3025, n2875, n3408);
nor  g3836 (n3883, n2782, n3623, n3658, n3413);
and  g3837 (n3860, n3377, n3222, n3646, n2765);
or   g3838 (n3728, n3487, n3233, n3485, n2761);
xor  g3839 (n3881, n3077, n3361, n3026, n3656);
nor  g3840 (n3845, n3399, n2748, n2708, n2927);
and  g3841 (n3937, n3103, n2867, n3170, n3651);
nor  g3842 (n3743, n2846, n2823, n2929, n2725);
and  g3843 (n3944, n3344, n3177, n2816, n3688);
xnor g3844 (n3855, n3433, n2971, n3165, n3607);
nor  g3845 (n3940, n3189, n2738, n2674, n3416);
and  g3846 (n3849, n3571, n3535, n3537, n3403);
xor  g3847 (n3701, n2796, n3343, n3027, n3311);
xor  g3848 (n3857, n3074, n3597, n3276, n3538);
or   g3849 (n3812, n2914, n2840, n3044, n2859);
xor  g3850 (n3933, n3532, n2848, n2723, n3070);
nor  g3851 (n3889, n3549, n2759, n3370, n3212);
xnor g3852 (n3925, n2955, n3455, n3417, n3179);
nor  g3853 (n3810, n3659, n3494, n2827, n3033);
and  g3854 (n3930, n3123, n3202, n3236, n3620);
nand g3855 (n3802, n2967, n3611, n2944, n3441);
nor  g3856 (n3928, n3230, n3498, n3209, n3042);
or   g3857 (n3733, n3068, n3676, n3135, n3600);
nor  g3858 (n3780, n3374, n2985, n3599, n2704);
or   g3859 (n3792, n3023, n3309, n2806, n2820);
and  g3860 (n3840, n3250, n3261, n2884, n3255);
or   g3861 (n3945, n3322, n3028, n3245, n3016);
xnor g3862 (n3924, n3326, n2703, n3337, n3196);
or   g3863 (n3907, n3368, n3580, n2886, n3615);
nand g3864 (n3762, n3159, n3167, n3102, n3589);
xnor g3865 (n3751, n3340, n2992, n2869, n3468);
xnor g3866 (n3704, n3474, n3502, n3666, n3292);
xor  g3867 (n3772, n2845, n3681, n3086, n2837);
xor  g3868 (n3789, n3226, n3426, n3562, n3115);
xor  g3869 (n3799, n3004, n3166, n2852, n2961);
xnor g3870 (n3941, n3149, n3220, n3447, n2932);
xor  g3871 (n3936, n3574, n3353, n3117, n3195);
and  g3872 (n3750, n2785, n3055, n3020, n3636);
xor  g3873 (n3898, n2809, n3640, n2778, n2726);
xor  g3874 (n3829, n3014, n3217, n3459, n3572);
nand g3875 (n3876, n3501, n3071, n3674, n3242);
xor  g3876 (n3777, n3316, n3632, n1157, n3409);
or   g3877 (n3843, n3425, n2756, n3483, n2724);
nand g3878 (n3707, n3175, n3254, n3400, n3325);
xor  g3879 (n3759, n3453, n2716, n2865, n3451);
xor  g3880 (n3747, n2679, n2787, n3251, n3093);
nor  g3881 (n3894, n2788, n3511, n3581, n3575);
nor  g3882 (n3864, n3056, n2812, n2996, n2776);
xor  g3883 (n3866, n2721, n3155, n3192, n2819);
xor  g3884 (n3877, n3520, n3691, n3090, n2957);
nand g3885 (n3794, n3606, n2856, n3479, n3320);
xnor g3886 (n3699, n2844, n3387, n3338, n3373);
nor  g3887 (n3785, n2742, n2939, n2903, n3246);
or   g3888 (n3834, n2758, n3533, n3631, n3057);
xnor g3889 (n3939, n2737, n2676, n3207, n3087);
and  g3890 (n3833, n2695, n2968, n3577, n3420);
xnor g3891 (n3929, n3342, n3329, n2735, n3428);
or   g3892 (n3926, n3684, n3354, n2705, n2878);
xor  g3893 (n3820, n3029, n2750, n3133, n2917);
xor  g3894 (n3918, n2946, n2952, n3680, n3355);
xnor g3895 (n3854, n2974, n2887, n2746, n3099);
xnor g3896 (n3694, n2972, n3544, n3210, n3516);
nor  g3897 (n3811, n3630, n3591, n2866, n3050);
and  g3898 (n3758, n2811, n2760, n3054, n2832);
nor  g3899 (n3879, n3069, n3381, n3008, n3392);
or   g3900 (n3756, n3414, n3199, n3348, n3394);
or   g3901 (n3722, n2718, n3476, n2810, n2959);
or   g3902 (n3838, n3401, n3301, n3273, n3121);
nor  g3903 (n3714, n3443, n2805, n3208, n2847);
and  g3904 (n3888, n3096, n2685, n2851, n3095);
nor  g3905 (n3917, n2976, n2900, n3448, n3610);
xor  g3906 (n3798, n3379, n3002, n2863, n2857);
xnor g3907 (n3863, n2762, n2798, n2907, n3098);
and  g3908 (n3790, n2879, n3522, n3380, n2918);
xnor g3909 (n3856, n3239, n3282, n3523, n2969);
nand g3910 (n3748, n3481, n2767, n3560, n3393);
xor  g3911 (n3844, n3397, n3559, n3512, n3191);
nand g3912 (n3878, n3269, n2953, n2908, n3006);
xor  g3913 (n3757, n2979, n3690, n3637, n3565);
or   g3914 (n3848, n3492, n2945, n3066, n2698);
nand g3915 (n3971, n3750, n3920, n3935, n3832);
nand g3916 (n3950, n3835, n3918, n3851, n3890);
nand g3917 (n3978, n3849, n3757, n3824, n3933);
and  g3918 (n3958, n3836, n3705, n3777, n3816);
nand g3919 (n3998, n3938, n3780, n3891, n3895);
nand g3920 (n4002, n3826, n3742, n3919, n3857);
nand g3921 (n3962, n3697, n3756, n3866, n3788);
or   g3922 (n3973, n3894, n3865, n3770, n3765);
xor  g3923 (n3994, n3696, n3781, n3889, n3707);
xnor g3924 (n3997, n3872, n3898, n3809, n3787);
xnor g3925 (n3975, n3734, n3699, n3821, n3860);
nand g3926 (n3948, n3846, n3772, n3917, n3764);
xnor g3927 (n3949, n3875, n3928, n3897, n3701);
or   g3928 (n3951, n3910, n3845, n3758, n3747);
xnor g3929 (n3979, n3873, n3947, n3899, n3823);
or   g3930 (n3974, n3753, n3830, n3859, n3703);
or   g3931 (n3982, n3794, n3829, n3804, n3748);
xnor g3932 (n3990, n3706, n3901, n3905, n3762);
nor  g3933 (n3986, n3767, n3833, n3736, n3793);
or   g3934 (n3989, n3730, n3783, n3911, n3914);
nand g3935 (n3963, n3774, n3896, n3912, n3800);
nor  g3936 (n4004, n3798, n3723, n3749, n3863);
nor  g3937 (n4010, n3884, n3881, n3892, n3729);
or   g3938 (n3985, n3864, n3796, n3805, n3942);
or   g3939 (n4003, n3934, n3907, n3871, n3822);
xor  g3940 (n3996, n3808, n3944, n3848, n3810);
xnor g3941 (n3961, n3817, n3751, n3925, n3778);
xor  g3942 (n3968, n3718, n3888, n3819, n3929);
nand g3943 (n3952, n3714, n3802, n3876, n3930);
and  g3944 (n3955, n3874, n3710, n3854, n3923);
nor  g3945 (n3959, n3728, n3885, n3725, n3791);
nand g3946 (n3987, n3715, n3939, n3921, n3893);
or   g3947 (n4000, n3784, n3858, n3775, n3702);
nand g3948 (n3969, n3763, n3735, n3932, n3722);
or   g3949 (n4001, n3838, n3856, n3904, n3852);
nand g3950 (n3970, n3877, n3727, n3806, n3946);
nor  g3951 (n3995, n3744, n3713, n3732, n3708);
xnor g3952 (n4006, n3766, n3882, n3692, n3769);
xor  g3953 (n4009, n3746, n3868, n3820, n3878);
nand g3954 (n4008, n3719, n3782, n3731, n3711);
and  g3955 (n3954, n3724, n3937, n3790, n3799);
nand g3956 (n3965, n3717, n3936, n3844, n3902);
xor  g3957 (n3984, n3839, n3721, n3903, n3738);
xnor g3958 (n3999, n3698, n3807, n3842, n3789);
nor  g3959 (n3957, n3941, n3900, n3726, n3869);
nand g3960 (n3964, n3841, n3908, n3840, n3818);
nor  g3961 (n3966, n3827, n3879, n3915, n3834);
nor  g3962 (n3988, n3931, n3814, n3704, n3922);
xnor g3963 (n4011, n3940, n3752, n3795, n3924);
xor  g3964 (n3960, n3855, n3825, n3786, n3880);
nand g3965 (n3980, n3755, n3740, n3785, n3733);
or   g3966 (n3977, n3712, n3813, n3760, n3926);
xnor g3967 (n3992, n3745, n3803, n3837, n3945);
nor  g3968 (n3993, n3916, n3709, n3870, n3913);
xor  g3969 (n3991, n3847, n3853, n3759, n3861);
or   g3970 (n3981, n3797, n3883, n3815, n3720);
xnor g3971 (n3967, n3850, n3743, n3828, n3862);
or   g3972 (n3983, n3754, n3739, n3779, n3700);
xnor g3973 (n4007, n3843, n3906, n3887, n3801);
xor  g3974 (n3976, n3773, n3792, n3693, n3695);
and  g3975 (n3956, n3886, n3741, n3694, n3776);
xnor g3976 (n3953, n3867, n3927, n3811, n3909);
xnor g3977 (n4005, n3831, n3943, n3812, n3771);
or   g3978 (n3972, n3716, n3761, n3737, n3768);
nor  g3979 (n4013, n3992, n3991, n4010, n3966);
xor  g3980 (n4025, n4005, n3965, n3950, n4011);
or   g3981 (n4012, n4002, n3974, n3997, n3964);
and  g3982 (n4018, n3988, n3998, n3952, n3956);
and  g3983 (n4024, n3973, n3979, n3986, n4008);
xor  g3984 (n4021, n3962, n3954, n3983, n3949);
nor  g3985 (n4022, n3959, n3957, n3978, n3996);
nor  g3986 (n4027, n3955, n3984, n3977, n3963);
xor  g3987 (n4014, n3995, n3980, n3953, n3967);
nand g3988 (n4015, n3960, n3972, n4001, n4003);
and  g3989 (n4019, n3971, n3975, n3982, n3970);
nor  g3990 (n4017, n3951, n4006, n3976, n4004);
xnor g3991 (n4020, n3999, n4009, n3969, n3985);
nor  g3992 (n4016, n3994, n4007, n3989, n3993);
xor  g3993 (n4023, n3990, n3958, n3987, n3968);
xor  g3994 (n4026, n3948, n3961, n3981, n4000);
nor  g3995 (n4030, n4013, n4026, n4021, n4018);
nand g3996 (n4031, n4016, n4022, n4024, n4015);
xnor g3997 (n4029, n4014, n4019, n4023, n4027);
and  g3998 (n4028, n4025, n4017, n4020, n4012);
and  g3999 (n4032, n4028, n4029, n4030, n4031);
endmodule
