

module Stat_2000_226
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n739,
  n715,
  n1183,
  n1173,
  n1169,
  n1179,
  n1175,
  n1194,
  n1188,
  n1196,
  n1177,
  n1185,
  n1167,
  n1187,
  n1408,
  n1424,
  n1412,
  n1418,
  n1423,
  n1395,
  n1425,
  n1403,
  n1396,
  n1401,
  n1397,
  n1393,
  n1426,
  n1415,
  n1411,
  n1406,
  n2031,
  n2032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n739;
  output n715;
  output n1183;
  output n1173;
  output n1169;
  output n1179;
  output n1175;
  output n1194;
  output n1188;
  output n1196;
  output n1177;
  output n1185;
  output n1167;
  output n1187;
  output n1408;
  output n1424;
  output n1412;
  output n1418;
  output n1423;
  output n1395;
  output n1425;
  output n1403;
  output n1396;
  output n1401;
  output n1397;
  output n1393;
  output n1426;
  output n1415;
  output n1411;
  output n1406;
  output n2031;
  output n2032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1168;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1174;
  wire n1176;
  wire n1178;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1184;
  wire n1186;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1195;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1394;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1402;
  wire n1404;
  wire n1405;
  wire n1407;
  wire n1409;
  wire n1410;
  wire n1413;
  wire n1414;
  wire n1416;
  wire n1417;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n80,
    n32
  );


  buf
  g1
  (
    n36,
    n4
  );


  not
  g2
  (
    n35,
    n20
  );


  not
  g3
  (
    n92,
    n28
  );


  buf
  g4
  (
    n34,
    n15
  );


  buf
  g5
  (
    n58,
    n23
  );


  buf
  g6
  (
    n67,
    n7
  );


  not
  g7
  (
    n123,
    n16
  );


  not
  g8
  (
    n158,
    n1
  );


  buf
  g9
  (
    KeyWire_0_11,
    n6
  );


  buf
  g10
  (
    n127,
    n32
  );


  not
  g11
  (
    n82,
    n10
  );


  not
  g12
  (
    n39,
    n12
  );


  not
  g13
  (
    KeyWire_0_0,
    n1
  );


  not
  g14
  (
    n68,
    n8
  );


  buf
  g15
  (
    n33,
    n22
  );


  not
  g16
  (
    n156,
    n17
  );


  not
  g17
  (
    n72,
    n10
  );


  buf
  g18
  (
    n97,
    n24
  );


  not
  g19
  (
    n77,
    n14
  );


  buf
  g20
  (
    n154,
    n11
  );


  buf
  g21
  (
    n87,
    n11
  );


  buf
  g22
  (
    n139,
    n3
  );


  not
  g23
  (
    n116,
    n2
  );


  buf
  g24
  (
    n69,
    n19
  );


  not
  g25
  (
    n151,
    n29
  );


  not
  g26
  (
    n132,
    n16
  );


  not
  g27
  (
    n101,
    n3
  );


  buf
  g28
  (
    n88,
    n7
  );


  buf
  g29
  (
    n38,
    n20
  );


  buf
  g30
  (
    n118,
    n24
  );


  not
  g31
  (
    n112,
    n3
  );


  buf
  g32
  (
    n145,
    n25
  );


  not
  g33
  (
    n100,
    n26
  );


  buf
  g34
  (
    n138,
    n12
  );


  not
  g35
  (
    n147,
    n20
  );


  not
  g36
  (
    n81,
    n5
  );


  buf
  g37
  (
    n129,
    n31
  );


  buf
  g38
  (
    n160,
    n9
  );


  not
  g39
  (
    n61,
    n14
  );


  not
  g40
  (
    n109,
    n27
  );


  buf
  g41
  (
    n78,
    n2
  );


  buf
  g42
  (
    n65,
    n7
  );


  buf
  g43
  (
    n89,
    n9
  );


  not
  g44
  (
    n152,
    n8
  );


  not
  g45
  (
    n55,
    n21
  );


  not
  g46
  (
    n153,
    n10
  );


  not
  g47
  (
    n108,
    n17
  );


  buf
  g48
  (
    n90,
    n25
  );


  not
  g49
  (
    n50,
    n23
  );


  not
  g50
  (
    n121,
    n29
  );


  buf
  g51
  (
    n111,
    n19
  );


  not
  g52
  (
    n45,
    n17
  );


  not
  g53
  (
    n110,
    n28
  );


  buf
  g54
  (
    n122,
    n31
  );


  not
  g55
  (
    n49,
    n9
  );


  buf
  g56
  (
    n75,
    n31
  );


  buf
  g57
  (
    n143,
    n25
  );


  not
  g58
  (
    n119,
    n5
  );


  not
  g59
  (
    n157,
    n26
  );


  not
  g60
  (
    n128,
    n14
  );


  not
  g61
  (
    n98,
    n22
  );


  not
  g62
  (
    n148,
    n4
  );


  not
  g63
  (
    n79,
    n24
  );


  buf
  g64
  (
    n76,
    n15
  );


  buf
  g65
  (
    n142,
    n18
  );


  not
  g66
  (
    n43,
    n21
  );


  not
  g67
  (
    n117,
    n10
  );


  buf
  g68
  (
    n94,
    n22
  );


  buf
  g69
  (
    n124,
    n28
  );


  not
  g70
  (
    n113,
    n32
  );


  buf
  g71
  (
    n74,
    n2
  );


  not
  g72
  (
    n93,
    n24
  );


  not
  g73
  (
    n115,
    n29
  );


  buf
  g74
  (
    n137,
    n26
  );


  not
  g75
  (
    n114,
    n14
  );


  not
  g76
  (
    n63,
    n18
  );


  not
  g77
  (
    n99,
    n13
  );


  buf
  g78
  (
    n103,
    n26
  );


  not
  g79
  (
    n107,
    n11
  );


  not
  g80
  (
    n136,
    n5
  );


  not
  g81
  (
    n125,
    n18
  );


  not
  g82
  (
    n85,
    n4
  );


  buf
  g83
  (
    n53,
    n29
  );


  buf
  g84
  (
    n149,
    n9
  );


  buf
  g85
  (
    n71,
    n4
  );


  buf
  g86
  (
    n130,
    n6
  );


  buf
  g87
  (
    n84,
    n23
  );


  not
  g88
  (
    n54,
    n15
  );


  buf
  g89
  (
    n150,
    n1
  );


  buf
  g90
  (
    n83,
    n32
  );


  buf
  g91
  (
    n140,
    n7
  );


  buf
  g92
  (
    n70,
    n16
  );


  buf
  g93
  (
    n41,
    n28
  );


  not
  g94
  (
    n133,
    n12
  );


  not
  g95
  (
    n59,
    n19
  );


  not
  g96
  (
    n47,
    n13
  );


  buf
  g97
  (
    n52,
    n11
  );


  not
  g98
  (
    n56,
    n6
  );


  buf
  g99
  (
    n51,
    n15
  );


  not
  g100
  (
    n126,
    n30
  );


  not
  g101
  (
    n106,
    n2
  );


  not
  g102
  (
    n96,
    n21
  );


  buf
  g103
  (
    n134,
    n19
  );


  not
  g104
  (
    n46,
    n8
  );


  buf
  g105
  (
    n44,
    n13
  );


  not
  g106
  (
    n42,
    n30
  );


  not
  g107
  (
    n104,
    n22
  );


  not
  g108
  (
    n91,
    n5
  );


  buf
  g109
  (
    n73,
    n1
  );


  buf
  g110
  (
    n135,
    n3
  );


  not
  g111
  (
    n64,
    n21
  );


  not
  g112
  (
    n105,
    n25
  );


  not
  g113
  (
    n48,
    n18
  );


  not
  g114
  (
    n120,
    n16
  );


  not
  g115
  (
    n141,
    n12
  );


  buf
  g116
  (
    n131,
    n27
  );


  not
  g117
  (
    n57,
    n30
  );


  not
  g118
  (
    n37,
    n20
  );


  not
  g119
  (
    n95,
    n30
  );


  not
  g120
  (
    n60,
    n17
  );


  buf
  g121
  (
    n40,
    n6
  );


  buf
  g122
  (
    n144,
    n23
  );


  buf
  g123
  (
    n159,
    n8
  );


  buf
  g124
  (
    n66,
    n31
  );


  buf
  g125
  (
    n155,
    n27
  );


  buf
  g126
  (
    n102,
    n27
  );


  not
  g127
  (
    n86,
    n13
  );


  not
  g128
  (
    n292,
    n97
  );


  not
  g129
  (
    n227,
    n143
  );


  not
  g130
  (
    n652,
    n36
  );


  not
  g131
  (
    n593,
    n46
  );


  not
  g132
  (
    n226,
    n33
  );


  buf
  g133
  (
    n286,
    n58
  );


  buf
  g134
  (
    n208,
    n113
  );


  not
  g135
  (
    n329,
    n39
  );


  not
  g136
  (
    n231,
    n50
  );


  buf
  g137
  (
    n243,
    n119
  );


  buf
  g138
  (
    n238,
    n76
  );


  buf
  g139
  (
    n449,
    n123
  );


  buf
  g140
  (
    n589,
    n147
  );


  buf
  g141
  (
    n366,
    n65
  );


  not
  g142
  (
    n453,
    n66
  );


  not
  g143
  (
    n300,
    n151
  );


  not
  g144
  (
    n585,
    n33
  );


  buf
  g145
  (
    n565,
    n153
  );


  buf
  g146
  (
    n483,
    n77
  );


  buf
  g147
  (
    n256,
    n159
  );


  not
  g148
  (
    n628,
    n60
  );


  buf
  g149
  (
    n202,
    n47
  );


  not
  g150
  (
    n295,
    n37
  );


  buf
  g151
  (
    n450,
    n114
  );


  not
  g152
  (
    n595,
    n100
  );


  not
  g153
  (
    n323,
    n101
  );


  buf
  g154
  (
    n327,
    n113
  );


  not
  g155
  (
    n291,
    n110
  );


  not
  g156
  (
    n415,
    n126
  );


  not
  g157
  (
    n284,
    n73
  );


  buf
  g158
  (
    n165,
    n66
  );


  buf
  g159
  (
    n599,
    n152
  );


  not
  g160
  (
    n426,
    n124
  );


  not
  g161
  (
    n511,
    n156
  );


  not
  g162
  (
    n161,
    n146
  );


  not
  g163
  (
    n663,
    n105
  );


  not
  g164
  (
    n220,
    n157
  );


  not
  g165
  (
    n367,
    n53
  );


  buf
  g166
  (
    n425,
    n108
  );


  buf
  g167
  (
    n169,
    n56
  );


  not
  g168
  (
    n413,
    n95
  );


  not
  g169
  (
    n167,
    n137
  );


  buf
  g170
  (
    n640,
    n130
  );


  not
  g171
  (
    n390,
    n131
  );


  not
  g172
  (
    n513,
    n128
  );


  not
  g173
  (
    n478,
    n126
  );


  not
  g174
  (
    n424,
    n152
  );


  buf
  g175
  (
    n171,
    n149
  );


  not
  g176
  (
    n358,
    n44
  );


  buf
  g177
  (
    n222,
    n50
  );


  buf
  g178
  (
    n351,
    n70
  );


  not
  g179
  (
    n214,
    n51
  );


  buf
  g180
  (
    n297,
    n83
  );


  buf
  g181
  (
    n491,
    n89
  );


  not
  g182
  (
    n409,
    n45
  );


  not
  g183
  (
    n439,
    n88
  );


  not
  g184
  (
    n287,
    n94
  );


  not
  g185
  (
    n645,
    n119
  );


  not
  g186
  (
    n400,
    n118
  );


  buf
  g187
  (
    n320,
    n120
  );


  buf
  g188
  (
    n257,
    n47
  );


  buf
  g189
  (
    n401,
    n154
  );


  buf
  g190
  (
    n641,
    n100
  );


  buf
  g191
  (
    n268,
    n146
  );


  not
  g192
  (
    n212,
    n144
  );


  not
  g193
  (
    n592,
    n130
  );


  not
  g194
  (
    n606,
    n74
  );


  not
  g195
  (
    n211,
    n93
  );


  buf
  g196
  (
    n228,
    n72
  );


  buf
  g197
  (
    n532,
    n72
  );


  not
  g198
  (
    n411,
    n74
  );


  buf
  g199
  (
    n482,
    n132
  );


  buf
  g200
  (
    n240,
    n111
  );


  not
  g201
  (
    n210,
    n84
  );


  buf
  g202
  (
    n234,
    n36
  );


  not
  g203
  (
    n190,
    n135
  );


  not
  g204
  (
    n246,
    n79
  );


  buf
  g205
  (
    n551,
    n44
  );


  buf
  g206
  (
    n617,
    n97
  );


  not
  g207
  (
    n388,
    n60
  );


  buf
  g208
  (
    n659,
    n139
  );


  not
  g209
  (
    n379,
    n154
  );


  buf
  g210
  (
    n340,
    n74
  );


  not
  g211
  (
    n625,
    n125
  );


  buf
  g212
  (
    n492,
    n108
  );


  buf
  g213
  (
    n163,
    n53
  );


  buf
  g214
  (
    n229,
    n160
  );


  buf
  g215
  (
    n441,
    n54
  );


  buf
  g216
  (
    n455,
    n160
  );


  not
  g217
  (
    n376,
    n80
  );


  not
  g218
  (
    n354,
    n45
  );


  not
  g219
  (
    n555,
    n106
  );


  not
  g220
  (
    n255,
    n106
  );


  buf
  g221
  (
    n578,
    n56
  );


  buf
  g222
  (
    n557,
    n58
  );


  not
  g223
  (
    n414,
    n42
  );


  not
  g224
  (
    n462,
    n141
  );


  buf
  g225
  (
    n536,
    n105
  );


  not
  g226
  (
    n573,
    n115
  );


  not
  g227
  (
    n479,
    n85
  );


  not
  g228
  (
    n363,
    n135
  );


  not
  g229
  (
    n259,
    n143
  );


  not
  g230
  (
    n473,
    n99
  );


  buf
  g231
  (
    n359,
    n72
  );


  buf
  g232
  (
    n576,
    n131
  );


  not
  g233
  (
    n647,
    n45
  );


  not
  g234
  (
    n371,
    n41
  );


  buf
  g235
  (
    n331,
    n114
  );


  buf
  g236
  (
    n584,
    n70
  );


  buf
  g237
  (
    n525,
    n157
  );


  not
  g238
  (
    n362,
    n121
  );


  buf
  g239
  (
    n270,
    n82
  );


  not
  g240
  (
    n260,
    n92
  );


  not
  g241
  (
    n446,
    n123
  );


  not
  g242
  (
    n199,
    n122
  );


  buf
  g243
  (
    n189,
    n64
  );


  buf
  g244
  (
    n375,
    n101
  );


  not
  g245
  (
    n484,
    n86
  );


  buf
  g246
  (
    n445,
    n95
  );


  buf
  g247
  (
    n644,
    n135
  );


  not
  g248
  (
    n530,
    n100
  );


  not
  g249
  (
    n187,
    n33
  );


  buf
  g250
  (
    n466,
    n101
  );


  not
  g251
  (
    n296,
    n117
  );


  not
  g252
  (
    n254,
    n109
  );


  not
  g253
  (
    n216,
    n54
  );


  buf
  g254
  (
    n539,
    n36
  );


  not
  g255
  (
    n407,
    n57
  );


  buf
  g256
  (
    n468,
    n63
  );


  not
  g257
  (
    n316,
    n61
  );


  not
  g258
  (
    n274,
    n85
  );


  buf
  g259
  (
    n639,
    n78
  );


  buf
  g260
  (
    n381,
    n132
  );


  buf
  g261
  (
    n281,
    n116
  );


  buf
  g262
  (
    n408,
    n46
  );


  not
  g263
  (
    n612,
    n54
  );


  buf
  g264
  (
    n634,
    n120
  );


  not
  g265
  (
    n494,
    n83
  );


  buf
  g266
  (
    n197,
    n38
  );


  buf
  g267
  (
    n633,
    n52
  );


  not
  g268
  (
    n501,
    n81
  );


  not
  g269
  (
    n609,
    n61
  );


  not
  g270
  (
    n604,
    n49
  );


  not
  g271
  (
    n384,
    n98
  );


  not
  g272
  (
    n527,
    n42
  );


  not
  g273
  (
    n572,
    n142
  );


  not
  g274
  (
    n267,
    n121
  );


  buf
  g275
  (
    n389,
    n133
  );


  not
  g276
  (
    n334,
    n84
  );


  not
  g277
  (
    n614,
    n158
  );


  buf
  g278
  (
    n568,
    n155
  );


  not
  g279
  (
    n613,
    n34
  );


  not
  g280
  (
    n324,
    n156
  );


  buf
  g281
  (
    n518,
    n46
  );


  not
  g282
  (
    n338,
    n91
  );


  buf
  g283
  (
    n514,
    n138
  );


  not
  g284
  (
    n396,
    n98
  );


  buf
  g285
  (
    n248,
    n110
  );


  buf
  g286
  (
    n404,
    n56
  );


  not
  g287
  (
    n262,
    n159
  );


  not
  g288
  (
    n556,
    n40
  );


  not
  g289
  (
    n610,
    n41
  );


  not
  g290
  (
    n304,
    n102
  );


  not
  g291
  (
    n350,
    n141
  );


  not
  g292
  (
    n183,
    n123
  );


  buf
  g293
  (
    n538,
    n127
  );


  buf
  g294
  (
    n658,
    n121
  );


  buf
  g295
  (
    n526,
    n41
  );


  buf
  g296
  (
    n637,
    n55
  );


  not
  g297
  (
    n280,
    n129
  );


  not
  g298
  (
    n176,
    n114
  );


  not
  g299
  (
    n269,
    n60
  );


  buf
  g300
  (
    n651,
    n48
  );


  buf
  g301
  (
    n193,
    n103
  );


  not
  g302
  (
    n213,
    n144
  );


  not
  g303
  (
    n397,
    n81
  );


  not
  g304
  (
    n469,
    n150
  );


  not
  g305
  (
    n326,
    n57
  );


  buf
  g306
  (
    n600,
    n58
  );


  buf
  g307
  (
    n310,
    n129
  );


  buf
  g308
  (
    n422,
    n62
  );


  buf
  g309
  (
    n219,
    n100
  );


  not
  g310
  (
    n186,
    n97
  );


  not
  g311
  (
    n205,
    n97
  );


  not
  g312
  (
    n626,
    n49
  );


  not
  g313
  (
    n447,
    n45
  );


  buf
  g314
  (
    n412,
    n43
  );


  buf
  g315
  (
    n416,
    n92
  );


  not
  g316
  (
    n662,
    n59
  );


  not
  g317
  (
    n464,
    n116
  );


  buf
  g318
  (
    n622,
    n118
  );


  not
  g319
  (
    n596,
    n95
  );


  buf
  g320
  (
    n583,
    n75
  );


  buf
  g321
  (
    n571,
    n131
  );


  not
  g322
  (
    n488,
    n68
  );


  buf
  g323
  (
    n548,
    n92
  );


  not
  g324
  (
    n430,
    n82
  );


  not
  g325
  (
    n343,
    n148
  );


  buf
  g326
  (
    n545,
    n77
  );


  not
  g327
  (
    n522,
    n34
  );


  buf
  g328
  (
    n177,
    n133
  );


  not
  g329
  (
    n303,
    n113
  );


  buf
  g330
  (
    n348,
    n153
  );


  not
  g331
  (
    n289,
    n52
  );


  not
  g332
  (
    n239,
    n111
  );


  buf
  g333
  (
    n458,
    n151
  );


  not
  g334
  (
    n657,
    n65
  );


  not
  g335
  (
    n448,
    n71
  );


  buf
  g336
  (
    n503,
    n67
  );


  buf
  g337
  (
    n519,
    n96
  );


  buf
  g338
  (
    n523,
    n77
  );


  not
  g339
  (
    n423,
    n109
  );


  not
  g340
  (
    n386,
    n125
  );


  not
  g341
  (
    n436,
    n74
  );


  buf
  g342
  (
    n339,
    n75
  );


  not
  g343
  (
    n504,
    n51
  );


  not
  g344
  (
    n342,
    n34
  );


  buf
  g345
  (
    n271,
    n93
  );


  buf
  g346
  (
    n623,
    n39
  );


  buf
  g347
  (
    n475,
    n88
  );


  buf
  g348
  (
    n463,
    n114
  );


  buf
  g349
  (
    n299,
    n147
  );


  buf
  g350
  (
    n322,
    n111
  );


  buf
  g351
  (
    n654,
    n35
  );


  not
  g352
  (
    n452,
    n81
  );


  not
  g353
  (
    n586,
    n94
  );


  buf
  g354
  (
    n290,
    n69
  );


  buf
  g355
  (
    n636,
    n63
  );


  buf
  g356
  (
    n166,
    n57
  );


  buf
  g357
  (
    n627,
    n38
  );


  buf
  g358
  (
    n170,
    n109
  );


  buf
  g359
  (
    n670,
    n115
  );


  not
  g360
  (
    n440,
    n136
  );


  buf
  g361
  (
    n629,
    n78
  );


  buf
  g362
  (
    n650,
    n78
  );


  buf
  g363
  (
    n476,
    n76
  );


  not
  g364
  (
    n500,
    n64
  );


  buf
  g365
  (
    n582,
    n63
  );


  buf
  g366
  (
    n454,
    n89
  );


  buf
  g367
  (
    n498,
    n87
  );


  buf
  g368
  (
    n417,
    n90
  );


  not
  g369
  (
    n508,
    n102
  );


  buf
  g370
  (
    n383,
    n136
  );


  not
  g371
  (
    n451,
    n117
  );


  not
  g372
  (
    n369,
    n140
  );


  buf
  g373
  (
    n567,
    n59
  );


  not
  g374
  (
    n574,
    n70
  );


  buf
  g375
  (
    n587,
    n104
  );


  buf
  g376
  (
    n217,
    n86
  );


  buf
  g377
  (
    n509,
    n124
  );


  buf
  g378
  (
    n378,
    n71
  );


  buf
  g379
  (
    n672,
    n148
  );


  buf
  g380
  (
    n178,
    n36
  );


  buf
  g381
  (
    n370,
    n64
  );


  buf
  g382
  (
    n624,
    n144
  );


  not
  g383
  (
    n631,
    n72
  );


  not
  g384
  (
    n361,
    n106
  );


  buf
  g385
  (
    n353,
    n53
  );


  not
  g386
  (
    n546,
    n49
  );


  buf
  g387
  (
    n278,
    n130
  );


  not
  g388
  (
    n428,
    n150
  );


  buf
  g389
  (
    n314,
    n133
  );


  not
  g390
  (
    n225,
    n67
  );


  not
  g391
  (
    n258,
    n108
  );


  buf
  g392
  (
    n543,
    n89
  );


  buf
  g393
  (
    n288,
    n88
  );


  buf
  g394
  (
    n360,
    n110
  );


  buf
  g395
  (
    n605,
    n119
  );


  buf
  g396
  (
    n620,
    n91
  );


  not
  g397
  (
    n632,
    n137
  );


  not
  g398
  (
    n419,
    n107
  );


  buf
  g399
  (
    n549,
    n159
  );


  not
  g400
  (
    n434,
    n35
  );


  not
  g401
  (
    n251,
    n94
  );


  not
  g402
  (
    n164,
    n132
  );


  not
  g403
  (
    n666,
    n67
  );


  buf
  g404
  (
    n664,
    n121
  );


  buf
  g405
  (
    n431,
    n149
  );


  buf
  g406
  (
    n497,
    n104
  );


  buf
  g407
  (
    n520,
    n124
  );


  not
  g408
  (
    n279,
    n96
  );


  not
  g409
  (
    n201,
    n145
  );


  not
  g410
  (
    n465,
    n87
  );


  buf
  g411
  (
    n250,
    n157
  );


  buf
  g412
  (
    n328,
    n145
  );


  buf
  g413
  (
    n560,
    n93
  );


  buf
  g414
  (
    n275,
    n69
  );


  buf
  g415
  (
    n437,
    n62
  );


  not
  g416
  (
    n444,
    n71
  );


  not
  g417
  (
    n649,
    n39
  );


  not
  g418
  (
    n380,
    n84
  );


  not
  g419
  (
    n377,
    n91
  );


  buf
  g420
  (
    n182,
    n151
  );


  not
  g421
  (
    n398,
    n107
  );


  not
  g422
  (
    n364,
    n146
  );


  buf
  g423
  (
    n619,
    n68
  );


  buf
  g424
  (
    n427,
    n126
  );


  buf
  g425
  (
    n387,
    n69
  );


  not
  g426
  (
    n559,
    n80
  );


  not
  g427
  (
    n318,
    n124
  );


  not
  g428
  (
    n661,
    n101
  );


  buf
  g429
  (
    n198,
    n112
  );


  not
  g430
  (
    n655,
    n59
  );


  not
  g431
  (
    n438,
    n83
  );


  buf
  g432
  (
    n588,
    n55
  );


  not
  g433
  (
    n341,
    n151
  );


  not
  g434
  (
    n347,
    n134
  );


  buf
  g435
  (
    n306,
    n90
  );


  not
  g436
  (
    n276,
    n75
  );


  buf
  g437
  (
    n204,
    n70
  );


  not
  g438
  (
    n352,
    n96
  );


  buf
  g439
  (
    n506,
    n145
  );


  buf
  g440
  (
    n293,
    n35
  );


  buf
  g441
  (
    n495,
    n87
  );


  buf
  g442
  (
    n315,
    n34
  );


  not
  g443
  (
    n597,
    n57
  );


  buf
  g444
  (
    n537,
    n155
  );


  buf
  g445
  (
    n496,
    n110
  );


  buf
  g446
  (
    n313,
    n153
  );


  not
  g447
  (
    n611,
    n140
  );


  buf
  g448
  (
    n577,
    n85
  );


  not
  g449
  (
    n528,
    n112
  );


  buf
  g450
  (
    n552,
    n62
  );


  buf
  g451
  (
    n547,
    n47
  );


  not
  g452
  (
    n311,
    n128
  );


  not
  g453
  (
    n391,
    n122
  );


  not
  g454
  (
    n206,
    n55
  );


  not
  g455
  (
    n283,
    n73
  );


  not
  g456
  (
    n590,
    n103
  );


  not
  g457
  (
    n481,
    n105
  );


  not
  g458
  (
    n249,
    n119
  );


  buf
  g459
  (
    n245,
    n145
  );


  buf
  g460
  (
    n180,
    n132
  );


  not
  g461
  (
    n667,
    n135
  );


  not
  g462
  (
    n235,
    n102
  );


  not
  g463
  (
    n515,
    n125
  );


  not
  g464
  (
    n172,
    n128
  );


  buf
  g465
  (
    n418,
    n50
  );


  not
  g466
  (
    n173,
    n61
  );


  buf
  g467
  (
    n194,
    n98
  );


  not
  g468
  (
    n221,
    n75
  );


  buf
  g469
  (
    KeyWire_0_8,
    n152
  );


  not
  g470
  (
    n233,
    n37
  );


  not
  g471
  (
    n558,
    n83
  );


  buf
  g472
  (
    n541,
    n80
  );


  not
  g473
  (
    n207,
    n60
  );


  not
  g474
  (
    n247,
    n42
  );


  not
  g475
  (
    n472,
    n94
  );


  not
  g476
  (
    n564,
    n86
  );


  not
  g477
  (
    n325,
    n65
  );


  not
  g478
  (
    n184,
    n76
  );


  not
  g479
  (
    n531,
    n87
  );


  buf
  g480
  (
    n507,
    n84
  );


  buf
  g481
  (
    n365,
    n103
  );


  buf
  g482
  (
    n668,
    n115
  );


  not
  g483
  (
    n385,
    n40
  );


  not
  g484
  (
    n242,
    n40
  );


  buf
  g485
  (
    n540,
    n138
  );


  not
  g486
  (
    n332,
    n159
  );


  buf
  g487
  (
    n648,
    n155
  );


  buf
  g488
  (
    n550,
    n56
  );


  not
  g489
  (
    n357,
    n108
  );


  buf
  g490
  (
    n218,
    n139
  );


  not
  g491
  (
    n298,
    n106
  );


  buf
  g492
  (
    n456,
    n157
  );


  buf
  g493
  (
    n580,
    n143
  );


  buf
  g494
  (
    n485,
    n107
  );


  not
  g495
  (
    n554,
    n156
  );


  not
  g496
  (
    n224,
    n150
  );


  not
  g497
  (
    n669,
    n149
  );


  buf
  g498
  (
    n253,
    n127
  );


  buf
  g499
  (
    n534,
    n129
  );


  not
  g500
  (
    n282,
    n120
  );


  not
  g501
  (
    n294,
    n96
  );


  not
  g502
  (
    n591,
    n141
  );


  buf
  g503
  (
    n467,
    n141
  );


  not
  g504
  (
    n368,
    n78
  );


  not
  g505
  (
    n460,
    n128
  );


  not
  g506
  (
    n330,
    n147
  );


  buf
  g507
  (
    n374,
    n154
  );


  not
  g508
  (
    n581,
    n133
  );


  not
  g509
  (
    n312,
    n77
  );


  not
  g510
  (
    n616,
    n149
  );


  not
  g511
  (
    n337,
    n38
  );


  not
  g512
  (
    n579,
    n109
  );


  not
  g513
  (
    n191,
    n104
  );


  buf
  g514
  (
    n575,
    n158
  );


  buf
  g515
  (
    n471,
    n160
  );


  buf
  g516
  (
    n356,
    n143
  );


  buf
  g517
  (
    n470,
    n127
  );


  not
  g518
  (
    n307,
    n93
  );


  buf
  g519
  (
    n459,
    n61
  );


  buf
  g520
  (
    n232,
    n137
  );


  buf
  g521
  (
    n516,
    n118
  );


  not
  g522
  (
    n236,
    n115
  );


  not
  g523
  (
    n477,
    n127
  );


  buf
  g524
  (
    n403,
    n66
  );


  not
  g525
  (
    n244,
    n79
  );


  buf
  g526
  (
    n521,
    n125
  );


  not
  g527
  (
    n223,
    n140
  );


  not
  g528
  (
    n429,
    n79
  );


  buf
  g529
  (
    n480,
    n59
  );


  not
  g530
  (
    n542,
    n134
  );


  buf
  g531
  (
    n630,
    n44
  );


  buf
  g532
  (
    n474,
    n91
  );


  not
  g533
  (
    n336,
    n90
  );


  buf
  g534
  (
    n569,
    n47
  );


  buf
  g535
  (
    n486,
    n136
  );


  buf
  g536
  (
    n175,
    n33
  );


  not
  g537
  (
    n395,
    n160
  );


  not
  g538
  (
    n435,
    n51
  );


  not
  g539
  (
    KeyWire_0_1,
    n82
  );


  buf
  g540
  (
    n461,
    n118
  );


  not
  g541
  (
    n443,
    n48
  );


  buf
  g542
  (
    n344,
    n123
  );


  not
  g543
  (
    n192,
    n44
  );


  not
  g544
  (
    n349,
    n65
  );


  buf
  g545
  (
    n535,
    n107
  );


  buf
  g546
  (
    n372,
    n117
  );


  not
  g547
  (
    n544,
    n92
  );


  not
  g548
  (
    n671,
    n68
  );


  not
  g549
  (
    n602,
    n85
  );


  buf
  g550
  (
    n188,
    n136
  );


  buf
  g551
  (
    n355,
    n142
  );


  not
  g552
  (
    n502,
    n62
  );


  not
  g553
  (
    n643,
    n81
  );


  not
  g554
  (
    n512,
    n41
  );


  not
  g555
  (
    n524,
    n131
  );


  not
  g556
  (
    n493,
    n43
  );


  not
  g557
  (
    n264,
    n49
  );


  not
  g558
  (
    n392,
    n95
  );


  not
  g559
  (
    n215,
    n52
  );


  not
  g560
  (
    n301,
    n52
  );


  not
  g561
  (
    n561,
    n88
  );


  buf
  g562
  (
    n346,
    n39
  );


  not
  g563
  (
    n570,
    n116
  );


  not
  g564
  (
    n263,
    n73
  );


  buf
  g565
  (
    n421,
    n148
  );


  buf
  g566
  (
    n638,
    n105
  );


  not
  g567
  (
    n162,
    n99
  );


  not
  g568
  (
    n209,
    n154
  );


  not
  g569
  (
    n406,
    n122
  );


  buf
  g570
  (
    n457,
    n138
  );


  not
  g571
  (
    n230,
    n158
  );


  buf
  g572
  (
    n642,
    n35
  );


  not
  g573
  (
    n308,
    n76
  );


  not
  g574
  (
    n345,
    n102
  );


  not
  g575
  (
    n399,
    n67
  );


  buf
  g576
  (
    n252,
    n43
  );


  buf
  g577
  (
    n394,
    n144
  );


  buf
  g578
  (
    n487,
    n150
  );


  buf
  g579
  (
    n319,
    n64
  );


  not
  g580
  (
    n517,
    n46
  );


  not
  g581
  (
    n553,
    n86
  );


  not
  g582
  (
    n317,
    n153
  );


  buf
  g583
  (
    n510,
    n148
  );


  not
  g584
  (
    n373,
    n43
  );


  buf
  g585
  (
    n665,
    n147
  );


  not
  g586
  (
    n608,
    n82
  );


  buf
  g587
  (
    n566,
    n58
  );


  buf
  g588
  (
    n203,
    n142
  );


  buf
  g589
  (
    n433,
    n69
  );


  not
  g590
  (
    n272,
    n146
  );


  buf
  g591
  (
    n174,
    n38
  );


  not
  g592
  (
    n402,
    n139
  );


  not
  g593
  (
    n200,
    n129
  );


  not
  g594
  (
    n603,
    n99
  );


  not
  g595
  (
    n533,
    n54
  );


  buf
  g596
  (
    n181,
    n37
  );


  not
  g597
  (
    n195,
    n48
  );


  not
  g598
  (
    n405,
    n50
  );


  buf
  g599
  (
    n185,
    n111
  );


  not
  g600
  (
    n305,
    n152
  );


  not
  g601
  (
    n382,
    n90
  );


  buf
  g602
  (
    n179,
    n53
  );


  buf
  g603
  (
    n273,
    n139
  );


  buf
  g604
  (
    n333,
    n37
  );


  buf
  g605
  (
    n285,
    n134
  );


  buf
  g606
  (
    n266,
    n120
  );


  not
  g607
  (
    n635,
    n155
  );


  buf
  g608
  (
    n615,
    n112
  );


  buf
  g609
  (
    n660,
    n103
  );


  not
  g610
  (
    n499,
    n116
  );


  buf
  g611
  (
    n420,
    n122
  );


  buf
  g612
  (
    n410,
    n48
  );


  not
  g613
  (
    n277,
    n113
  );


  buf
  g614
  (
    n618,
    n55
  );


  not
  g615
  (
    n594,
    n80
  );


  not
  g616
  (
    n237,
    n40
  );


  buf
  g617
  (
    n505,
    n63
  );


  buf
  g618
  (
    KeyWire_0_5,
    n73
  );


  not
  g619
  (
    n563,
    n137
  );


  not
  g620
  (
    n442,
    n142
  );


  buf
  g621
  (
    n241,
    n138
  );


  buf
  g622
  (
    n335,
    n130
  );


  buf
  g623
  (
    n302,
    n140
  );


  not
  g624
  (
    n656,
    n79
  );


  buf
  g625
  (
    n321,
    n51
  );


  not
  g626
  (
    n601,
    n66
  );


  not
  g627
  (
    n265,
    n42
  );


  buf
  g628
  (
    n432,
    n156
  );


  buf
  g629
  (
    n607,
    n68
  );


  buf
  g630
  (
    n621,
    n117
  );


  buf
  g631
  (
    n489,
    n158
  );


  not
  g632
  (
    n646,
    n112
  );


  buf
  g633
  (
    n196,
    n104
  );


  buf
  g634
  (
    n562,
    n99
  );


  not
  g635
  (
    n309,
    n89
  );


  not
  g636
  (
    n598,
    n71
  );


  not
  g637
  (
    n490,
    n126
  );


  buf
  g638
  (
    n261,
    n134
  );


  not
  g639
  (
    n529,
    n98
  );


  xnor
  g640
  (
    n845,
    n430,
    n456,
    n333,
    n486
  );


  nor
  g641
  (
    n685,
    n280,
    n461,
    n353,
    n357
  );


  nand
  g642
  (
    n814,
    n380,
    n332,
    n272,
    n378
  );


  and
  g643
  (
    n851,
    n438,
    n407,
    n363,
    n423
  );


  or
  g644
  (
    n903,
    n264,
    n484,
    n375,
    n369
  );


  nand
  g645
  (
    n726,
    n186,
    n319,
    n447,
    n303
  );


  nand
  g646
  (
    n746,
    n327,
    n233,
    n277,
    n426
  );


  xor
  g647
  (
    n773,
    n167,
    n266,
    n442,
    n344
  );


  xor
  g648
  (
    n843,
    n497,
    n459,
    n489,
    n417
  );


  xor
  g649
  (
    n751,
    n348,
    n378,
    n398,
    n488
  );


  nand
  g650
  (
    n922,
    n367,
    n314,
    n269,
    n303
  );


  xnor
  g651
  (
    n800,
    n202,
    n282,
    n382,
    n266
  );


  nand
  g652
  (
    n863,
    n306,
    n344,
    n362,
    n229
  );


  and
  g653
  (
    n693,
    n489,
    n386,
    n189,
    n480
  );


  xor
  g654
  (
    n927,
    n165,
    n473,
    n287,
    n279
  );


  nor
  g655
  (
    n912,
    n381,
    n322,
    n473,
    n428
  );


  and
  g656
  (
    n749,
    n330,
    n244,
    n471,
    n478
  );


  or
  g657
  (
    n870,
    n364,
    n381,
    n389,
    n383
  );


  xor
  g658
  (
    n899,
    n409,
    n295,
    n274,
    n456
  );


  or
  g659
  (
    n756,
    n446,
    n399,
    n313,
    n428
  );


  nand
  g660
  (
    n929,
    n387,
    n465,
    n406,
    n445
  );


  and
  g661
  (
    n784,
    n452,
    n445,
    n314,
    n308
  );


  or
  g662
  (
    n677,
    n348,
    n313,
    n300,
    n356
  );


  xor
  g663
  (
    n824,
    n171,
    n410,
    n414,
    n369
  );


  xnor
  g664
  (
    n766,
    n297,
    n371,
    n434,
    n396
  );


  and
  g665
  (
    n806,
    n230,
    n491,
    n351,
    n435
  );


  and
  g666
  (
    n879,
    n334,
    n482,
    n312,
    n359
  );


  nand
  g667
  (
    n911,
    n255,
    n466,
    n352,
    n465
  );


  or
  g668
  (
    n902,
    n416,
    n304,
    n450,
    n267
  );


  xor
  g669
  (
    n859,
    n258,
    n311,
    n335,
    n461
  );


  xor
  g670
  (
    n872,
    n385,
    n224,
    n377,
    n370
  );


  or
  g671
  (
    n778,
    n422,
    n339,
    n408,
    n318
  );


  xor
  g672
  (
    n865,
    n287,
    n260,
    n266,
    n269
  );


  xnor
  g673
  (
    n837,
    n445,
    n277,
    n205,
    n370
  );


  or
  g674
  (
    n812,
    n425,
    n400,
    n417,
    n284
  );


  nand
  g675
  (
    n886,
    n274,
    n411,
    n290,
    n370
  );


  and
  g676
  (
    n679,
    n345,
    n405,
    n421,
    n387
  );


  nand
  g677
  (
    n836,
    n309,
    n356,
    n444,
    n292
  );


  nor
  g678
  (
    n890,
    n198,
    n372,
    n435
  );


  and
  g679
  (
    n847,
    n330,
    n174,
    n380,
    n484
  );


  nand
  g680
  (
    n901,
    n423,
    n325,
    n289,
    n474
  );


  xnor
  g681
  (
    n690,
    n354,
    n446,
    n261,
    n176
  );


  or
  g682
  (
    n793,
    n319,
    n338,
    n206,
    n342
  );


  xor
  g683
  (
    n737,
    n490,
    n262,
    n449,
    n483
  );


  xnor
  g684
  (
    n834,
    n195,
    n355,
    n333,
    n484
  );


  and
  g685
  (
    n842,
    n335,
    n460,
    n336,
    n326
  );


  xor
  g686
  (
    n937,
    n398,
    n297,
    n481,
    n498
  );


  xnor
  g687
  (
    n909,
    n375,
    n315,
    n340,
    n390
  );


  and
  g688
  (
    n700,
    n498,
    n307,
    n356,
    n455
  );


  or
  g689
  (
    n704,
    n263,
    n361,
    n300,
    n420
  );


  nand
  g690
  (
    n829,
    n353,
    n259,
    n344,
    n245
  );


  xnor
  g691
  (
    n792,
    n390,
    n384,
    n161,
    n258
  );


  and
  g692
  (
    n880,
    n295,
    n425,
    n163,
    n298
  );


  or
  g693
  (
    n893,
    n367,
    n391,
    n458,
    n314
  );


  xor
  g694
  (
    n817,
    n256,
    n493,
    n397,
    n360
  );


  xnor
  g695
  (
    n802,
    n472,
    n468,
    n414,
    n393
  );


  xor
  g696
  (
    n908,
    n350,
    n178,
    n271,
    n427
  );


  and
  g697
  (
    n830,
    n315,
    n187,
    n405,
    n376
  );


  and
  g698
  (
    n915,
    n381,
    n359,
    n219,
    n291
  );


  xnor
  g699
  (
    n720,
    n434,
    n439,
    n416,
    n366
  );


  nand
  g700
  (
    n831,
    n475,
    n223,
    n409,
    n406
  );


  and
  g701
  (
    n673,
    n379,
    n270,
    n448,
    n298
  );


  xor
  g702
  (
    n796,
    n192,
    n265,
    n456,
    n293
  );


  xor
  g703
  (
    n684,
    n427,
    n378,
    n443,
    n301
  );


  xor
  g704
  (
    n926,
    n388,
    n373,
    n261,
    n291
  );


  xnor
  g705
  (
    n736,
    n331,
    n488,
    n411,
    n251
  );


  and
  g706
  (
    n885,
    n292,
    n492,
    n455,
    n349
  );


  nor
  g707
  (
    n846,
    n440,
    n336,
    n319,
    n307
  );


  and
  g708
  (
    n923,
    n485,
    n418,
    n177,
    n326
  );


  nand
  g709
  (
    n730,
    n310,
    n388,
    n396,
    n458
  );


  or
  g710
  (
    n891,
    n354,
    n375,
    n304,
    n267
  );


  or
  g711
  (
    n686,
    n397,
    n469,
    n259,
    n472
  );


  nand
  g712
  (
    n921,
    n275,
    n299,
    n278
  );


  or
  g713
  (
    n713,
    n431,
    n431,
    n443,
    n412
  );


  nor
  g714
  (
    n876,
    n457,
    n166,
    n391,
    n276
  );


  xor
  g715
  (
    n810,
    n489,
    n364,
    n493,
    n325
  );


  or
  g716
  (
    n883,
    n388,
    n384,
    n261,
    n211
  );


  and
  g717
  (
    n873,
    n359,
    n438,
    n296,
    n243
  );


  xor
  g718
  (
    n848,
    n474,
    n276,
    n494,
    n280
  );


  xor
  g719
  (
    n898,
    n342,
    n281,
    n370,
    n312
  );


  xor
  g720
  (
    n887,
    n183,
    n465,
    n347,
    n381
  );


  and
  g721
  (
    n930,
    n490,
    n448,
    n409,
    n469
  );


  nand
  g722
  (
    n764,
    n300,
    n345,
    n306,
    n318
  );


  nor
  g723
  (
    n725,
    n466,
    n330,
    n394,
    n372
  );


  nor
  g724
  (
    n884,
    n277,
    n419,
    n262,
    n497
  );


  nor
  g725
  (
    n676,
    n321,
    n280,
    n413,
    n439
  );


  xnor
  g726
  (
    n680,
    n373,
    n424,
    n271,
    n391
  );


  or
  g727
  (
    n900,
    n435,
    n497,
    n282,
    n321
  );


  nor
  g728
  (
    KeyWire_0_12,
    n284,
    n225,
    n464,
    n345
  );


  xor
  g729
  (
    n743,
    n423,
    n216,
    n270,
    n353
  );


  xor
  g730
  (
    n731,
    n291,
    n374,
    n433
  );


  xor
  g731
  (
    n904,
    n308,
    n179,
    n313,
    n397
  );


  nor
  g732
  (
    n894,
    n253,
    n494,
    n364,
    n487
  );


  xnor
  g733
  (
    n925,
    n326,
    n263,
    n324,
    n463
  );


  xor
  g734
  (
    n933,
    n485,
    n320,
    n352,
    n309
  );


  nand
  g735
  (
    n809,
    n271,
    n459,
    n440,
    n443
  );


  and
  g736
  (
    n758,
    n310,
    n287,
    n196,
    n355
  );


  or
  g737
  (
    n936,
    n283,
    n279,
    n286,
    n449
  );


  nand
  g738
  (
    KeyWire_0_13,
    n349,
    n386,
    n309,
    n318
  );


  or
  g739
  (
    n807,
    n418,
    n348,
    n376,
    n337
  );


  nor
  g740
  (
    n896,
    n297,
    n411,
    n435,
    n445
  );


  xor
  g741
  (
    n708,
    n468,
    n252,
    n460,
    n422
  );


  xnor
  g742
  (
    n828,
    n356,
    n371,
    n485,
    n412
  );


  and
  g743
  (
    n775,
    n317,
    n340,
    n305,
    n498
  );


  or
  g744
  (
    n695,
    n403,
    n392,
    n408,
    n469
  );


  xnor
  g745
  (
    n740,
    n410,
    n263,
    n374,
    n349
  );


  and
  g746
  (
    n729,
    n392,
    n376,
    n478,
    n258
  );


  nand
  g747
  (
    n808,
    n402,
    n348,
    n499,
    n281
  );


  nand
  g748
  (
    n741,
    n496,
    n301,
    n315,
    n324
  );


  and
  g749
  (
    n748,
    n430,
    n443,
    n463,
    n254
  );


  and
  g750
  (
    n785,
    n479,
    n295,
    n301,
    n382
  );


  xnor
  g751
  (
    n889,
    n184,
    n416,
    n349,
    n358
  );


  and
  g752
  (
    n682,
    n441,
    n476,
    n492,
    n334
  );


  and
  g753
  (
    n854,
    n282,
    n293,
    n241,
    n329
  );


  nor
  g754
  (
    n783,
    n273,
    n362,
    n412,
    n299
  );


  nor
  g755
  (
    n850,
    n494,
    n471,
    n221
  );


  xor
  g756
  (
    n888,
    n302,
    n496,
    n374,
    n285
  );


  xnor
  g757
  (
    n935,
    n170,
    n427,
    n321,
    n473
  );


  nand
  g758
  (
    n739,
    n332,
    n437,
    n220,
    n260
  );


  and
  g759
  (
    n841,
    n482,
    n457,
    n350,
    n360
  );


  xnor
  g760
  (
    n771,
    n315,
    n389,
    n199,
    n360
  );


  nor
  g761
  (
    n916,
    n404,
    n368,
    n346,
    n292
  );


  xnor
  g762
  (
    n857,
    n320,
    n429,
    n188,
    n453
  );


  nand
  g763
  (
    n789,
    n289,
    n392,
    n433,
    n272
  );


  nand
  g764
  (
    n795,
    n465,
    n405,
    n375,
    n172
  );


  nor
  g765
  (
    n815,
    n442,
    n391,
    n331,
    n288
  );


  and
  g766
  (
    n849,
    n386,
    n493,
    n437,
    n477
  );


  nand
  g767
  (
    n840,
    n404,
    n401,
    n407,
    n384
  );


  nor
  g768
  (
    n907,
    n397,
    n325,
    n327,
    n363
  );


  or
  g769
  (
    n786,
    n246,
    n451,
    n311,
    n300
  );


  or
  g770
  (
    n924,
    n294,
    n463,
    n407,
    n308
  );


  xor
  g771
  (
    n747,
    n424,
    n351,
    n339,
    n438
  );


  xor
  g772
  (
    n728,
    n386,
    n294,
    n353,
    n303
  );


  xnor
  g773
  (
    n701,
    n341,
    n477,
    n307,
    n476
  );


  nand
  g774
  (
    n691,
    n302,
    n434,
    n454,
    n476
  );


  xor
  g775
  (
    n852,
    n331,
    n269,
    n413,
    n395
  );


  nand
  g776
  (
    n733,
    n310,
    n404,
    n342,
    n359
  );


  xnor
  g777
  (
    n860,
    n264,
    n478,
    n222,
    n447
  );


  nor
  g778
  (
    n895,
    n268,
    n434,
    n487,
    n405
  );


  nor
  g779
  (
    n750,
    n476,
    n290,
    n383,
    n436
  );


  xor
  g780
  (
    n820,
    n265,
    n428,
    n292,
    n193
  );


  xor
  g781
  (
    n727,
    n310,
    n483,
    n467,
    n323
  );


  or
  g782
  (
    n787,
    n340,
    n257,
    n283,
    n273
  );


  nand
  g783
  (
    n913,
    n486,
    n411,
    n413,
    n340
  );


  xnor
  g784
  (
    n897,
    n347,
    n232,
    n432,
    n346
  );


  and
  g785
  (
    KeyWire_0_14,
    n417,
    n470,
    n446,
    n326
  );


  xor
  g786
  (
    n735,
    n256,
    n460,
    n369,
    n164
  );


  and
  g787
  (
    n791,
    n294,
    n361,
    n328,
    n362
  );


  or
  g788
  (
    n801,
    n439,
    n472,
    n488,
    n461
  );


  or
  g789
  (
    n772,
    n319,
    n485,
    n368,
    n395
  );


  and
  g790
  (
    n892,
    n373,
    n406,
    n347,
    n366
  );


  or
  g791
  (
    n878,
    n484,
    n431,
    n332,
    n317
  );


  nand
  g792
  (
    n774,
    n427,
    n453,
    n496,
    n328
  );


  nand
  g793
  (
    n753,
    n288,
    n328,
    n383,
    n217
  );


  xor
  g794
  (
    n714,
    n346,
    n379,
    n248,
    n314
  );


  nand
  g795
  (
    n871,
    n255,
    n421,
    n268,
    n290
  );


  xor
  g796
  (
    n855,
    n304,
    n238,
    n456,
    n479
  );


  xnor
  g797
  (
    n862,
    n384,
    n256,
    n415,
    n226
  );


  nor
  g798
  (
    n813,
    n491,
    n471,
    n480,
    n369
  );


  nor
  g799
  (
    n763,
    n394,
    n296,
    n444,
    n461
  );


  xnor
  g800
  (
    n853,
    n323,
    n210,
    n403,
    n285
  );


  or
  g801
  (
    n767,
    n262,
    n267,
    n482,
    n338
  );


  nand
  g802
  (
    n805,
    n347,
    n422,
    n277,
    n256
  );


  or
  g803
  (
    n719,
    n312,
    n185,
    n399,
    n306
  );


  xor
  g804
  (
    n864,
    n394,
    n436,
    n459,
    n255
  );


  nand
  g805
  (
    n877,
    n316,
    n200,
    n288,
    n416
  );


  nand
  g806
  (
    n711,
    n367,
    n454,
    n285,
    n439
  );


  or
  g807
  (
    n867,
    n260,
    n335,
    n323,
    n295
  );


  and
  g808
  (
    n822,
    n467,
    n474,
    n379,
    n260
  );


  xor
  g809
  (
    n868,
    n424,
    n237,
    n469,
    n406
  );


  xor
  g810
  (
    n689,
    n488,
    n432,
    n451,
    n258
  );


  xnor
  g811
  (
    n705,
    n354,
    n377,
    n357,
    n432
  );


  or
  g812
  (
    n914,
    n453,
    n190,
    n316,
    n419
  );


  nand
  g813
  (
    n882,
    n371,
    n395,
    n454,
    n472
  );


  nand
  g814
  (
    n825,
    n396,
    n440,
    n290,
    n419
  );


  or
  g815
  (
    n939,
    n402,
    n351,
    n429,
    n274
  );


  and
  g816
  (
    n917,
    n479,
    n312,
    n418,
    n452
  );


  or
  g817
  (
    n938,
    n382,
    n388,
    n491,
    n430
  );


  nor
  g818
  (
    n827,
    n392,
    n408,
    n478,
    n407
  );


  nor
  g819
  (
    n832,
    n430,
    n380,
    n462,
    n343
  );


  xnor
  g820
  (
    n823,
    n257,
    n338,
    n400,
    n448
  );


  nand
  g821
  (
    n707,
    n389,
    n259,
    n417,
    n316
  );


  xor
  g822
  (
    n715,
    n259,
    n242,
    n280,
    n376
  );


  or
  g823
  (
    n782,
    n212,
    n420,
    n273,
    n352
  );


  nand
  g824
  (
    n724,
    n486,
    n483,
    n466,
    n283
  );


  nand
  g825
  (
    n717,
    n236,
    n180,
    n475,
    n234
  );


  nor
  g826
  (
    n752,
    n361,
    n385,
    n366,
    n401
  );


  xnor
  g827
  (
    n770,
    n305,
    n299,
    n486,
    n425
  );


  nand
  g828
  (
    n797,
    n480,
    n284,
    n468,
    n350
  );


  and
  g829
  (
    n838,
    n436,
    n325,
    n495,
    n366
  );


  nand
  g830
  (
    n745,
    n377,
    n449,
    n264,
    n477
  );


  or
  g831
  (
    n780,
    n470,
    n304,
    n377,
    n331
  );


  or
  g832
  (
    n702,
    n317,
    n448,
    n327,
    n399
  );


  or
  g833
  (
    n755,
    n250,
    n308,
    n418,
    n487
  );


  xnor
  g834
  (
    n688,
    n313,
    n367,
    n181,
    n403
  );


  nand
  g835
  (
    n768,
    n473,
    n285,
    n275,
    n432
  );


  nor
  g836
  (
    n732,
    n274,
    n169,
    n379,
    n477
  );


  xnor
  g837
  (
    n940,
    n311,
    n415,
    n235,
    n284
  );


  and
  g838
  (
    n765,
    n362,
    n231,
    n303,
    n364
  );


  nand
  g839
  (
    n811,
    n335,
    n276,
    n299,
    n296
  );


  nand
  g840
  (
    n918,
    n344,
    n378,
    n341,
    n365
  );


  or
  g841
  (
    n696,
    n329,
    n455,
    n343,
    n197
  );


  xor
  g842
  (
    n716,
    n247,
    n336,
    n327,
    n447
  );


  nor
  g843
  (
    n721,
    n426,
    n293,
    n492,
    n257
  );


  nor
  g844
  (
    n826,
    n446,
    n428,
    n333,
    n429
  );


  xnor
  g845
  (
    n776,
    n275,
    n480,
    n475,
    n287
  );


  nor
  g846
  (
    n881,
    n382,
    n227,
    n393,
    n279
  );


  xor
  g847
  (
    n905,
    n400,
    n404,
    n263,
    n479
  );


  and
  g848
  (
    n712,
    n426,
    n275,
    n361,
    n468
  );


  and
  g849
  (
    n687,
    n270,
    n368,
    n398,
    n301
  );


  nor
  g850
  (
    n866,
    n499,
    n393,
    n293,
    n289
  );


  and
  g851
  (
    n803,
    n272,
    n462,
    n433,
    n239
  );


  xnor
  g852
  (
    n694,
    n398,
    n450,
    n481,
    n298
  );


  nor
  g853
  (
    n760,
    n463,
    n306,
    n395,
    n339
  );


  nor
  g854
  (
    n722,
    n341,
    n342,
    n286
  );


  xor
  g855
  (
    n839,
    n288,
    n329,
    n441,
    n334
  );


  xor
  g856
  (
    n761,
    n408,
    n459,
    n168,
    n401
  );


  xnor
  g857
  (
    n804,
    n324,
    n337,
    n368,
    n390
  );


  xnor
  g858
  (
    n920,
    n458,
    n266,
    n278,
    n457
  );


  xnor
  g859
  (
    n931,
    n447,
    n496,
    n466,
    n339
  );


  nor
  g860
  (
    n906,
    n419,
    n423,
    n267,
    n318
  );


  xor
  g861
  (
    n875,
    n414,
    n268,
    n352,
    n207
  );


  nand
  g862
  (
    n706,
    n302,
    n268,
    n357,
    n208
  );


  or
  g863
  (
    n681,
    n402,
    n358,
    n265,
    n322
  );


  and
  g864
  (
    n697,
    n271,
    n343,
    n283,
    n470
  );


  and
  g865
  (
    n742,
    n452,
    n341,
    n444,
    n495
  );


  or
  g866
  (
    n754,
    n457,
    n330,
    n354,
    n494
  );


  or
  g867
  (
    n799,
    n355,
    n218,
    n422,
    n390
  );


  and
  g868
  (
    n794,
    n426,
    n402,
    n444,
    n396
  );


  nor
  g869
  (
    n819,
    n452,
    n328,
    n462,
    n357
  );


  xnor
  g870
  (
    n779,
    n297,
    n316,
    n450,
    n203
  );


  nand
  g871
  (
    n777,
    n191,
    n436,
    n294,
    n334
  );


  and
  g872
  (
    n856,
    n333,
    n194,
    n403,
    n400
  );


  xor
  g873
  (
    n757,
    n464,
    n482,
    n454,
    n249
  );


  xor
  g874
  (
    n932,
    n305,
    n175,
    n324,
    n264
  );


  nand
  g875
  (
    n692,
    n449,
    n393,
    n498,
    n346
  );


  xnor
  g876
  (
    n861,
    n255,
    n410,
    n329,
    n495
  );


  nor
  g877
  (
    n790,
    n336,
    n286,
    n414,
    n385
  );


  or
  g878
  (
    n844,
    n358,
    n343,
    n491,
    n365
  );


  xnor
  g879
  (
    n821,
    n209,
    n279,
    n272,
    n438
  );


  xnor
  g880
  (
    n816,
    n481,
    n173,
    n490,
    n451
  );


  or
  g881
  (
    n683,
    n464,
    n240,
    n273,
    n421
  );


  or
  g882
  (
    n723,
    n317,
    n338,
    n497,
    n363
  );


  or
  g883
  (
    n674,
    n453,
    n321,
    n311,
    n410
  );


  nor
  g884
  (
    n734,
    n412,
    n276,
    n455,
    n467
  );


  xnor
  g885
  (
    n675,
    n495,
    n320,
    n214,
    n383
  );


  and
  g886
  (
    n781,
    n490,
    n257,
    n302,
    n380
  );


  xnor
  g887
  (
    n703,
    n322,
    n365,
    n358,
    n269
  );


  or
  g888
  (
    n718,
    n363,
    n481,
    n487,
    n442
  );


  and
  g889
  (
    n798,
    n355,
    n182,
    n421,
    n270
  );


  nor
  g890
  (
    n919,
    n483,
    n278,
    n281
  );


  nor
  g891
  (
    n738,
    n429,
    n332,
    n467,
    n442
  );


  nand
  g892
  (
    n858,
    n373,
    n470,
    n282,
    n372
  );


  and
  g893
  (
    n678,
    n415,
    n433,
    n460,
    n387
  );


  nand
  g894
  (
    n910,
    n493,
    n450,
    n320,
    n474
  );


  xor
  g895
  (
    n769,
    n437,
    n424,
    n296,
    n289
  );


  or
  g896
  (
    n818,
    n401,
    n213,
    n204,
    n420
  );


  xnor
  g897
  (
    n833,
    n489,
    n298,
    n441,
    n265
  );


  xor
  g898
  (
    n788,
    n309,
    n399,
    n389,
    n323
  );


  nand
  g899
  (
    n709,
    n337,
    n440,
    n322,
    n351
  );


  xor
  g900
  (
    n699,
    n492,
    n431,
    n387,
    n360
  );


  xnor
  g901
  (
    n762,
    n437,
    n420,
    n415,
    n215
  );


  nand
  g902
  (
    n710,
    n291,
    n307,
    n441,
    n458
  );


  nor
  g903
  (
    n928,
    n451,
    n385,
    n337,
    n425
  );


  or
  g904
  (
    n934,
    n464,
    n262,
    n462,
    n394
  );


  xnor
  g905
  (
    n698,
    n345,
    n371,
    n365,
    n261
  );


  nand
  g906
  (
    n874,
    n201,
    n409,
    n350,
    n228
  );


  nand
  g907
  (
    n835,
    n162,
    n475,
    n413,
    n305
  );


  or
  g908
  (
    n1148,
    n640,
    n605,
    n569,
    n887
  );


  nand
  g909
  (
    n982,
    n638,
    n536,
    n515,
    n636
  );


  xnor
  g910
  (
    n1041,
    n592,
    n631,
    n500,
    n572
  );


  xnor
  g911
  (
    n1070,
    n704,
    n749,
    n620,
    n518
  );


  nand
  g912
  (
    n1149,
    n560,
    n529,
    n615,
    n587
  );


  or
  g913
  (
    n1046,
    n502,
    n574,
    n659,
    n549
  );


  xnor
  g914
  (
    n1098,
    n630,
    n514,
    n622,
    n886
  );


  and
  g915
  (
    n1133,
    n512,
    n641,
    n647,
    n607
  );


  xor
  g916
  (
    n1107,
    n601,
    n659,
    n756,
    n658
  );


  nand
  g917
  (
    n1109,
    n534,
    n666,
    n632,
    n686
  );


  or
  g918
  (
    n1152,
    n864,
    n551,
    n611,
    n733
  );


  nor
  g919
  (
    n1075,
    n718,
    n654,
    n594,
    n633
  );


  or
  g920
  (
    n963,
    n646,
    n503,
    n530,
    n578
  );


  nand
  g921
  (
    n1092,
    n593,
    n521,
    n586,
    n509
  );


  xor
  g922
  (
    n1037,
    n577,
    n649,
    n595,
    n548
  );


  and
  g923
  (
    n956,
    n600,
    n598,
    n627,
    n893
  );


  nor
  g924
  (
    n1047,
    n667,
    n602,
    n800,
    n590
  );


  or
  g925
  (
    n1159,
    n505,
    n649,
    n598,
    n645
  );


  xor
  g926
  (
    n1134,
    n820,
    n668,
    n859,
    n727
  );


  xnor
  g927
  (
    n988,
    n506,
    n755,
    n678,
    n510
  );


  xnor
  g928
  (
    n977,
    n602,
    n603,
    n528,
    n648
  );


  nand
  g929
  (
    n1061,
    n639,
    n525,
    n837,
    n599
  );


  and
  g930
  (
    n1150,
    n597,
    n843,
    n762,
    n620
  );


  xnor
  g931
  (
    n979,
    n879,
    n809,
    n556,
    n836
  );


  xor
  g932
  (
    n1043,
    n806,
    n657,
    n882,
    n808
  );


  xor
  g933
  (
    n1019,
    n878,
    n650,
    n831,
    n517
  );


  and
  g934
  (
    n1027,
    n612,
    n518,
    n770,
    n594
  );


  nand
  g935
  (
    n1062,
    n615,
    n612,
    n601,
    n510
  );


  xor
  g936
  (
    n1066,
    n509,
    n612,
    n703,
    n782
  );


  nand
  g937
  (
    n1079,
    n559,
    n580,
    n603,
    n554
  );


  nor
  g938
  (
    n1108,
    n614,
    n547,
    n648,
    n661
  );


  and
  g939
  (
    KeyWire_0_15,
    n559,
    n504,
    n766,
    n853
  );


  and
  g940
  (
    n966,
    n538,
    n534,
    n740,
    n846
  );


  xnor
  g941
  (
    n1165,
    n544,
    n535,
    n790,
    n632
  );


  and
  g942
  (
    n1063,
    n589,
    n659,
    n550,
    n665
  );


  and
  g943
  (
    n1073,
    n535,
    n513,
    n574,
    n503
  );


  xor
  g944
  (
    n1031,
    n714,
    n529,
    n516,
    n628
  );


  xnor
  g945
  (
    n1124,
    n657,
    n757,
    n812,
    n538
  );


  xor
  g946
  (
    n1033,
    n538,
    n675,
    n735,
    n665
  );


  xor
  g947
  (
    n952,
    n532,
    n590,
    n639,
    n585
  );


  or
  g948
  (
    n1096,
    n610,
    n619,
    n581,
    n695
  );


  xnor
  g949
  (
    n1029,
    n642,
    n616,
    n537,
    n676
  );


  nor
  g950
  (
    n980,
    n515,
    n765,
    n510,
    n728
  );


  xnor
  g951
  (
    n1086,
    n842,
    n521,
    n643,
    n701
  );


  nor
  g952
  (
    n1099,
    n573,
    n604,
    n779,
    n521
  );


  nor
  g953
  (
    n954,
    n577,
    n869,
    n618,
    n657
  );


  nor
  g954
  (
    n984,
    n506,
    n594,
    n571,
    n513
  );


  nand
  g955
  (
    n1163,
    n553,
    n629,
    n562,
    n517
  );


  nor
  g956
  (
    n969,
    n531,
    n691,
    n710,
    n620
  );


  xor
  g957
  (
    n983,
    n635,
    n738,
    n645,
    n816
  );


  or
  g958
  (
    n1128,
    n606,
    n900,
    n777,
    n797
  );


  xor
  g959
  (
    n1007,
    n641,
    n507,
    n570,
    n523
  );


  nor
  g960
  (
    n1009,
    n559,
    n776,
    n530,
    n641
  );


  xor
  g961
  (
    n1156,
    n586,
    n668,
    n561,
    n522
  );


  nor
  g962
  (
    n1054,
    n511,
    n606,
    n567,
    n637
  );


  nor
  g963
  (
    n949,
    n538,
    n519,
    n540,
    n520
  );


  and
  g964
  (
    n987,
    n665,
    n616,
    n888,
    n516
  );


  nor
  g965
  (
    n1008,
    n519,
    n600,
    n612,
    n635
  );


  xor
  g966
  (
    n955,
    n528,
    n590,
    n608,
    n663
  );


  xor
  g967
  (
    n944,
    n659,
    n614,
    n767,
    n543
  );


  xnor
  g968
  (
    n1132,
    n744,
    n505,
    n646,
    n563
  );


  xor
  g969
  (
    KeyWire_0_9,
    n663,
    n535,
    n504,
    n698
  );


  xor
  g970
  (
    n989,
    n817,
    n634,
    n522,
    n615
  );


  or
  g971
  (
    n981,
    n523,
    n562,
    n617,
    n582
  );


  xor
  g972
  (
    n1042,
    n536,
    n699,
    n575,
    n500
  );


  xor
  g973
  (
    n1144,
    n527,
    n608,
    n603,
    n563
  );


  xnor
  g974
  (
    n1069,
    n533,
    n655,
    n540,
    n568
  );


  and
  g975
  (
    n959,
    n717,
    n605,
    n543,
    n683
  );


  nor
  g976
  (
    n960,
    n720,
    n566,
    n531,
    n557
  );


  nor
  g977
  (
    n994,
    n619,
    n752,
    n662,
    n898
  );


  or
  g978
  (
    n1064,
    n589,
    n645,
    n581,
    n793
  );


  xor
  g979
  (
    n1111,
    n653,
    n540,
    n833,
    n579
  );


  or
  g980
  (
    n1091,
    n753,
    n617,
    n630,
    n524
  );


  or
  g981
  (
    n1089,
    n880,
    n636,
    n628,
    n525
  );


  or
  g982
  (
    n1038,
    n841,
    n845,
    n550
  );


  xnor
  g983
  (
    n1093,
    n537,
    n871,
    n571,
    n541
  );


  xor
  g984
  (
    n1074,
    n618,
    n613,
    n614,
    n642
  );


  nand
  g985
  (
    n992,
    n828,
    n608,
    n537,
    n680
  );


  and
  g986
  (
    n999,
    n515,
    n629,
    n599,
    n607
  );


  xor
  g987
  (
    n942,
    n874,
    n811,
    n835,
    n677
  );


  xnor
  g988
  (
    n1115,
    n660,
    n656,
    n629,
    n534
  );


  xor
  g989
  (
    n1100,
    n741,
    n666,
    n590,
    n622
  );


  xor
  g990
  (
    n1157,
    n876,
    n570,
    n526,
    n865
  );


  nand
  g991
  (
    n1114,
    n583,
    n600,
    n601,
    n517
  );


  or
  g992
  (
    n1013,
    n575,
    n604,
    n527,
    n715
  );


  xor
  g993
  (
    n1000,
    n644,
    n507,
    n891,
    n557
  );


  or
  g994
  (
    n1143,
    n568,
    n557,
    n664,
    n592
  );


  and
  g995
  (
    n1095,
    n546,
    n613,
    n625,
    n595
  );


  or
  g996
  (
    n1056,
    n520,
    n839,
    n791,
    n635
  );


  or
  g997
  (
    n1105,
    n587,
    n524,
    n774,
    n775
  );


  and
  g998
  (
    n976,
    n636,
    n652,
    n544,
    n586
  );


  xor
  g999
  (
    KeyWire_0_7,
    n539,
    n564,
    n730,
    n649
  );


  nor
  g1000
  (
    n993,
    n586,
    n826,
    n642,
    n796
  );


  and
  g1001
  (
    n1022,
    n854,
    n892,
    n631,
    n834
  );


  nor
  g1002
  (
    n1080,
    n705,
    n618,
    n515,
    n801
  );


  nand
  g1003
  (
    n1025,
    n795,
    n579,
    n502,
    n522
  );


  and
  g1004
  (
    n1094,
    n576,
    n589,
    n688,
    n747
  );


  or
  g1005
  (
    n1118,
    n610,
    n638,
    n783,
    n643
  );


  nand
  g1006
  (
    KeyWire_0_2,
    n664,
    n549,
    n622,
    n588
  );


  and
  g1007
  (
    n1001,
    n585,
    n499,
    n535,
    n639
  );


  nor
  g1008
  (
    n1034,
    n870,
    n823,
    n521,
    n504
  );


  or
  g1009
  (
    n1136,
    n550,
    n792,
    n598,
    n542
  );


  xnor
  g1010
  (
    n1116,
    n514,
    n637,
    n570,
    n739
  );


  xor
  g1011
  (
    n1015,
    n519,
    n868,
    n615,
    n732
  );


  nor
  g1012
  (
    n968,
    n555,
    n580,
    n664,
    n563
  );


  nor
  g1013
  (
    n1050,
    n802,
    n501,
    n573,
    n863
  );


  xnor
  g1014
  (
    n1102,
    n611,
    n650,
    n531,
    n520
  );


  xor
  g1015
  (
    n1123,
    n789,
    n697,
    n799,
    n584
  );


  nor
  g1016
  (
    n1032,
    n662,
    n507,
    n501,
    n585
  );


  xor
  g1017
  (
    n1028,
    n760,
    n544,
    n606,
    n661
  );


  xor
  g1018
  (
    n1011,
    n584,
    n572,
    n518,
    n685
  );


  xnor
  g1019
  (
    n1018,
    n651,
    n707,
    n643,
    n655
  );


  nand
  g1020
  (
    n943,
    n528,
    n626,
    n623,
    n593
  );


  or
  g1021
  (
    n1067,
    n696,
    n548,
    n651,
    n572
  );


  nand
  g1022
  (
    n1090,
    n556,
    n572,
    n566,
    n724
  );


  and
  g1023
  (
    n974,
    n588,
    n647,
    n627,
    n591
  );


  nor
  g1024
  (
    n1110,
    n508,
    n621,
    n526,
    n569
  );


  or
  g1025
  (
    n1164,
    n523,
    n541,
    n609,
    n575
  );


  xor
  g1026
  (
    n1087,
    n564,
    n646,
    n595,
    n848
  );


  xor
  g1027
  (
    n1048,
    n667,
    n524,
    n608,
    n540
  );


  and
  g1028
  (
    n1068,
    n784,
    n539,
    n578,
    n547
  );


  xor
  g1029
  (
    n1057,
    n661,
    n617,
    n885,
    n507
  );


  nand
  g1030
  (
    n1077,
    n838,
    n743,
    n596,
    n543
  );


  nor
  g1031
  (
    n1162,
    n682,
    n872,
    n599,
    n713
  );


  xnor
  g1032
  (
    n1076,
    n668,
    n509,
    n712,
    n532
  );


  nand
  g1033
  (
    n946,
    n579,
    n822,
    n561,
    n616
  );


  xnor
  g1034
  (
    n1160,
    n541,
    n821,
    n644,
    n624
  );


  or
  g1035
  (
    n1101,
    n585,
    n751,
    n645,
    n623
  );


  nand
  g1036
  (
    n1053,
    n679,
    n617,
    n810,
    n737
  );


  nand
  g1037
  (
    n1142,
    n505,
    n895,
    n654,
    n638
  );


  or
  g1038
  (
    n1131,
    n622,
    n580,
    n805,
    n537
  );


  xor
  g1039
  (
    n985,
    n716,
    n827,
    n505,
    n551
  );


  xor
  g1040
  (
    n1045,
    n544,
    n693,
    n546,
    n794
  );


  or
  g1041
  (
    n948,
    n897,
    n589,
    n706,
    n815
  );


  or
  g1042
  (
    n1005,
    n651,
    n639,
    n851,
    n502
  );


  nor
  g1043
  (
    n971,
    n662,
    n655,
    n736,
    n648
  );


  nor
  g1044
  (
    n986,
    n819,
    n640,
    n778,
    n502
  );


  nand
  g1045
  (
    n1039,
    n609,
    n554,
    n829,
    n624
  );


  nand
  g1046
  (
    n945,
    n654,
    n581,
    n588
  );


  xnor
  g1047
  (
    n947,
    n553,
    n519,
    n689,
    n652
  );


  nand
  g1048
  (
    n1121,
    n850,
    n875,
    n771,
    n619
  );


  xor
  g1049
  (
    n1104,
    n630,
    n648,
    n511,
    n745
  );


  and
  g1050
  (
    n1112,
    n576,
    n605,
    n656,
    n582
  );


  nand
  g1051
  (
    n1141,
    n577,
    n866,
    n553,
    n616
  );


  or
  g1052
  (
    n1036,
    n621,
    n532,
    n511,
    n559
  );


  xor
  g1053
  (
    n1072,
    n504,
    n514,
    n556,
    n552
  );


  xnor
  g1054
  (
    n1129,
    n877,
    n803,
    n595,
    n596
  );


  xor
  g1055
  (
    n1153,
    n726,
    n646,
    n644,
    n541
  );


  and
  g1056
  (
    n1154,
    n587,
    n536,
    n861,
    n746
  );


  nor
  g1057
  (
    n951,
    n692,
    n596,
    n593,
    n506
  );


  or
  g1058
  (
    n1017,
    n621,
    n856,
    n534,
    n840
  );


  and
  g1059
  (
    n1044,
    n578,
    n609,
    n619,
    n527
  );


  or
  g1060
  (
    n1055,
    n632,
    n641,
    n721,
    n552
  );


  and
  g1061
  (
    n1020,
    n501,
    n547,
    n530,
    n602
  );


  or
  g1062
  (
    n1125,
    n652,
    n526,
    n832,
    n633
  );


  nor
  g1063
  (
    n1051,
    n661,
    n763,
    n729,
    n665
  );


  xor
  g1064
  (
    n1016,
    n625,
    n798,
    n613,
    n830
  );


  or
  g1065
  (
    n1059,
    n565,
    n533,
    n660,
    n722
  );


  nand
  g1066
  (
    n1126,
    n786,
    n583,
    n633,
    n587
  );


  nor
  g1067
  (
    n1113,
    n542,
    n614,
    n658,
    n620
  );


  nand
  g1068
  (
    n995,
    n666,
    n857,
    n607,
    n564
  );


  nor
  g1069
  (
    n1030,
    n600,
    n700,
    n862,
    n621
  );


  xor
  g1070
  (
    n997,
    n558,
    n643,
    n690,
    n660
  );


  xor
  g1071
  (
    n970,
    n593,
    n569,
    n561,
    n528
  );


  nor
  g1072
  (
    n1085,
    n825,
    n525,
    n899,
    n663
  );


  xnor
  g1073
  (
    n961,
    n579,
    n558,
    n543
  );


  nor
  g1074
  (
    n1127,
    n889,
    n884,
    n626,
    n630
  );


  nand
  g1075
  (
    n973,
    n582,
    n855,
    n568,
    n633
  );


  xor
  g1076
  (
    n975,
    n570,
    n653,
    n545,
    n580
  );


  nand
  g1077
  (
    n1010,
    n552,
    n613,
    n631,
    n635
  );


  nor
  g1078
  (
    n1146,
    n516,
    n571,
    n634,
    n847
  );


  and
  g1079
  (
    n1103,
    n546,
    n560,
    n500,
    n708
  );


  and
  g1080
  (
    n957,
    n522,
    n627,
    n601,
    n781
  );


  xnor
  g1081
  (
    n1012,
    n571,
    n629,
    n567,
    n563
  );


  nand
  g1082
  (
    n1122,
    n592,
    n561,
    n558,
    n565
  );


  xor
  g1083
  (
    n991,
    n583,
    n551,
    n636,
    n759
  );


  xor
  g1084
  (
    n1014,
    n574,
    n573,
    n638,
    n582
  );


  xor
  g1085
  (
    n1151,
    n557,
    n512,
    n666,
    n576
  );


  and
  g1086
  (
    n1097,
    n512,
    n533,
    n529,
    n642
  );


  xor
  g1087
  (
    n1155,
    n725,
    n625,
    n592,
    n742
  );


  and
  g1088
  (
    n1052,
    n653,
    n539,
    n511,
    n702
  );


  nor
  g1089
  (
    n962,
    n577,
    n548,
    n723,
    n536
  );


  nor
  g1090
  (
    n1166,
    n644,
    n560,
    n552,
    n525
  );


  and
  g1091
  (
    n998,
    n598,
    n576,
    n768,
    n656
  );


  nor
  g1092
  (
    n1023,
    n566,
    n565,
    n769,
    n508
  );


  and
  g1093
  (
    n1065,
    n611,
    n547,
    n849,
    n605
  );


  nor
  g1094
  (
    n958,
    n750,
    n780,
    n660,
    n664
  );


  xnor
  g1095
  (
    n1049,
    n551,
    n883,
    n628,
    n556
  );


  xor
  g1096
  (
    n996,
    n637,
    n567,
    n658,
    n545
  );


  xor
  g1097
  (
    n1083,
    n518,
    n647,
    n533,
    n549
  );


  and
  g1098
  (
    n1006,
    n787,
    n567,
    n609,
    n542
  );


  nor
  g1099
  (
    n1002,
    n632,
    n640,
    n748,
    n503
  );


  nand
  g1100
  (
    n1140,
    n555,
    n553,
    n554,
    n734
  );


  or
  g1101
  (
    n1040,
    n896,
    n509,
    n584,
    n627
  );


  nand
  g1102
  (
    n990,
    n532,
    n510,
    n555,
    n512
  );


  and
  g1103
  (
    n1139,
    n529,
    n565,
    n623,
    n596
  );


  or
  g1104
  (
    n978,
    n545,
    n813,
    n890,
    n574
  );


  xnor
  g1105
  (
    n1078,
    n618,
    n731,
    n514,
    n761
  );


  nand
  g1106
  (
    n1119,
    n562,
    n852,
    n591,
    n773
  );


  and
  g1107
  (
    n1145,
    n545,
    n807,
    n814,
    n662
  );


  nor
  g1108
  (
    n1060,
    n555,
    n597,
    n566,
    n611
  );


  xor
  g1109
  (
    n1120,
    n684,
    n594,
    n573,
    n531
  );


  xor
  g1110
  (
    n953,
    n569,
    n772,
    n513,
    n719
  );


  or
  g1111
  (
    n1082,
    n578,
    n597,
    n560,
    n658
  );


  and
  g1112
  (
    n1003,
    n568,
    n562,
    n881,
    n709
  );


  or
  g1113
  (
    n1161,
    n610,
    n575,
    n524,
    n694
  );


  xnor
  g1114
  (
    n1035,
    n526,
    n506,
    n508,
    n818
  );


  nor
  g1115
  (
    n941,
    n804,
    n867,
    n824,
    n523
  );


  and
  g1116
  (
    n1084,
    n501,
    n656,
    n764,
    n650
  );


  and
  g1117
  (
    n964,
    n623,
    n626,
    n583
  );


  and
  g1118
  (
    n1137,
    n548,
    n651,
    n508,
    n527
  );


  or
  g1119
  (
    n1088,
    n711,
    n844,
    n637,
    n647
  );


  xnor
  g1120
  (
    n972,
    n591,
    n624,
    n681,
    n606
  );


  xor
  g1121
  (
    n1130,
    n530,
    n663,
    n894,
    n599
  );


  xor
  g1122
  (
    n1106,
    n858,
    n517,
    n754,
    n652
  );


  xor
  g1123
  (
    n1117,
    n542,
    n650,
    n624,
    n667
  );


  and
  g1124
  (
    n965,
    n657,
    n785,
    n520,
    n499
  );


  and
  g1125
  (
    n1058,
    n539,
    n607,
    n549,
    n602
  );


  nand
  g1126
  (
    n1135,
    n634,
    n653,
    n655,
    n604
  );


  nand
  g1127
  (
    n1004,
    n581,
    n654,
    n610,
    n513
  );


  and
  g1128
  (
    n1138,
    n667,
    n788,
    n500,
    n860
  );


  nand
  g1129
  (
    n1147,
    n516,
    n649,
    n640,
    n564
  );


  xnor
  g1130
  (
    n950,
    n634,
    n628,
    n604,
    n584
  );


  or
  g1131
  (
    n1026,
    n687,
    n591,
    n668,
    n631
  );


  nor
  g1132
  (
    n1081,
    n546,
    n873,
    n758,
    n503
  );


  nand
  g1133
  (
    n1158,
    n603,
    n625,
    n554,
    n597
  );


  or
  g1134
  (
    n1194,
    n933,
    n1004,
    n960,
    n916
  );


  xor
  g1135
  (
    n1168,
    n1015,
    n1049,
    n943,
    n1013
  );


  xor
  g1136
  (
    n1171,
    n911,
    n932,
    n1063,
    n1068
  );


  xor
  g1137
  (
    n1176,
    n907,
    n915,
    n1054,
    n957
  );


  or
  g1138
  (
    n1172,
    n1023,
    n924,
    n920,
    n972
  );


  xnor
  g1139
  (
    n1202,
    n927,
    n1017,
    n1011,
    n1066
  );


  nand
  g1140
  (
    n1197,
    n1067,
    n903,
    n925,
    n975
  );


  nor
  g1141
  (
    n1186,
    n948,
    n968,
    n1032,
    n1069
  );


  and
  g1142
  (
    KeyWire_0_3,
    n1018,
    n1074,
    n909,
    n1061
  );


  nor
  g1143
  (
    n1196,
    n934,
    n964,
    n990,
    n996
  );


  nand
  g1144
  (
    n1169,
    n1012,
    n984,
    n917,
    n1019
  );


  nor
  g1145
  (
    n1195,
    n1031,
    n985,
    n904,
    n978
  );


  nand
  g1146
  (
    n1207,
    n1036,
    n1059,
    n918,
    n1041
  );


  and
  g1147
  (
    n1187,
    n1008,
    n1046,
    n914,
    n1070
  );


  xor
  g1148
  (
    n1184,
    n999,
    n1025,
    n912,
    n988
  );


  nor
  g1149
  (
    n1191,
    n1053,
    n1035,
    n1052,
    n942
  );


  nor
  g1150
  (
    n1204,
    n958,
    n1022,
    n928,
    n902
  );


  or
  g1151
  (
    n1201,
    n1006,
    n908,
    n950,
    n997
  );


  or
  g1152
  (
    n1181,
    n1062,
    n959,
    n966,
    n973
  );


  or
  g1153
  (
    n1173,
    n1065,
    n923,
    n989,
    n1047
  );


  or
  g1154
  (
    n1175,
    n986,
    n1021,
    n952,
    n969
  );


  xor
  g1155
  (
    n1208,
    n1034,
    n1030,
    n1027,
    n955
  );


  nand
  g1156
  (
    n1189,
    n1003,
    n1029,
    n998,
    n1073
  );


  and
  g1157
  (
    n1200,
    n944,
    n971,
    n1064,
    n1039
  );


  xor
  g1158
  (
    n1180,
    n1048,
    n931,
    n947,
    n921
  );


  or
  g1159
  (
    n1177,
    n981,
    n995,
    n1009,
    n976
  );


  or
  g1160
  (
    n1182,
    n929,
    n919,
    n974,
    n953
  );


  xnor
  g1161
  (
    n1206,
    n930,
    n956,
    n946,
    n1055
  );


  xnor
  g1162
  (
    n1185,
    n901,
    n1057,
    n991,
    n1010
  );


  or
  g1163
  (
    n1179,
    n1038,
    n1040,
    n951,
    n1028
  );


  and
  g1164
  (
    n1167,
    n1005,
    n906,
    n1037,
    n1002
  );


  xor
  g1165
  (
    n1190,
    n967,
    n970,
    n1051,
    n1020
  );


  and
  g1166
  (
    n1192,
    n1000,
    n1043,
    n1058,
    n941
  );


  or
  g1167
  (
    n1178,
    n1042,
    n1044,
    n949,
    n926
  );


  xnor
  g1168
  (
    n1193,
    n910,
    n1026,
    n980,
    n1016
  );


  and
  g1169
  (
    n1203,
    n1007,
    n983,
    n945,
    n994
  );


  nor
  g1170
  (
    n1174,
    n987,
    n913,
    n905,
    n922
  );


  nand
  g1171
  (
    n1188,
    n993,
    n1056,
    n1024,
    n1050
  );


  xor
  g1172
  (
    n1170,
    n982,
    n992,
    n1071,
    n1014
  );


  or
  g1173
  (
    n1198,
    n954,
    n979,
    n1001,
    n977
  );


  or
  g1174
  (
    n1199,
    n1033,
    n1060,
    n961,
    n962
  );


  xor
  g1175
  (
    n1205,
    n1072,
    n965,
    n1045,
    n963
  );


  nand
  g1176
  (
    n1222,
    n1079,
    n1145,
    n1195
  );


  nand
  g1177
  (
    n1214,
    n1098,
    n1119,
    n1189
  );


  nor
  g1178
  (
    n1211,
    n1107,
    n1133,
    n1150,
    n1132
  );


  xor
  g1179
  (
    n1212,
    n1105,
    n1193,
    n1115,
    n1096
  );


  nor
  g1180
  (
    n1220,
    n1087,
    n1192,
    n1139,
    n1086
  );


  nor
  g1181
  (
    n1226,
    n1116,
    n1190,
    n1184,
    n1185
  );


  xnor
  g1182
  (
    n1218,
    n1117,
    n1147,
    n1148,
    n1089
  );


  and
  g1183
  (
    n1227,
    n1095,
    n1099,
    n1138,
    n1202
  );


  xor
  g1184
  (
    n1217,
    n1142,
    n1084,
    n1194,
    n1088
  );


  xnor
  g1185
  (
    n1234,
    n1091,
    n1094,
    n1082,
    n1125
  );


  xnor
  g1186
  (
    n1230,
    n1141,
    n1118,
    n1093,
    n1108
  );


  xor
  g1187
  (
    n1213,
    n1104,
    n1123,
    n1114,
    n1078
  );


  xnor
  g1188
  (
    n1219,
    n1129,
    n1201,
    n1090,
    n1134
  );


  xor
  g1189
  (
    n1210,
    n1181,
    n1077,
    n1198,
    n1200
  );


  or
  g1190
  (
    n1223,
    n1186,
    n1113,
    n1203,
    n1110
  );


  nand
  g1191
  (
    n1216,
    n1146,
    n1140,
    n1076,
    n1191
  );


  nor
  g1192
  (
    n1232,
    n1135,
    n1130,
    n1122,
    n1187
  );


  nor
  g1193
  (
    n1225,
    n1182,
    n1083,
    n1131,
    n1106
  );


  and
  g1194
  (
    n1209,
    n1097,
    n1124,
    n1197,
    n1128
  );


  nor
  g1195
  (
    n1228,
    n1112,
    n1188,
    n1137,
    n1111
  );


  xnor
  g1196
  (
    n1231,
    n1136,
    n1075,
    n1101,
    n1103
  );


  and
  g1197
  (
    n1215,
    n1179,
    n1143,
    n1127,
    n1183
  );


  and
  g1198
  (
    n1224,
    n1092,
    n1085,
    n1126,
    n1081
  );


  xor
  g1199
  (
    KeyWire_0_6,
    n1180,
    n1120,
    n1199,
    n1121
  );


  xor
  g1200
  (
    n1233,
    n1204,
    n1196,
    n1109,
    n1080
  );


  nand
  g1201
  (
    n1229,
    n1102,
    n1149,
    n1144,
    n1100
  );


  not
  g1202
  (
    n1258,
    n1154
  );


  not
  g1203
  (
    n1256,
    n1233
  );


  buf
  g1204
  (
    n1240,
    n1225
  );


  buf
  g1205
  (
    n1238,
    n1151
  );


  not
  g1206
  (
    n1248,
    n1222
  );


  not
  g1207
  (
    n1247,
    n1152
  );


  not
  g1208
  (
    n1235,
    n1219
  );


  not
  g1209
  (
    n1242,
    n1223
  );


  buf
  g1210
  (
    n1237,
    n1210
  );


  not
  g1211
  (
    n1236,
    n1215
  );


  not
  g1212
  (
    n1252,
    n1226
  );


  buf
  g1213
  (
    n1253,
    n1221
  );


  buf
  g1214
  (
    n1260,
    n1212
  );


  not
  g1215
  (
    n1239,
    n1214
  );


  buf
  g1216
  (
    n1250,
    n1153
  );


  buf
  g1217
  (
    n1254,
    n1216
  );


  not
  g1218
  (
    n1241,
    n1227
  );


  not
  g1219
  (
    n1246,
    n1234
  );


  not
  g1220
  (
    n1245,
    n1211
  );


  buf
  g1221
  (
    n1251,
    n1232
  );


  not
  g1222
  (
    n1244,
    n1220
  );


  not
  g1223
  (
    n1255,
    n1218
  );


  nand
  g1224
  (
    n1257,
    n1224,
    n1230
  );


  and
  g1225
  (
    n1249,
    n1228,
    n1234
  );


  and
  g1226
  (
    n1243,
    n1229,
    n1217
  );


  nor
  g1227
  (
    n1259,
    n1209,
    n1155
  );


  xnor
  g1228
  (
    n1261,
    n1231,
    n1213
  );


  not
  g1229
  (
    n1302,
    n1243
  );


  not
  g1230
  (
    n1312,
    n1235
  );


  not
  g1231
  (
    n1325,
    n1249
  );


  buf
  g1232
  (
    n1262,
    n1250
  );


  not
  g1233
  (
    n1275,
    n1242
  );


  buf
  g1234
  (
    n1267,
    n1240
  );


  not
  g1235
  (
    n1335,
    n1248
  );


  not
  g1236
  (
    n1276,
    n1248
  );


  not
  g1237
  (
    n1310,
    n1253
  );


  not
  g1238
  (
    n1296,
    n1251
  );


  not
  g1239
  (
    n1271,
    n1238
  );


  not
  g1240
  (
    n1332,
    n1254
  );


  not
  g1241
  (
    n1265,
    n1247
  );


  buf
  g1242
  (
    n1334,
    n1240
  );


  not
  g1243
  (
    n1329,
    n1254
  );


  not
  g1244
  (
    n1294,
    n1248
  );


  buf
  g1245
  (
    n1311,
    n1236
  );


  buf
  g1246
  (
    n1322,
    n1242
  );


  not
  g1247
  (
    n1326,
    n1235
  );


  buf
  g1248
  (
    n1331,
    n1247
  );


  not
  g1249
  (
    n1338,
    n1242
  );


  buf
  g1250
  (
    n1297,
    n1252
  );


  buf
  g1251
  (
    n1288,
    n1241
  );


  buf
  g1252
  (
    n1336,
    n1237
  );


  not
  g1253
  (
    n1289,
    n1239
  );


  buf
  g1254
  (
    n1304,
    n1241
  );


  not
  g1255
  (
    n1290,
    n1237
  );


  not
  g1256
  (
    n1284,
    n1246
  );


  not
  g1257
  (
    n1274,
    n1247
  );


  buf
  g1258
  (
    n1317,
    n1243
  );


  not
  g1259
  (
    n1330,
    n1241
  );


  buf
  g1260
  (
    n1269,
    n1237
  );


  buf
  g1261
  (
    n1318,
    n1237
  );


  buf
  g1262
  (
    n1295,
    n1244
  );


  not
  g1263
  (
    n1301,
    n1254
  );


  not
  g1264
  (
    n1314,
    n1235
  );


  not
  g1265
  (
    n1263,
    n1253
  );


  not
  g1266
  (
    n1278,
    n1249
  );


  not
  g1267
  (
    n1327,
    n1249
  );


  buf
  g1268
  (
    n1292,
    n1243
  );


  buf
  g1269
  (
    n1266,
    n1253
  );


  not
  g1270
  (
    n1293,
    n1240
  );


  not
  g1271
  (
    n1291,
    n1246
  );


  not
  g1272
  (
    n1287,
    n1251
  );


  buf
  g1273
  (
    n1303,
    n1236
  );


  not
  g1274
  (
    n1300,
    n1252
  );


  buf
  g1275
  (
    n1321,
    n1238
  );


  buf
  g1276
  (
    n1299,
    n1246
  );


  not
  g1277
  (
    n1283,
    n1244
  );


  buf
  g1278
  (
    n1273,
    n1238
  );


  buf
  g1279
  (
    n1340,
    n1249
  );


  not
  g1280
  (
    n1333,
    n1241
  );


  not
  g1281
  (
    n1268,
    n1250
  );


  buf
  g1282
  (
    n1324,
    n1246
  );


  buf
  g1283
  (
    n1308,
    n1254
  );


  buf
  g1284
  (
    n1341,
    n1238
  );


  buf
  g1285
  (
    n1313,
    n1239
  );


  not
  g1286
  (
    n1315,
    n1245
  );


  buf
  g1287
  (
    n1272,
    n1244
  );


  buf
  g1288
  (
    n1279,
    n1240
  );


  buf
  g1289
  (
    n1282,
    n1250
  );


  buf
  g1290
  (
    n1264,
    n1253
  );


  not
  g1291
  (
    n1316,
    n1242
  );


  buf
  g1292
  (
    n1277,
    n1235
  );


  not
  g1293
  (
    n1319,
    n1239
  );


  not
  g1294
  (
    n1320,
    n1251
  );


  not
  g1295
  (
    n1281,
    n1252
  );


  buf
  g1296
  (
    n1339,
    n1239
  );


  not
  g1297
  (
    n1309,
    n1251
  );


  not
  g1298
  (
    n1328,
    n1245
  );


  buf
  g1299
  (
    n1270,
    n1245
  );


  not
  g1300
  (
    n1337,
    n1250
  );


  buf
  g1301
  (
    n1280,
    n1248
  );


  buf
  g1302
  (
    n1306,
    n1245
  );


  not
  g1303
  (
    n1286,
    n1236
  );


  not
  g1304
  (
    n1307,
    n1247
  );


  buf
  g1305
  (
    n1305,
    n1244
  );


  buf
  g1306
  (
    n1323,
    n1236
  );


  not
  g1307
  (
    n1298,
    n1243
  );


  not
  g1308
  (
    n1285,
    n1252
  );


  xnor
  g1309
  (
    n1353,
    n1255,
    n1261,
    n1288,
    n1272
  );


  nand
  g1310
  (
    n1376,
    n1284,
    n1273,
    n1298,
    n1264
  );


  xnor
  g1311
  (
    n1346,
    n1293,
    n1269,
    n1291,
    n1264
  );


  nor
  g1312
  (
    n1364,
    n1290,
    n1276,
    n1299,
    n1257
  );


  and
  g1313
  (
    n1350,
    n1288,
    n1272,
    n1259,
    n1290
  );


  nand
  g1314
  (
    n1382,
    n1292,
    n1263,
    n1287,
    n1268
  );


  and
  g1315
  (
    n1361,
    n1284,
    n1301,
    n1265,
    n1283
  );


  xnor
  g1316
  (
    n1374,
    n1267,
    n1275,
    n1281,
    n1263
  );


  xnor
  g1317
  (
    n1383,
    n1262,
    n1270
  );


  xnor
  g1318
  (
    n1375,
    n1285,
    n1272,
    n1260,
    n1281
  );


  or
  g1319
  (
    n1363,
    n1274,
    n1269,
    n1278,
    n1277
  );


  and
  g1320
  (
    n1343,
    n1278,
    n1287,
    n1304,
    n1282
  );


  xor
  g1321
  (
    n1344,
    n1281,
    n1290,
    n1292,
    n1274
  );


  nand
  g1322
  (
    n1351,
    n1279,
    n1260,
    n1289,
    n1286
  );


  nand
  g1323
  (
    n1372,
    n1264,
    n1294,
    n1265,
    n1295
  );


  and
  g1324
  (
    n1370,
    n1276,
    n1275,
    n1289,
    n1260
  );


  xor
  g1325
  (
    n1391,
    n1301,
    n1294,
    n1258,
    n1302
  );


  or
  g1326
  (
    n1387,
    n1268,
    n1267,
    n1258,
    n1295
  );


  or
  g1327
  (
    n1362,
    n1298,
    n1271,
    n1264,
    n1289
  );


  or
  g1328
  (
    n1356,
    n1282,
    n1277,
    n1255,
    n1298
  );


  nand
  g1329
  (
    n1388,
    n1301,
    n1277,
    n1260,
    n1287
  );


  xor
  g1330
  (
    n1373,
    n1289,
    n1257,
    n1297,
    n1274
  );


  nor
  g1331
  (
    n1366,
    n1294,
    n1273,
    n1259,
    n1300
  );


  nor
  g1332
  (
    n1354,
    n1293,
    n1276,
    n1302,
    n1280
  );


  xnor
  g1333
  (
    n1378,
    n1266,
    n1271,
    n1270
  );


  nor
  g1334
  (
    n1347,
    n1303,
    n1295,
    n1262,
    n1256
  );


  nand
  g1335
  (
    n1385,
    n1285,
    n1276,
    n1274,
    n1265
  );


  and
  g1336
  (
    n1359,
    n1303,
    n1266,
    n1283,
    n1286
  );


  nand
  g1337
  (
    n1380,
    n1297,
    n1300,
    n1257
  );


  nor
  g1338
  (
    n1355,
    n1297,
    n1255,
    n1270,
    n1263
  );


  xor
  g1339
  (
    n1371,
    n1293,
    n1303,
    n1298,
    n1256
  );


  nand
  g1340
  (
    n1367,
    n1275,
    n1257,
    n1285,
    n1286
  );


  and
  g1341
  (
    n1384,
    n1256,
    n1266,
    n1285,
    n1296
  );


  nand
  g1342
  (
    n1357,
    n1299,
    n1303,
    n1258,
    n1291
  );


  and
  g1343
  (
    n1358,
    n1268,
    n1259,
    n1301,
    n1299
  );


  and
  g1344
  (
    n1368,
    n1255,
    n1280,
    n1279,
    n1261
  );


  or
  g1345
  (
    n1348,
    n1279,
    n1291,
    n1283,
    n1272
  );


  and
  g1346
  (
    n1379,
    n1282,
    n1290,
    n1267,
    n1291
  );


  nand
  g1347
  (
    n1381,
    n1273,
    n1271,
    n1302,
    n1284
  );


  and
  g1348
  (
    n1345,
    n1278,
    n1299,
    n1261,
    n1296
  );


  xor
  g1349
  (
    n1365,
    n1269,
    n1265,
    n1278,
    n1296
  );


  or
  g1350
  (
    n1352,
    n1280,
    n1268,
    n1273,
    n1284
  );


  xor
  g1351
  (
    n1386,
    n1288,
    n1287,
    n1304,
    n1261
  );


  or
  g1352
  (
    n1349,
    n1293,
    n1294,
    n1256,
    n1277
  );


  or
  g1353
  (
    n1369,
    n1258,
    n1269,
    n1292,
    n1295
  );


  and
  g1354
  (
    n1342,
    n1304,
    n1292,
    n1266,
    n1283
  );


  nor
  g1355
  (
    n1389,
    n1296,
    n1275,
    n1286,
    n1262
  );


  nand
  g1356
  (
    n1360,
    n1259,
    n1288,
    n1263,
    n1297
  );


  nand
  g1357
  (
    n1377,
    n1302,
    n1281,
    n1282,
    n1300
  );


  xor
  g1358
  (
    n1390,
    n1304,
    n1267,
    n1279,
    n1280
  );


  buf
  g1359
  (
    n1398,
    n1306
  );


  buf
  g1360
  (
    n1412,
    n1311
  );


  not
  g1361
  (
    n1414,
    n1305
  );


  not
  g1362
  (
    n1419,
    n1308
  );


  buf
  g1363
  (
    n1410,
    n1347
  );


  not
  g1364
  (
    n1400,
    n1313
  );


  buf
  g1365
  (
    n1406,
    n1312
  );


  not
  g1366
  (
    n1417,
    n1365
  );


  not
  g1367
  (
    n1422,
    n1358
  );


  not
  g1368
  (
    n1404,
    n1343
  );


  buf
  g1369
  (
    n1408,
    n1369
  );


  not
  g1370
  (
    n1403,
    n1315
  );


  buf
  g1371
  (
    n1423,
    n1313
  );


  not
  g1372
  (
    n1415,
    n1367
  );


  not
  g1373
  (
    n1394,
    n1346
  );


  buf
  g1374
  (
    n1407,
    n1307
  );


  buf
  g1375
  (
    n1418,
    n1315
  );


  not
  g1376
  (
    n1401,
    n1313
  );


  not
  g1377
  (
    n1420,
    n1310
  );


  buf
  g1378
  (
    n1413,
    n1316
  );


  xnor
  g1379
  (
    n1393,
    n1352,
    n1307,
    n1362,
    n1305
  );


  xor
  g1380
  (
    n1425,
    n1309,
    n1363,
    n1311,
    n1306
  );


  nand
  g1381
  (
    n1421,
    n1309,
    n1351,
    n1370,
    n1345
  );


  nand
  g1382
  (
    n1409,
    n1356,
    n1364,
    n1312,
    n1355
  );


  xnor
  g1383
  (
    n1405,
    n1308,
    n1305,
    n1376
  );


  or
  g1384
  (
    n1411,
    n1361,
    n1312,
    n1315,
    n1307
  );


  nor
  g1385
  (
    n1426,
    n1307,
    n1310,
    n1374,
    n1371
  );


  xor
  g1386
  (
    n1399,
    n1350,
    n1308,
    n1306,
    n1314
  );


  and
  g1387
  (
    n1416,
    n1344,
    n1309,
    n1357,
    n1375
  );


  nand
  g1388
  (
    n1397,
    n1349,
    n1308,
    n1314,
    n1372
  );


  xnor
  g1389
  (
    n1392,
    n1312,
    n1310,
    n1309
  );


  xnor
  g1390
  (
    n1424,
    n1315,
    n1314,
    n1313
  );


  nor
  g1391
  (
    n1395,
    n1353,
    n1359,
    n1311,
    n1342
  );


  xor
  g1392
  (
    n1396,
    n1373,
    n1311,
    n1354,
    n1348
  );


  xor
  g1393
  (
    n1402,
    n1368,
    n1306,
    n1366,
    n1360
  );


  not
  g1394
  (
    n1434,
    n1394
  );


  not
  g1395
  (
    n1429,
    n1393
  );


  not
  g1396
  (
    n1431,
    n1317
  );


  buf
  g1397
  (
    n1427,
    n1397
  );


  buf
  g1398
  (
    n1433,
    n1397
  );


  buf
  g1399
  (
    n1436,
    n1398
  );


  buf
  g1400
  (
    n1428,
    n1396
  );


  buf
  g1401
  (
    n1437,
    n1316
  );


  buf
  g1402
  (
    n1432,
    n1397
  );


  xnor
  g1403
  (
    n1430,
    n1398,
    n1317
  );


  nand
  g1404
  (
    n1435,
    n1395,
    n1398,
    n1316
  );


  xnor
  g1405
  (
    n1438,
    n1436,
    n1328,
    n1326,
    n1320
  );


  or
  g1406
  (
    n1479,
    n1379,
    n1389,
    n1321,
    n1399
  );


  nor
  g1407
  (
    n1461,
    n1435,
    n1427,
    n1329,
    n1431
  );


  and
  g1408
  (
    n1452,
    n1436,
    n1378,
    n1389,
    n1433
  );


  and
  g1409
  (
    n1476,
    n1381,
    n1431,
    n1325,
    n1388
  );


  xnor
  g1410
  (
    n1456,
    n1318,
    n1434,
    n1382,
    n1329
  );


  nor
  g1411
  (
    n1450,
    n1401,
    n1332,
    n1382,
    n1387
  );


  nand
  g1412
  (
    n1444,
    n1390,
    n1386,
    n1431,
    n1327
  );


  nor
  g1413
  (
    n1465,
    n1317,
    n1326,
    n1385,
    n1321
  );


  nand
  g1414
  (
    n1448,
    n1433,
    n1398,
    n1377,
    n1383
  );


  and
  g1415
  (
    n1453,
    n1434,
    n1430,
    n1323,
    n1386
  );


  and
  g1416
  (
    n1470,
    n1384,
    n1388,
    n1387,
    n1381
  );


  or
  g1417
  (
    n1441,
    n1324,
    n1319,
    n1318,
    n1331
  );


  and
  g1418
  (
    n1463,
    n1437,
    n1427,
    n1428,
    n1323
  );


  or
  g1419
  (
    n1462,
    n1327,
    n1379,
    n1329,
    n1428
  );


  xor
  g1420
  (
    n1478,
    n1432,
    n1391,
    n1325,
    n1427
  );


  or
  g1421
  (
    n1471,
    n1320,
    n1428,
    n1387,
    n1324
  );


  or
  g1422
  (
    n1455,
    n1391,
    n1400,
    n1434,
    n1331
  );


  xor
  g1423
  (
    n1445,
    n1379,
    n1437,
    n1385,
    n1319
  );


  nand
  g1424
  (
    n1472,
    n1432,
    n1384,
    n1399,
    n1386
  );


  nand
  g1425
  (
    n1443,
    n1320,
    n1330,
    n1325,
    n1326
  );


  xnor
  g1426
  (
    n1440,
    n1328,
    n1434,
    n1321,
    n1317
  );


  nor
  g1427
  (
    n1439,
    n1388,
    n1429,
    n1330
  );


  nand
  g1428
  (
    n1457,
    n1331,
    n1326,
    n1432,
    n1319
  );


  nor
  g1429
  (
    n1449,
    n1430,
    n1383,
    n1323,
    n1321
  );


  xnor
  g1430
  (
    n1477,
    n1377,
    n1320,
    n1386,
    n1322
  );


  xnor
  g1431
  (
    n1469,
    n1400,
    n1389,
    n1430,
    n1380
  );


  nand
  g1432
  (
    n1468,
    n1390,
    n1437,
    n1436,
    n1378
  );


  nor
  g1433
  (
    n1480,
    n1322,
    n1385,
    n1376,
    n1433
  );


  nor
  g1434
  (
    n1474,
    n1330,
    n1322,
    n1325,
    n1327
  );


  xnor
  g1435
  (
    n1473,
    n1427,
    n1377,
    n1379,
    n1385
  );


  and
  g1436
  (
    n1466,
    n1383,
    n1388,
    n1400,
    n1435
  );


  or
  g1437
  (
    n1460,
    n1430,
    n1328,
    n1378
  );


  xor
  g1438
  (
    n1442,
    n1428,
    n1431,
    n1389,
    n1429
  );


  or
  g1439
  (
    n1451,
    n1436,
    n1384,
    n1327,
    n1399
  );


  nor
  g1440
  (
    n1475,
    n1380,
    n1381,
    n1376
  );


  xor
  g1441
  (
    n1454,
    n1323,
    n1390,
    n1380,
    n1382
  );


  nor
  g1442
  (
    n1467,
    n1319,
    n1429,
    n1435,
    n1376
  );


  or
  g1443
  (
    n1459,
    n1384,
    n1437,
    n1383,
    n1324
  );


  nand
  g1444
  (
    n1446,
    n1400,
    n1390,
    n1318,
    n1387
  );


  or
  g1445
  (
    KeyWire_0_10,
    n1391,
    n1433,
    n1382,
    n1328
  );


  or
  g1446
  (
    n1464,
    n1380,
    n1399,
    n1377,
    n1432
  );


  xnor
  g1447
  (
    n1447,
    n1329,
    n1429,
    n1391,
    n1318
  );


  nor
  g1448
  (
    n1458,
    n1331,
    n1435,
    n1324,
    n1322
  );


  not
  g1449
  (
    n1486,
    n1452
  );


  not
  g1450
  (
    n1491,
    n1448
  );


  buf
  g1451
  (
    n1484,
    n1450
  );


  not
  g1452
  (
    n1485,
    n1439
  );


  not
  g1453
  (
    n1496,
    n1449
  );


  buf
  g1454
  (
    n1488,
    n1440
  );


  buf
  g1455
  (
    n1492,
    n1438
  );


  not
  g1456
  (
    n1483,
    n1446
  );


  not
  g1457
  (
    n1482,
    n1444
  );


  buf
  g1458
  (
    n1495,
    n1443
  );


  buf
  g1459
  (
    n1490,
    n1442
  );


  buf
  g1460
  (
    n1494,
    n1441
  );


  not
  g1461
  (
    n1493,
    n1453
  );


  not
  g1462
  (
    n1489,
    n1447
  );


  not
  g1463
  (
    n1487,
    n1451
  );


  not
  g1464
  (
    n1497,
    n1445
  );


  or
  g1465
  (
    n1502,
    n1415,
    n1455,
    n1411,
    n1488
  );


  nand
  g1466
  (
    n1511,
    n1401,
    n1416,
    n1403,
    n1404
  );


  xnor
  g1467
  (
    n1528,
    n1490,
    n1404,
    n1418
  );


  nor
  g1468
  (
    n1526,
    n1335,
    n1409,
    n1333,
    n1417
  );


  xor
  g1469
  (
    n1514,
    n1413,
    n1489,
    n1409,
    n1421
  );


  nor
  g1470
  (
    n1503,
    n1411,
    n1335,
    n1416,
    n1401
  );


  xnor
  g1471
  (
    n1504,
    n1410,
    n1408,
    n1418,
    n1484
  );


  and
  g1472
  (
    n1523,
    n1418,
    n1334,
    n1485,
    n1409
  );


  and
  g1473
  (
    n1529,
    n1413,
    n1411,
    n1409,
    n1484
  );


  or
  g1474
  (
    n1507,
    n1421,
    n1406,
    n1412,
    n1414
  );


  xnor
  g1475
  (
    n1516,
    n1485,
    n1402,
    n1334,
    n1457
  );


  nand
  g1476
  (
    n1499,
    n1414,
    n1410,
    n1419,
    n1408
  );


  and
  g1477
  (
    n1531,
    n1401,
    n1336,
    n1402,
    n1405
  );


  nand
  g1478
  (
    n1518,
    n1406,
    n1415,
    n1410,
    n1420
  );


  and
  g1479
  (
    n1519,
    n1484,
    n1417,
    n1415,
    n1413
  );


  nand
  g1480
  (
    n1525,
    n1454,
    n1485,
    n1417,
    n1414
  );


  xnor
  g1481
  (
    n1532,
    n1417,
    n1404,
    n1403,
    n1407
  );


  and
  g1482
  (
    n1501,
    n1407,
    n1490,
    n1333,
    n1484
  );


  nor
  g1483
  (
    n1505,
    n1482,
    n1405,
    n1488,
    n1489
  );


  xor
  g1484
  (
    n1521,
    n1487,
    n1482,
    n1411,
    n1332
  );


  or
  g1485
  (
    n1522,
    n1487,
    n1482,
    n1334,
    n1485
  );


  xor
  g1486
  (
    n1500,
    n1488,
    n1403,
    n1486,
    n1332
  );


  xnor
  g1487
  (
    n1513,
    n1489,
    n1419,
    n1416,
    n1487
  );


  and
  g1488
  (
    n1509,
    n1483,
    n1420
  );


  or
  g1489
  (
    n1510,
    n1334,
    n1482,
    n1406,
    n1413
  );


  or
  g1490
  (
    n1506,
    n1490,
    n1408,
    n1488,
    n1483
  );


  xor
  g1491
  (
    n1530,
    n1419,
    n1412,
    n1422,
    n1487
  );


  and
  g1492
  (
    n1508,
    n1405,
    n1422,
    n1333
  );


  xor
  g1493
  (
    n1512,
    n1414,
    n1406,
    n1486,
    n1420
  );


  nand
  g1494
  (
    n1524,
    n1419,
    n1489,
    n1335,
    n1402
  );


  and
  g1495
  (
    n1520,
    n1486,
    n1405,
    n1402,
    n1416
  );


  xnor
  g1496
  (
    n1517,
    n1412,
    n1412,
    n1407,
    n1403
  );


  xnor
  g1497
  (
    n1515,
    n1421,
    n1418,
    n1332,
    n1486
  );


  or
  g1498
  (
    n1498,
    n1483,
    n1407,
    n1410,
    n1421
  );


  nand
  g1499
  (
    n1527,
    n1408,
    n1456,
    n1335,
    n1415
  );


  buf
  g1500
  (
    n1543,
    n1513
  );


  not
  g1501
  (
    n1549,
    n1516
  );


  buf
  g1502
  (
    n1546,
    n1504
  );


  buf
  g1503
  (
    n1534,
    n1521
  );


  not
  g1504
  (
    n1541,
    n1505
  );


  buf
  g1505
  (
    n1545,
    n1515
  );


  not
  g1506
  (
    n1560,
    n1509
  );


  buf
  g1507
  (
    n1544,
    n1510
  );


  not
  g1508
  (
    n1552,
    n1524
  );


  not
  g1509
  (
    n1559,
    n1498
  );


  not
  g1510
  (
    n1538,
    n1525
  );


  not
  g1511
  (
    n1556,
    n1517
  );


  not
  g1512
  (
    n1548,
    n1523
  );


  not
  g1513
  (
    n1539,
    n1512
  );


  not
  g1514
  (
    n1535,
    n1506
  );


  not
  g1515
  (
    n1542,
    n1520
  );


  buf
  g1516
  (
    n1540,
    n1522
  );


  not
  g1517
  (
    n1557,
    n1503
  );


  not
  g1518
  (
    n1537,
    n1499
  );


  buf
  g1519
  (
    n1554,
    n1508
  );


  not
  g1520
  (
    n1536,
    n1518
  );


  buf
  g1521
  (
    n1547,
    n1514
  );


  not
  g1522
  (
    n1553,
    n1511
  );


  not
  g1523
  (
    n1551,
    n1507
  );


  not
  g1524
  (
    n1533,
    n1519
  );


  not
  g1525
  (
    n1558,
    n1500
  );


  not
  g1526
  (
    n1550,
    n1502
  );


  not
  g1527
  (
    n1555,
    n1501
  );


  not
  g1528
  (
    n1587,
    n1534
  );


  buf
  g1529
  (
    n1593,
    n1471
  );


  buf
  g1530
  (
    n1632,
    n1475
  );


  not
  g1531
  (
    n1597,
    n1543
  );


  not
  g1532
  (
    n1608,
    n1492
  );


  buf
  g1533
  (
    n1581,
    n1538
  );


  not
  g1534
  (
    n1616,
    n1337
  );


  not
  g1535
  (
    n1621,
    n1467
  );


  not
  g1536
  (
    n1627,
    n1547
  );


  not
  g1537
  (
    n1561,
    n1550
  );


  buf
  g1538
  (
    n1572,
    n1546
  );


  buf
  g1539
  (
    n1623,
    n1472
  );


  not
  g1540
  (
    n1574,
    n1461
  );


  buf
  g1541
  (
    n1595,
    n1475
  );


  not
  g1542
  (
    n1626,
    n1538
  );


  buf
  g1543
  (
    n1609,
    n1471
  );


  buf
  g1544
  (
    n1594,
    n1474
  );


  buf
  g1545
  (
    n1604,
    n1546
  );


  not
  g1546
  (
    n1585,
    n1491
  );


  buf
  g1547
  (
    n1619,
    n1495
  );


  not
  g1548
  (
    n1598,
    n1544
  );


  buf
  g1549
  (
    n1592,
    n1475
  );


  buf
  g1550
  (
    n1566,
    n1468
  );


  not
  g1551
  (
    n1596,
    n1462
  );


  buf
  g1552
  (
    n1602,
    n1542
  );


  not
  g1553
  (
    n1607,
    n1536
  );


  buf
  g1554
  (
    n1611,
    n1541
  );


  buf
  g1555
  (
    n1575,
    n1544
  );


  buf
  g1556
  (
    n1631,
    n1544
  );


  buf
  g1557
  (
    n1606,
    n1493
  );


  not
  g1558
  (
    n1568,
    n1543
  );


  buf
  g1559
  (
    n1599,
    n1465
  );


  buf
  g1560
  (
    n1618,
    n1493
  );


  not
  g1561
  (
    n1586,
    n1495
  );


  not
  g1562
  (
    n1580,
    n1545
  );


  not
  g1563
  (
    n1565,
    n1534
  );


  not
  g1564
  (
    n1603,
    n1471
  );


  buf
  g1565
  (
    n1590,
    n1459
  );


  not
  g1566
  (
    n1630,
    n1535
  );


  not
  g1567
  (
    n1576,
    n1541
  );


  buf
  g1568
  (
    n1578,
    n1539
  );


  buf
  g1569
  (
    n1615,
    n1536
  );


  buf
  g1570
  (
    n1589,
    n1550
  );


  not
  g1571
  (
    n1567,
    n1473
  );


  buf
  g1572
  (
    n1613,
    n1464
  );


  buf
  g1573
  (
    n1563,
    n1545
  );


  buf
  g1574
  (
    n1617,
    n1161
  );


  not
  g1575
  (
    n1583,
    n1470
  );


  nand
  g1576
  (
    n1569,
    n1469,
    n1472
  );


  or
  g1577
  (
    n1573,
    n1494,
    n1460
  );


  or
  g1578
  (
    n1610,
    n1472,
    n1540,
    n1539,
    n1474
  );


  nand
  g1579
  (
    n1564,
    n1492,
    n1156,
    n1160,
    n1336
  );


  and
  g1580
  (
    n1625,
    n1548,
    n1538,
    n1533,
    n1549
  );


  or
  g1581
  (
    n1612,
    n1550,
    n1548,
    n1541,
    n1492
  );


  or
  g1582
  (
    n1628,
    n1472,
    n1458,
    n1473,
    n1542
  );


  and
  g1583
  (
    n1571,
    n1537,
    n1491,
    n1549
  );


  nand
  g1584
  (
    n1562,
    n1159,
    n1158,
    n1539,
    n1543
  );


  nand
  g1585
  (
    n1570,
    n1539,
    n1537,
    n1336
  );


  xnor
  g1586
  (
    n1629,
    n1540,
    n1536,
    n1545,
    n1544
  );


  xor
  g1587
  (
    n1588,
    n1474,
    n1547,
    n1491,
    n1538
  );


  xnor
  g1588
  (
    n1579,
    n1546,
    n1545,
    n1493,
    n1535
  );


  nand
  g1589
  (
    n1584,
    n1549,
    n1548,
    n1543,
    n1534
  );


  or
  g1590
  (
    n1605,
    n1533,
    n1337,
    n1495,
    n1537
  );


  and
  g1591
  (
    n1582,
    n1541,
    n1490,
    n1542,
    n1547
  );


  and
  g1592
  (
    n1614,
    n1493,
    n1534,
    n1494
  );


  or
  g1593
  (
    n1622,
    n1536,
    n1535,
    n1540,
    n1473
  );


  nor
  g1594
  (
    n1591,
    n1336,
    n1337,
    n1474,
    n1495
  );


  nor
  g1595
  (
    n1624,
    n1548,
    n1533,
    n1337,
    n1547
  );


  xor
  g1596
  (
    n1620,
    n1533,
    n1494,
    n1471,
    n1546
  );


  or
  g1597
  (
    n1577,
    n1492,
    n1542,
    n1473,
    n1491
  );


  and
  g1598
  (
    n1601,
    n1475,
    n1535,
    n1550,
    n1466
  );


  and
  g1599
  (
    n1600,
    n1157,
    n1463,
    n1540,
    n1496
  );


  buf
  g1600
  (
    n1834,
    n1612
  );


  not
  g1601
  (
    n1794,
    n1566
  );


  not
  g1602
  (
    n1769,
    n1568
  );


  buf
  g1603
  (
    n1793,
    n1582
  );


  buf
  g1604
  (
    n1705,
    n1618
  );


  buf
  g1605
  (
    n1844,
    n1555
  );


  not
  g1606
  (
    n1784,
    n1593
  );


  not
  g1607
  (
    n1648,
    n1621
  );


  buf
  g1608
  (
    n1791,
    n1559
  );


  not
  g1609
  (
    n1811,
    n1619
  );


  not
  g1610
  (
    n1847,
    n1567
  );


  not
  g1611
  (
    n1782,
    n1594
  );


  not
  g1612
  (
    n1816,
    n1616
  );


  buf
  g1613
  (
    n1693,
    n1341
  );


  buf
  g1614
  (
    n1674,
    n1555
  );


  not
  g1615
  (
    n1854,
    n1561
  );


  buf
  g1616
  (
    n1742,
    n1579
  );


  not
  g1617
  (
    n1747,
    n1573
  );


  not
  g1618
  (
    n1745,
    n1594
  );


  not
  g1619
  (
    n1827,
    n1602
  );


  buf
  g1620
  (
    n1634,
    n1614
  );


  not
  g1621
  (
    n1649,
    n669
  );


  not
  g1622
  (
    n1800,
    n1586
  );


  buf
  g1623
  (
    n1741,
    n1560
  );


  not
  g1624
  (
    n1727,
    n1592
  );


  not
  g1625
  (
    n1746,
    n1572
  );


  not
  g1626
  (
    n1732,
    n1559
  );


  buf
  g1627
  (
    n1828,
    n1603
  );


  not
  g1628
  (
    n1724,
    n1611
  );


  buf
  g1629
  (
    n1787,
    n1570
  );


  not
  g1630
  (
    n1721,
    n1630
  );


  buf
  g1631
  (
    n1848,
    n671
  );


  not
  g1632
  (
    n1846,
    n1551
  );


  buf
  g1633
  (
    n1754,
    n1589
  );


  not
  g1634
  (
    n1717,
    n1592
  );


  buf
  g1635
  (
    n1734,
    n1561
  );


  not
  g1636
  (
    n1678,
    n1206
  );


  buf
  g1637
  (
    n1756,
    n1584
  );


  not
  g1638
  (
    n1819,
    n1621
  );


  not
  g1639
  (
    n1656,
    n1608
  );


  not
  g1640
  (
    n1707,
    n1565
  );


  not
  g1641
  (
    n1663,
    n1558
  );


  not
  g1642
  (
    n1807,
    n1608
  );


  not
  g1643
  (
    n1825,
    n1606
  );


  buf
  g1644
  (
    n1633,
    n1628
  );


  not
  g1645
  (
    n1808,
    n1552
  );


  buf
  g1646
  (
    n1760,
    n1604
  );


  buf
  g1647
  (
    n1651,
    n1624
  );


  not
  g1648
  (
    n1829,
    n1610
  );


  buf
  g1649
  (
    n1691,
    n1588
  );


  not
  g1650
  (
    n1711,
    n1615
  );


  buf
  g1651
  (
    n1713,
    n1581
  );


  not
  g1652
  (
    n1655,
    n1628
  );


  buf
  g1653
  (
    n1753,
    n1584
  );


  buf
  g1654
  (
    n1752,
    n1164
  );


  buf
  g1655
  (
    n1809,
    n672
  );


  not
  g1656
  (
    n1720,
    n1339
  );


  buf
  g1657
  (
    n1641,
    n1626
  );


  buf
  g1658
  (
    n1698,
    n1589
  );


  not
  g1659
  (
    n1695,
    n1632
  );


  buf
  g1660
  (
    n1817,
    n1601
  );


  buf
  g1661
  (
    n1673,
    n1601
  );


  not
  g1662
  (
    n1687,
    n1617
  );


  buf
  g1663
  (
    n1843,
    n1586
  );


  not
  g1664
  (
    n1798,
    n1602
  );


  buf
  g1665
  (
    n1683,
    n1585
  );


  buf
  g1666
  (
    n1778,
    n1480
  );


  not
  g1667
  (
    n1661,
    n1165
  );


  not
  g1668
  (
    n1676,
    n1625
  );


  buf
  g1669
  (
    n1670,
    n1340
  );


  not
  g1670
  (
    n1708,
    n1558
  );


  not
  g1671
  (
    n1726,
    n1616
  );


  buf
  g1672
  (
    n1772,
    n1593
  );


  buf
  g1673
  (
    n1743,
    n1605
  );


  not
  g1674
  (
    n1758,
    n1571
  );


  not
  g1675
  (
    n1709,
    n1566
  );


  not
  g1676
  (
    n1737,
    n1599
  );


  buf
  g1677
  (
    n1842,
    n1426
  );


  buf
  g1678
  (
    n1728,
    n1630
  );


  not
  g1679
  (
    n1637,
    n1581
  );


  not
  g1680
  (
    n1749,
    n1559
  );


  buf
  g1681
  (
    n1820,
    n1340
  );


  buf
  g1682
  (
    n1660,
    n1163
  );


  buf
  g1683
  (
    n1821,
    n1607
  );


  buf
  g1684
  (
    n1738,
    n1598
  );


  not
  g1685
  (
    n1748,
    n1480
  );


  buf
  g1686
  (
    n1849,
    n672
  );


  not
  g1687
  (
    n1804,
    n1617
  );


  not
  g1688
  (
    n1740,
    n1593
  );


  not
  g1689
  (
    n1723,
    n1569
  );


  buf
  g1690
  (
    n1658,
    n1477
  );


  not
  g1691
  (
    n1725,
    n1628
  );


  buf
  g1692
  (
    n1715,
    n1597
  );


  not
  g1693
  (
    n1764,
    n1621
  );


  buf
  g1694
  (
    n1735,
    n1560
  );


  not
  g1695
  (
    n1642,
    n1574
  );


  not
  g1696
  (
    n1763,
    n1562
  );


  not
  g1697
  (
    n1675,
    n1588
  );


  buf
  g1698
  (
    n1806,
    n1631
  );


  buf
  g1699
  (
    n1671,
    n1587
  );


  not
  g1700
  (
    n1704,
    n1612
  );


  buf
  g1701
  (
    n1694,
    n1574
  );


  not
  g1702
  (
    n1759,
    n1622
  );


  not
  g1703
  (
    n1803,
    n1570
  );


  buf
  g1704
  (
    n1799,
    n1162
  );


  not
  g1705
  (
    n1666,
    n1579
  );


  not
  g1706
  (
    n1700,
    n1584
  );


  buf
  g1707
  (
    n1852,
    n1627
  );


  buf
  g1708
  (
    n1767,
    n1424
  );


  buf
  g1709
  (
    n1639,
    n1423
  );


  not
  g1710
  (
    n1668,
    n1596
  );


  buf
  g1711
  (
    n1647,
    n1592
  );


  not
  g1712
  (
    n1680,
    n1611
  );


  buf
  g1713
  (
    n1783,
    n1578
  );


  not
  g1714
  (
    n1839,
    n1572
  );


  buf
  g1715
  (
    n1835,
    n1605
  );


  not
  g1716
  (
    n1719,
    n1565
  );


  not
  g1717
  (
    n1654,
    n1478
  );


  buf
  g1718
  (
    n1822,
    n1166
  );


  not
  g1719
  (
    n1712,
    n1629
  );


  buf
  g1720
  (
    n1686,
    n1166
  );


  buf
  g1721
  (
    n1810,
    n1607
  );


  not
  g1722
  (
    n1797,
    n1527
  );


  buf
  g1723
  (
    n1688,
    n1600
  );


  not
  g1724
  (
    n1792,
    n1426
  );


  not
  g1725
  (
    n1702,
    n1562
  );


  buf
  g1726
  (
    n1770,
    n1579
  );


  buf
  g1727
  (
    n1774,
    n1529
  );


  not
  g1728
  (
    n1850,
    n940
  );


  not
  g1729
  (
    n1714,
    n1629
  );


  buf
  g1730
  (
    n1853,
    n1586
  );


  not
  g1731
  (
    n1801,
    n1425
  );


  not
  g1732
  (
    n1729,
    n1551
  );


  not
  g1733
  (
    n1766,
    n1596
  );


  buf
  g1734
  (
    n1833,
    n1632
  );


  buf
  g1735
  (
    n1730,
    n1599
  );


  not
  g1736
  (
    n1744,
    n1605
  );


  not
  g1737
  (
    n1771,
    n671
  );


  buf
  g1738
  (
    n1699,
    n1564
  );


  buf
  g1739
  (
    n1796,
    n1476
  );


  not
  g1740
  (
    n1635,
    n1574
  );


  not
  g1741
  (
    n1838,
    n1558
  );


  buf
  g1742
  (
    n1775,
    n1594
  );


  not
  g1743
  (
    n1837,
    n1581
  );


  buf
  g1744
  (
    n1731,
    n1583
  );


  buf
  g1745
  (
    n1773,
    n1424
  );


  buf
  g1746
  (
    n1710,
    n1338
  );


  not
  g1747
  (
    n1795,
    n1585
  );


  buf
  g1748
  (
    n1823,
    n1562
  );


  buf
  g1749
  (
    n1768,
    n1481
  );


  and
  g1750
  (
    n1640,
    n1624,
    n1577,
    n1553
  );


  and
  g1751
  (
    n1813,
    n1166,
    n1598,
    n1614,
    n1339
  );


  xor
  g1752
  (
    n1659,
    n1599,
    n1565,
    n1617,
    n1556
  );


  or
  g1753
  (
    n1677,
    n1557,
    n1592,
    n1496,
    n1607
  );


  nor
  g1754
  (
    n1664,
    n1425,
    n1563,
    n1480,
    n1554
  );


  xnor
  g1755
  (
    n1669,
    n1557,
    n1426,
    n1621,
    n1423
  );


  xor
  g1756
  (
    n1785,
    n1163,
    n1567,
    n1424,
    n1582
  );


  xnor
  g1757
  (
    n1718,
    n1164,
    n1479,
    n1531,
    n1555
  );


  nor
  g1758
  (
    n1644,
    n1590,
    n1580,
    n1604,
    n1340
  );


  xor
  g1759
  (
    n1780,
    n1165,
    n1341,
    n1563,
    n1616
  );


  nor
  g1760
  (
    n1781,
    n1574,
    n1569,
    n1564,
    n1619
  );


  or
  g1761
  (
    n1814,
    n1625,
    n1589,
    n1594,
    n1617
  );


  nand
  g1762
  (
    n1751,
    n1573,
    n1573,
    n1600,
    n1165
  );


  or
  g1763
  (
    n1831,
    n1570,
    n1426,
    n1622,
    n1587
  );


  nor
  g1764
  (
    n1681,
    n1532,
    n1568,
    n1497,
    n1612
  );


  xnor
  g1765
  (
    n1696,
    n1563,
    n1578,
    n1613,
    n1163
  );


  xor
  g1766
  (
    n1697,
    n1570,
    n1568,
    n1575,
    n1609
  );


  xnor
  g1767
  (
    n1812,
    n1476,
    n1338,
    n1623,
    n1552
  );


  or
  g1768
  (
    n1650,
    n1575,
    n1590,
    n1583,
    n1609
  );


  xnor
  g1769
  (
    n1706,
    n1576,
    n1618,
    n1554,
    n1591
  );


  nand
  g1770
  (
    n1845,
    n1595,
    n1575,
    n1615,
    n1497
  );


  and
  g1771
  (
    n1638,
    n1632,
    n1207,
    n1477,
    n1580
  );


  xnor
  g1772
  (
    n1762,
    n1496,
    n1627,
    n670,
    n1618
  );


  and
  g1773
  (
    n1750,
    n1564,
    n1580,
    n1551,
    n1582
  );


  and
  g1774
  (
    n1739,
    n1620,
    n1627,
    n1586,
    n1619
  );


  nand
  g1775
  (
    n1851,
    n1611,
    n1476,
    n1571,
    n1596
  );


  or
  g1776
  (
    n1777,
    n936,
    n670,
    n1163,
    n1554
  );


  and
  g1777
  (
    n1805,
    n1620,
    n1571,
    n1607,
    n1557
  );


  or
  g1778
  (
    n1645,
    n1591,
    n1563,
    n670,
    n1425
  );


  nand
  g1779
  (
    n1662,
    n1619,
    n1591,
    n1479,
    n1578
  );


  and
  g1780
  (
    n1682,
    n1583,
    n1557,
    n1208,
    n1553
  );


  or
  g1781
  (
    n1643,
    n1578,
    n1631,
    n1479,
    n1590
  );


  nor
  g1782
  (
    n1840,
    n1165,
    n1559,
    n1604,
    n1576
  );


  xor
  g1783
  (
    n1786,
    n1587,
    n1338,
    n1606,
    n1610
  );


  and
  g1784
  (
    n1646,
    n1589,
    n1597,
    n1422,
    n1581
  );


  xor
  g1785
  (
    n1689,
    n1614,
    n1613,
    n1477,
    n1424
  );


  and
  g1786
  (
    n1701,
    n1590,
    n1596,
    n1624,
    n1601
  );


  nand
  g1787
  (
    n1672,
    n1600,
    n1553,
    n1588,
    n1625
  );


  or
  g1788
  (
    n1755,
    n1591,
    n1579,
    n1477,
    n1595
  );


  xnor
  g1789
  (
    n1733,
    n670,
    n1497,
    n1599,
    n1587
  );


  or
  g1790
  (
    n1790,
    n1609,
    n1624,
    n1585,
    n1628
  );


  xor
  g1791
  (
    n1761,
    n1561,
    n1609,
    n669,
    n1564
  );


  or
  g1792
  (
    n1665,
    n939,
    n1340,
    n1630,
    n1569
  );


  xnor
  g1793
  (
    n1636,
    n1608,
    n1476,
    n1598,
    n1595
  );


  and
  g1794
  (
    n1779,
    n1580,
    n1595,
    n1603,
    n1481
  );


  and
  g1795
  (
    n1832,
    n1603,
    n1571,
    n1584,
    n1588
  );


  xnor
  g1796
  (
    n1685,
    n935,
    n1602,
    n1629,
    n1577
  );


  and
  g1797
  (
    n1855,
    n1569,
    n1585,
    n938,
    n1603
  );


  nand
  g1798
  (
    n1788,
    n671,
    n1478,
    n1597,
    n1630
  );


  xnor
  g1799
  (
    n1824,
    n1341,
    n1602,
    n1601,
    n1572
  );


  or
  g1800
  (
    n1841,
    n1629,
    n1164,
    n1606,
    n1338
  );


  nor
  g1801
  (
    n1692,
    n1593,
    n669,
    n1558,
    n1423
  );


  xnor
  g1802
  (
    n1703,
    n1481,
    n1166,
    n1339,
    n1613
  );


  xnor
  g1803
  (
    n1765,
    n1613,
    n1598,
    n1605,
    n1576
  );


  xnor
  g1804
  (
    n1836,
    n1610,
    n1626,
    n1631
  );


  or
  g1805
  (
    n1818,
    n1615,
    n1425,
    n1556,
    n1528
  );


  or
  g1806
  (
    n1716,
    n1339,
    n1422,
    n1572,
    n1555
  );


  xnor
  g1807
  (
    n1667,
    n1618,
    n1608,
    n1556,
    n1497
  );


  and
  g1808
  (
    n1802,
    n1205,
    n1164,
    n1620,
    n1631
  );


  and
  g1809
  (
    n1789,
    n1341,
    n1610,
    n1552,
    n1480
  );


  nor
  g1810
  (
    n1815,
    n1479,
    n1623,
    n671,
    n669
  );


  xor
  g1811
  (
    n1757,
    n1582,
    n1560,
    n1562,
    n1632
  );


  nor
  g1812
  (
    n1830,
    n1627,
    n1481,
    n1614,
    n1478
  );


  and
  g1813
  (
    n1657,
    n1600,
    n1626,
    n1576,
    n1622
  );


  nor
  g1814
  (
    n1679,
    n1611,
    n1423,
    n1573,
    n1597
  );


  or
  g1815
  (
    n1722,
    n1577,
    n1526,
    n1623,
    n1530
  );


  and
  g1816
  (
    n1690,
    n1551,
    n1583,
    n1561,
    n1625
  );


  xnor
  g1817
  (
    n1684,
    n1554,
    n1567,
    n1568,
    n1604
  );


  nor
  g1818
  (
    n1826,
    n1556,
    n1622,
    n1567,
    n1566
  );


  nor
  g1819
  (
    n1776,
    n1612,
    n1552,
    n1566,
    n1553
  );


  nand
  g1820
  (
    n1736,
    n672,
    n1616,
    n1606,
    n1496
  );


  xnor
  g1821
  (
    n1653,
    n1623,
    n937,
    n1620,
    n1615
  );


  xor
  g1822
  (
    n1652,
    n1478,
    n1575,
    n1560,
    n1565
  );


  nor
  g1823
  (
    n1937,
    n1785,
    n1659,
    n1791,
    n1798
  );


  xnor
  g1824
  (
    n1857,
    n1769,
    n1749,
    n1846,
    n1817
  );


  nand
  g1825
  (
    n1875,
    n1817,
    n1800,
    n1734,
    n1827
  );


  or
  g1826
  (
    n1960,
    n1683,
    n1823,
    n1810,
    n1674
  );


  nand
  g1827
  (
    n1963,
    n1818,
    n1850,
    n1783,
    n1777
  );


  nand
  g1828
  (
    n1982,
    n1773,
    n1708,
    n1770,
    n1836
  );


  and
  g1829
  (
    n1914,
    n1715,
    n1778,
    n1795,
    n1757
  );


  xnor
  g1830
  (
    n1978,
    n1836,
    n1820,
    n1822,
    n1748
  );


  xnor
  g1831
  (
    n1905,
    n1707,
    n1824,
    n1852,
    n1780
  );


  xnor
  g1832
  (
    n1896,
    n1808,
    n1712,
    n1737,
    n1849
  );


  nand
  g1833
  (
    n1923,
    n1825,
    n1742,
    n1759,
    n1807
  );


  xor
  g1834
  (
    n1931,
    n1749,
    n1790,
    n1838,
    n1762
  );


  nand
  g1835
  (
    n1908,
    n1842,
    n1810,
    n1831,
    n1837
  );


  or
  g1836
  (
    n1885,
    n1797,
    n1832,
    n1660,
    n1779
  );


  nor
  g1837
  (
    n1911,
    n1850,
    n1847,
    n1830,
    n1826
  );


  xnor
  g1838
  (
    n1915,
    n1817,
    n1842,
    n1652,
    n1725
  );


  nor
  g1839
  (
    n1866,
    n1804,
    n1665,
    n1774,
    n1756
  );


  nor
  g1840
  (
    n1930,
    n1781,
    n1648,
    n1798,
    n1760
  );


  xnor
  g1841
  (
    n1864,
    n1687,
    n1801,
    n1851,
    n1793
  );


  nor
  g1842
  (
    n1925,
    n1785,
    n1761,
    n1830,
    n1788
  );


  or
  g1843
  (
    n1918,
    n1816,
    n1705,
    n1719,
    n1855
  );


  and
  g1844
  (
    n1901,
    n1826,
    n1664,
    n1776,
    n1787
  );


  xor
  g1845
  (
    n1883,
    n1819,
    n1783,
    n1851,
    n1784
  );


  xor
  g1846
  (
    n1909,
    n1853,
    n1788,
    n1699,
    n1786
  );


  or
  g1847
  (
    KeyWire_0_4,
    n1841,
    n1789,
    n1851,
    n1744
  );


  xnor
  g1848
  (
    n1942,
    n1838,
    n1828,
    n1786,
    n1780
  );


  xnor
  g1849
  (
    n1859,
    n1807,
    n1662,
    n1789,
    n1803
  );


  nand
  g1850
  (
    n1916,
    n1783,
    n1827,
    n1677,
    n1705
  );


  nand
  g1851
  (
    n1939,
    n1824,
    n1852,
    n1771,
    n1818
  );


  xor
  g1852
  (
    n1959,
    n1757,
    n1761,
    n1710,
    n1810
  );


  and
  g1853
  (
    n1878,
    n1754,
    n1754,
    n1823,
    n1814
  );


  nand
  g1854
  (
    n1902,
    n1784,
    n1737,
    n1845,
    n1841
  );


  xor
  g1855
  (
    n1904,
    n1713,
    n1821,
    n1779,
    n1800
  );


  and
  g1856
  (
    n1961,
    n1736,
    n1739,
    n1786,
    n1721
  );


  nor
  g1857
  (
    n1858,
    n1673,
    n1649,
    n1813,
    n1812
  );


  nor
  g1858
  (
    n1899,
    n1773,
    n1684,
    n1730,
    n1780
  );


  xor
  g1859
  (
    n1867,
    n1690,
    n1822,
    n1728,
    n1782
  );


  nand
  g1860
  (
    n1919,
    n1806,
    n1845,
    n1679,
    n1810
  );


  and
  g1861
  (
    n1889,
    n1718,
    n1831,
    n1802,
    n1676
  );


  nand
  g1862
  (
    n1881,
    n1835,
    n1829,
    n1682,
    n1772
  );


  nor
  g1863
  (
    n1862,
    n1655,
    n1650,
    n1852,
    n1809
  );


  nor
  g1864
  (
    n1892,
    n1837,
    n1805,
    n1835,
    n1840
  );


  or
  g1865
  (
    n1922,
    n1828,
    n1815,
    n1692
  );


  xnor
  g1866
  (
    n1967,
    n1829,
    n1709,
    n1818,
    n1775
  );


  and
  g1867
  (
    n1893,
    n1803,
    n1846,
    n1755,
    n1784
  );


  nand
  g1868
  (
    n1983,
    n1747,
    n1724,
    n1833
  );


  nor
  g1869
  (
    n1980,
    n1731,
    n1832,
    n1654,
    n1822
  );


  nor
  g1870
  (
    n1962,
    n1796,
    n1732,
    n1731,
    n1704
  );


  or
  g1871
  (
    n1928,
    n1694,
    n1789,
    n1779,
    n1806
  );


  nor
  g1872
  (
    n1977,
    n1672,
    n1792,
    n1712,
    n1796
  );


  or
  g1873
  (
    n1964,
    n1762,
    n1831,
    n1855,
    n1790
  );


  and
  g1874
  (
    n1870,
    n1787,
    n1675,
    n1726,
    n1729
  );


  xnor
  g1875
  (
    n1953,
    n1847,
    n1719,
    n1803,
    n1741
  );


  xnor
  g1876
  (
    n1865,
    n1841,
    n1752,
    n1742,
    n1738
  );


  xor
  g1877
  (
    n1884,
    n1793,
    n1748,
    n1693,
    n1667
  );


  xnor
  g1878
  (
    n1907,
    n1834,
    n1839,
    n1668
  );


  nor
  g1879
  (
    n1880,
    n1835,
    n1815,
    n1799,
    n1670
  );


  xnor
  g1880
  (
    n1946,
    n1780,
    n1855,
    n1788,
    n1797
  );


  and
  g1881
  (
    n1932,
    n1720,
    n1822,
    n1782,
    n1763
  );


  nand
  g1882
  (
    n1948,
    n1722,
    n672,
    n1814,
    n1807
  );


  nand
  g1883
  (
    n1936,
    n1854,
    n1771,
    n1849,
    n1697
  );


  xor
  g1884
  (
    n1945,
    n1813,
    n1811,
    n1847,
    n1735
  );


  or
  g1885
  (
    n1888,
    n1707,
    n1824,
    n1821,
    n1784
  );


  or
  g1886
  (
    n1876,
    n1714,
    n1766,
    n1691,
    n1743
  );


  or
  g1887
  (
    n1934,
    n1702,
    n1853,
    n1729,
    n1799
  );


  xnor
  g1888
  (
    n1981,
    n1808,
    n1826,
    n1829,
    n1811
  );


  or
  g1889
  (
    n1951,
    n1750,
    n1767,
    n1755,
    n1723
  );


  nand
  g1890
  (
    n1920,
    n1788,
    n1850,
    n1710,
    n1686
  );


  or
  g1891
  (
    n1898,
    n1815,
    n1803,
    n1769,
    n1844
  );


  nor
  g1892
  (
    n1906,
    n1842,
    n1739,
    n1651,
    n1703
  );


  nand
  g1893
  (
    n1944,
    n1772,
    n1841,
    n1812,
    n1848
  );


  xnor
  g1894
  (
    n1974,
    n1658,
    n1838,
    n1805,
    n1745
  );


  or
  g1895
  (
    n1968,
    n1701,
    n1794,
    n1795,
    n1793
  );


  or
  g1896
  (
    n1900,
    n1801,
    n1730,
    n1716,
    n1802
  );


  and
  g1897
  (
    n1891,
    n1718,
    n1753,
    n1818,
    n1775
  );


  or
  g1898
  (
    n1860,
    n1843,
    n1816,
    n1758,
    n1751
  );


  nand
  g1899
  (
    n1926,
    n1740,
    n1819,
    n1760,
    n1720
  );


  xnor
  g1900
  (
    n1933,
    n1848,
    n1804,
    n1727,
    n1809
  );


  and
  g1901
  (
    n1938,
    n1825,
    n1827,
    n1799,
    n1661
  );


  and
  g1902
  (
    n1950,
    n1798,
    n1768,
    n1716,
    n1844
  );


  nand
  g1903
  (
    n1913,
    n1721,
    n1787,
    n1774,
    n1843
  );


  xnor
  g1904
  (
    n1975,
    n1656,
    n1826,
    n1767,
    n1795
  );


  nor
  g1905
  (
    n1887,
    n1725,
    n1843,
    n1806,
    n1756
  );


  nand
  g1906
  (
    n1869,
    n1819,
    n1820,
    n1698,
    n1778
  );


  or
  g1907
  (
    n1965,
    n1765,
    n1759,
    n1681,
    n1744
  );


  xnor
  g1908
  (
    n1856,
    n1800,
    n1834,
    n1835,
    n1746
  );


  xnor
  g1909
  (
    n1976,
    n1752,
    n1777,
    n1852,
    n1740
  );


  or
  g1910
  (
    n1903,
    n1847,
    n1838,
    n1798,
    n1781
  );


  xnor
  g1911
  (
    n1895,
    n1824,
    n1845,
    n1827,
    n1792
  );


  or
  g1912
  (
    n1873,
    n1823,
    n1669,
    n1854,
    n1829
  );


  xnor
  g1913
  (
    n1863,
    n1703,
    n1790,
    n1836,
    n1746
  );


  and
  g1914
  (
    n1958,
    n1816,
    n1840,
    n1854,
    n1741
  );


  xnor
  g1915
  (
    n1890,
    n1808,
    n1783,
    n1776,
    n1657
  );


  nand
  g1916
  (
    n1971,
    n1817,
    n1821,
    n1695
  );


  and
  g1917
  (
    n1868,
    n1723,
    n1671,
    n1764,
    n1728
  );


  nor
  g1918
  (
    n1955,
    n1846,
    n1732,
    n1850,
    n1830
  );


  xor
  g1919
  (
    n1877,
    n1706,
    n1825,
    n1805,
    n1804
  );


  and
  g1920
  (
    n1979,
    n1794,
    n1834,
    n1704,
    n1848
  );


  nor
  g1921
  (
    n1947,
    n1717,
    n1666,
    n1812,
    n1696
  );


  xor
  g1922
  (
    n1966,
    n1711,
    n1766,
    n1724,
    n1688
  );


  and
  g1923
  (
    n1897,
    n1796,
    n1751,
    n1753,
    n1781
  );


  nand
  g1924
  (
    n1874,
    n1765,
    n1782,
    n1853,
    n1792
  );


  and
  g1925
  (
    n1935,
    n1812,
    n1828,
    n1685,
    n1813
  );


  or
  g1926
  (
    n1910,
    n1809,
    n1787,
    n1792,
    n1848
  );


  or
  g1927
  (
    n1894,
    n1770,
    n1709,
    n1830,
    n1717
  );


  xor
  g1928
  (
    n1929,
    n1777,
    n1804,
    n1811,
    n1789
  );


  or
  g1929
  (
    n1957,
    n1785,
    n1796,
    n1708,
    n1700
  );


  xnor
  g1930
  (
    n1984,
    n1745,
    n1747,
    n1791,
    n1823
  );


  xor
  g1931
  (
    n1886,
    n1797,
    n1779,
    n1813,
    n1849
  );


  xnor
  g1932
  (
    n1924,
    n1734,
    n1736,
    n1786,
    n1842
  );


  nor
  g1933
  (
    n1940,
    n1778,
    n1722,
    n1794,
    n1833
  );


  nor
  g1934
  (
    n1969,
    n1689,
    n1836,
    n1840,
    n1839
  );


  xor
  g1935
  (
    n1927,
    n1678,
    n1844,
    n1849,
    n1743
  );


  nand
  g1936
  (
    n1941,
    n1844,
    n1811,
    n1807,
    n1733
  );


  or
  g1937
  (
    n1871,
    n1834,
    n1768,
    n1819,
    n1790
  );


  and
  g1938
  (
    n1861,
    n1843,
    n1750,
    n1820,
    n1833
  );


  nor
  g1939
  (
    n1912,
    n1663,
    n1738,
    n1714,
    n1764
  );


  nor
  g1940
  (
    n1970,
    n1801,
    n1735,
    n1797,
    n1799
  );


  nor
  g1941
  (
    n1985,
    n1832,
    n1837,
    n1733,
    n1706
  );


  xnor
  g1942
  (
    n1949,
    n1854,
    n1653,
    n1828,
    n1846
  );


  xnor
  g1943
  (
    n1879,
    n1777,
    n1713,
    n1781,
    n1839
  );


  nor
  g1944
  (
    n1872,
    n1809,
    n1851,
    n1727,
    n1831
  );


  or
  g1945
  (
    n1956,
    n1806,
    n1845,
    n1715,
    n1711
  );


  and
  g1946
  (
    n1973,
    n1795,
    n1853,
    n1802,
    n1832
  );


  nand
  g1947
  (
    n1921,
    n1808,
    n1782,
    n1814,
    n1794
  );


  or
  g1948
  (
    n1972,
    n1778,
    n1802,
    n1801,
    n1800
  );


  xor
  g1949
  (
    n1882,
    n1840,
    n1758,
    n1814,
    n1805
  );


  and
  g1950
  (
    n1954,
    n1785,
    n1816,
    n1680,
    n1820
  );


  nor
  g1951
  (
    n1943,
    n1763,
    n1825,
    n1793,
    n1855
  );


  nand
  g1952
  (
    n1952,
    n1837,
    n1791,
    n1726
  );


  xor
  g1953
  (
    n2013,
    n1896,
    n1912,
    n1931,
    n1902
  );


  or
  g1954
  (
    n2004,
    n1978,
    n1939,
    n1895,
    n1893
  );


  and
  g1955
  (
    n2007,
    n1944,
    n1905,
    n1900,
    n1907
  );


  nor
  g1956
  (
    n2015,
    n1954,
    n1929,
    n1947,
    n1867
  );


  nor
  g1957
  (
    n1998,
    n1903,
    n1878,
    n1924,
    n1964
  );


  or
  g1958
  (
    n1996,
    n1973,
    n1914,
    n1983,
    n1962
  );


  or
  g1959
  (
    n2012,
    n1937,
    n1943,
    n1934,
    n1857
  );


  xor
  g1960
  (
    n1988,
    n1864,
    n1955,
    n1891,
    n1872
  );


  or
  g1961
  (
    n2017,
    n1927,
    n1894,
    n1909,
    n1963
  );


  xor
  g1962
  (
    n2016,
    n1925,
    n1911,
    n1877,
    n1887
  );


  xnor
  g1963
  (
    n2011,
    n1948,
    n1960,
    n1921,
    n1976
  );


  xor
  g1964
  (
    n1994,
    n1908,
    n1886,
    n1979,
    n1951
  );


  xnor
  g1965
  (
    n2005,
    n1888,
    n1901,
    n1946,
    n1974
  );


  nand
  g1966
  (
    n1993,
    n1889,
    n1860,
    n1862,
    n1972
  );


  nand
  g1967
  (
    n1986,
    n1874,
    n1922,
    n1869,
    n1910
  );


  or
  g1968
  (
    n2000,
    n1950,
    n1885,
    n1861,
    n1923
  );


  xnor
  g1969
  (
    n2006,
    n1980,
    n1898,
    n1906,
    n1875
  );


  or
  g1970
  (
    n1991,
    n1913,
    n1904,
    n1949,
    n1940
  );


  nor
  g1971
  (
    n2008,
    n1965,
    n1871,
    n1881,
    n1932
  );


  xnor
  g1972
  (
    n1989,
    n1868,
    n1956,
    n1942,
    n1866
  );


  xnor
  g1973
  (
    n1992,
    n1953,
    n1897,
    n1941,
    n1967
  );


  nand
  g1974
  (
    n1995,
    n1938,
    n1982,
    n1945,
    n1933
  );


  or
  g1975
  (
    n2009,
    n1926,
    n1957,
    n1918,
    n1928
  );


  or
  g1976
  (
    n2002,
    n1879,
    n1920,
    n1961,
    n1890
  );


  nand
  g1977
  (
    n2014,
    n1970,
    n1892,
    n1884,
    n1975
  );


  nor
  g1978
  (
    n2010,
    n1880,
    n1856,
    n1968,
    n1916
  );


  nand
  g1979
  (
    n2001,
    n1876,
    n1873,
    n1959,
    n1883
  );


  nand
  g1980
  (
    n2003,
    n1935,
    n1958,
    n1882,
    n1870
  );


  and
  g1981
  (
    n1997,
    n1952,
    n1930,
    n1859,
    n1971
  );


  xor
  g1982
  (
    n1987,
    n1917,
    n1915,
    n1865,
    n1899
  );


  xor
  g1983
  (
    n1999,
    n1981,
    n1919,
    n1977,
    n1863
  );


  nand
  g1984
  (
    n1990,
    n1969,
    n1936,
    n1966,
    n1858
  );


  not
  g1985
  (
    n2020,
    n1988
  );


  not
  g1986
  (
    n2018,
    n1993
  );


  xnor
  g1987
  (
    n2021,
    n1985,
    n1986
  );


  xnor
  g1988
  (
    n2022,
    n1990,
    n1984
  );


  nor
  g1989
  (
    n2019,
    n1992,
    n1987,
    n1989,
    n1991
  );


  nor
  g1990
  (
    n2025,
    n2022,
    n1999,
    n2010,
    n1998
  );


  or
  g1991
  (
    n2026,
    n2001,
    n2017,
    n2011,
    n2003
  );


  xnor
  g1992
  (
    n2024,
    n2007,
    n2020,
    n2009,
    n2021
  );


  xnor
  g1993
  (
    n2027,
    n1996,
    n2004,
    n2022,
    n2019
  );


  nand
  g1994
  (
    n2029,
    n2016,
    n1997,
    n2014,
    n2006
  );


  xnor
  g1995
  (
    n2023,
    n2013,
    n2022,
    n2000,
    n2008
  );


  nand
  g1996
  (
    n2030,
    n2015,
    n2018,
    n2012,
    n1994
  );


  and
  g1997
  (
    n2028,
    n2022,
    n1995,
    n2005,
    n2002
  );


  nand
  g1998
  (
    n2032,
    n2026,
    n2023,
    n2027,
    n2030
  );


  xnor
  g1999
  (
    n2031,
    n2028,
    n2029,
    n2024,
    n2025
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n62,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n653,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n1024,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1183,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1917,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n168,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1221,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n967,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n393,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1021,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1481,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n146,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n744,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n869,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n759,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1071,
    KeyNOTWire_0_15
  );


endmodule

