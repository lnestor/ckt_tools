

module Stat_1120_14_8
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n1108,
  n1097,
  n1103,
  n1098,
  n1104,
  n1099,
  n1100,
  n1086,
  n1101,
  n1089,
  n1106,
  n1091,
  n1134,
  n1136,
  n1140,
  n1142,
  n1141,
  n1143,
  n1144,
  n1145,
  n1139,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n1108;
  output n1097;
  output n1103;
  output n1098;
  output n1104;
  output n1099;
  output n1100;
  output n1086;
  output n1101;
  output n1089;
  output n1106;
  output n1091;
  output n1134;
  output n1136;
  output n1140;
  output n1142;
  output n1141;
  output n1143;
  output n1144;
  output n1145;
  output n1139;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1087;
  wire n1088;
  wire n1090;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1102;
  wire n1105;
  wire n1107;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1135;
  wire n1137;
  wire n1138;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n28,
    n2
  );


  not
  g1
  (
    n27,
    n3
  );


  not
  g2
  (
    n34,
    n7
  );


  not
  g3
  (
    n33,
    n3
  );


  not
  g4
  (
    n30,
    n1
  );


  buf
  g5
  (
    n36,
    n8
  );


  not
  g6
  (
    n35,
    n2
  );


  buf
  g7
  (
    n32,
    n5
  );


  buf
  g8
  (
    n29,
    n6
  );


  not
  g9
  (
    n37,
    n2
  );


  not
  g10
  (
    n31,
    n4
  );


  or
  g11
  (
    n39,
    n6,
    n4,
    n7,
    n5
  );


  xor
  g12
  (
    n38,
    n3,
    n7,
    n6,
    n4
  );


  xnor
  g13
  (
    n26,
    n5,
    n8,
    n1
  );


  not
  g14
  (
    n43,
    n32
  );


  buf
  g15
  (
    n40,
    n27
  );


  not
  g16
  (
    n49,
    n28
  );


  buf
  g17
  (
    n51,
    n31
  );


  buf
  g18
  (
    n41,
    n34
  );


  buf
  g19
  (
    n52,
    n28
  );


  buf
  g20
  (
    n53,
    n37
  );


  buf
  g21
  (
    n57,
    n29
  );


  nand
  g22
  (
    n42,
    n26,
    n30
  );


  and
  g23
  (
    KeyWire_0_41,
    n33,
    n32,
    n29
  );


  and
  g24
  (
    n55,
    n36,
    n26,
    n27
  );


  and
  g25
  (
    n54,
    n34,
    n36,
    n30,
    n33
  );


  and
  g26
  (
    n44,
    n32,
    n28,
    n35,
    n31
  );


  or
  g27
  (
    n58,
    n28,
    n36,
    n35
  );


  nand
  g28
  (
    n48,
    n34,
    n27,
    n30,
    n35
  );


  nor
  g29
  (
    n46,
    n30,
    n35,
    n27,
    n31
  );


  or
  g30
  (
    n45,
    n33,
    n31,
    n26,
    n37
  );


  or
  g31
  (
    n50,
    n34,
    n29,
    n32,
    n33
  );


  nor
  g32
  (
    n56,
    n37,
    n38
  );


  or
  g33
  (
    n64,
    n42,
    n50,
    n55,
    n56
  );


  xnor
  g34
  (
    n62,
    n40,
    n53,
    n54,
    n49
  );


  nor
  g35
  (
    n61,
    n51,
    n50,
    n53,
    n41
  );


  or
  g36
  (
    n63,
    n43,
    n48,
    n54,
    n44
  );


  xor
  g37
  (
    n60,
    n47,
    n55,
    n51
  );


  xor
  g38
  (
    n59,
    n45,
    n52,
    n46
  );


  buf
  g39
  (
    n74,
    n59
  );


  not
  g40
  (
    n73,
    n38
  );


  not
  g41
  (
    n67,
    n38
  );


  buf
  g42
  (
    n70,
    n64
  );


  buf
  g43
  (
    n65,
    n9
  );


  not
  g44
  (
    n72,
    n9
  );


  buf
  g45
  (
    n71,
    n8
  );


  not
  g46
  (
    n68,
    n63
  );


  not
  g47
  (
    n66,
    n63
  );


  not
  g48
  (
    n79,
    n60
  );


  buf
  g49
  (
    n77,
    n62
  );


  buf
  g50
  (
    n69,
    n59
  );


  and
  g51
  (
    n75,
    n62,
    n64,
    n9,
    n63
  );


  nand
  g52
  (
    n76,
    n62,
    n61,
    n64,
    n9
  );


  nand
  g53
  (
    n78,
    n63,
    n60,
    n10,
    n59
  );


  or
  g54
  (
    n80,
    n60,
    n61,
    n64
  );


  not
  g55
  (
    n90,
    n70
  );


  buf
  g56
  (
    n100,
    n13
  );


  not
  g57
  (
    KeyWire_0_7,
    n73
  );


  not
  g58
  (
    KeyWire_0_53,
    n56
  );


  buf
  g59
  (
    n102,
    n13
  );


  buf
  g60
  (
    n91,
    n68
  );


  xor
  g61
  (
    n96,
    n14,
    n77
  );


  or
  g62
  (
    n95,
    n71,
    n78
  );


  nand
  g63
  (
    n83,
    n78,
    n77
  );


  nand
  g64
  (
    n110,
    n76,
    n11
  );


  nand
  g65
  (
    n101,
    n14,
    n11
  );


  xnor
  g66
  (
    n87,
    n75,
    n77
  );


  or
  g67
  (
    n93,
    n65,
    n74
  );


  and
  g68
  (
    n92,
    n80,
    n14
  );


  and
  g69
  (
    n107,
    n15,
    n72
  );


  xnor
  g70
  (
    n85,
    n79,
    n76
  );


  xor
  g71
  (
    n109,
    n12,
    n73
  );


  and
  g72
  (
    n111,
    n10,
    n66
  );


  and
  g73
  (
    n89,
    n15,
    n67
  );


  or
  g74
  (
    n97,
    n11,
    n12
  );


  buf
  g75
  (
    n104,
    n79
  );


  and
  g76
  (
    n112,
    n16,
    n80
  );


  nor
  g77
  (
    KeyWire_0_15,
    n13,
    n16
  );


  nand
  g78
  (
    n84,
    n69,
    n75
  );


  nor
  g79
  (
    n98,
    n15,
    n12
  );


  and
  g80
  (
    KeyWire_0_45,
    n75,
    n74
  );


  and
  g81
  (
    n106,
    n78,
    n73
  );


  xor
  g82
  (
    n105,
    n14,
    n13
  );


  or
  g83
  (
    n108,
    n12,
    n15
  );


  or
  g84
  (
    n94,
    n10,
    n74
  );


  or
  g85
  (
    n103,
    n10,
    n11
  );


  nand
  g86
  (
    n99,
    n80,
    n76
  );


  not
  g87
  (
    n117,
    n81
  );


  not
  g88
  (
    n205,
    n92
  );


  buf
  g89
  (
    n148,
    n87
  );


  buf
  g90
  (
    n214,
    n106
  );


  buf
  g91
  (
    n139,
    n97
  );


  not
  g92
  (
    n136,
    n101
  );


  buf
  g93
  (
    n125,
    n101
  );


  not
  g94
  (
    n113,
    n93
  );


  not
  g95
  (
    n239,
    n88
  );


  buf
  g96
  (
    n198,
    n90
  );


  not
  g97
  (
    n114,
    n104
  );


  buf
  g98
  (
    n206,
    n98
  );


  buf
  g99
  (
    n119,
    n111
  );


  buf
  g100
  (
    n210,
    n112
  );


  not
  g101
  (
    n132,
    n102
  );


  buf
  g102
  (
    n202,
    n83
  );


  buf
  g103
  (
    n207,
    n93
  );


  not
  g104
  (
    n153,
    n82
  );


  not
  g105
  (
    n219,
    n102
  );


  not
  g106
  (
    n134,
    n88
  );


  buf
  g107
  (
    n116,
    n89
  );


  not
  g108
  (
    n222,
    n112
  );


  buf
  g109
  (
    n124,
    n107
  );


  not
  g110
  (
    n221,
    n103
  );


  buf
  g111
  (
    n179,
    n101
  );


  not
  g112
  (
    n181,
    n104
  );


  not
  g113
  (
    n204,
    n85
  );


  not
  g114
  (
    n176,
    n81
  );


  buf
  g115
  (
    n175,
    n103
  );


  not
  g116
  (
    n232,
    n106
  );


  buf
  g117
  (
    n201,
    n95
  );


  buf
  g118
  (
    n229,
    n89
  );


  buf
  g119
  (
    n190,
    n94
  );


  not
  g120
  (
    n140,
    n89
  );


  buf
  g121
  (
    n200,
    n111
  );


  not
  g122
  (
    n189,
    n110
  );


  buf
  g123
  (
    n171,
    n99
  );


  buf
  g124
  (
    n185,
    n89
  );


  not
  g125
  (
    n195,
    n97
  );


  buf
  g126
  (
    n180,
    n82
  );


  not
  g127
  (
    n162,
    n90
  );


  not
  g128
  (
    n143,
    n85
  );


  not
  g129
  (
    KeyWire_0_4,
    n86
  );


  not
  g130
  (
    n235,
    n100
  );


  buf
  g131
  (
    n147,
    n109
  );


  buf
  g132
  (
    n127,
    n108
  );


  buf
  g133
  (
    n126,
    n99
  );


  not
  g134
  (
    n160,
    n102
  );


  buf
  g135
  (
    n217,
    n106
  );


  buf
  g136
  (
    n178,
    n97
  );


  not
  g137
  (
    n224,
    n86
  );


  buf
  g138
  (
    n120,
    n97
  );


  buf
  g139
  (
    n118,
    n81
  );


  not
  g140
  (
    n166,
    n94
  );


  not
  g141
  (
    n233,
    n90
  );


  buf
  g142
  (
    n177,
    n110
  );


  not
  g143
  (
    n228,
    n96
  );


  buf
  g144
  (
    n142,
    n95
  );


  buf
  g145
  (
    n129,
    n84
  );


  buf
  g146
  (
    n169,
    n95
  );


  not
  g147
  (
    n155,
    n92
  );


  buf
  g148
  (
    n216,
    n83
  );


  not
  g149
  (
    n208,
    n87
  );


  not
  g150
  (
    n130,
    n81
  );


  buf
  g151
  (
    n141,
    n95
  );


  buf
  g152
  (
    n227,
    n107
  );


  not
  g153
  (
    n193,
    n84
  );


  not
  g154
  (
    n240,
    n108
  );


  not
  g155
  (
    n225,
    n92
  );


  not
  g156
  (
    n203,
    n93
  );


  not
  g157
  (
    n196,
    n99
  );


  buf
  g158
  (
    n123,
    n98
  );


  buf
  g159
  (
    n150,
    n82
  );


  buf
  g160
  (
    n213,
    n106
  );


  buf
  g161
  (
    n223,
    n87
  );


  not
  g162
  (
    n212,
    n105
  );


  not
  g163
  (
    n154,
    n98
  );


  not
  g164
  (
    n194,
    n109
  );


  not
  g165
  (
    n236,
    n105
  );


  buf
  g166
  (
    n135,
    n93
  );


  not
  g167
  (
    n220,
    n108
  );


  buf
  g168
  (
    n133,
    n107
  );


  not
  g169
  (
    n173,
    n96
  );


  buf
  g170
  (
    n174,
    n92
  );


  buf
  g171
  (
    KeyWire_0_30,
    n85
  );


  not
  g172
  (
    KeyWire_0_33,
    n100
  );


  not
  g173
  (
    n152,
    n111
  );


  not
  g174
  (
    KeyWire_0_29,
    n91
  );


  not
  g175
  (
    KeyWire_0_20,
    n82
  );


  buf
  g176
  (
    KeyWire_0_38,
    n100
  );


  not
  g177
  (
    n158,
    n112
  );


  buf
  g178
  (
    n151,
    n101
  );


  not
  g179
  (
    n167,
    n84
  );


  buf
  g180
  (
    n209,
    n98
  );


  buf
  g181
  (
    n161,
    n102
  );


  buf
  g182
  (
    n156,
    n85
  );


  buf
  g183
  (
    n168,
    n105
  );


  not
  g184
  (
    n226,
    n91
  );


  not
  g185
  (
    n192,
    n90
  );


  not
  g186
  (
    n163,
    n87
  );


  buf
  g187
  (
    n186,
    n91
  );


  not
  g188
  (
    n231,
    n86
  );


  buf
  g189
  (
    n211,
    n111
  );


  not
  g190
  (
    KeyWire_0_26,
    n100
  );


  buf
  g191
  (
    n182,
    n88
  );


  buf
  g192
  (
    n157,
    n103
  );


  not
  g193
  (
    n137,
    n96
  );


  not
  g194
  (
    n165,
    n96
  );


  not
  g195
  (
    n115,
    n83
  );


  buf
  g196
  (
    n146,
    n110
  );


  not
  g197
  (
    n183,
    n104
  );


  buf
  g198
  (
    n184,
    n112
  );


  not
  g199
  (
    n149,
    n84
  );


  buf
  g200
  (
    n121,
    n94
  );


  not
  g201
  (
    n170,
    n109
  );


  buf
  g202
  (
    n138,
    n91
  );


  buf
  g203
  (
    KeyWire_0_31,
    n103
  );


  buf
  g204
  (
    n197,
    n94
  );


  buf
  g205
  (
    n128,
    n86
  );


  buf
  g206
  (
    n187,
    n99
  );


  buf
  g207
  (
    n218,
    n110
  );


  buf
  g208
  (
    n144,
    n83
  );


  not
  g209
  (
    n131,
    n88
  );


  not
  g210
  (
    n172,
    n108
  );


  buf
  g211
  (
    n188,
    n109
  );


  buf
  g212
  (
    n199,
    n107
  );


  not
  g213
  (
    n145,
    n104
  );


  buf
  g214
  (
    n191,
    n105
  );


  not
  g215
  (
    n406,
    n116
  );


  buf
  g216
  (
    n452,
    n120
  );


  buf
  g217
  (
    n372,
    n220
  );


  not
  g218
  (
    n414,
    n236
  );


  buf
  g219
  (
    n428,
    n196
  );


  not
  g220
  (
    KeyWire_0_13,
    n127
  );


  not
  g221
  (
    n479,
    n173
  );


  not
  g222
  (
    n285,
    n189
  );


  not
  g223
  (
    n358,
    n228
  );


  buf
  g224
  (
    n312,
    n213
  );


  buf
  g225
  (
    n346,
    n184
  );


  not
  g226
  (
    n331,
    n214
  );


  buf
  g227
  (
    n337,
    n151
  );


  not
  g228
  (
    n326,
    n208
  );


  not
  g229
  (
    n419,
    n157
  );


  buf
  g230
  (
    n482,
    n154
  );


  buf
  g231
  (
    n332,
    n178
  );


  not
  g232
  (
    n304,
    n178
  );


  not
  g233
  (
    n311,
    n207
  );


  buf
  g234
  (
    n274,
    n224
  );


  buf
  g235
  (
    n437,
    n220
  );


  not
  g236
  (
    n261,
    n202
  );


  buf
  g237
  (
    n328,
    n228
  );


  buf
  g238
  (
    n383,
    n179
  );


  not
  g239
  (
    n499,
    n206
  );


  not
  g240
  (
    n457,
    n134
  );


  buf
  g241
  (
    n402,
    n176
  );


  not
  g242
  (
    n266,
    n227
  );


  buf
  g243
  (
    n315,
    n178
  );


  not
  g244
  (
    n434,
    n197
  );


  buf
  g245
  (
    n345,
    n157
  );


  buf
  g246
  (
    n470,
    n238
  );


  not
  g247
  (
    n291,
    n126
  );


  buf
  g248
  (
    n405,
    n181
  );


  not
  g249
  (
    n483,
    n144
  );


  buf
  g250
  (
    n333,
    n143
  );


  not
  g251
  (
    n458,
    n183
  );


  buf
  g252
  (
    n469,
    n125
  );


  not
  g253
  (
    n427,
    n163
  );


  buf
  g254
  (
    n282,
    n179
  );


  buf
  g255
  (
    n362,
    n159
  );


  not
  g256
  (
    n490,
    n155
  );


  buf
  g257
  (
    n276,
    n153
  );


  not
  g258
  (
    n454,
    n129
  );


  buf
  g259
  (
    n410,
    n117
  );


  buf
  g260
  (
    n342,
    n122
  );


  not
  g261
  (
    n415,
    n233
  );


  buf
  g262
  (
    n356,
    n132
  );


  not
  g263
  (
    n330,
    n174
  );


  not
  g264
  (
    n303,
    n195
  );


  buf
  g265
  (
    n322,
    n215
  );


  not
  g266
  (
    n382,
    n135
  );


  not
  g267
  (
    n387,
    n161
  );


  not
  g268
  (
    n253,
    n158
  );


  not
  g269
  (
    n249,
    n177
  );


  not
  g270
  (
    n471,
    n169
  );


  buf
  g271
  (
    n307,
    n227
  );


  not
  g272
  (
    n497,
    n161
  );


  not
  g273
  (
    KeyWire_0_16,
    n128
  );


  buf
  g274
  (
    n318,
    n212
  );


  not
  g275
  (
    n306,
    n133
  );


  buf
  g276
  (
    n302,
    n211
  );


  buf
  g277
  (
    n334,
    n149
  );


  buf
  g278
  (
    n280,
    n237
  );


  buf
  g279
  (
    n338,
    n193
  );


  buf
  g280
  (
    n461,
    n177
  );


  buf
  g281
  (
    n329,
    n149
  );


  not
  g282
  (
    n412,
    n199
  );


  buf
  g283
  (
    n289,
    n148
  );


  buf
  g284
  (
    n449,
    n223
  );


  buf
  g285
  (
    n409,
    n131
  );


  buf
  g286
  (
    n258,
    n184
  );


  buf
  g287
  (
    n354,
    n231
  );


  not
  g288
  (
    n250,
    n176
  );


  not
  g289
  (
    n324,
    n176
  );


  not
  g290
  (
    n456,
    n234
  );


  buf
  g291
  (
    n448,
    n130
  );


  not
  g292
  (
    n468,
    n118
  );


  buf
  g293
  (
    n502,
    n156
  );


  not
  g294
  (
    n259,
    n207
  );


  buf
  g295
  (
    n496,
    n178
  );


  not
  g296
  (
    n385,
    n129
  );


  buf
  g297
  (
    n264,
    n194
  );


  not
  g298
  (
    n283,
    n204
  );


  not
  g299
  (
    n263,
    n222
  );


  not
  g300
  (
    n341,
    n237
  );


  not
  g301
  (
    n284,
    n209
  );


  buf
  g302
  (
    n265,
    n132
  );


  not
  g303
  (
    n391,
    n234
  );


  buf
  g304
  (
    n316,
    n126
  );


  buf
  g305
  (
    KeyWire_0_57,
    n196
  );


  not
  g306
  (
    n435,
    n199
  );


  not
  g307
  (
    n487,
    n228
  );


  not
  g308
  (
    n492,
    n233
  );


  buf
  g309
  (
    n393,
    n201
  );


  not
  g310
  (
    n270,
    n200
  );


  not
  g311
  (
    n277,
    n159
  );


  buf
  g312
  (
    n422,
    n56
  );


  buf
  g313
  (
    n371,
    n215
  );


  buf
  g314
  (
    n272,
    n168
  );


  not
  g315
  (
    n464,
    n197
  );


  buf
  g316
  (
    n401,
    n136
  );


  buf
  g317
  (
    n426,
    n164
  );


  buf
  g318
  (
    n295,
    n239
  );


  not
  g319
  (
    n474,
    n161
  );


  not
  g320
  (
    n369,
    n196
  );


  buf
  g321
  (
    n467,
    n114
  );


  buf
  g322
  (
    KeyWire_0_63,
    n140
  );


  not
  g323
  (
    n488,
    n156
  );


  buf
  g324
  (
    n460,
    n122
  );


  not
  g325
  (
    n248,
    n159
  );


  not
  g326
  (
    n439,
    n115
  );


  not
  g327
  (
    n299,
    n218
  );


  not
  g328
  (
    n273,
    n170
  );


  not
  g329
  (
    n494,
    n164
  );


  buf
  g330
  (
    n376,
    n165
  );


  not
  g331
  (
    n363,
    n136
  );


  buf
  g332
  (
    n357,
    n172
  );


  buf
  g333
  (
    n486,
    n156
  );


  buf
  g334
  (
    n404,
    n236
  );


  not
  g335
  (
    n374,
    n216
  );


  not
  g336
  (
    n390,
    n212
  );


  not
  g337
  (
    n394,
    n149
  );


  buf
  g338
  (
    n375,
    n157
  );


  not
  g339
  (
    n498,
    n234
  );


  not
  g340
  (
    n466,
    n217
  );


  buf
  g341
  (
    n472,
    n132
  );


  not
  g342
  (
    n365,
    n167
  );


  buf
  g343
  (
    n313,
    n165
  );


  not
  g344
  (
    n429,
    n152
  );


  buf
  g345
  (
    n335,
    n174
  );


  not
  g346
  (
    n484,
    n145
  );


  not
  g347
  (
    n290,
    n166
  );


  not
  g348
  (
    n396,
    n153
  );


  buf
  g349
  (
    n244,
    n240
  );


  buf
  g350
  (
    n389,
    n150
  );


  not
  g351
  (
    n267,
    n113
  );


  buf
  g352
  (
    n325,
    n116
  );


  buf
  g353
  (
    n453,
    n123
  );


  buf
  g354
  (
    n241,
    n120
  );


  buf
  g355
  (
    n355,
    n181
  );


  not
  g356
  (
    n441,
    n163
  );


  not
  g357
  (
    n403,
    n128
  );


  buf
  g358
  (
    n443,
    n195
  );


  not
  g359
  (
    n243,
    n232
  );


  buf
  g360
  (
    n408,
    n240
  );


  buf
  g361
  (
    n268,
    n193
  );


  buf
  g362
  (
    n336,
    n224
  );


  not
  g363
  (
    n378,
    n138
  );


  buf
  g364
  (
    n432,
    n206
  );


  buf
  g365
  (
    n257,
    n122
  );


  buf
  g366
  (
    n278,
    n118
  );


  buf
  g367
  (
    n339,
    n186
  );


  buf
  g368
  (
    KeyWire_0_14,
    n177
  );


  not
  g369
  (
    n310,
    n172
  );


  buf
  g370
  (
    KeyWire_0_55,
    n188
  );


  buf
  g371
  (
    n301,
    n130
  );


  not
  g372
  (
    n397,
    n138
  );


  not
  g373
  (
    n424,
    n141
  );


  not
  g374
  (
    n478,
    n230
  );


  not
  g375
  (
    n379,
    n224
  );


  buf
  g376
  (
    KeyWire_0_3,
    n233
  );


  buf
  g377
  (
    KeyWire_0_46,
    n187
  );


  buf
  g378
  (
    n481,
    n114
  );


  buf
  g379
  (
    n451,
    n223
  );


  not
  g380
  (
    n377,
    n182
  );


  buf
  g381
  (
    n392,
    n123
  );


  buf
  g382
  (
    n317,
    n142
  );


  buf
  g383
  (
    n308,
    n230
  );


  not
  g384
  (
    n400,
    n135
  );


  not
  g385
  (
    n254,
    n129
  );


  buf
  g386
  (
    KeyWire_0_39,
    n162
  );


  not
  g387
  (
    n319,
    n222
  );


  not
  g388
  (
    n373,
    n224
  );


  not
  g389
  (
    n347,
    n191
  );


  buf
  g390
  (
    n288,
    n125
  );


  buf
  g391
  (
    n349,
    n239
  );


  buf
  g392
  (
    n294,
    n238
  );


  and
  g393
  (
    n361,
    n182,
    n127,
    n218
  );


  nor
  g394
  (
    n269,
    n194,
    n133,
    n236,
    n128
  );


  xnor
  g395
  (
    n298,
    n157,
    n193,
    n137,
    n139
  );


  and
  g396
  (
    n255,
    n232,
    n126,
    n217,
    n196
  );


  xnor
  g397
  (
    n446,
    n183,
    n148,
    n180,
    n121
  );


  nor
  g398
  (
    n380,
    n197,
    n225,
    n173,
    n162
  );


  xnor
  g399
  (
    n245,
    n201,
    n211,
    n210,
    n161
  );


  xor
  g400
  (
    n501,
    n189,
    n226,
    n152,
    n160
  );


  or
  g401
  (
    n242,
    n173,
    n205,
    n235,
    n127
  );


  xnor
  g402
  (
    n351,
    n229,
    n135,
    n190,
    n221
  );


  xor
  g403
  (
    n275,
    n165,
    n212,
    n185,
    n215
  );


  and
  g404
  (
    n251,
    n183,
    n206,
    n154,
    n150
  );


  xnor
  g405
  (
    n411,
    n131,
    n141,
    n119,
    n221
  );


  xor
  g406
  (
    n309,
    n166,
    n210,
    n174,
    n170
  );


  or
  g407
  (
    n416,
    n147,
    n147,
    n159,
    n152
  );


  xor
  g408
  (
    n366,
    n185,
    n203,
    n115,
    n163
  );


  and
  g409
  (
    n381,
    n235,
    n188,
    n184,
    n216
  );


  or
  g410
  (
    n413,
    n191,
    n232,
    n210,
    n144
  );


  nor
  g411
  (
    n386,
    n203,
    n167,
    n143,
    n151
  );


  and
  g412
  (
    n297,
    n134,
    n208,
    n204,
    n215
  );


  nor
  g413
  (
    n440,
    n237,
    n198,
    n131,
    n136
  );


  nand
  g414
  (
    n340,
    n194,
    n170,
    n190,
    n216
  );


  or
  g415
  (
    n477,
    n184,
    n119,
    n221,
    n118
  );


  or
  g416
  (
    n485,
    n164,
    n199,
    n183,
    n181
  );


  or
  g417
  (
    n450,
    n192,
    n238,
    n171,
    n239
  );


  xor
  g418
  (
    n463,
    n218,
    n162,
    n202,
    n131
  );


  xor
  g419
  (
    n252,
    n180,
    n129,
    n229,
    n182
  );


  or
  g420
  (
    n465,
    n137,
    n237,
    n192,
    n115
  );


  or
  g421
  (
    KeyWire_0_27,
    n190,
    n197,
    n121,
    n217
  );


  nand
  g422
  (
    n292,
    n122,
    n226,
    n181,
    n177
  );


  and
  g423
  (
    KeyWire_0_25,
    n195,
    n113,
    n185,
    n182
  );


  and
  g424
  (
    n370,
    n227,
    n154,
    n155,
    n124
  );


  nand
  g425
  (
    n430,
    n160,
    n155,
    n192,
    n240
  );


  or
  g426
  (
    n442,
    n146,
    n142,
    n164,
    n219
  );


  or
  g427
  (
    n279,
    n175,
    n175,
    n231,
    n128
  );


  or
  g428
  (
    n271,
    n198,
    n230,
    n186,
    n225
  );


  nand
  g429
  (
    n438,
    n141,
    n145,
    n125,
    n205
  );


  nor
  g430
  (
    n359,
    n123,
    n124,
    n216,
    n205
  );


  and
  g431
  (
    n348,
    n133,
    n141,
    n226,
    n235
  );


  and
  g432
  (
    n462,
    n179,
    n170,
    n140,
    n199
  );


  and
  g433
  (
    n360,
    n174,
    n117,
    n234,
    n213
  );


  xnor
  g434
  (
    n398,
    n211,
    n120,
    n143,
    n166
  );


  xor
  g435
  (
    n491,
    n180,
    n139,
    n144
  );


  and
  g436
  (
    n480,
    n114,
    n185,
    n162,
    n207
  );


  nor
  g437
  (
    n489,
    n145,
    n172,
    n168,
    n142
  );


  nand
  g438
  (
    n495,
    n232,
    n190,
    n225,
    n220
  );


  nor
  g439
  (
    n321,
    n201,
    n228,
    n203,
    n167
  );


  nor
  g440
  (
    n445,
    n125,
    n186,
    n147,
    n146
  );


  xor
  g441
  (
    n327,
    n113,
    n158,
    n222,
    n203
  );


  xor
  g442
  (
    n305,
    n124,
    n238,
    n139,
    n116
  );


  and
  g443
  (
    n473,
    n193,
    n113,
    n172,
    n192
  );


  and
  g444
  (
    n395,
    n213,
    n117,
    n223,
    n187
  );


  or
  g445
  (
    n323,
    n163,
    n188,
    n155,
    n239
  );


  xor
  g446
  (
    n476,
    n175,
    n133,
    n200,
    n209
  );


  or
  g447
  (
    n417,
    n219,
    n143,
    n189,
    n168
  );


  and
  g448
  (
    n350,
    n117,
    n227,
    n231,
    n142
  );


  or
  g449
  (
    n344,
    n119,
    n160,
    n231,
    n114
  );


  and
  g450
  (
    n455,
    n158,
    n145,
    n147,
    n171
  );


  or
  g451
  (
    n384,
    n194,
    n121,
    n201,
    n195
  );


  xor
  g452
  (
    n256,
    n209,
    n212,
    n167,
    n225
  );


  xnor
  g453
  (
    n320,
    n189,
    n153,
    n198,
    n148
  );


  nor
  g454
  (
    KeyWire_0_42,
    n138,
    n148,
    n134,
    n136
  );


  xnor
  g455
  (
    n444,
    n205,
    n169,
    n208,
    n175
  );


  or
  g456
  (
    n500,
    n149,
    n176,
    n200,
    n150
  );


  nand
  g457
  (
    n364,
    n121,
    n130,
    n191,
    n187
  );


  and
  g458
  (
    n433,
    n156,
    n119,
    n166,
    n168
  );


  or
  g459
  (
    n493,
    n206,
    n204,
    n217,
    n137
  );


  or
  g460
  (
    n293,
    n218,
    n140,
    n132,
    n207
  );


  or
  g461
  (
    n447,
    n229,
    n219,
    n151,
    n126
  );


  xnor
  g462
  (
    n423,
    n116,
    n169,
    n230,
    n118
  );


  and
  g463
  (
    n247,
    n115,
    n214,
    n135,
    n236
  );


  xnor
  g464
  (
    n388,
    n139,
    n233,
    n208,
    n153
  );


  xnor
  g465
  (
    KeyWire_0_50,
    n179,
    n140,
    n214,
    n165
  );


  nor
  g466
  (
    n425,
    n180,
    n200,
    n123,
    n198
  );


  nand
  g467
  (
    n418,
    n146,
    n226,
    n187,
    n210
  );


  and
  g468
  (
    n421,
    n150,
    n219,
    n154,
    n146
  );


  or
  g469
  (
    n260,
    n169,
    n120,
    n202,
    n173
  );


  xor
  g470
  (
    n343,
    n188,
    n152,
    n240,
    n221
  );


  xnor
  g471
  (
    n281,
    n171,
    n151,
    n204,
    n186
  );


  nand
  g472
  (
    n436,
    n211,
    n220,
    n158,
    n127
  );


  or
  g473
  (
    n399,
    n222,
    n137,
    n130,
    n171
  );


  or
  g474
  (
    n368,
    n191,
    n214,
    n202,
    n124
  );


  xor
  g475
  (
    KeyWire_0_2,
    n138,
    n213,
    n229,
    n209
  );


  or
  g476
  (
    n286,
    n134,
    n223,
    n160,
    n235
  );


  not
  g477
  (
    n762,
    n337
  );


  buf
  g478
  (
    n673,
    n402
  );


  buf
  g479
  (
    n682,
    n456
  );


  not
  g480
  (
    n534,
    n279
  );


  not
  g481
  (
    n845,
    n348
  );


  buf
  g482
  (
    n590,
    n299
  );


  not
  g483
  (
    n528,
    n344
  );


  buf
  g484
  (
    n747,
    n18
  );


  not
  g485
  (
    n823,
    n320
  );


  not
  g486
  (
    n776,
    n483
  );


  not
  g487
  (
    n899,
    n374
  );


  not
  g488
  (
    n721,
    n477
  );


  not
  g489
  (
    n654,
    n259
  );


  buf
  g490
  (
    n798,
    n303
  );


  buf
  g491
  (
    n792,
    n312
  );


  buf
  g492
  (
    n810,
    n374
  );


  not
  g493
  (
    n584,
    n376
  );


  buf
  g494
  (
    n724,
    n345
  );


  buf
  g495
  (
    n917,
    n403
  );


  buf
  g496
  (
    n913,
    n323
  );


  not
  g497
  (
    n729,
    n273
  );


  buf
  g498
  (
    n872,
    n441
  );


  buf
  g499
  (
    n780,
    n461
  );


  buf
  g500
  (
    n625,
    n475
  );


  not
  g501
  (
    n617,
    n389
  );


  buf
  g502
  (
    n740,
    n409
  );


  buf
  g503
  (
    n681,
    n57
  );


  not
  g504
  (
    n831,
    n482
  );


  not
  g505
  (
    n766,
    n337
  );


  not
  g506
  (
    n954,
    n390
  );


  buf
  g507
  (
    n842,
    n411
  );


  not
  g508
  (
    n542,
    n360
  );


  not
  g509
  (
    n609,
    n417
  );


  not
  g510
  (
    n870,
    n443
  );


  buf
  g511
  (
    n518,
    n18
  );


  not
  g512
  (
    n647,
    n417
  );


  not
  g513
  (
    n770,
    n446
  );


  not
  g514
  (
    n697,
    n329
  );


  not
  g515
  (
    n962,
    n245
  );


  buf
  g516
  (
    KeyWire_0_5,
    n485
  );


  buf
  g517
  (
    n541,
    n469
  );


  not
  g518
  (
    n514,
    n281
  );


  buf
  g519
  (
    KeyWire_0_23,
    n495
  );


  not
  g520
  (
    n704,
    n476
  );


  not
  g521
  (
    n649,
    n283
  );


  not
  g522
  (
    n614,
    n344
  );


  not
  g523
  (
    n522,
    n272
  );


  buf
  g524
  (
    n765,
    n267
  );


  buf
  g525
  (
    n841,
    n452
  );


  not
  g526
  (
    n540,
    n296
  );


  buf
  g527
  (
    n879,
    n423
  );


  not
  g528
  (
    n675,
    n300
  );


  not
  g529
  (
    n888,
    n302
  );


  not
  g530
  (
    n859,
    n299
  );


  not
  g531
  (
    n858,
    n368
  );


  not
  g532
  (
    n607,
    n380
  );


  not
  g533
  (
    n904,
    n342
  );


  not
  g534
  (
    n964,
    n458
  );


  buf
  g535
  (
    n887,
    n471
  );


  not
  g536
  (
    n662,
    n472
  );


  not
  g537
  (
    n652,
    n341
  );


  buf
  g538
  (
    n574,
    n248
  );


  not
  g539
  (
    n703,
    n250
  );


  buf
  g540
  (
    n644,
    n248
  );


  buf
  g541
  (
    n808,
    n479
  );


  buf
  g542
  (
    n637,
    n411
  );


  buf
  g543
  (
    n725,
    n277
  );


  not
  g544
  (
    n559,
    n313
  );


  not
  g545
  (
    n728,
    n413
  );


  not
  g546
  (
    n757,
    n400
  );


  buf
  g547
  (
    n715,
    n367
  );


  buf
  g548
  (
    n612,
    n251
  );


  not
  g549
  (
    n633,
    n382
  );


  buf
  g550
  (
    n796,
    n308
  );


  buf
  g551
  (
    n783,
    n241
  );


  buf
  g552
  (
    n691,
    n488
  );


  not
  g553
  (
    n670,
    n408
  );


  not
  g554
  (
    n549,
    n312
  );


  not
  g555
  (
    n521,
    n338
  );


  not
  g556
  (
    n961,
    n397
  );


  buf
  g557
  (
    n722,
    n498
  );


  buf
  g558
  (
    n925,
    n421
  );


  not
  g559
  (
    n854,
    n317
  );


  not
  g560
  (
    n733,
    n454
  );


  buf
  g561
  (
    n579,
    n419
  );


  buf
  g562
  (
    n587,
    n363
  );


  buf
  g563
  (
    n867,
    n265
  );


  not
  g564
  (
    n717,
    n430
  );


  not
  g565
  (
    n640,
    n461
  );


  buf
  g566
  (
    n832,
    n454
  );


  buf
  g567
  (
    n865,
    n311
  );


  buf
  g568
  (
    n892,
    n308
  );


  buf
  g569
  (
    n509,
    n362
  );


  buf
  g570
  (
    n695,
    n296
  );


  not
  g571
  (
    n781,
    n490
  );


  not
  g572
  (
    n850,
    n387
  );


  buf
  g573
  (
    n575,
    n365
  );


  buf
  g574
  (
    n567,
    n279
  );


  not
  g575
  (
    KeyWire_0_40,
    n325
  );


  not
  g576
  (
    n802,
    n354
  );


  buf
  g577
  (
    n804,
    n260
  );


  buf
  g578
  (
    KeyWire_0_28,
    n267
  );


  not
  g579
  (
    n545,
    n326
  );


  not
  g580
  (
    n539,
    n251
  );


  buf
  g581
  (
    n576,
    n491
  );


  not
  g582
  (
    n566,
    n426
  );


  buf
  g583
  (
    KeyWire_0_18,
    n334
  );


  buf
  g584
  (
    n634,
    n481
  );


  buf
  g585
  (
    n864,
    n289
  );


  not
  g586
  (
    n732,
    n310
  );


  buf
  g587
  (
    n905,
    n385
  );


  not
  g588
  (
    KeyWire_0_11,
    n380
  );


  not
  g589
  (
    n684,
    n379
  );


  not
  g590
  (
    n818,
    n442
  );


  not
  g591
  (
    n583,
    n289
  );


  buf
  g592
  (
    KeyWire_0_9,
    n318
  );


  not
  g593
  (
    n746,
    n365
  );


  not
  g594
  (
    n943,
    n338
  );


  not
  g595
  (
    n803,
    n280
  );


  buf
  g596
  (
    n606,
    n308
  );


  buf
  g597
  (
    n742,
    n364
  );


  not
  g598
  (
    n581,
    n375
  );


  not
  g599
  (
    n713,
    n348
  );


  buf
  g600
  (
    n585,
    n271
  );


  buf
  g601
  (
    n743,
    n413
  );


  buf
  g602
  (
    n779,
    n297
  );


  not
  g603
  (
    n761,
    n328
  );


  not
  g604
  (
    n886,
    n375
  );


  buf
  g605
  (
    n772,
    n309
  );


  not
  g606
  (
    n941,
    n464
  );


  not
  g607
  (
    n608,
    n266
  );


  not
  g608
  (
    n690,
    n389
  );


  not
  g609
  (
    n664,
    n279
  );


  buf
  g610
  (
    n526,
    n378
  );


  not
  g611
  (
    n699,
    n335
  );


  buf
  g612
  (
    n786,
    n374
  );


  not
  g613
  (
    n828,
    n306
  );


  not
  g614
  (
    n829,
    n255
  );


  not
  g615
  (
    n693,
    n488
  );


  buf
  g616
  (
    n598,
    n485
  );


  buf
  g617
  (
    KeyWire_0_62,
    n502
  );


  buf
  g618
  (
    n951,
    n482
  );


  buf
  g619
  (
    KeyWire_0_21,
    n309
  );


  buf
  g620
  (
    n689,
    n323
  );


  buf
  g621
  (
    n914,
    n487
  );


  buf
  g622
  (
    n911,
    n491
  );


  not
  g623
  (
    n705,
    n383
  );


  buf
  g624
  (
    n618,
    n398
  );


  not
  g625
  (
    n718,
    n308
  );


  buf
  g626
  (
    n927,
    n276
  );


  buf
  g627
  (
    n727,
    n295
  );


  buf
  g628
  (
    n547,
    n254
  );


  buf
  g629
  (
    KeyWire_0_47,
    n307
  );


  buf
  g630
  (
    n702,
    n492
  );


  buf
  g631
  (
    n696,
    n435
  );


  not
  g632
  (
    n550,
    n344
  );


  not
  g633
  (
    n855,
    n315
  );


  buf
  g634
  (
    n869,
    n18
  );


  not
  g635
  (
    KeyWire_0_8,
    n379
  );


  buf
  g636
  (
    n834,
    n17
  );


  not
  g637
  (
    n745,
    n270
  );


  buf
  g638
  (
    n931,
    n268
  );


  buf
  g639
  (
    n853,
    n386
  );


  buf
  g640
  (
    n674,
    n252
  );


  not
  g641
  (
    n785,
    n340
  );


  not
  g642
  (
    n846,
    n16
  );


  not
  g643
  (
    n656,
    n356
  );


  buf
  g644
  (
    n592,
    n322
  );


  buf
  g645
  (
    n885,
    n249
  );


  not
  g646
  (
    n738,
    n254
  );


  buf
  g647
  (
    KeyWire_0_56,
    n405
  );


  buf
  g648
  (
    n597,
    n391
  );


  buf
  g649
  (
    n601,
    n356
  );


  buf
  g650
  (
    n908,
    n263
  );


  buf
  g651
  (
    n963,
    n282
  );


  buf
  g652
  (
    n833,
    n478
  );


  buf
  g653
  (
    n760,
    n404
  );


  buf
  g654
  (
    n815,
    n492
  );


  not
  g655
  (
    n852,
    n345
  );


  not
  g656
  (
    n525,
    n378
  );


  buf
  g657
  (
    n700,
    n355
  );


  buf
  g658
  (
    n944,
    n399
  );


  not
  g659
  (
    n657,
    n294
  );


  not
  g660
  (
    n929,
    n442
  );


  buf
  g661
  (
    n671,
    n242
  );


  not
  g662
  (
    n650,
    n464
  );


  buf
  g663
  (
    n873,
    n290
  );


  not
  g664
  (
    n685,
    n304
  );


  not
  g665
  (
    n714,
    n17
  );


  not
  g666
  (
    n755,
    n459
  );


  not
  g667
  (
    n897,
    n440
  );


  buf
  g668
  (
    n767,
    n441
  );


  not
  g669
  (
    n805,
    n388
  );


  buf
  g670
  (
    n558,
    n264
  );


  not
  g671
  (
    n701,
    n422
  );


  not
  g672
  (
    n748,
    n352
  );


  buf
  g673
  (
    n641,
    n365
  );


  not
  g674
  (
    n546,
    n448
  );


  not
  g675
  (
    n946,
    n478
  );


  buf
  g676
  (
    n639,
    n288
  );


  buf
  g677
  (
    n953,
    n325
  );


  not
  g678
  (
    n898,
    n17
  );


  not
  g679
  (
    n847,
    n447
  );


  buf
  g680
  (
    n512,
    n309
  );


  buf
  g681
  (
    n933,
    n463
  );


  buf
  g682
  (
    n555,
    n405
  );


  buf
  g683
  (
    KeyWire_0_22,
    n306
  );


  not
  g684
  (
    n775,
    n459
  );


  buf
  g685
  (
    n744,
    n498
  );


  not
  g686
  (
    n942,
    n323
  );


  buf
  g687
  (
    n794,
    n463
  );


  buf
  g688
  (
    n616,
    n450
  );


  buf
  g689
  (
    n874,
    n39
  );


  buf
  g690
  (
    n809,
    n347
  );


  not
  g691
  (
    n688,
    n352
  );


  buf
  g692
  (
    n615,
    n462
  );


  not
  g693
  (
    n825,
    n320
  );


  not
  g694
  (
    n720,
    n442
  );


  not
  g695
  (
    n707,
    n295
  );


  not
  g696
  (
    n737,
    n256
  );


  not
  g697
  (
    n503,
    n350
  );


  not
  g698
  (
    n920,
    n246
  );


  buf
  g699
  (
    n838,
    n317
  );


  not
  g700
  (
    n570,
    n294
  );


  not
  g701
  (
    KeyWire_0_49,
    n386
  );


  buf
  g702
  (
    n921,
    n476
  );


  buf
  g703
  (
    n891,
    n294
  );


  not
  g704
  (
    n800,
    n304
  );


  not
  g705
  (
    n948,
    n396
  );


  not
  g706
  (
    n824,
    n490
  );


  buf
  g707
  (
    n513,
    n423
  );


  not
  g708
  (
    n749,
    n293
  );


  not
  g709
  (
    n949,
    n450
  );


  buf
  g710
  (
    n679,
    n355
  );


  buf
  g711
  (
    n940,
    n458
  );


  not
  g712
  (
    n790,
    n292
  );


  not
  g713
  (
    n677,
    n413
  );


  buf
  g714
  (
    n843,
    n415
  );


  not
  g715
  (
    n645,
    n385
  );


  buf
  g716
  (
    KeyWire_0_59,
    n333
  );


  buf
  g717
  (
    KeyWire_0_32,
    n331
  );


  not
  g718
  (
    n698,
    n362
  );


  not
  g719
  (
    n814,
    n499
  );


  not
  g720
  (
    n706,
    n18
  );


  buf
  g721
  (
    n894,
    n282
  );


  not
  g722
  (
    n939,
    n492
  );


  not
  g723
  (
    n906,
    n493
  );


  not
  g724
  (
    n777,
    n342
  );


  buf
  g725
  (
    n801,
    n452
  );


  buf
  g726
  (
    n900,
    n490
  );


  buf
  g727
  (
    n957,
    n501
  );


  not
  g728
  (
    n840,
    n19
  );


  not
  g729
  (
    n519,
    n432
  );


  buf
  g730
  (
    n544,
    n290
  );


  buf
  g731
  (
    n543,
    n253
  );


  buf
  g732
  (
    n537,
    n377
  );


  buf
  g733
  (
    n508,
    n343
  );


  buf
  g734
  (
    n907,
    n486
  );


  buf
  g735
  (
    n789,
    n332
  );


  buf
  g736
  (
    n924,
    n324
  );


  not
  g737
  (
    n646,
    n484
  );


  buf
  g738
  (
    n569,
    n367
  );


  not
  g739
  (
    n915,
    n431
  );


  not
  g740
  (
    n868,
    n323
  );


  not
  g741
  (
    n588,
    n443
  );


  xnor
  g742
  (
    KeyWire_0_52,
    n298,
    n348
  );


  nand
  g743
  (
    n936,
    n368,
    n357,
    n341,
    n356
  );


  nand
  g744
  (
    n602,
    n410,
    n493,
    n370,
    n325
  );


  xor
  g745
  (
    n626,
    n400,
    n366,
    n363,
    n359
  );


  nor
  g746
  (
    n932,
    n424,
    n435,
    n247,
    n482
  );


  and
  g747
  (
    KeyWire_0_43,
    n425,
    n281,
    n346,
    n242
  );


  nand
  g748
  (
    n667,
    n331,
    n366,
    n336,
    n496
  );


  xor
  g749
  (
    n551,
    n262,
    n457,
    n388,
    n479
  );


  nor
  g750
  (
    n883,
    n350,
    n421,
    n414,
    n392
  );


  xnor
  g751
  (
    n938,
    n259,
    n422,
    n429,
    n257
  );


  and
  g752
  (
    n826,
    n375,
    n270,
    n420,
    n429
  );


  and
  g753
  (
    n912,
    n415,
    n500,
    n361,
    n377
  );


  xnor
  g754
  (
    n511,
    n438,
    n405,
    n39,
    n428
  );


  and
  g755
  (
    n945,
    n336,
    n486,
    n360,
    n418
  );


  nor
  g756
  (
    n532,
    n351,
    n291,
    n253,
    n274
  );


  and
  g757
  (
    n935,
    n301,
    n276,
    n395,
    n488
  );


  and
  g758
  (
    n764,
    n440,
    n387,
    n343,
    n363
  );


  xnor
  g759
  (
    n716,
    n257,
    n466,
    n480,
    n370
  );


  and
  g760
  (
    n788,
    n305,
    n320,
    n424,
    n278
  );


  and
  g761
  (
    n622,
    n380,
    n252,
    n495,
    n17
  );


  and
  g762
  (
    n758,
    n272,
    n430,
    n368,
    n392
  );


  nor
  g763
  (
    n750,
    n342,
    n357,
    n437,
    n355
  );


  nand
  g764
  (
    n564,
    n439,
    n241,
    n484,
    n483
  );


  and
  g765
  (
    n510,
    n401,
    n502,
    n305,
    n416
  );


  xnor
  g766
  (
    n910,
    n371,
    n433,
    n243,
    n400
  );


  or
  g767
  (
    n821,
    n427,
    n299,
    n485,
    n278
  );


  xor
  g768
  (
    n861,
    n307,
    n384,
    n321,
    n427
  );


  or
  g769
  (
    n571,
    n429,
    n493,
    n398
  );


  or
  g770
  (
    n604,
    n295,
    n340,
    n302,
    n258
  );


  nand
  g771
  (
    n605,
    n291,
    n487,
    n277,
    n501
  );


  or
  g772
  (
    n552,
    n334,
    n329,
    n371,
    n495
  );


  nand
  g773
  (
    n860,
    n440,
    n263,
    n393,
    n500
  );


  nor
  g774
  (
    n603,
    n290,
    n252,
    n269,
    n258
  );


  nand
  g775
  (
    n623,
    n412,
    n428,
    n335,
    n367
  );


  nor
  g776
  (
    KeyWire_0_58,
    n359,
    n245,
    n447,
    n329
  );


  nand
  g777
  (
    n934,
    n286,
    n462,
    n403,
    n371
  );


  nand
  g778
  (
    n782,
    n353,
    n465,
    n268,
    n285
  );


  nand
  g779
  (
    KeyWire_0_1,
    n407,
    n305,
    n446,
    n462
  );


  nand
  g780
  (
    n735,
    n474,
    n354,
    n477,
    n351
  );


  and
  g781
  (
    n531,
    n445,
    n258,
    n491,
    n343
  );


  or
  g782
  (
    n620,
    n465,
    n401,
    n427,
    n246
  );


  xor
  g783
  (
    n902,
    n319,
    n341,
    n387,
    n490
  );


  nor
  g784
  (
    n573,
    n473,
    n481,
    n393,
    n461
  );


  and
  g785
  (
    n947,
    n451,
    n367,
    n352,
    n260
  );


  and
  g786
  (
    n527,
    n322,
    n395,
    n423,
    n460
  );


  nand
  g787
  (
    n769,
    n409,
    n424,
    n410,
    n342
  );


  xnor
  g788
  (
    n928,
    n251,
    n261,
    n466,
    n285
  );


  and
  g789
  (
    n816,
    n287,
    n281,
    n494,
    n316
  );


  xnor
  g790
  (
    KeyWire_0_61,
    n498,
    n425,
    n386,
    n369
  );


  xor
  g791
  (
    n635,
    n482,
    n468,
    n285,
    n280
  );


  nor
  g792
  (
    n572,
    n262,
    n309,
    n340,
    n440
  );


  xor
  g793
  (
    n889,
    n284,
    n287,
    n419,
    n426
  );


  xnor
  g794
  (
    n880,
    n477,
    n385,
    n283,
    n404
  );


  and
  g795
  (
    n683,
    n286,
    n481,
    n349,
    n288
  );


  and
  g796
  (
    n965,
    n393,
    n480,
    n477,
    n470
  );


  nand
  g797
  (
    n669,
    n273,
    n409,
    n394,
    n470
  );


  xor
  g798
  (
    KeyWire_0_19,
    n306,
    n354,
    n313,
    n345
  );


  nand
  g799
  (
    n580,
    n288,
    n470,
    n417,
    n497
  );


  nand
  g800
  (
    n844,
    n288,
    n303,
    n439,
    n275
  );


  xor
  g801
  (
    n771,
    n337,
    n273,
    n326,
    n500
  );


  xor
  g802
  (
    n866,
    n412,
    n311,
    n262,
    n270
  );


  or
  g803
  (
    n565,
    n435,
    n411,
    n473,
    n331
  );


  and
  g804
  (
    n751,
    n461,
    n349,
    n329,
    n366
  );


  xor
  g805
  (
    n586,
    n349,
    n416,
    n265,
    n418
  );


  nand
  g806
  (
    n563,
    n394,
    n256,
    n258,
    n415
  );


  xnor
  g807
  (
    n875,
    n424,
    n491,
    n352,
    n414
  );


  or
  g808
  (
    n589,
    n468,
    n460,
    n343,
    n313
  );


  or
  g809
  (
    n708,
    n406,
    n405,
    n332,
    n336
  );


  or
  g810
  (
    n863,
    n416,
    n437,
    n403,
    n419
  );


  nor
  g811
  (
    n922,
    n330,
    n327,
    n277,
    n339
  );


  nand
  g812
  (
    n950,
    n271,
    n346,
    n318,
    n410
  );


  or
  g813
  (
    n797,
    n267,
    n396,
    n334,
    n353
  );


  and
  g814
  (
    n515,
    n437,
    n472,
    n257,
    n391
  );


  or
  g815
  (
    n806,
    n250,
    n486,
    n398,
    n358
  );


  nand
  g816
  (
    n817,
    n255,
    n331,
    n303,
    n423
  );


  nor
  g817
  (
    n595,
    n407,
    n264,
    n313,
    n426
  );


  nor
  g818
  (
    KeyWire_0_37,
    n260,
    n397,
    n243,
    n422
  );


  xnor
  g819
  (
    n791,
    n292,
    n328,
    n448,
    n314
  );


  xor
  g820
  (
    n877,
    n251,
    n254,
    n249,
    n322
  );


  xor
  g821
  (
    n960,
    n432,
    n357,
    n389,
    n449
  );


  nor
  g822
  (
    n636,
    n381,
    n341,
    n407,
    n496
  );


  nor
  g823
  (
    n600,
    n421,
    n446,
    n346,
    n403
  );


  or
  g824
  (
    n582,
    n397,
    n452,
    n484,
    n383
  );


  nor
  g825
  (
    KeyWire_0_54,
    n457,
    n319,
    n434,
    n360
  );


  nand
  g826
  (
    n837,
    n500,
    n428,
    n442,
    n411
  );


  xor
  g827
  (
    n561,
    n391,
    n453,
    n378,
    n298
  );


  and
  g828
  (
    n666,
    n377,
    n454,
    n374,
    n381
  );


  nand
  g829
  (
    n710,
    n362,
    n335,
    n372,
    n497
  );


  nand
  g830
  (
    n878,
    n373,
    n274,
    n291,
    n471
  );


  or
  g831
  (
    n711,
    n269,
    n456,
    n262,
    n266
  );


  and
  g832
  (
    n752,
    n447,
    n276,
    n271,
    n468
  );


  xnor
  g833
  (
    n857,
    n432,
    n253,
    n324,
    n314
  );


  nor
  g834
  (
    n517,
    n315,
    n321,
    n299,
    n479
  );


  xnor
  g835
  (
    n958,
    n282,
    n419,
    n346,
    n370
  );


  and
  g836
  (
    n773,
    n416,
    n466,
    n301,
    n383
  );


  or
  g837
  (
    n807,
    n363,
    n489,
    n360,
    n268
  );


  nand
  g838
  (
    n651,
    n383,
    n320,
    n418,
    n420
  );


  nor
  g839
  (
    n734,
    n255,
    n364,
    n347,
    n289
  );


  nand
  g840
  (
    n520,
    n297,
    n449,
    n314,
    n379
  );


  or
  g841
  (
    n668,
    n487,
    n441,
    n443,
    n369
  );


  nand
  g842
  (
    n630,
    n316,
    n380,
    n353,
    n399
  );


  or
  g843
  (
    n754,
    n444,
    n270,
    n430,
    n389
  );


  xnor
  g844
  (
    n655,
    n499,
    n387,
    n324,
    n275
  );


  xnor
  g845
  (
    n903,
    n265,
    n437,
    n469,
    n285
  );


  and
  g846
  (
    n632,
    n420,
    n464,
    n485,
    n399
  );


  nor
  g847
  (
    n909,
    n354,
    n489,
    n396,
    n317
  );


  xor
  g848
  (
    n562,
    n470,
    n496,
    n349,
    n361
  );


  or
  g849
  (
    n741,
    n439,
    n263,
    n372,
    n394
  );


  xor
  g850
  (
    n918,
    n444,
    n487,
    n295,
    n368
  );


  xor
  g851
  (
    n660,
    n376,
    n286,
    n254,
    n492
  );


  and
  g852
  (
    KeyWire_0_17,
    n384,
    n333,
    n350,
    n361
  );


  nand
  g853
  (
    n610,
    n330,
    n404,
    n436,
    n336
  );


  nand
  g854
  (
    n836,
    n460,
    n372,
    n392,
    n248
  );


  or
  g855
  (
    n624,
    n444,
    n333,
    n496,
    n322
  );


  nor
  g856
  (
    n694,
    n16,
    n358,
    n244,
    n401
  );


  nand
  g857
  (
    n901,
    n473,
    n307,
    n373,
    n406
  );


  and
  g858
  (
    n768,
    n436,
    n431,
    n330,
    n402
  );


  xor
  g859
  (
    n523,
    n245,
    n266,
    n296,
    n450
  );


  and
  g860
  (
    n553,
    n438,
    n364,
    n479,
    n388
  );


  or
  g861
  (
    n505,
    n339,
    n465,
    n247,
    n451
  );


  xnor
  g862
  (
    n822,
    n328,
    n445,
    n427,
    n391
  );


  and
  g863
  (
    n628,
    n327,
    n364,
    n301,
    n247
  );


  or
  g864
  (
    n952,
    n356,
    n351,
    n337,
    n481
  );


  xor
  g865
  (
    n648,
    n425,
    n256,
    n414,
    n249
  );


  and
  g866
  (
    n611,
    n319,
    n422,
    n438,
    n358
  );


  nand
  g867
  (
    n956,
    n292,
    n448,
    n269,
    n497
  );


  xor
  g868
  (
    n638,
    n373,
    n501,
    n311,
    n280
  );


  xnor
  g869
  (
    n529,
    n328,
    n456,
    n399,
    n256
  );


  xnor
  g870
  (
    n930,
    n426,
    n494,
    n264,
    n448
  );


  xnor
  g871
  (
    n778,
    n459,
    n303,
    n434,
    n339
  );


  or
  g872
  (
    n507,
    n296,
    n402,
    n287,
    n289
  );


  nand
  g873
  (
    n723,
    n472,
    n272,
    n277,
    n244
  );


  xor
  g874
  (
    n524,
    n483,
    n369,
    n480,
    n283
  );


  nand
  g875
  (
    n663,
    n443,
    n459,
    n316,
    n445
  );


  xor
  g876
  (
    n557,
    n460,
    n259,
    n395,
    n474
  );


  nor
  g877
  (
    n937,
    n458,
    n347,
    n281,
    n400
  );


  or
  g878
  (
    KeyWire_0_12,
    n455,
    n408,
    n465,
    n499
  );


  or
  g879
  (
    n848,
    n304,
    n351,
    n392,
    n488
  );


  xnor
  g880
  (
    n882,
    n318,
    n259,
    n269,
    n475
  );


  nand
  g881
  (
    n759,
    n475,
    n39,
    n406,
    n489
  );


  nand
  g882
  (
    n820,
    n338,
    n432,
    n433,
    n483
  );


  nor
  g883
  (
    KeyWire_0_36,
    n287,
    n311,
    n332,
    n330
  );


  nor
  g884
  (
    n813,
    n434,
    n494,
    n464,
    n446
  );


  or
  g885
  (
    n736,
    n453,
    n271,
    n457,
    n340
  );


  xor
  g886
  (
    n812,
    n292,
    n257,
    n324,
    n314
  );


  xor
  g887
  (
    n659,
    n407,
    n293,
    n390,
    n333
  );


  nor
  g888
  (
    n916,
    n300,
    n347,
    n406,
    n371
  );


  or
  g889
  (
    n680,
    n434,
    n325,
    n372,
    n267
  );


  xnor
  g890
  (
    n658,
    n307,
    n458,
    n462,
    n265
  );


  xor
  g891
  (
    n896,
    n456,
    n286,
    n431,
    n344
  );


  xnor
  g892
  (
    n763,
    n421,
    n498,
    n19,
    n469
  );


  xnor
  g893
  (
    n795,
    n410,
    n495,
    n381,
    n279
  );


  xor
  g894
  (
    n678,
    n348,
    n291,
    n260,
    n390
  );


  and
  g895
  (
    n774,
    n476,
    n316,
    n359,
    n350
  );


  nor
  g896
  (
    KeyWire_0_0,
    n429,
    n358,
    n420,
    n390
  );


  nand
  g897
  (
    n692,
    n384,
    n318,
    n275,
    n430
  );


  nand
  g898
  (
    n811,
    n317,
    n357,
    n474,
    n370
  );


  nor
  g899
  (
    n506,
    n475,
    n376,
    n339,
    n402
  );


  xor
  g900
  (
    n793,
    n353,
    n297,
    n451,
    n369
  );


  xor
  g901
  (
    n881,
    n293,
    n282,
    n396,
    n244
  );


  xnor
  g902
  (
    n726,
    n393,
    n398,
    n304,
    n335
  );


  or
  g903
  (
    n687,
    n274,
    n438,
    n253,
    n453
  );


  nand
  g904
  (
    n535,
    n376,
    n327,
    n263,
    n284
  );


  nand
  g905
  (
    n672,
    n241,
    n417,
    n382,
    n455
  );


  xnor
  g906
  (
    n835,
    n468,
    n312,
    n294,
    n321
  );


  and
  g907
  (
    n893,
    n319,
    n455,
    n290,
    n471
  );


  nand
  g908
  (
    n621,
    n467,
    n473,
    n478,
    n302
  );


  xor
  g909
  (
    n577,
    n261,
    n457,
    n409,
    n441
  );


  xor
  g910
  (
    n686,
    n243,
    n361,
    n272,
    n449
  );


  nand
  g911
  (
    n862,
    n486,
    n408,
    n268
  );


  nor
  g912
  (
    KeyWire_0_44,
    n480,
    n433,
    n418,
    n300
  );


  nor
  g913
  (
    n890,
    n315,
    n401,
    n366,
    n502
  );


  xnor
  g914
  (
    n876,
    n332,
    n280,
    n278,
    n467
  );


  or
  g915
  (
    n554,
    n474,
    n450,
    n255,
    n246
  );


  nand
  g916
  (
    n578,
    n453,
    n306,
    n463,
    n394
  );


  xor
  g917
  (
    n665,
    n471,
    n310,
    n447,
    n428
  );


  and
  g918
  (
    n784,
    n365,
    n415,
    n355,
    n466
  );


  xor
  g919
  (
    n849,
    n362,
    n375,
    n382,
    n435
  );


  nor
  g920
  (
    n619,
    n454,
    n312,
    n39,
    n310
  );


  xor
  g921
  (
    n871,
    n359,
    n274,
    n300,
    n242
  );


  xnor
  g922
  (
    n504,
    n463,
    n382,
    n297,
    n439
  );


  nand
  g923
  (
    KeyWire_0_34,
    n378,
    n326,
    n452,
    n436
  );


  nor
  g924
  (
    n959,
    n326,
    n472,
    n388,
    n444
  );


  and
  g925
  (
    n787,
    n315,
    n502,
    n455,
    n478
  );


  and
  g926
  (
    n923,
    n467,
    n449,
    n381,
    n278
  );


  or
  g927
  (
    n856,
    n275,
    n250,
    n264,
    n298
  );


  xor
  g928
  (
    n753,
    n377,
    n501,
    n436,
    n397
  );


  xnor
  g929
  (
    n538,
    n261,
    n425,
    n445,
    n284
  );


  xor
  g930
  (
    n819,
    n412,
    n476,
    n384,
    n413
  );


  nand
  g931
  (
    n599,
    n284,
    n433,
    n310,
    n261
  );


  xor
  g932
  (
    n731,
    n489,
    n385,
    n414,
    n494
  );


  xnor
  g933
  (
    n719,
    n252,
    n412,
    n386,
    n298
  );


  xnor
  g934
  (
    n676,
    n404,
    n302,
    n334,
    n338
  );


  nor
  g935
  (
    n653,
    n379,
    n266,
    n345,
    n431
  );


  or
  g936
  (
    n629,
    n321,
    n373,
    n467,
    n283
  );


  or
  g937
  (
    n756,
    n293,
    n276,
    n484,
    n273
  );


  nor
  g938
  (
    n709,
    n497,
    n499,
    n327,
    n469
  );


  xnor
  g939
  (
    n594,
    n395,
    n305,
    n451,
    n301
  );


  xnor
  g940
  (
    n1065,
    n964,
    n676,
    n796,
    n761
  );


  xnor
  g941
  (
    n1015,
    n520,
    n632,
    n963,
    n829
  );


  xnor
  g942
  (
    n1011,
    n954,
    n755,
    n546,
    n771
  );


  or
  g943
  (
    n966,
    n673,
    n619,
    n898,
    n798
  );


  nand
  g944
  (
    n1071,
    n887,
    n958,
    n665,
    n578
  );


  xnor
  g945
  (
    n1080,
    n651,
    n772,
    n835,
    n960
  );


  nor
  g946
  (
    n1035,
    n884,
    n911,
    n720,
    n633
  );


  xor
  g947
  (
    n1009,
    n932,
    n569,
    n856,
    n737
  );


  xor
  g948
  (
    n1068,
    n740,
    n641,
    n852,
    n838
  );


  xnor
  g949
  (
    n1063,
    n751,
    n645,
    n853,
    n843
  );


  and
  g950
  (
    n1000,
    n913,
    n867,
    n515,
    n945
  );


  or
  g951
  (
    n986,
    n809,
    n621,
    n612,
    n953
  );


  nor
  g952
  (
    n968,
    n734,
    n817,
    n943,
    n821
  );


  nand
  g953
  (
    n1029,
    n560,
    n675,
    n758,
    n618
  );


  xor
  g954
  (
    n970,
    n699,
    n568,
    n797,
    n636
  );


  nor
  g955
  (
    n1053,
    n875,
    n625,
    n775,
    n731
  );


  xor
  g956
  (
    n1008,
    n959,
    n929,
    n643,
    n690
  );


  nor
  g957
  (
    n1023,
    n837,
    n869,
    n537,
    n539
  );


  xnor
  g958
  (
    n1039,
    n600,
    n886,
    n890,
    n799
  );


  or
  g959
  (
    n1042,
    n519,
    n629,
    n790,
    n933
  );


  nand
  g960
  (
    n1046,
    n710,
    n698,
    n759,
    n601
  );


  or
  g961
  (
    KeyWire_0_10,
    n942,
    n963,
    n711,
    n514
  );


  or
  g962
  (
    n1005,
    n536,
    n604,
    n779,
    n727
  );


  xnor
  g963
  (
    n1075,
    n679,
    n575,
    n635,
    n952
  );


  and
  g964
  (
    n1062,
    n693,
    n926,
    n548,
    n683
  );


  xor
  g965
  (
    n1041,
    n812,
    n895,
    n824,
    n791
  );


  xnor
  g966
  (
    n1051,
    n879,
    n605,
    n940,
    n802
  );


  xor
  g967
  (
    n1048,
    n844,
    n863,
    n777,
    n792
  );


  nand
  g968
  (
    n981,
    n544,
    n707,
    n960,
    n881
  );


  and
  g969
  (
    n1001,
    n672,
    n860,
    n505,
    n961
  );


  nor
  g970
  (
    n1074,
    n834,
    n658,
    n778,
    n573
  );


  and
  g971
  (
    n1076,
    n677,
    n717,
    n756,
    n745
  );


  nor
  g972
  (
    n1081,
    n598,
    n811,
    n893,
    n752
  );


  nand
  g973
  (
    n1037,
    n694,
    n614,
    n748,
    n735
  );


  nand
  g974
  (
    n987,
    n814,
    n706,
    n764,
    n511
  );


  xor
  g975
  (
    n974,
    n905,
    n956,
    n729,
    n701
  );


  and
  g976
  (
    n980,
    n522,
    n868,
    n800,
    n883
  );


  xnor
  g977
  (
    n994,
    n577,
    n934,
    n552,
    n957
  );


  xnor
  g978
  (
    n998,
    n921,
    n611,
    n521,
    n682
  );


  xnor
  g979
  (
    n1034,
    n718,
    n902,
    n785,
    n702
  );


  or
  g980
  (
    n1020,
    n556,
    n565,
    n857,
    n832
  );


  nand
  g981
  (
    n989,
    n557,
    n849,
    n616,
    n951
  );


  xor
  g982
  (
    n1047,
    n649,
    n958,
    n674,
    n566
  );


  and
  g983
  (
    n977,
    n874,
    n916,
    n952,
    n613
  );


  xnor
  g984
  (
    n1066,
    n754,
    n965,
    n610,
    n789
  );


  xnor
  g985
  (
    n1018,
    n864,
    n634,
    n862,
    n527
  );


  nand
  g986
  (
    n973,
    n769,
    n762,
    n508,
    n586
  );


  nor
  g987
  (
    n991,
    n558,
    n816,
    n554,
    n861
  );


  xnor
  g988
  (
    n1033,
    n736,
    n591,
    n647,
    n846
  );


  nand
  g989
  (
    n1030,
    n813,
    n962,
    n786,
    n865
  );


  or
  g990
  (
    n992,
    n845,
    n903,
    n750,
    n631
  );


  nand
  g991
  (
    n1043,
    n794,
    n908,
    n526,
    n739
  );


  or
  g992
  (
    n978,
    n741,
    n842,
    n815,
    n776
  );


  xnor
  g993
  (
    n1010,
    n553,
    n551,
    n766,
    n582
  );


  xnor
  g994
  (
    n1038,
    n770,
    n581,
    n545,
    n685
  );


  nor
  g995
  (
    n995,
    n839,
    n939,
    n567,
    n744
  );


  xor
  g996
  (
    n1070,
    n584,
    n650,
    n697,
    n946
  );


  xnor
  g997
  (
    n1024,
    n962,
    n877,
    n858,
    n657
  );


  or
  g998
  (
    n997,
    n836,
    n851,
    n607,
    n914
  );


  nand
  g999
  (
    n1077,
    n524,
    n894,
    n725,
    n507
  );


  nand
  g1000
  (
    n1028,
    n630,
    n904,
    n572,
    n746
  );


  nor
  g1001
  (
    n975,
    n749,
    n826,
    n922,
    n543
  );


  or
  g1002
  (
    n976,
    n724,
    n555,
    n599,
    n804
  );


  xnor
  g1003
  (
    n1002,
    n823,
    n620,
    n708,
    n907
  );


  xnor
  g1004
  (
    n999,
    n892,
    n660,
    n924,
    n954
  );


  nand
  g1005
  (
    n1049,
    n533,
    n955,
    n885,
    n589
  );


  xnor
  g1006
  (
    n1016,
    n595,
    n623,
    n918,
    n965
  );


  or
  g1007
  (
    n1055,
    n678,
    n882,
    n803,
    n901
  );


  nand
  g1008
  (
    n1058,
    n726,
    n959,
    n593,
    n767
  );


  nor
  g1009
  (
    n1012,
    n615,
    n663,
    n847,
    n506
  );


  or
  g1010
  (
    n1027,
    n805,
    n587,
    n897,
    n841
  );


  and
  g1011
  (
    n1054,
    n850,
    n757,
    n919,
    n900
  );


  xor
  g1012
  (
    n1013,
    n656,
    n781,
    n912,
    n585
  );


  or
  g1013
  (
    n1006,
    n529,
    n733,
    n662,
    n906
  );


  and
  g1014
  (
    n1064,
    n518,
    n563,
    n872,
    n655
  );


  nor
  g1015
  (
    n1079,
    n628,
    n878,
    n760,
    n590
  );


  xor
  g1016
  (
    n1044,
    n580,
    n542,
    n525,
    n915
  );


  or
  g1017
  (
    n1007,
    n592,
    n859,
    n899,
    n774
  );


  and
  g1018
  (
    n1014,
    n602,
    n531,
    n541,
    n828
  );


  xor
  g1019
  (
    n1040,
    n889,
    n719,
    n747,
    n638
  );


  xor
  g1020
  (
    n1073,
    n583,
    n920,
    n876,
    n936
  );


  or
  g1021
  (
    n1082,
    n705,
    n830,
    n788,
    n855
  );


  and
  g1022
  (
    n1022,
    n848,
    n709,
    n671,
    n571
  );


  xor
  g1023
  (
    n988,
    n528,
    n696,
    n576,
    n550
  );


  xor
  g1024
  (
    n1067,
    n715,
    n941,
    n810,
    n742
  );


  nor
  g1025
  (
    n1069,
    n603,
    n723,
    n646,
    n949
  );


  nor
  g1026
  (
    n1057,
    n637,
    n819,
    n686,
    n820
  );


  xor
  g1027
  (
    n971,
    n961,
    n948,
    n609,
    n784
  );


  xnor
  g1028
  (
    n996,
    n668,
    n654,
    n714,
    n669
  );


  or
  g1029
  (
    n1031,
    n753,
    n938,
    n713,
    n688
  );


  nor
  g1030
  (
    n1004,
    n953,
    n806,
    n680,
    n574
  );


  xnor
  g1031
  (
    n1050,
    n763,
    n930,
    n866,
    n523
  );


  nor
  g1032
  (
    n993,
    n666,
    n642,
    n597,
    n831
  );


  nand
  g1033
  (
    n1036,
    n570,
    n712,
    n782,
    n854
  );


  xnor
  g1034
  (
    n1017,
    n716,
    n738,
    n684,
    n722
  );


  and
  g1035
  (
    n1072,
    n562,
    n691,
    n925,
    n703
  );


  or
  g1036
  (
    n984,
    n670,
    n534,
    n937,
    n549
  );


  or
  g1037
  (
    n967,
    n957,
    n822,
    n639,
    n773
  );


  and
  g1038
  (
    n990,
    n840,
    n516,
    n743,
    n538
  );


  xnor
  g1039
  (
    n985,
    n730,
    n692,
    n644,
    n765
  );


  xor
  g1040
  (
    n1003,
    n659,
    n917,
    n513,
    n579
  );


  xor
  g1041
  (
    n1026,
    n624,
    n667,
    n808,
    n928
  );


  nor
  g1042
  (
    KeyWire_0_35,
    n880,
    n964,
    n653,
    n947
  );


  and
  g1043
  (
    n972,
    n732,
    n594,
    n910,
    n956
  );


  nand
  g1044
  (
    n969,
    n931,
    n768,
    n535,
    n661
  );


  or
  g1045
  (
    n979,
    n721,
    n695,
    n681,
    n728
  );


  nor
  g1046
  (
    n1032,
    n873,
    n532,
    n807,
    n588
  );


  and
  g1047
  (
    n982,
    n564,
    n617,
    n783,
    n793
  );


  xor
  g1048
  (
    n1045,
    n935,
    n627,
    n704,
    n801
  );


  xor
  g1049
  (
    n1060,
    n606,
    n825,
    n795,
    n559
  );


  xor
  g1050
  (
    n1056,
    n787,
    n504,
    n871,
    n512
  );


  or
  g1051
  (
    n1021,
    n664,
    n944,
    n780,
    n626
  );


  nor
  g1052
  (
    n1084,
    n608,
    n888,
    n510,
    n540
  );


  nand
  g1053
  (
    n1052,
    n640,
    n833,
    n909,
    n517
  );


  or
  g1054
  (
    n1078,
    n891,
    n927,
    n870,
    n530
  );


  xnor
  g1055
  (
    n1061,
    n955,
    n827,
    n547,
    n596
  );


  nor
  g1056
  (
    n1059,
    n509,
    n622,
    n648,
    n923
  );


  xnor
  g1057
  (
    KeyWire_0_6,
    n818,
    n689,
    n896,
    n561
  );


  or
  g1058
  (
    n1019,
    n950,
    n700,
    n652,
    n687
  );


  nand
  g1059
  (
    n1111,
    n990,
    n1051,
    n1079,
    n1015
  );


  xnor
  g1060
  (
    n1110,
    n1040,
    n1034,
    n1035,
    n974
  );


  xor
  g1061
  (
    n1091,
    n1066,
    n1064,
    n1020,
    n1014
  );


  nand
  g1062
  (
    n1101,
    n1003,
    n1000,
    n1036,
    n1056
  );


  or
  g1063
  (
    n1106,
    n1065,
    n1010,
    n1026,
    n1002
  );


  or
  g1064
  (
    n1100,
    n994,
    n1012,
    n979,
    n1021
  );


  nand
  g1065
  (
    n1094,
    n1080,
    n1068,
    n1075,
    n1022
  );


  nor
  g1066
  (
    n1109,
    n1057,
    n1071,
    n1006,
    n986
  );


  xor
  g1067
  (
    n1112,
    n969,
    n995,
    n1031,
    n1039
  );


  or
  g1068
  (
    n1095,
    n968,
    n981,
    n1044,
    n1053
  );


  or
  g1069
  (
    n1087,
    n1050,
    n989,
    n996,
    n966
  );


  xor
  g1070
  (
    n1108,
    n1063,
    n1058,
    n1009,
    n988
  );


  xor
  g1071
  (
    n1104,
    n1073,
    n1016,
    n1025,
    n1052
  );


  and
  g1072
  (
    n1092,
    n978,
    n997,
    n1061,
    n1028
  );


  xor
  g1073
  (
    n1088,
    n1024,
    n980,
    n1011,
    n1019
  );


  nor
  g1074
  (
    n1090,
    n973,
    n1005,
    n1042,
    n971
  );


  nand
  g1075
  (
    n1085,
    n1017,
    n972,
    n1033,
    n1077
  );


  nor
  g1076
  (
    n1089,
    n998,
    n1037,
    n1008,
    n967
  );


  xnor
  g1077
  (
    n1096,
    n1067,
    n1004,
    n991,
    n1018
  );


  nor
  g1078
  (
    n1093,
    n1007,
    n1046,
    n985,
    n1001
  );


  nand
  g1079
  (
    n1097,
    n1072,
    n970,
    n1029,
    n1070
  );


  xnor
  g1080
  (
    n1105,
    n1043,
    n1060,
    n987,
    n1048
  );


  xnor
  g1081
  (
    KeyWire_0_48,
    n983,
    n1013,
    n993,
    n984
  );


  xnor
  g1082
  (
    n1102,
    n992,
    n1059,
    n1030,
    n976
  );


  xor
  g1083
  (
    n1113,
    n1081,
    n1078,
    n1049,
    n975
  );


  and
  g1084
  (
    n1107,
    n1076,
    n977,
    n1027,
    n1069
  );


  nor
  g1085
  (
    n1099,
    n1045,
    n1047,
    n1032,
    n1062
  );


  nor
  g1086
  (
    n1086,
    n999,
    n1023,
    n982,
    n1041
  );


  nand
  g1087
  (
    n1098,
    n1054,
    n1038,
    n1055,
    n1074
  );


  xor
  g1088
  (
    n1123,
    n24,
    n58,
    n25,
    n1111
  );


  or
  g1089
  (
    n1121,
    n21,
    n21,
    n25,
    n20
  );


  and
  g1090
  (
    n1125,
    n23,
    n22,
    n57
  );


  nor
  g1091
  (
    n1122,
    n1110,
    n23,
    n20,
    n24
  );


  xor
  g1092
  (
    n1119,
    n1097,
    n1102,
    n1107,
    n19
  );


  nand
  g1093
  (
    n1118,
    n1105,
    n58,
    n1104,
    n1098
  );


  nand
  g1094
  (
    n1117,
    n1100,
    n23,
    n19
  );


  nand
  g1095
  (
    n1115,
    n1103,
    n22,
    n57
  );


  nand
  g1096
  (
    n1120,
    n25,
    n20,
    n58,
    n1099
  );


  xnor
  g1097
  (
    n1116,
    n21,
    n1112,
    n1108,
    n25
  );


  xnor
  g1098
  (
    n1124,
    n1106,
    n1109,
    n24,
    n1101
  );


  xnor
  g1099
  (
    KeyWire_0_51,
    n21,
    n20,
    n1113,
    n24
  );


  buf
  g1100
  (
    n1129,
    n1114
  );


  not
  g1101
  (
    n1127,
    n1115
  );


  or
  g1102
  (
    n1128,
    n1118,
    n1117,
    n1115,
    n1114
  );


  xnor
  g1103
  (
    n1130,
    n1118,
    n1115,
    n1116,
    n1117
  );


  xor
  g1104
  (
    n1126,
    n1114,
    n1116,
    n1117
  );


  and
  g1105
  (
    n1132,
    n1119,
    n1127,
    n1118
  );


  and
  g1106
  (
    n1138,
    n1128,
    n1127,
    n1084,
    n1126
  );


  xnor
  g1107
  (
    n1136,
    n1130,
    n1126,
    n1129,
    n1127
  );


  nor
  g1108
  (
    n1133,
    n1126,
    n1128,
    n1129,
    n1118
  );


  nor
  g1109
  (
    n1135,
    n1120,
    n1129,
    n1130
  );


  nor
  g1110
  (
    KeyWire_0_24,
    n1128,
    n1119,
    n1083
  );


  xor
  g1111
  (
    n1137,
    n1120,
    n1119,
    n1082,
    n1126
  );


  or
  g1112
  (
    n1134,
    n1130,
    n1129,
    n1120,
    n1128
  );


  xor
  g1113
  (
    n1139,
    n1120,
    n1123,
    n1122,
    n1121
  );


  xor
  g1114
  (
    n1141,
    n1123,
    n1122,
    n1121
  );


  or
  g1115
  (
    n1142,
    n1121,
    n1122,
    n1137,
    n1125
  );


  xor
  g1116
  (
    n1144,
    n1121,
    n1124,
    n1125
  );


  or
  g1117
  (
    n1140,
    n1123,
    n1134,
    n1125,
    n1133
  );


  nor
  g1118
  (
    n1145,
    n1125,
    n1136,
    n1124,
    n1123
  );


  and
  g1119
  (
    KeyWire_0_60,
    n1135,
    n1132,
    n1138,
    n1124
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n560,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n730,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n262,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n352,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n122,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n613,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1025,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n82,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n593,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n839,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n1083,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n799,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n919,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n367,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n296,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n81,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n246,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n884,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n631,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n568,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n234,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n530,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n591,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n895,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1131,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n407,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n237,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n287,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n536,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n238,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n215,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n230,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n643,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n164,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n851,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n983,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n627,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n926,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n159,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n431,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n642,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n47,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n459,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n827,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n661,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n88,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n314,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n548,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n1103,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n533,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n300,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n1114,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n596,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n86,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n516,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n353,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n830,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n420,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n556,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n739,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n1143,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n712,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n955,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n475,
    KeyNOTWire_0_63
  );


endmodule

