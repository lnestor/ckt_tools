

module Stat_3512_42_5
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n779,
  n796,
  n949,
  n940,
  n945,
  n938,
  n941,
  n947,
  n946,
  n934,
  n943,
  n3543,
  n3546,
  n3544,
  n3541,
  n3547,
  n3542,
  n3545,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n779;output n796;output n949;output n940;output n945;output n938;output n941;output n947;output n946;output n934;output n943;output n3543;output n3546;output n3544;output n3541;output n3547;output n3542;output n3545;
  wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n935;wire n936;wire n937;wire n939;wire n942;wire n944;wire n948;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire n3011;wire n3012;wire n3013;wire n3014;wire n3015;wire n3016;wire n3017;wire n3018;wire n3019;wire n3020;wire n3021;wire n3022;wire n3023;wire n3024;wire n3025;wire n3026;wire n3027;wire n3028;wire n3029;wire n3030;wire n3031;wire n3032;wire n3033;wire n3034;wire n3035;wire n3036;wire n3037;wire n3038;wire n3039;wire n3040;wire n3041;wire n3042;wire n3043;wire n3044;wire n3045;wire n3046;wire n3047;wire n3048;wire n3049;wire n3050;wire n3051;wire n3052;wire n3053;wire n3054;wire n3055;wire n3056;wire n3057;wire n3058;wire n3059;wire n3060;wire n3061;wire n3062;wire n3063;wire n3064;wire n3065;wire n3066;wire n3067;wire n3068;wire n3069;wire n3070;wire n3071;wire n3072;wire n3073;wire n3074;wire n3075;wire n3076;wire n3077;wire n3078;wire n3079;wire n3080;wire n3081;wire n3082;wire n3083;wire n3084;wire n3085;wire n3086;wire n3087;wire n3088;wire n3089;wire n3090;wire n3091;wire n3092;wire n3093;wire n3094;wire n3095;wire n3096;wire n3097;wire n3098;wire n3099;wire n3100;wire n3101;wire n3102;wire n3103;wire n3104;wire n3105;wire n3106;wire n3107;wire n3108;wire n3109;wire n3110;wire n3111;wire n3112;wire n3113;wire n3114;wire n3115;wire n3116;wire n3117;wire n3118;wire n3119;wire n3120;wire n3121;wire n3122;wire n3123;wire n3124;wire n3125;wire n3126;wire n3127;wire n3128;wire n3129;wire n3130;wire n3131;wire n3132;wire n3133;wire n3134;wire n3135;wire n3136;wire n3137;wire n3138;wire n3139;wire n3140;wire n3141;wire n3142;wire n3143;wire n3144;wire n3145;wire n3146;wire n3147;wire n3148;wire n3149;wire n3150;wire n3151;wire n3152;wire n3153;wire n3154;wire n3155;wire n3156;wire n3157;wire n3158;wire n3159;wire n3160;wire n3161;wire n3162;wire n3163;wire n3164;wire n3165;wire n3166;wire n3167;wire n3168;wire n3169;wire n3170;wire n3171;wire n3172;wire n3173;wire n3174;wire n3175;wire n3176;wire n3177;wire n3178;wire n3179;wire n3180;wire n3181;wire n3182;wire n3183;wire n3184;wire n3185;wire n3186;wire n3187;wire n3188;wire n3189;wire n3190;wire n3191;wire n3192;wire n3193;wire n3194;wire n3195;wire n3196;wire n3197;wire n3198;wire n3199;wire n3200;wire n3201;wire n3202;wire n3203;wire n3204;wire n3205;wire n3206;wire n3207;wire n3208;wire n3209;wire n3210;wire n3211;wire n3212;wire n3213;wire n3214;wire n3215;wire n3216;wire n3217;wire n3218;wire n3219;wire n3220;wire n3221;wire n3222;wire n3223;wire n3224;wire n3225;wire n3226;wire n3227;wire n3228;wire n3229;wire n3230;wire n3231;wire n3232;wire n3233;wire n3234;wire n3235;wire n3236;wire n3237;wire n3238;wire n3239;wire n3240;wire n3241;wire n3242;wire n3243;wire n3244;wire n3245;wire n3246;wire n3247;wire n3248;wire n3249;wire n3250;wire n3251;wire n3252;wire n3253;wire n3254;wire n3255;wire n3256;wire n3257;wire n3258;wire n3259;wire n3260;wire n3261;wire n3262;wire n3263;wire n3264;wire n3265;wire n3266;wire n3267;wire n3268;wire n3269;wire n3270;wire n3271;wire n3272;wire n3273;wire n3274;wire n3275;wire n3276;wire n3277;wire n3278;wire n3279;wire n3280;wire n3281;wire n3282;wire n3283;wire n3284;wire n3285;wire n3286;wire n3287;wire n3288;wire n3289;wire n3290;wire n3291;wire n3292;wire n3293;wire n3294;wire n3295;wire n3296;wire n3297;wire n3298;wire n3299;wire n3300;wire n3301;wire n3302;wire n3303;wire n3304;wire n3305;wire n3306;wire n3307;wire n3308;wire n3309;wire n3310;wire n3311;wire n3312;wire n3313;wire n3314;wire n3315;wire n3316;wire n3317;wire n3318;wire n3319;wire n3320;wire n3321;wire n3322;wire n3323;wire n3324;wire n3325;wire n3326;wire n3327;wire n3328;wire n3329;wire n3330;wire n3331;wire n3332;wire n3333;wire n3334;wire n3335;wire n3336;wire n3337;wire n3338;wire n3339;wire n3340;wire n3341;wire n3342;wire n3343;wire n3344;wire n3345;wire n3346;wire n3347;wire n3348;wire n3349;wire n3350;wire n3351;wire n3352;wire n3353;wire n3354;wire n3355;wire n3356;wire n3357;wire n3358;wire n3359;wire n3360;wire n3361;wire n3362;wire n3363;wire n3364;wire n3365;wire n3366;wire n3367;wire n3368;wire n3369;wire n3370;wire n3371;wire n3372;wire n3373;wire n3374;wire n3375;wire n3376;wire n3377;wire n3378;wire n3379;wire n3380;wire n3381;wire n3382;wire n3383;wire n3384;wire n3385;wire n3386;wire n3387;wire n3388;wire n3389;wire n3390;wire n3391;wire n3392;wire n3393;wire n3394;wire n3395;wire n3396;wire n3397;wire n3398;wire n3399;wire n3400;wire n3401;wire n3402;wire n3403;wire n3404;wire n3405;wire n3406;wire n3407;wire n3408;wire n3409;wire n3410;wire n3411;wire n3412;wire n3413;wire n3414;wire n3415;wire n3416;wire n3417;wire n3418;wire n3419;wire n3420;wire n3421;wire n3422;wire n3423;wire n3424;wire n3425;wire n3426;wire n3427;wire n3428;wire n3429;wire n3430;wire n3431;wire n3432;wire n3433;wire n3434;wire n3435;wire n3436;wire n3437;wire n3438;wire n3439;wire n3440;wire n3441;wire n3442;wire n3443;wire n3444;wire n3445;wire n3446;wire n3447;wire n3448;wire n3449;wire n3450;wire n3451;wire n3452;wire n3453;wire n3454;wire n3455;wire n3456;wire n3457;wire n3458;wire n3459;wire n3460;wire n3461;wire n3462;wire n3463;wire n3464;wire n3465;wire n3466;wire n3467;wire n3468;wire n3469;wire n3470;wire n3471;wire n3472;wire n3473;wire n3474;wire n3475;wire n3476;wire n3477;wire n3478;wire n3479;wire n3480;wire n3481;wire n3482;wire n3483;wire n3484;wire n3485;wire n3486;wire n3487;wire n3488;wire n3489;wire n3490;wire n3491;wire n3492;wire n3493;wire n3494;wire n3495;wire n3496;wire n3497;wire n3498;wire n3499;wire n3500;wire n3501;wire n3502;wire n3503;wire n3504;wire n3505;wire n3506;wire n3507;wire n3508;wire n3509;wire n3510;wire n3511;wire n3512;wire n3513;wire n3514;wire n3515;wire n3516;wire n3517;wire n3518;wire n3519;wire n3520;wire n3521;wire n3522;wire n3523;wire n3524;wire n3525;wire n3526;wire n3527;wire n3528;wire n3529;wire n3530;wire n3531;wire n3532;wire n3533;wire n3534;wire n3535;wire n3536;wire n3537;wire n3538;wire n3539;wire n3540;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n52,
    n30
  );


  buf
  g1
  (
    n56,
    n17
  );


  buf
  g2
  (
    n74,
    n18
  );


  buf
  g3
  (
    n143,
    n29
  );


  not
  g4
  (
    n72,
    n10
  );


  buf
  g5
  (
    n60,
    n2
  );


  not
  g6
  (
    n57,
    n26
  );


  not
  g7
  (
    n123,
    n32
  );


  buf
  g8
  (
    n78,
    n21
  );


  buf
  g9
  (
    n163,
    n19
  );


  not
  g10
  (
    n101,
    n20
  );


  not
  g11
  (
    n133,
    n31
  );


  buf
  g12
  (
    n140,
    n31
  );


  buf
  g13
  (
    n112,
    n16
  );


  not
  g14
  (
    n50,
    n11
  );


  buf
  g15
  (
    n145,
    n1
  );


  not
  g16
  (
    n142,
    n7
  );


  not
  g17
  (
    n161,
    n7
  );


  buf
  g18
  (
    n164,
    n32
  );


  buf
  g19
  (
    n68,
    n9
  );


  not
  g20
  (
    n95,
    n1
  );


  buf
  g21
  (
    n90,
    n11
  );


  buf
  g22
  (
    n137,
    n24
  );


  not
  g23
  (
    n171,
    n26
  );


  not
  g24
  (
    n138,
    n23
  );


  buf
  g25
  (
    n41,
    n4
  );


  buf
  g26
  (
    n169,
    n10
  );


  buf
  g27
  (
    n126,
    n35
  );


  not
  g28
  (
    n38,
    n6
  );


  buf
  g29
  (
    n61,
    n7
  );


  not
  g30
  (
    n122,
    n21
  );


  not
  g31
  (
    n108,
    n18
  );


  buf
  g32
  (
    n160,
    n13
  );


  not
  g33
  (
    n144,
    n14
  );


  not
  g34
  (
    n81,
    n20
  );


  buf
  g35
  (
    n59,
    n33
  );


  not
  g36
  (
    n152,
    n32
  );


  buf
  g37
  (
    n106,
    n18
  );


  buf
  g38
  (
    n149,
    n13
  );


  not
  g39
  (
    n127,
    n6
  );


  buf
  g40
  (
    n135,
    n29
  );


  not
  g41
  (
    n54,
    n17
  );


  buf
  g42
  (
    n116,
    n1
  );


  buf
  g43
  (
    n173,
    n30
  );


  not
  g44
  (
    n139,
    n5
  );


  not
  g45
  (
    n45,
    n15
  );


  buf
  g46
  (
    n113,
    n9
  );


  buf
  g47
  (
    n55,
    n29
  );


  buf
  g48
  (
    n159,
    n16
  );


  buf
  g49
  (
    n174,
    n35
  );


  buf
  g50
  (
    n44,
    n34
  );


  not
  g51
  (
    n51,
    n6
  );


  buf
  g52
  (
    n94,
    n24
  );


  not
  g53
  (
    n79,
    n12
  );


  not
  g54
  (
    n53,
    n30
  );


  buf
  g55
  (
    n166,
    n19
  );


  buf
  g56
  (
    n70,
    n23
  );


  buf
  g57
  (
    n80,
    n12
  );


  not
  g58
  (
    n100,
    n34
  );


  buf
  g59
  (
    n46,
    n29
  );


  buf
  g60
  (
    n65,
    n2
  );


  buf
  g61
  (
    n40,
    n22
  );


  not
  g62
  (
    n75,
    n18
  );


  not
  g63
  (
    n119,
    n4
  );


  buf
  g64
  (
    n47,
    n6
  );


  buf
  g65
  (
    n162,
    n14
  );


  buf
  g66
  (
    n141,
    n9
  );


  not
  g67
  (
    n157,
    n24
  );


  buf
  g68
  (
    n49,
    n22
  );


  buf
  g69
  (
    n124,
    n28
  );


  buf
  g70
  (
    n89,
    n13
  );


  buf
  g71
  (
    n110,
    n3
  );


  buf
  g72
  (
    n87,
    n20
  );


  buf
  g73
  (
    n132,
    n8
  );


  not
  g74
  (
    n58,
    n1
  );


  buf
  g75
  (
    n73,
    n14
  );


  buf
  g76
  (
    n129,
    n3
  );


  not
  g77
  (
    n62,
    n24
  );


  buf
  g78
  (
    n84,
    n13
  );


  not
  g79
  (
    n158,
    n28
  );


  not
  g80
  (
    n118,
    n9
  );


  buf
  g81
  (
    n48,
    n8
  );


  not
  g82
  (
    n86,
    n34
  );


  not
  g83
  (
    n114,
    n26
  );


  buf
  g84
  (
    n130,
    n21
  );


  not
  g85
  (
    n105,
    n15
  );


  buf
  g86
  (
    n102,
    n2
  );


  buf
  g87
  (
    n39,
    n15
  );


  buf
  g88
  (
    n170,
    n30
  );


  not
  g89
  (
    n150,
    n12
  );


  buf
  g90
  (
    n134,
    n31
  );


  not
  g91
  (
    n109,
    n10
  );


  buf
  g92
  (
    n64,
    n27
  );


  buf
  g93
  (
    n77,
    n16
  );


  not
  g94
  (
    n153,
    n2
  );


  not
  g95
  (
    n168,
    n5
  );


  buf
  g96
  (
    n63,
    n19
  );


  buf
  g97
  (
    n128,
    n27
  );


  not
  g98
  (
    n67,
    n25
  );


  not
  g99
  (
    n131,
    n27
  );


  not
  g100
  (
    n93,
    n22
  );


  buf
  g101
  (
    n103,
    n25
  );


  buf
  g102
  (
    n97,
    n10
  );


  buf
  g103
  (
    n172,
    n28
  );


  not
  g104
  (
    n111,
    n17
  );


  buf
  g105
  (
    n92,
    n5
  );


  not
  g106
  (
    n121,
    n21
  );


  not
  g107
  (
    n156,
    n20
  );


  not
  g108
  (
    n136,
    n26
  );


  not
  g109
  (
    n98,
    n32
  );


  not
  g110
  (
    n165,
    n23
  );


  buf
  g111
  (
    n107,
    n8
  );


  not
  g112
  (
    n71,
    n14
  );


  not
  g113
  (
    n125,
    n7
  );


  not
  g114
  (
    n115,
    n19
  );


  buf
  g115
  (
    n42,
    n25
  );


  buf
  g116
  (
    n147,
    n34
  );


  buf
  g117
  (
    n175,
    n12
  );


  buf
  g118
  (
    n88,
    n25
  );


  not
  g119
  (
    n85,
    n15
  );


  not
  g120
  (
    n104,
    n23
  );


  not
  g121
  (
    n120,
    n17
  );


  buf
  g122
  (
    n99,
    n33
  );


  buf
  g123
  (
    n155,
    n22
  );


  buf
  g124
  (
    n91,
    n8
  );


  buf
  g125
  (
    n66,
    n11
  );


  not
  g126
  (
    n83,
    n33
  );


  not
  g127
  (
    n37,
    n31
  );


  buf
  g128
  (
    n151,
    n28
  );


  buf
  g129
  (
    n43,
    n35
  );


  buf
  g130
  (
    n76,
    n27
  );


  not
  g131
  (
    n117,
    n4
  );


  buf
  g132
  (
    n82,
    n11
  );


  buf
  g133
  (
    n146,
    n5
  );


  buf
  g134
  (
    n36,
    n3
  );


  buf
  g135
  (
    n96,
    n35
  );


  buf
  g136
  (
    n167,
    n4
  );


  buf
  g137
  (
    n154,
    n16
  );


  not
  g138
  (
    n148,
    n33
  );


  buf
  g139
  (
    n69,
    n3
  );


  buf
  g140
  (
    n406,
    n145
  );


  not
  g141
  (
    n249,
    n106
  );


  not
  g142
  (
    n660,
    n134
  );


  not
  g143
  (
    n624,
    n160
  );


  buf
  g144
  (
    n394,
    n65
  );


  not
  g145
  (
    n191,
    n110
  );


  buf
  g146
  (
    n392,
    n143
  );


  buf
  g147
  (
    n314,
    n81
  );


  buf
  g148
  (
    n450,
    n142
  );


  not
  g149
  (
    n488,
    n119
  );


  buf
  g150
  (
    n486,
    n51
  );


  buf
  g151
  (
    n310,
    n133
  );


  buf
  g152
  (
    n495,
    n121
  );


  not
  g153
  (
    n319,
    n124
  );


  buf
  g154
  (
    n227,
    n171
  );


  buf
  g155
  (
    n557,
    n164
  );


  buf
  g156
  (
    n251,
    n38
  );


  buf
  g157
  (
    n533,
    n113
  );


  buf
  g158
  (
    n590,
    n50
  );


  not
  g159
  (
    n492,
    n54
  );


  buf
  g160
  (
    n320,
    n115
  );


  buf
  g161
  (
    n291,
    n75
  );


  not
  g162
  (
    n252,
    n57
  );


  buf
  g163
  (
    n654,
    n84
  );


  buf
  g164
  (
    n321,
    n73
  );


  not
  g165
  (
    n532,
    n77
  );


  buf
  g166
  (
    n703,
    n130
  );


  not
  g167
  (
    n579,
    n82
  );


  buf
  g168
  (
    n403,
    n64
  );


  not
  g169
  (
    n538,
    n158
  );


  buf
  g170
  (
    n539,
    n72
  );


  not
  g171
  (
    n339,
    n116
  );


  buf
  g172
  (
    n678,
    n105
  );


  not
  g173
  (
    n199,
    n133
  );


  not
  g174
  (
    n513,
    n171
  );


  buf
  g175
  (
    n286,
    n142
  );


  not
  g176
  (
    n720,
    n165
  );


  not
  g177
  (
    n418,
    n54
  );


  buf
  g178
  (
    n573,
    n74
  );


  buf
  g179
  (
    n574,
    n151
  );


  not
  g180
  (
    n243,
    n77
  );


  not
  g181
  (
    n679,
    n78
  );


  not
  g182
  (
    n411,
    n105
  );


  buf
  g183
  (
    n299,
    n157
  );


  buf
  g184
  (
    n652,
    n97
  );


  buf
  g185
  (
    n318,
    n139
  );


  buf
  g186
  (
    n276,
    n85
  );


  buf
  g187
  (
    n494,
    n57
  );


  buf
  g188
  (
    n201,
    n106
  );


  not
  g189
  (
    n666,
    n88
  );


  not
  g190
  (
    n663,
    n111
  );


  buf
  g191
  (
    n448,
    n90
  );


  not
  g192
  (
    n307,
    n88
  );


  not
  g193
  (
    n689,
    n70
  );


  not
  g194
  (
    n472,
    n59
  );


  buf
  g195
  (
    n219,
    n161
  );


  not
  g196
  (
    n331,
    n159
  );


  buf
  g197
  (
    n504,
    n118
  );


  not
  g198
  (
    n537,
    n49
  );


  not
  g199
  (
    n554,
    n131
  );


  not
  g200
  (
    n675,
    n116
  );


  not
  g201
  (
    n717,
    n56
  );


  buf
  g202
  (
    n711,
    n59
  );


  buf
  g203
  (
    n522,
    n39
  );


  not
  g204
  (
    n461,
    n121
  );


  not
  g205
  (
    n715,
    n121
  );


  not
  g206
  (
    n563,
    n42
  );


  not
  g207
  (
    n233,
    n141
  );


  not
  g208
  (
    n503,
    n103
  );


  not
  g209
  (
    n226,
    n50
  );


  buf
  g210
  (
    n306,
    n54
  );


  not
  g211
  (
    n259,
    n149
  );


  buf
  g212
  (
    n655,
    n110
  );


  buf
  g213
  (
    n343,
    n97
  );


  not
  g214
  (
    n214,
    n40
  );


  buf
  g215
  (
    n681,
    n58
  );


  not
  g216
  (
    n561,
    n132
  );


  buf
  g217
  (
    n661,
    n42
  );


  buf
  g218
  (
    n628,
    n162
  );


  buf
  g219
  (
    n673,
    n146
  );


  buf
  g220
  (
    n351,
    n84
  );


  not
  g221
  (
    n302,
    n130
  );


  buf
  g222
  (
    n519,
    n53
  );


  buf
  g223
  (
    n440,
    n149
  );


  buf
  g224
  (
    n405,
    n112
  );


  not
  g225
  (
    n723,
    n172
  );


  not
  g226
  (
    n308,
    n120
  );


  buf
  g227
  (
    n433,
    n65
  );


  not
  g228
  (
    n386,
    n163
  );


  not
  g229
  (
    n508,
    n44
  );


  not
  g230
  (
    n580,
    n98
  );


  buf
  g231
  (
    n208,
    n45
  );


  buf
  g232
  (
    n225,
    n116
  );


  buf
  g233
  (
    n360,
    n153
  );


  buf
  g234
  (
    n721,
    n56
  );


  not
  g235
  (
    n650,
    n86
  );


  buf
  g236
  (
    n460,
    n83
  );


  buf
  g237
  (
    n281,
    n110
  );


  buf
  g238
  (
    n415,
    n82
  );


  not
  g239
  (
    n551,
    n132
  );


  not
  g240
  (
    n707,
    n84
  );


  buf
  g241
  (
    n667,
    n170
  );


  buf
  g242
  (
    n190,
    n47
  );


  buf
  g243
  (
    n327,
    n127
  );


  buf
  g244
  (
    n204,
    n90
  );


  not
  g245
  (
    n582,
    n159
  );


  buf
  g246
  (
    n454,
    n169
  );


  buf
  g247
  (
    n328,
    n148
  );


  buf
  g248
  (
    n670,
    n168
  );


  buf
  g249
  (
    n512,
    n128
  );


  not
  g250
  (
    n569,
    n153
  );


  not
  g251
  (
    n303,
    n74
  );


  buf
  g252
  (
    n184,
    n46
  );


  not
  g253
  (
    n410,
    n138
  );


  buf
  g254
  (
    n435,
    n109
  );


  not
  g255
  (
    n188,
    n139
  );


  buf
  g256
  (
    n490,
    n138
  );


  not
  g257
  (
    n627,
    n147
  );


  buf
  g258
  (
    n271,
    n147
  );


  not
  g259
  (
    n591,
    n71
  );


  not
  g260
  (
    n357,
    n165
  );


  buf
  g261
  (
    n336,
    n43
  );


  not
  g262
  (
    n546,
    n38
  );


  not
  g263
  (
    n297,
    n83
  );


  buf
  g264
  (
    n217,
    n95
  );


  buf
  g265
  (
    n457,
    n53
  );


  buf
  g266
  (
    n425,
    n136
  );


  not
  g267
  (
    n366,
    n130
  );


  not
  g268
  (
    n431,
    n72
  );


  not
  g269
  (
    n282,
    n102
  );


  not
  g270
  (
    n547,
    n87
  );


  buf
  g271
  (
    n260,
    n159
  );


  not
  g272
  (
    n672,
    n141
  );


  buf
  g273
  (
    n493,
    n113
  );


  buf
  g274
  (
    n189,
    n68
  );


  not
  g275
  (
    n211,
    n80
  );


  buf
  g276
  (
    n255,
    n39
  );


  buf
  g277
  (
    n378,
    n91
  );


  buf
  g278
  (
    n657,
    n166
  );


  buf
  g279
  (
    n706,
    n47
  );


  buf
  g280
  (
    n633,
    n114
  );


  not
  g281
  (
    n467,
    n37
  );


  not
  g282
  (
    n432,
    n168
  );


  not
  g283
  (
    n334,
    n128
  );


  buf
  g284
  (
    n589,
    n79
  );


  not
  g285
  (
    n640,
    n86
  );


  not
  g286
  (
    n423,
    n36
  );


  buf
  g287
  (
    n617,
    n145
  );


  not
  g288
  (
    n210,
    n133
  );


  not
  g289
  (
    n384,
    n62
  );


  buf
  g290
  (
    n412,
    n96
  );


  not
  g291
  (
    n629,
    n65
  );


  buf
  g292
  (
    n258,
    n164
  );


  not
  g293
  (
    n498,
    n111
  );


  not
  g294
  (
    n604,
    n122
  );


  buf
  g295
  (
    n453,
    n90
  );


  not
  g296
  (
    n383,
    n43
  );


  buf
  g297
  (
    n593,
    n134
  );


  buf
  g298
  (
    n434,
    n50
  );


  buf
  g299
  (
    n581,
    n97
  );


  buf
  g300
  (
    n480,
    n77
  );


  not
  g301
  (
    n525,
    n101
  );


  buf
  g302
  (
    n283,
    n102
  );


  buf
  g303
  (
    n602,
    n115
  );


  buf
  g304
  (
    n216,
    n59
  );


  not
  g305
  (
    n280,
    n125
  );


  not
  g306
  (
    n585,
    n137
  );


  buf
  g307
  (
    n583,
    n160
  );


  not
  g308
  (
    n300,
    n50
  );


  buf
  g309
  (
    n441,
    n136
  );


  buf
  g310
  (
    n228,
    n120
  );


  not
  g311
  (
    n301,
    n117
  );


  not
  g312
  (
    n407,
    n149
  );


  buf
  g313
  (
    n342,
    n86
  );


  buf
  g314
  (
    n674,
    n131
  );


  buf
  g315
  (
    n177,
    n157
  );


  buf
  g316
  (
    n474,
    n170
  );


  buf
  g317
  (
    n608,
    n71
  );


  not
  g318
  (
    n716,
    n93
  );


  buf
  g319
  (
    n240,
    n155
  );


  buf
  g320
  (
    n263,
    n40
  );


  buf
  g321
  (
    n618,
    n154
  );


  not
  g322
  (
    n196,
    n38
  );


  not
  g323
  (
    n298,
    n103
  );


  buf
  g324
  (
    n489,
    n127
  );


  not
  g325
  (
    n659,
    n98
  );


  buf
  g326
  (
    n375,
    n113
  );


  buf
  g327
  (
    n344,
    n104
  );


  buf
  g328
  (
    n700,
    n156
  );


  buf
  g329
  (
    n183,
    n129
  );


  buf
  g330
  (
    n195,
    n78
  );


  not
  g331
  (
    n267,
    n127
  );


  buf
  g332
  (
    n718,
    n112
  );


  buf
  g333
  (
    n290,
    n170
  );


  not
  g334
  (
    n468,
    n80
  );


  not
  g335
  (
    n595,
    n155
  );


  not
  g336
  (
    n288,
    n41
  );


  buf
  g337
  (
    n178,
    n52
  );


  buf
  g338
  (
    n612,
    n119
  );


  not
  g339
  (
    n324,
    n47
  );


  buf
  g340
  (
    n680,
    n41
  );


  buf
  g341
  (
    n284,
    n62
  );


  not
  g342
  (
    n649,
    n66
  );


  buf
  g343
  (
    n295,
    n142
  );


  not
  g344
  (
    n197,
    n44
  );


  buf
  g345
  (
    n400,
    n162
  );


  buf
  g346
  (
    n364,
    n88
  );


  not
  g347
  (
    n540,
    n37
  );


  not
  g348
  (
    n443,
    n153
  );


  buf
  g349
  (
    n510,
    n152
  );


  buf
  g350
  (
    n568,
    n89
  );


  not
  g351
  (
    n352,
    n166
  );


  not
  g352
  (
    n428,
    n129
  );


  not
  g353
  (
    n577,
    n140
  );


  not
  g354
  (
    n662,
    n46
  );


  buf
  g355
  (
    n322,
    n66
  );


  not
  g356
  (
    n279,
    n126
  );


  buf
  g357
  (
    n714,
    n127
  );


  buf
  g358
  (
    n424,
    n136
  );


  buf
  g359
  (
    n213,
    n102
  );


  buf
  g360
  (
    n393,
    n135
  );


  not
  g361
  (
    n576,
    n143
  );


  buf
  g362
  (
    n187,
    n112
  );


  not
  g363
  (
    n545,
    n125
  );


  buf
  g364
  (
    n241,
    n79
  );


  buf
  g365
  (
    n239,
    n165
  );


  buf
  g366
  (
    n359,
    n74
  );


  buf
  g367
  (
    n311,
    n154
  );


  buf
  g368
  (
    n683,
    n55
  );


  buf
  g369
  (
    n684,
    n102
  );


  buf
  g370
  (
    n549,
    n117
  );


  not
  g371
  (
    n611,
    n90
  );


  buf
  g372
  (
    n382,
    n77
  );


  not
  g373
  (
    n520,
    n60
  );


  buf
  g374
  (
    n610,
    n39
  );


  not
  g375
  (
    n592,
    n59
  );


  buf
  g376
  (
    n643,
    n98
  );


  not
  g377
  (
    n194,
    n128
  );


  not
  g378
  (
    n558,
    n117
  );


  not
  g379
  (
    n523,
    n85
  );


  buf
  g380
  (
    n264,
    n95
  );


  not
  g381
  (
    n698,
    n70
  );


  not
  g382
  (
    n388,
    n72
  );


  not
  g383
  (
    n570,
    n123
  );


  buf
  g384
  (
    n636,
    n65
  );


  not
  g385
  (
    n456,
    n100
  );


  not
  g386
  (
    n401,
    n99
  );


  not
  g387
  (
    n245,
    n148
  );


  buf
  g388
  (
    n621,
    n94
  );


  not
  g389
  (
    n565,
    n49
  );


  buf
  g390
  (
    n292,
    n100
  );


  not
  g391
  (
    n373,
    n150
  );


  not
  g392
  (
    n598,
    n100
  );


  not
  g393
  (
    n452,
    n68
  );


  buf
  g394
  (
    n552,
    n132
  );


  buf
  g395
  (
    n349,
    n140
  );


  not
  g396
  (
    n597,
    n46
  );


  not
  g397
  (
    n497,
    n64
  );


  not
  g398
  (
    n505,
    n71
  );


  buf
  g399
  (
    n413,
    n53
  );


  buf
  g400
  (
    n614,
    n104
  );


  not
  g401
  (
    n417,
    n135
  );


  not
  g402
  (
    n230,
    n122
  );


  not
  g403
  (
    n688,
    n62
  );


  not
  g404
  (
    n466,
    n61
  );


  not
  g405
  (
    n555,
    n73
  );


  buf
  g406
  (
    n398,
    n57
  );


  not
  g407
  (
    n571,
    n134
  );


  not
  g408
  (
    n690,
    n93
  );


  not
  g409
  (
    n556,
    n44
  );


  not
  g410
  (
    n390,
    n158
  );


  not
  g411
  (
    n202,
    n48
  );


  buf
  g412
  (
    n644,
    n101
  );


  not
  g413
  (
    n603,
    n78
  );


  not
  g414
  (
    n222,
    n68
  );


  not
  g415
  (
    n514,
    n141
  );


  not
  g416
  (
    n346,
    n152
  );


  not
  g417
  (
    n309,
    n58
  );


  not
  g418
  (
    n528,
    n144
  );


  not
  g419
  (
    n368,
    n107
  );


  not
  g420
  (
    n600,
    n86
  );


  buf
  g421
  (
    n181,
    n139
  );


  not
  g422
  (
    n693,
    n37
  );


  buf
  g423
  (
    n250,
    n104
  );


  not
  g424
  (
    n442,
    n165
  );


  not
  g425
  (
    n518,
    n64
  );


  buf
  g426
  (
    KeyWire_0_10,
    n52
  );


  not
  g427
  (
    n491,
    n108
  );


  buf
  g428
  (
    n594,
    n43
  );


  not
  g429
  (
    n408,
    n164
  );


  not
  g430
  (
    n658,
    n63
  );


  not
  g431
  (
    n507,
    n107
  );


  buf
  g432
  (
    n370,
    n154
  );


  buf
  g433
  (
    n399,
    n76
  );


  not
  g434
  (
    n362,
    n129
  );


  buf
  g435
  (
    n464,
    n172
  );


  buf
  g436
  (
    n502,
    n87
  );


  not
  g437
  (
    n316,
    n135
  );


  buf
  g438
  (
    n664,
    n170
  );


  not
  g439
  (
    n395,
    n144
  );


  buf
  g440
  (
    n587,
    n81
  );


  buf
  g441
  (
    n607,
    n145
  );


  not
  g442
  (
    n444,
    n76
  );


  not
  g443
  (
    n526,
    n161
  );


  buf
  g444
  (
    n176,
    n67
  );


  not
  g445
  (
    n478,
    n41
  );


  not
  g446
  (
    n462,
    n36
  );


  not
  g447
  (
    n548,
    n81
  );


  not
  g448
  (
    n256,
    n151
  );


  buf
  g449
  (
    n285,
    n150
  );


  not
  g450
  (
    n377,
    n56
  );


  buf
  g451
  (
    n686,
    n52
  );


  not
  g452
  (
    n294,
    n71
  );


  not
  g453
  (
    n416,
    n122
  );


  buf
  g454
  (
    n358,
    n131
  );


  buf
  g455
  (
    n606,
    n80
  );


  not
  g456
  (
    n235,
    n109
  );


  buf
  g457
  (
    n185,
    n108
  );


  not
  g458
  (
    n638,
    n146
  );


  buf
  g459
  (
    n631,
    n123
  );


  not
  g460
  (
    n315,
    n133
  );


  buf
  g461
  (
    n430,
    n79
  );


  buf
  g462
  (
    n380,
    n58
  );


  not
  g463
  (
    n348,
    n101
  );


  not
  g464
  (
    n304,
    n141
  );


  not
  g465
  (
    n634,
    n75
  );


  buf
  g466
  (
    n332,
    n83
  );


  not
  g467
  (
    n685,
    n94
  );


  buf
  g468
  (
    n708,
    n36
  );


  buf
  g469
  (
    n374,
    n66
  );


  buf
  g470
  (
    n365,
    n113
  );


  buf
  g471
  (
    n566,
    n156
  );


  not
  g472
  (
    n429,
    n152
  );


  not
  g473
  (
    n317,
    n91
  );


  buf
  g474
  (
    n553,
    n69
  );


  not
  g475
  (
    n699,
    n115
  );


  buf
  g476
  (
    n426,
    n92
  );


  not
  g477
  (
    n458,
    n150
  );


  not
  g478
  (
    n312,
    n111
  );


  not
  g479
  (
    n275,
    n128
  );


  not
  g480
  (
    n355,
    n130
  );


  not
  g481
  (
    n653,
    n48
  );


  buf
  g482
  (
    n268,
    n119
  );


  not
  g483
  (
    n330,
    n111
  );


  buf
  g484
  (
    n500,
    n163
  );


  not
  g485
  (
    n427,
    n137
  );


  buf
  g486
  (
    n381,
    n53
  );


  not
  g487
  (
    n209,
    n73
  );


  buf
  g488
  (
    n712,
    n122
  );


  buf
  g489
  (
    n620,
    n114
  );


  not
  g490
  (
    n623,
    n60
  );


  not
  g491
  (
    n182,
    n75
  );


  not
  g492
  (
    n709,
    n124
  );


  buf
  g493
  (
    n677,
    n76
  );


  buf
  g494
  (
    n445,
    n103
  );


  not
  g495
  (
    KeyWire_0_19,
    n151
  );


  not
  g496
  (
    n449,
    n49
  );


  not
  g497
  (
    n626,
    n67
  );


  buf
  g498
  (
    n536,
    n36
  );


  buf
  g499
  (
    n361,
    n146
  );


  not
  g500
  (
    n527,
    n63
  );


  buf
  g501
  (
    n578,
    n158
  );


  buf
  g502
  (
    n261,
    n60
  );


  buf
  g503
  (
    n630,
    n136
  );


  buf
  g504
  (
    n421,
    n162
  );


  buf
  g505
  (
    n385,
    n57
  );


  buf
  g506
  (
    n722,
    n168
  );


  buf
  g507
  (
    n220,
    n92
  );


  not
  g508
  (
    n326,
    n61
  );


  buf
  g509
  (
    n534,
    n166
  );


  not
  g510
  (
    n616,
    n154
  );


  buf
  g511
  (
    n323,
    n48
  );


  not
  g512
  (
    n371,
    n89
  );


  buf
  g513
  (
    n272,
    n108
  );


  buf
  g514
  (
    n476,
    n109
  );


  not
  g515
  (
    n719,
    n69
  );


  buf
  g516
  (
    n710,
    n157
  );


  buf
  g517
  (
    n237,
    n151
  );


  not
  g518
  (
    n588,
    n37
  );


  not
  g519
  (
    n645,
    n73
  );


  buf
  g520
  (
    n637,
    n88
  );


  not
  g521
  (
    n193,
    n124
  );


  buf
  g522
  (
    n704,
    n96
  );


  not
  g523
  (
    n186,
    n169
  );


  buf
  g524
  (
    n584,
    n156
  );


  buf
  g525
  (
    n236,
    n126
  );


  not
  g526
  (
    n287,
    n55
  );


  not
  g527
  (
    n257,
    n120
  );


  not
  g528
  (
    n363,
    n143
  );


  buf
  g529
  (
    n482,
    n172
  );


  buf
  g530
  (
    n234,
    n95
  );


  buf
  g531
  (
    n572,
    n85
  );


  buf
  g532
  (
    n379,
    n41
  );


  not
  g533
  (
    n487,
    n40
  );


  buf
  g534
  (
    n671,
    n148
  );


  not
  g535
  (
    n596,
    n56
  );


  not
  g536
  (
    n376,
    n171
  );


  buf
  g537
  (
    n437,
    n156
  );


  buf
  g538
  (
    n296,
    n100
  );


  not
  g539
  (
    n560,
    n125
  );


  buf
  g540
  (
    n496,
    n120
  );


  buf
  g541
  (
    n419,
    n42
  );


  not
  g542
  (
    n529,
    n82
  );


  not
  g543
  (
    n389,
    n60
  );


  buf
  g544
  (
    n481,
    n138
  );


  not
  g545
  (
    n516,
    n172
  );


  buf
  g546
  (
    n479,
    n47
  );


  not
  g547
  (
    n229,
    n91
  );


  buf
  g548
  (
    n485,
    n153
  );


  buf
  g549
  (
    n397,
    n97
  );


  not
  g550
  (
    n223,
    n103
  );


  not
  g551
  (
    n273,
    n74
  );


  buf
  g552
  (
    n337,
    n79
  );


  not
  g553
  (
    n483,
    n159
  );


  buf
  g554
  (
    n278,
    n38
  );


  not
  g555
  (
    n696,
    n81
  );


  not
  g556
  (
    n289,
    n66
  );


  buf
  g557
  (
    n648,
    n58
  );


  not
  g558
  (
    n499,
    n119
  );


  not
  g559
  (
    n509,
    n166
  );


  not
  g560
  (
    n248,
    n94
  );


  not
  g561
  (
    n218,
    n62
  );


  not
  g562
  (
    n391,
    n123
  );


  not
  g563
  (
    n446,
    n54
  );


  not
  g564
  (
    n484,
    n80
  );


  not
  g565
  (
    n609,
    n139
  );


  buf
  g566
  (
    n207,
    n157
  );


  not
  g567
  (
    n369,
    n96
  );


  buf
  g568
  (
    n501,
    n99
  );


  not
  g569
  (
    n586,
    n42
  );


  buf
  g570
  (
    n459,
    n67
  );


  buf
  g571
  (
    n224,
    n72
  );


  buf
  g572
  (
    n697,
    n163
  );


  not
  g573
  (
    n463,
    n126
  );


  buf
  g574
  (
    n713,
    n149
  );


  not
  g575
  (
    n646,
    n142
  );


  not
  g576
  (
    n269,
    n64
  );


  buf
  g577
  (
    n447,
    n162
  );


  not
  g578
  (
    n451,
    n39
  );


  not
  g579
  (
    n203,
    n98
  );


  not
  g580
  (
    n682,
    n51
  );


  buf
  g581
  (
    n262,
    n158
  );


  buf
  g582
  (
    n402,
    n105
  );


  buf
  g583
  (
    n215,
    n105
  );


  buf
  g584
  (
    n562,
    n101
  );


  not
  g585
  (
    n277,
    n123
  );


  not
  g586
  (
    n477,
    n84
  );


  not
  g587
  (
    n635,
    n44
  );


  not
  g588
  (
    n438,
    n45
  );


  buf
  g589
  (
    n254,
    n160
  );


  buf
  g590
  (
    n266,
    n144
  );


  buf
  g591
  (
    n619,
    n78
  );


  buf
  g592
  (
    n232,
    n92
  );


  buf
  g593
  (
    n656,
    n146
  );


  not
  g594
  (
    n615,
    n129
  );


  buf
  g595
  (
    n613,
    n85
  );


  not
  g596
  (
    n541,
    n48
  );


  not
  g597
  (
    n641,
    n115
  );


  not
  g598
  (
    n471,
    n106
  );


  not
  g599
  (
    n270,
    n94
  );


  buf
  g600
  (
    n694,
    n55
  );


  buf
  g601
  (
    n205,
    n148
  );


  not
  g602
  (
    n559,
    n110
  );


  buf
  g603
  (
    n511,
    n45
  );


  not
  g604
  (
    n246,
    n135
  );


  not
  g605
  (
    n473,
    n124
  );


  buf
  g606
  (
    n198,
    n46
  );


  not
  g607
  (
    n550,
    n125
  );


  buf
  g608
  (
    n347,
    n40
  );


  buf
  g609
  (
    n543,
    n61
  );


  buf
  g610
  (
    n702,
    n83
  );


  not
  g611
  (
    n535,
    n109
  );


  buf
  g612
  (
    n691,
    n131
  );


  buf
  g613
  (
    n354,
    n155
  );


  not
  g614
  (
    n325,
    n114
  );


  buf
  g615
  (
    n305,
    n160
  );


  not
  g616
  (
    n564,
    n167
  );


  not
  g617
  (
    n345,
    n169
  );


  not
  g618
  (
    n221,
    n167
  );


  buf
  g619
  (
    n231,
    n171
  );


  not
  g620
  (
    n639,
    n137
  );


  not
  g621
  (
    n524,
    n107
  );


  not
  g622
  (
    n530,
    n137
  );


  buf
  g623
  (
    n335,
    n118
  );


  buf
  g624
  (
    n387,
    n99
  );


  not
  g625
  (
    n192,
    n161
  );


  not
  g626
  (
    n506,
    n95
  );


  buf
  g627
  (
    n180,
    n126
  );


  buf
  g628
  (
    n701,
    n76
  );


  not
  g629
  (
    n353,
    n43
  );


  not
  g630
  (
    n599,
    n114
  );


  buf
  g631
  (
    n206,
    n93
  );


  not
  g632
  (
    n293,
    n168
  );


  not
  g633
  (
    n341,
    n118
  );


  buf
  g634
  (
    n313,
    n147
  );


  buf
  g635
  (
    n521,
    n52
  );


  buf
  g636
  (
    n244,
    n106
  );


  buf
  g637
  (
    n542,
    n145
  );


  buf
  g638
  (
    n265,
    n87
  );


  buf
  g639
  (
    n338,
    n51
  );


  buf
  g640
  (
    n469,
    n155
  );


  not
  g641
  (
    n531,
    n82
  );


  buf
  g642
  (
    n647,
    n167
  );


  buf
  g643
  (
    n179,
    n75
  );


  buf
  g644
  (
    n372,
    n143
  );


  not
  g645
  (
    n515,
    n147
  );


  not
  g646
  (
    n356,
    n150
  );


  not
  g647
  (
    n695,
    n152
  );


  not
  g648
  (
    n575,
    n70
  );


  not
  g649
  (
    n692,
    n91
  );


  not
  g650
  (
    n420,
    n118
  );


  not
  g651
  (
    n396,
    n68
  );


  buf
  g652
  (
    n455,
    n112
  );


  buf
  g653
  (
    n622,
    n89
  );


  buf
  g654
  (
    n651,
    n163
  );


  buf
  g655
  (
    n567,
    n140
  );


  not
  g656
  (
    n668,
    n51
  );


  not
  g657
  (
    n642,
    n121
  );


  buf
  g658
  (
    n422,
    n164
  );


  buf
  g659
  (
    n238,
    n96
  );


  buf
  g660
  (
    n436,
    n69
  );


  buf
  g661
  (
    n669,
    n63
  );


  buf
  g662
  (
    n517,
    n107
  );


  buf
  g663
  (
    n367,
    n49
  );


  not
  g664
  (
    n439,
    n63
  );


  not
  g665
  (
    n404,
    n116
  );


  not
  g666
  (
    n605,
    n104
  );


  buf
  g667
  (
    n465,
    n169
  );


  buf
  g668
  (
    n475,
    n70
  );


  buf
  g669
  (
    n676,
    n161
  );


  buf
  g670
  (
    n665,
    n140
  );


  buf
  g671
  (
    n632,
    n144
  );


  not
  g672
  (
    n409,
    n134
  );


  not
  g673
  (
    n705,
    n45
  );


  not
  g674
  (
    n470,
    n69
  );


  buf
  g675
  (
    n274,
    n108
  );


  not
  g676
  (
    n212,
    n92
  );


  not
  g677
  (
    n601,
    n99
  );


  buf
  g678
  (
    n333,
    n55
  );


  buf
  g679
  (
    n253,
    n89
  );


  not
  g680
  (
    n687,
    n138
  );


  not
  g681
  (
    n200,
    n93
  );


  buf
  g682
  (
    n625,
    n61
  );


  not
  g683
  (
    n329,
    n87
  );


  buf
  g684
  (
    n414,
    n132
  );


  not
  g685
  (
    n242,
    n67
  );


  buf
  g686
  (
    n247,
    n117
  );


  buf
  g687
  (
    n340,
    n167
  );


  buf
  g688
  (
    n725,
    n177
  );


  not
  g689
  (
    n724,
    n176
  );


  nand
  g690
  (
    n726,
    n725,
    n724
  );


  nand
  g691
  (
    n727,
    n178,
    n726
  );


  buf
  g692
  (
    n730,
    n727
  );


  buf
  g693
  (
    n731,
    n727
  );


  buf
  g694
  (
    n728,
    n727
  );


  buf
  g695
  (
    n729,
    n727
  );


  buf
  g696
  (
    n737,
    n730
  );


  not
  g697
  (
    n736,
    n730
  );


  not
  g698
  (
    n732,
    n731
  );


  buf
  g699
  (
    n733,
    n179
  );


  buf
  g700
  (
    n734,
    n731
  );


  not
  g701
  (
    n741,
    n187
  );


  xor
  g702
  (
    n739,
    n729,
    n730
  );


  or
  g703
  (
    n738,
    n183,
    n186,
    n184,
    n185
  );


  xor
  g704
  (
    n735,
    n188,
    n731,
    n728
  );


  xor
  g705
  (
    n740,
    n180,
    n182,
    n181,
    n730
  );


  not
  g706
  (
    n742,
    n738
  );


  buf
  g707
  (
    n752,
    n193
  );


  not
  g708
  (
    n746,
    n199
  );


  buf
  g709
  (
    n754,
    n734
  );


  not
  g710
  (
    n758,
    n737
  );


  buf
  g711
  (
    n748,
    n736
  );


  not
  g712
  (
    n759,
    n737
  );


  buf
  g713
  (
    n750,
    n734
  );


  not
  g714
  (
    n743,
    n736
  );


  buf
  g715
  (
    n756,
    n195
  );


  buf
  g716
  (
    n749,
    n189
  );


  nand
  g717
  (
    n751,
    n732,
    n191,
    n733
  );


  xnor
  g718
  (
    n757,
    n200,
    n198,
    n202
  );


  xor
  g719
  (
    n747,
    n192,
    n196,
    n735
  );


  xor
  g720
  (
    n744,
    n738,
    n739,
    n190
  );


  xnor
  g721
  (
    n753,
    n737,
    n735
  );


  and
  g722
  (
    n755,
    n736,
    n197,
    n201
  );


  xnor
  g723
  (
    n745,
    n194,
    n738,
    n734
  );


  nor
  g724
  (
    n760,
    n742,
    n204,
    n203,
    n205
  );


  or
  g725
  (
    n762,
    n210,
    n207,
    n208,
    n211
  );


  nand
  g726
  (
    n761,
    n206,
    n760,
    n209
  );


  not
  g727
  (
    n763,
    n761
  );


  buf
  g728
  (
    n765,
    n763
  );


  buf
  g729
  (
    n764,
    n763
  );


  buf
  g730
  (
    n768,
    n764
  );


  not
  g731
  (
    n771,
    n764
  );


  buf
  g732
  (
    n767,
    n764
  );


  buf
  g733
  (
    n770,
    n765
  );


  not
  g734
  (
    n766,
    n765
  );


  not
  g735
  (
    n772,
    n765
  );


  not
  g736
  (
    n769,
    n765
  );


  not
  g737
  (
    n775,
    n766
  );


  buf
  g738
  (
    n773,
    n767
  );


  not
  g739
  (
    n774,
    n767
  );


  and
  g740
  (
    n776,
    n213,
    n212,
    n773,
    n214
  );


  and
  g741
  (
    n778,
    n725,
    n776
  );


  xor
  g742
  (
    n777,
    n767,
    n768,
    n725,
    n776
  );


  buf
  g743
  (
    n780,
    n778
  );


  buf
  g744
  (
    n779,
    n777
  );


  nand
  g745
  (
    n781,
    n762,
    n780
  );


  or
  g746
  (
    n783,
    n217,
    n219,
    n215,
    n220
  );


  nor
  g747
  (
    n782,
    n216,
    n781,
    n218
  );


  nand
  g748
  (
    n784,
    n768,
    n782
  );


  buf
  g749
  (
    n785,
    n784
  );


  buf
  g750
  (
    n786,
    n784
  );


  xnor
  g751
  (
    n792,
    n778,
    n785
  );


  xor
  g752
  (
    n788,
    n775,
    n768,
    n770,
    n760
  );


  or
  g753
  (
    n794,
    n786,
    n769,
    n783,
    n770
  );


  xnor
  g754
  (
    n790,
    n778,
    n769,
    n774,
    n785
  );


  xnor
  g755
  (
    n789,
    n786,
    n786,
    n783,
    n775
  );


  xor
  g756
  (
    n791,
    n773,
    n783,
    n785,
    n775
  );


  nand
  g757
  (
    n793,
    n771,
    n769,
    n770,
    n774
  );


  xnor
  g758
  (
    n787,
    n774,
    n773,
    n786,
    n785
  );


  buf
  g759
  (
    n795,
    n787
  );


  not
  g760
  (
    n796,
    n787
  );


  xnor
  g761
  (
    n797,
    n739,
    n796
  );


  not
  g762
  (
    n798,
    n797
  );


  not
  g763
  (
    n799,
    n797
  );


  buf
  g764
  (
    n800,
    n798
  );


  not
  g765
  (
    n801,
    n798
  );


  not
  g766
  (
    n802,
    n798
  );


  not
  g767
  (
    n804,
    n802
  );


  buf
  g768
  (
    n805,
    n802
  );


  buf
  g769
  (
    n807,
    n800
  );


  not
  g770
  (
    n806,
    n802
  );


  buf
  g771
  (
    n803,
    n801
  );


  not
  g772
  (
    n808,
    n802
  );


  nor
  g773
  (
    n830,
    n792,
    n788
  );


  nand
  g774
  (
    n823,
    n174,
    n173
  );


  nor
  g775
  (
    n818,
    n803,
    n790
  );


  and
  g776
  (
    n813,
    n794,
    n788
  );


  xor
  g777
  (
    n820,
    n175,
    n797
  );


  nor
  g778
  (
    n815,
    n799,
    n174
  );


  and
  g779
  (
    n826,
    n175,
    n771
  );


  nand
  g780
  (
    n816,
    n808,
    n804
  );


  and
  g781
  (
    n821,
    n806,
    n807
  );


  and
  g782
  (
    n824,
    n790,
    n807
  );


  nand
  g783
  (
    n809,
    n804,
    n808
  );


  xor
  g784
  (
    n814,
    n799,
    n789
  );


  and
  g785
  (
    n811,
    n805,
    n789,
    n808,
    n792
  );


  nand
  g786
  (
    n810,
    n789,
    n807,
    n793
  );


  xnor
  g787
  (
    n832,
    n794,
    n791,
    n173
  );


  nor
  g788
  (
    n819,
    n804,
    n808,
    n794,
    n174
  );


  xor
  g789
  (
    n827,
    n788,
    n174,
    n792,
    n175
  );


  and
  g790
  (
    n822,
    n791,
    n803,
    n804,
    n799
  );


  xnor
  g791
  (
    n825,
    n805,
    n790,
    n787
  );


  and
  g792
  (
    n817,
    n173,
    n793,
    n776,
    n806
  );


  and
  g793
  (
    n828,
    n793,
    n794,
    n789,
    n805
  );


  or
  g794
  (
    n831,
    n806,
    n173,
    n792,
    n788
  );


  xnor
  g795
  (
    n812,
    n793,
    n790,
    n175,
    n806
  );


  and
  g796
  (
    n829,
    n803,
    n803,
    n805,
    n791
  );


  nor
  g797
  (
    n905,
    n489,
    n348,
    n819,
    n827
  );


  nand
  g798
  (
    n878,
    n421,
    n413,
    n824,
    n392
  );


  nor
  g799
  (
    n882,
    n328,
    n385,
    n810,
    n832
  );


  or
  g800
  (
    n850,
    n419,
    n809,
    n261
  );


  and
  g801
  (
    n917,
    n822,
    n431,
    n455,
    n227
  );


  nand
  g802
  (
    n880,
    n466,
    n820,
    n327,
    n376
  );


  nor
  g803
  (
    n888,
    n821,
    n384,
    n352,
    n829
  );


  nor
  g804
  (
    n914,
    n356,
    n248,
    n831,
    n461
  );


  xnor
  g805
  (
    n859,
    n241,
    n493,
    n333,
    n820
  );


  or
  g806
  (
    n912,
    n473,
    n222,
    n507,
    n821
  );


  nor
  g807
  (
    n858,
    n504,
    n818,
    n224,
    n445
  );


  xor
  g808
  (
    n889,
    n305,
    n828,
    n456,
    n820
  );


  nand
  g809
  (
    n835,
    n437,
    n231,
    n221,
    n810
  );


  or
  g810
  (
    n851,
    n374,
    n313,
    n433,
    n389
  );


  xnor
  g811
  (
    n843,
    n825,
    n294,
    n429,
    n502
  );


  xor
  g812
  (
    KeyWire_0_18,
    n255,
    n478,
    n372,
    n386
  );


  and
  g813
  (
    n845,
    n815,
    n828,
    n816,
    n447
  );


  or
  g814
  (
    n861,
    n298,
    n353,
    n309,
    n299
  );


  or
  g815
  (
    n913,
    n406,
    n393,
    n238,
    n278
  );


  or
  g816
  (
    n874,
    n306,
    n826,
    n815,
    n813
  );


  nand
  g817
  (
    n834,
    n382,
    n417,
    n831,
    n438
  );


  nand
  g818
  (
    n872,
    n826,
    n827,
    n246,
    n225
  );


  nand
  g819
  (
    n857,
    n271,
    n452,
    n492,
    n343
  );


  nor
  g820
  (
    n863,
    n810,
    n269,
    n317,
    n505
  );


  nand
  g821
  (
    n873,
    n373,
    n290,
    n342,
    n488
  );


  nand
  g822
  (
    n928,
    n288,
    n418,
    n256,
    n365
  );


  xor
  g823
  (
    n908,
    n239,
    n310,
    n816,
    n329
  );


  xnor
  g824
  (
    n879,
    n830,
    n812,
    n463,
    n486
  );


  or
  g825
  (
    n870,
    n415,
    n822,
    n811,
    n457
  );


  and
  g826
  (
    n910,
    n251,
    n427,
    n401,
    n366
  );


  nor
  g827
  (
    n846,
    n361,
    n816,
    n822,
    n321
  );


  nor
  g828
  (
    n838,
    n821,
    n380,
    n240,
    n474
  );


  nor
  g829
  (
    n885,
    n323,
    n282,
    n495,
    n812
  );


  xor
  g830
  (
    n848,
    n325,
    n407,
    n475,
    n249
  );


  nor
  g831
  (
    n925,
    n381,
    n399,
    n831,
    n402
  );


  nand
  g832
  (
    n915,
    n350,
    n345,
    n331,
    n387
  );


  or
  g833
  (
    n842,
    n295,
    n363,
    n276,
    n441
  );


  nand
  g834
  (
    n864,
    n454,
    n809,
    n815,
    n360
  );


  nand
  g835
  (
    n849,
    n496,
    n301,
    n228,
    n316
  );


  nor
  g836
  (
    n926,
    n275,
    n825,
    n405,
    n336
  );


  xnor
  g837
  (
    n918,
    n448,
    n330,
    n469,
    n395
  );


  xor
  g838
  (
    n867,
    n270,
    n824,
    n337,
    n817
  );


  xor
  g839
  (
    n833,
    n357,
    n390,
    n355,
    n824
  );


  xnor
  g840
  (
    n887,
    n422,
    n823,
    n237,
    n817
  );


  or
  g841
  (
    n898,
    n829,
    n257,
    n831,
    n811
  );


  xnor
  g842
  (
    n922,
    n230,
    n832,
    n829,
    n442
  );


  xor
  g843
  (
    n897,
    n281,
    n300,
    n308,
    n820
  );


  or
  g844
  (
    n920,
    n267,
    n388,
    n245,
    n440
  );


  nor
  g845
  (
    n903,
    n279,
    n825,
    n349,
    n259
  );


  xor
  g846
  (
    n852,
    n320,
    n268,
    n476,
    n483
  );


  nor
  g847
  (
    n891,
    n459,
    n414,
    n818,
    n425
  );


  nand
  g848
  (
    n862,
    n260,
    n508,
    n272,
    n443
  );


  and
  g849
  (
    n866,
    n368,
    n811,
    n464,
    n503
  );


  xnor
  g850
  (
    KeyWire_0_7,
    n335,
    n332,
    n500,
    n232
  );


  nor
  g851
  (
    n871,
    n304,
    n832,
    n428,
    n391
  );


  nand
  g852
  (
    n894,
    n340,
    n816,
    n293,
    n273
  );


  nor
  g853
  (
    n856,
    n811,
    n823,
    n311,
    n338
  );


  nor
  g854
  (
    n837,
    n346,
    n813,
    n827,
    n283
  );


  or
  g855
  (
    n883,
    n830,
    n487,
    n824,
    n462
  );


  or
  g856
  (
    n876,
    n400,
    n498,
    n814
  );


  xor
  g857
  (
    n901,
    n426,
    n253,
    n291,
    n813
  );


  xnor
  g858
  (
    n909,
    n303,
    n297,
    n817,
    n828
  );


  nand
  g859
  (
    n892,
    n809,
    n312,
    n286,
    n501
  );


  xnor
  g860
  (
    n923,
    n446,
    n817,
    n477,
    n497
  );


  nor
  g861
  (
    n884,
    n319,
    n344,
    n403,
    n409
  );


  and
  g862
  (
    n899,
    n416,
    n287,
    n449,
    n485
  );


  xnor
  g863
  (
    n924,
    n280,
    n810,
    n266,
    n814
  );


  nor
  g864
  (
    n868,
    n334,
    n296,
    n471,
    n819
  );


  nand
  g865
  (
    n900,
    n435,
    n247,
    n424,
    n412
  );


  xor
  g866
  (
    n890,
    n351,
    n818,
    n243,
    n264
  );


  xnor
  g867
  (
    n844,
    n460,
    n813,
    n307,
    n379
  );


  and
  g868
  (
    n853,
    n277,
    n827,
    n274,
    n358
  );


  xnor
  g869
  (
    n854,
    n284,
    n432,
    n490,
    n397
  );


  nand
  g870
  (
    n895,
    n472,
    n444,
    n491,
    n377
  );


  nor
  g871
  (
    n921,
    n430,
    n434,
    n819,
    n341
  );


  xor
  g872
  (
    n840,
    n458,
    n479,
    n223,
    n818
  );


  xnor
  g873
  (
    n869,
    n226,
    n359,
    n234,
    n318
  );


  or
  g874
  (
    n855,
    n347,
    n404,
    n812,
    n826
  );


  and
  g875
  (
    n927,
    n481,
    n439,
    n411,
    n450
  );


  xnor
  g876
  (
    n865,
    n375,
    n364,
    n258,
    n829
  );


  or
  g877
  (
    n886,
    n396,
    n812,
    n292,
    n339
  );


  nor
  g878
  (
    n911,
    n814,
    n823,
    n244,
    n378
  );


  and
  g879
  (
    n916,
    n826,
    n236,
    n410,
    n423
  );


  or
  g880
  (
    n847,
    n229,
    n383,
    n235,
    n825
  );


  nor
  g881
  (
    n836,
    n370,
    n482,
    n465,
    n285
  );


  and
  g882
  (
    n881,
    n314,
    n289,
    n242,
    n480
  );


  and
  g883
  (
    n919,
    n832,
    n467,
    n451,
    n315
  );


  or
  g884
  (
    n906,
    n815,
    n819,
    n302,
    n499
  );


  xor
  g885
  (
    n896,
    n394,
    n252,
    n408,
    n354
  );


  and
  g886
  (
    n904,
    n324,
    n436,
    n470,
    n398
  );


  or
  g887
  (
    n875,
    n828,
    n362,
    n250,
    n263
  );


  or
  g888
  (
    n893,
    n468,
    n822,
    n233,
    n367
  );


  or
  g889
  (
    n877,
    n484,
    n262,
    n265,
    n420
  );


  or
  g890
  (
    n841,
    n494,
    n506,
    n371,
    n322
  );


  nand
  g891
  (
    n902,
    n823,
    n830,
    n326,
    n369
  );


  xnor
  g892
  (
    n839,
    n821,
    n830,
    n254,
    n453
  );


  not
  g893
  (
    n929,
    n833
  );


  not
  g894
  (
    n932,
    n929
  );


  buf
  g895
  (
    n933,
    n929
  );


  not
  g896
  (
    n931,
    n929
  );


  buf
  g897
  (
    n930,
    n929
  );


  xor
  g898
  (
    n947,
    n551,
    n525,
    n533,
    n515
  );


  nor
  g899
  (
    n939,
    n532,
    n552,
    n932,
    n554
  );


  nand
  g900
  (
    n943,
    n553,
    n549,
    n931,
    n514
  );


  nor
  g901
  (
    n946,
    n512,
    n517,
    n933,
    n536
  );


  xnor
  g902
  (
    n937,
    n537,
    n527,
    n510,
    n516
  );


  nor
  g903
  (
    n944,
    n539,
    n932,
    n521,
    n529
  );


  xor
  g904
  (
    n948,
    n543,
    n545,
    n526,
    n931
  );


  and
  g905
  (
    n945,
    n933,
    n513,
    n522,
    n932
  );


  xor
  g906
  (
    n934,
    n548,
    n933,
    n509,
    n528
  );


  xnor
  g907
  (
    n936,
    n542,
    n556,
    n531,
    n511
  );


  xor
  g908
  (
    n949,
    n555,
    n930,
    n547
  );


  nand
  g909
  (
    n935,
    n524,
    n931,
    n518
  );


  nand
  g910
  (
    n942,
    n523,
    n538,
    n530,
    n930
  );


  and
  g911
  (
    n940,
    n933,
    n544,
    n932,
    n550
  );


  xnor
  g912
  (
    n938,
    n541,
    n546,
    n535,
    n540
  );


  and
  g913
  (
    n941,
    n930,
    n520,
    n534,
    n519
  );


  buf
  g914
  (
    n951,
    n943
  );


  not
  g915
  (
    n950,
    n944
  );


  buf
  g916
  (
    n957,
    n950
  );


  buf
  g917
  (
    n955,
    n950
  );


  buf
  g918
  (
    n953,
    n950
  );


  not
  g919
  (
    n952,
    n951
  );


  buf
  g920
  (
    n956,
    n951
  );


  not
  g921
  (
    n958,
    n951
  );


  not
  g922
  (
    n959,
    n950
  );


  not
  g923
  (
    n954,
    n951
  );


  buf
  g924
  (
    n971,
    n956
  );


  not
  g925
  (
    n985,
    n954
  );


  not
  g926
  (
    n977,
    n955
  );


  buf
  g927
  (
    n981,
    n954
  );


  not
  g928
  (
    n984,
    n955
  );


  buf
  g929
  (
    n982,
    n952
  );


  buf
  g930
  (
    n967,
    n956
  );


  buf
  g931
  (
    n969,
    n958
  );


  not
  g932
  (
    n979,
    n957
  );


  not
  g933
  (
    n983,
    n954
  );


  buf
  g934
  (
    n973,
    n957
  );


  buf
  g935
  (
    n968,
    n955
  );


  buf
  g936
  (
    n960,
    n952
  );


  buf
  g937
  (
    n970,
    n953
  );


  buf
  g938
  (
    n972,
    n956
  );


  not
  g939
  (
    n976,
    n952
  );


  not
  g940
  (
    n961,
    n953
  );


  buf
  g941
  (
    n975,
    n956
  );


  not
  g942
  (
    n965,
    n954
  );


  buf
  g943
  (
    n966,
    n957
  );


  buf
  g944
  (
    n974,
    n955
  );


  buf
  g945
  (
    n962,
    n953
  );


  buf
  g946
  (
    n978,
    n953
  );


  not
  g947
  (
    n963,
    n952
  );


  buf
  g948
  (
    n964,
    n958
  );


  buf
  g949
  (
    n980,
    n957
  );


  buf
  g950
  (
    n1059,
    n984
  );


  buf
  g951
  (
    n1084,
    n973
  );


  not
  g952
  (
    n988,
    n979
  );


  not
  g953
  (
    n1053,
    n962
  );


  not
  g954
  (
    n993,
    n967
  );


  not
  g955
  (
    n1012,
    n984
  );


  not
  g956
  (
    n1021,
    n965
  );


  buf
  g957
  (
    n1023,
    n982
  );


  buf
  g958
  (
    n1088,
    n978
  );


  buf
  g959
  (
    n1041,
    n981
  );


  buf
  g960
  (
    n1062,
    n963
  );


  not
  g961
  (
    n1057,
    n985
  );


  not
  g962
  (
    n986,
    n970
  );


  buf
  g963
  (
    n1086,
    n978
  );


  not
  g964
  (
    n1010,
    n981
  );


  not
  g965
  (
    n1081,
    n974
  );


  buf
  g966
  (
    n1066,
    n972
  );


  not
  g967
  (
    n1024,
    n971
  );


  not
  g968
  (
    n1003,
    n984
  );


  buf
  g969
  (
    n1031,
    n983
  );


  not
  g970
  (
    n1038,
    n971
  );


  buf
  g971
  (
    n995,
    n963
  );


  not
  g972
  (
    n1045,
    n984
  );


  buf
  g973
  (
    n1005,
    n966
  );


  buf
  g974
  (
    n1052,
    n982
  );


  buf
  g975
  (
    n997,
    n966
  );


  not
  g976
  (
    n1006,
    n971
  );


  not
  g977
  (
    n1067,
    n968
  );


  not
  g978
  (
    n1061,
    n982
  );


  not
  g979
  (
    n1042,
    n772
  );


  buf
  g980
  (
    n1002,
    n970
  );


  not
  g981
  (
    n992,
    n970
  );


  not
  g982
  (
    n1032,
    n962
  );


  not
  g983
  (
    n1025,
    n973
  );


  buf
  g984
  (
    n1078,
    n964
  );


  not
  g985
  (
    n1017,
    n970
  );


  not
  g986
  (
    n1026,
    n980
  );


  not
  g987
  (
    n1077,
    n969
  );


  buf
  g988
  (
    n1063,
    n958
  );


  not
  g989
  (
    n1001,
    n964
  );


  buf
  g990
  (
    n1051,
    n961
  );


  buf
  g991
  (
    n1035,
    n977
  );


  buf
  g992
  (
    n1019,
    n979
  );


  buf
  g993
  (
    n989,
    n967
  );


  buf
  g994
  (
    n1004,
    n964
  );


  buf
  g995
  (
    n991,
    n968
  );


  not
  g996
  (
    n1047,
    n969
  );


  buf
  g997
  (
    n1015,
    n968
  );


  not
  g998
  (
    n1075,
    n965
  );


  buf
  g999
  (
    n1056,
    n979
  );


  not
  g1000
  (
    n1036,
    n962
  );


  not
  g1001
  (
    n1043,
    n963
  );


  not
  g1002
  (
    n1071,
    n960
  );


  not
  g1003
  (
    n1022,
    n964
  );


  not
  g1004
  (
    n1039,
    n772
  );


  buf
  g1005
  (
    n1007,
    n969
  );


  buf
  g1006
  (
    n1085,
    n971
  );


  buf
  g1007
  (
    n1046,
    n976
  );


  buf
  g1008
  (
    n1054,
    n771
  );


  not
  g1009
  (
    n1087,
    n974
  );


  not
  g1010
  (
    n1011,
    n968
  );


  buf
  g1011
  (
    n1060,
    n973
  );


  not
  g1012
  (
    n1072,
    n975
  );


  not
  g1013
  (
    n1000,
    n979
  );


  not
  g1014
  (
    n1089,
    n972
  );


  buf
  g1015
  (
    n999,
    n985
  );


  not
  g1016
  (
    n1074,
    n977
  );


  buf
  g1017
  (
    n1034,
    n772
  );


  not
  g1018
  (
    n1058,
    n966
  );


  buf
  g1019
  (
    n1027,
    n967
  );


  buf
  g1020
  (
    n990,
    n772
  );


  buf
  g1021
  (
    n1064,
    n965
  );


  not
  g1022
  (
    n1044,
    n981
  );


  not
  g1023
  (
    n1050,
    n983
  );


  not
  g1024
  (
    n1049,
    n973
  );


  not
  g1025
  (
    n1048,
    n975
  );


  not
  g1026
  (
    n1009,
    n983
  );


  buf
  g1027
  (
    n1069,
    n976
  );


  buf
  g1028
  (
    KeyWire_0_30,
    n976
  );


  buf
  g1029
  (
    n1016,
    n965
  );


  buf
  g1030
  (
    n1079,
    n975
  );


  not
  g1031
  (
    n994,
    n980
  );


  buf
  g1032
  (
    n1030,
    n961
  );


  buf
  g1033
  (
    n1073,
    n975
  );


  not
  g1034
  (
    n1020,
    n983
  );


  not
  g1035
  (
    n1029,
    n974
  );


  not
  g1036
  (
    n1008,
    n985
  );


  buf
  g1037
  (
    n1080,
    n961
  );


  buf
  g1038
  (
    n998,
    n963
  );


  buf
  g1039
  (
    n1070,
    n960
  );


  not
  g1040
  (
    n1076,
    n961
  );


  not
  g1041
  (
    n987,
    n962
  );


  buf
  g1042
  (
    n1033,
    n974
  );


  not
  g1043
  (
    n1068,
    n969
  );


  buf
  g1044
  (
    n1082,
    n978
  );


  buf
  g1045
  (
    n1013,
    n967
  );


  buf
  g1046
  (
    n1065,
    n966
  );


  buf
  g1047
  (
    n1040,
    n960
  );


  buf
  g1048
  (
    n1037,
    n978
  );


  buf
  g1049
  (
    n1018,
    n980
  );


  buf
  g1050
  (
    n1028,
    n972
  );


  not
  g1051
  (
    n1055,
    n972
  );


  and
  g1052
  (
    n1014,
    n985,
    n977,
    n980
  );


  and
  g1053
  (
    n1083,
    n981,
    n976,
    n960,
    n982
  );


  not
  g1054
  (
    n1309,
    n740
  );


  not
  g1055
  (
    n1480,
    n1041
  );


  buf
  g1056
  (
    n1410,
    n1070
  );


  buf
  g1057
  (
    n1487,
    n1015
  );


  buf
  g1058
  (
    n1411,
    n838
  );


  not
  g1059
  (
    n1389,
    n861
  );


  buf
  g1060
  (
    n1297,
    n1024
  );


  buf
  g1061
  (
    n1245,
    n1008
  );


  buf
  g1062
  (
    n1357,
    n1026
  );


  not
  g1063
  (
    n1431,
    n1068
  );


  buf
  g1064
  (
    n1499,
    n891
  );


  buf
  g1065
  (
    n1208,
    n1013
  );


  not
  g1066
  (
    n1222,
    n1057
  );


  buf
  g1067
  (
    n1278,
    n853
  );


  not
  g1068
  (
    n1149,
    n868
  );


  buf
  g1069
  (
    n1285,
    n1002
  );


  buf
  g1070
  (
    n1127,
    n838
  );


  buf
  g1071
  (
    n1335,
    n1016
  );


  not
  g1072
  (
    n1488,
    n895
  );


  not
  g1073
  (
    n1383,
    n849
  );


  not
  g1074
  (
    n1144,
    n1046
  );


  not
  g1075
  (
    n1492,
    n1061
  );


  buf
  g1076
  (
    n1476,
    n1041
  );


  buf
  g1077
  (
    n1465,
    n1087
  );


  buf
  g1078
  (
    n1253,
    n1020
  );


  not
  g1079
  (
    n1240,
    n917
  );


  not
  g1080
  (
    n1132,
    n1074
  );


  not
  g1081
  (
    n1286,
    n1012
  );


  buf
  g1082
  (
    n1243,
    n891
  );


  not
  g1083
  (
    n1439,
    n1012
  );


  buf
  g1084
  (
    n1458,
    n1015
  );


  buf
  g1085
  (
    n1442,
    n882
  );


  buf
  g1086
  (
    n1112,
    n1079
  );


  buf
  g1087
  (
    n1348,
    n994
  );


  buf
  g1088
  (
    n1113,
    n1001
  );


  buf
  g1089
  (
    n1415,
    n924
  );


  not
  g1090
  (
    n1408,
    n851
  );


  buf
  g1091
  (
    n1427,
    n1069
  );


  not
  g1092
  (
    n1241,
    n908
  );


  buf
  g1093
  (
    n1198,
    n928
  );


  buf
  g1094
  (
    n1280,
    n849
  );


  not
  g1095
  (
    n1391,
    n1065
  );


  not
  g1096
  (
    n1138,
    n1000
  );


  not
  g1097
  (
    n1231,
    n1051
  );


  not
  g1098
  (
    n1261,
    n915
  );


  not
  g1099
  (
    n1294,
    n1068
  );


  not
  g1100
  (
    n1456,
    n989
  );


  buf
  g1101
  (
    n1232,
    n873
  );


  buf
  g1102
  (
    n1179,
    n1080
  );


  not
  g1103
  (
    n1327,
    n1081
  );


  not
  g1104
  (
    n1239,
    n901
  );


  buf
  g1105
  (
    n1402,
    n1072
  );


  buf
  g1106
  (
    n1299,
    n1013
  );


  buf
  g1107
  (
    n1190,
    n1014
  );


  not
  g1108
  (
    n1090,
    n834
  );


  not
  g1109
  (
    n1407,
    n913
  );


  not
  g1110
  (
    n1331,
    n1077
  );


  not
  g1111
  (
    n1466,
    n1046
  );


  buf
  g1112
  (
    n1305,
    n1086
  );


  buf
  g1113
  (
    n1369,
    n882
  );


  not
  g1114
  (
    n1249,
    n902
  );


  buf
  g1115
  (
    n1344,
    n905
  );


  buf
  g1116
  (
    n1443,
    n1026
  );


  buf
  g1117
  (
    n1459,
    n868
  );


  buf
  g1118
  (
    n1346,
    n1001
  );


  not
  g1119
  (
    n1436,
    n840
  );


  buf
  g1120
  (
    n1159,
    n1055
  );


  not
  g1121
  (
    n1171,
    n916
  );


  not
  g1122
  (
    n1306,
    n909
  );


  buf
  g1123
  (
    n1228,
    n959
  );


  buf
  g1124
  (
    n1312,
    n1062
  );


  buf
  g1125
  (
    n1233,
    n858
  );


  not
  g1126
  (
    n1468,
    n1079
  );


  buf
  g1127
  (
    n1255,
    n991
  );


  not
  g1128
  (
    n1098,
    n879
  );


  buf
  g1129
  (
    n1355,
    n1080
  );


  buf
  g1130
  (
    n1417,
    n923
  );


  buf
  g1131
  (
    n1258,
    n910
  );


  buf
  g1132
  (
    n1288,
    n1067
  );


  not
  g1133
  (
    n1289,
    n903
  );


  not
  g1134
  (
    n1191,
    n872
  );


  buf
  g1135
  (
    n1237,
    n881
  );


  buf
  g1136
  (
    n1244,
    n1079
  );


  buf
  g1137
  (
    n1152,
    n1000
  );


  not
  g1138
  (
    n1474,
    n879
  );


  buf
  g1139
  (
    n1446,
    n1084
  );


  not
  g1140
  (
    n1412,
    n1058
  );


  buf
  g1141
  (
    n1291,
    n1078
  );


  buf
  g1142
  (
    n1182,
    n1071
  );


  buf
  g1143
  (
    n1314,
    n877
  );


  buf
  g1144
  (
    n1100,
    n996
  );


  not
  g1145
  (
    n1192,
    n1031
  );


  buf
  g1146
  (
    n1096,
    n1085
  );


  buf
  g1147
  (
    n1102,
    n1053
  );


  not
  g1148
  (
    n1329,
    n877
  );


  not
  g1149
  (
    n1490,
    n863
  );


  buf
  g1150
  (
    n1178,
    n1087
  );


  not
  g1151
  (
    n1212,
    n1015
  );


  not
  g1152
  (
    n1393,
    n883
  );


  not
  g1153
  (
    n1359,
    n1006
  );


  not
  g1154
  (
    n1452,
    n1032
  );


  buf
  g1155
  (
    n1390,
    n1002
  );


  buf
  g1156
  (
    n1125,
    n898
  );


  buf
  g1157
  (
    n1143,
    n864
  );


  not
  g1158
  (
    n1366,
    n1047
  );


  buf
  g1159
  (
    n1284,
    n1019
  );


  not
  g1160
  (
    n1338,
    n834
  );


  buf
  g1161
  (
    n1223,
    n915
  );


  not
  g1162
  (
    n1221,
    n959
  );


  buf
  g1163
  (
    n1124,
    n1070
  );


  buf
  g1164
  (
    n1200,
    n835
  );


  buf
  g1165
  (
    n1328,
    n920
  );


  not
  g1166
  (
    n1292,
    n896
  );


  buf
  g1167
  (
    n1301,
    n859
  );


  buf
  g1168
  (
    n1129,
    n881
  );


  buf
  g1169
  (
    n1130,
    n884
  );


  buf
  g1170
  (
    n1247,
    n875
  );


  buf
  g1171
  (
    n1105,
    n844
  );


  buf
  g1172
  (
    n1375,
    n1013
  );


  not
  g1173
  (
    n1414,
    n918
  );


  buf
  g1174
  (
    n1091,
    n1056
  );


  not
  g1175
  (
    n1422,
    n927
  );


  buf
  g1176
  (
    n1265,
    n1027
  );


  not
  g1177
  (
    n1399,
    n1060
  );


  buf
  g1178
  (
    n1449,
    n846
  );


  not
  g1179
  (
    n1347,
    n1027
  );


  not
  g1180
  (
    n1116,
    n896
  );


  not
  g1181
  (
    n1336,
    n916
  );


  not
  g1182
  (
    n1404,
    n1012
  );


  not
  g1183
  (
    n1351,
    n993
  );


  not
  g1184
  (
    n1454,
    n1084
  );


  not
  g1185
  (
    n1093,
    n835
  );


  not
  g1186
  (
    n1106,
    n866
  );


  buf
  g1187
  (
    n1308,
    n894
  );


  not
  g1188
  (
    n1364,
    n1008
  );


  not
  g1189
  (
    n1406,
    n848
  );


  not
  g1190
  (
    n1498,
    n1000
  );


  buf
  g1191
  (
    n1101,
    n833
  );


  buf
  g1192
  (
    n1156,
    n878
  );


  not
  g1193
  (
    n1400,
    n1049
  );


  not
  g1194
  (
    n1464,
    n1051
  );


  buf
  g1195
  (
    n1425,
    n914
  );


  buf
  g1196
  (
    n1199,
    n1081
  );


  buf
  g1197
  (
    n1374,
    n860
  );


  buf
  g1198
  (
    n1227,
    n1075
  );


  buf
  g1199
  (
    n1111,
    n998
  );


  not
  g1200
  (
    n1413,
    n1044
  );


  not
  g1201
  (
    n1287,
    n991
  );


  not
  g1202
  (
    n1146,
    n843
  );


  not
  g1203
  (
    n1204,
    n851
  );


  buf
  g1204
  (
    n1438,
    n901
  );


  not
  g1205
  (
    n1453,
    n1034
  );


  buf
  g1206
  (
    n1254,
    n873
  );


  not
  g1207
  (
    n1259,
    n1059
  );


  buf
  g1208
  (
    n1320,
    n903
  );


  not
  g1209
  (
    n1447,
    n857
  );


  not
  g1210
  (
    n1173,
    n741
  );


  not
  g1211
  (
    n1209,
    n1019
  );


  buf
  g1212
  (
    n1372,
    n861
  );


  buf
  g1213
  (
    n1483,
    n921
  );


  buf
  g1214
  (
    n1142,
    n1066
  );


  buf
  g1215
  (
    n1358,
    n921
  );


  buf
  g1216
  (
    n1290,
    n1003
  );


  not
  g1217
  (
    n1441,
    n911
  );


  buf
  g1218
  (
    n1162,
    n1013
  );


  not
  g1219
  (
    n1360,
    n882
  );


  buf
  g1220
  (
    n1435,
    n833
  );


  not
  g1221
  (
    n1214,
    n1005
  );


  not
  g1222
  (
    n1371,
    n1041
  );


  not
  g1223
  (
    n1154,
    n837
  );


  not
  g1224
  (
    n1282,
    n1009
  );


  buf
  g1225
  (
    KeyWire_0_5,
    n1042
  );


  buf
  g1226
  (
    n1187,
    n741
  );


  not
  g1227
  (
    n1267,
    n1052
  );


  not
  g1228
  (
    n1386,
    n920
  );


  not
  g1229
  (
    n1275,
    n899
  );


  buf
  g1230
  (
    n1135,
    n918
  );


  not
  g1231
  (
    n1109,
    n855
  );


  buf
  g1232
  (
    n1201,
    n1047
  );


  buf
  g1233
  (
    n1317,
    n1061
  );


  buf
  g1234
  (
    n1445,
    n859
  );


  buf
  g1235
  (
    n1202,
    n893
  );


  not
  g1236
  (
    n1491,
    n1069
  );


  buf
  g1237
  (
    n1462,
    n1026
  );


  not
  g1238
  (
    n1450,
    n884
  );


  not
  g1239
  (
    n1107,
    n873
  );


  not
  g1240
  (
    n1170,
    n903
  );


  not
  g1241
  (
    n1172,
    n1080
  );


  not
  g1242
  (
    n1262,
    n836
  );


  buf
  g1243
  (
    n1455,
    n1021
  );


  not
  g1244
  (
    n1174,
    n839
  );


  not
  g1245
  (
    n1368,
    n870
  );


  buf
  g1246
  (
    n1242,
    n900
  );


  buf
  g1247
  (
    n1473,
    n1043
  );


  buf
  g1248
  (
    n1215,
    n1088
  );


  buf
  g1249
  (
    n1379,
    n1043
  );


  buf
  g1250
  (
    n1332,
    n876
  );


  buf
  g1251
  (
    KeyWire_0_11,
    n919
  );


  not
  g1252
  (
    n1424,
    n997
  );


  buf
  g1253
  (
    n1334,
    n1088
  );


  buf
  g1254
  (
    n1382,
    n1052
  );


  not
  g1255
  (
    n1185,
    n1053
  );


  buf
  g1256
  (
    n1225,
    n923
  );


  buf
  g1257
  (
    n1134,
    n841
  );


  buf
  g1258
  (
    n1457,
    n1003
  );


  not
  g1259
  (
    n1167,
    n904
  );


  buf
  g1260
  (
    n1429,
    n1058
  );


  buf
  g1261
  (
    n1356,
    n1072
  );


  buf
  g1262
  (
    n1363,
    n1067
  );


  not
  g1263
  (
    n1184,
    n1052
  );


  buf
  g1264
  (
    n1120,
    n879
  );


  buf
  g1265
  (
    n1307,
    n872
  );


  buf
  g1266
  (
    n1108,
    n904
  );


  not
  g1267
  (
    n1343,
    n1078
  );


  buf
  g1268
  (
    n1114,
    n1070
  );


  not
  g1269
  (
    n1396,
    n1022
  );


  not
  g1270
  (
    n1119,
    n846
  );


  buf
  g1271
  (
    n1145,
    n1036
  );


  not
  g1272
  (
    n1502,
    n882
  );


  buf
  g1273
  (
    n1104,
    n1089
  );


  buf
  g1274
  (
    n1342,
    n881
  );


  not
  g1275
  (
    n1256,
    n1078
  );


  buf
  g1276
  (
    n1181,
    n1040
  );


  buf
  g1277
  (
    n1218,
    n835
  );


  not
  g1278
  (
    n1207,
    n1011
  );


  buf
  g1279
  (
    n1479,
    n890
  );


  buf
  g1280
  (
    n1213,
    n1035
  );


  buf
  g1281
  (
    n1340,
    n1064
  );


  buf
  g1282
  (
    n1416,
    n922
  );


  buf
  g1283
  (
    n1180,
    n875
  );


  buf
  g1284
  (
    n1463,
    n1028
  );


  not
  g1285
  (
    n1230,
    n1059
  );


  buf
  g1286
  (
    n1423,
    n1084
  );


  not
  g1287
  (
    n1103,
    n1082
  );


  not
  g1288
  (
    n1197,
    n996
  );


  not
  g1289
  (
    n1151,
    n1082
  );


  buf
  g1290
  (
    n1354,
    n986
  );


  not
  g1291
  (
    n1270,
    n1083
  );


  buf
  g1292
  (
    n1216,
    n905
  );


  buf
  g1293
  (
    n1220,
    n1035
  );


  not
  g1294
  (
    n1401,
    n1061
  );


  not
  g1295
  (
    n1131,
    n1089
  );


  not
  g1296
  (
    n1426,
    n866
  );


  buf
  g1297
  (
    n1303,
    n1031
  );


  not
  g1298
  (
    n1398,
    n912
  );


  not
  g1299
  (
    n1210,
    n845
  );


  buf
  g1300
  (
    n1196,
    n1081
  );


  buf
  g1301
  (
    n1362,
    n834
  );


  not
  g1302
  (
    n1163,
    n1005
  );


  buf
  g1303
  (
    n1277,
    n885
  );


  not
  g1304
  (
    n1339,
    n838
  );


  not
  g1305
  (
    n1418,
    n897
  );


  buf
  g1306
  (
    n1248,
    n987
  );


  buf
  g1307
  (
    n1133,
    n900
  );


  not
  g1308
  (
    n1434,
    n1038
  );


  not
  g1309
  (
    n1161,
    n1054
  );


  buf
  g1310
  (
    n1295,
    n1083
  );


  not
  g1311
  (
    n1475,
    n862
  );


  buf
  g1312
  (
    n1318,
    n1085
  );


  buf
  g1313
  (
    n1503,
    n903
  );


  buf
  g1314
  (
    n1378,
    n1075
  );


  not
  g1315
  (
    n1341,
    n986
  );


  buf
  g1316
  (
    n1293,
    n1074
  );


  buf
  g1317
  (
    n1257,
    n1037
  );


  not
  g1318
  (
    n1150,
    n906
  );


  buf
  g1319
  (
    n1097,
    n1066
  );


  buf
  g1320
  (
    n1252,
    n1042
  );


  buf
  g1321
  (
    n1419,
    n901
  );


  buf
  g1322
  (
    n1121,
    n1056
  );


  not
  g1323
  (
    n1316,
    n1025
  );


  buf
  g1324
  (
    n1333,
    n927
  );


  buf
  g1325
  (
    n1251,
    n1043
  );


  buf
  g1326
  (
    n1319,
    n987
  );


  not
  g1327
  (
    n1166,
    n843
  );


  not
  g1328
  (
    n1183,
    n848
  );


  not
  g1329
  (
    n1203,
    n847
  );


  buf
  g1330
  (
    n1229,
    n1009
  );


  buf
  g1331
  (
    n1323,
    n1005
  );


  buf
  g1332
  (
    n1496,
    n1067
  );


  buf
  g1333
  (
    n1160,
    n1053
  );


  not
  g1334
  (
    n1164,
    n1024
  );


  not
  g1335
  (
    n1380,
    n991
  );


  not
  g1336
  (
    n1126,
    n863
  );


  not
  g1337
  (
    n1430,
    n1039
  );


  xor
  g1338
  (
    n1494,
    n888,
    n852,
    n922,
    n883
  );


  xnor
  g1339
  (
    n1193,
    n1082,
    n1018,
    n876,
    n1010
  );


  or
  g1340
  (
    n1272,
    n1044,
    n1012,
    n1070,
    n916
  );


  xnor
  g1341
  (
    n1186,
    n1064,
    n871,
    n879,
    n886
  );


  xor
  g1342
  (
    n1448,
    n841,
    n1041,
    n901,
    n891
  );


  nor
  g1343
  (
    n1409,
    n989,
    n1026,
    n1034,
    n880
  );


  and
  g1344
  (
    n1326,
    n897,
    n908,
    n918,
    n1044
  );


  or
  g1345
  (
    n1246,
    n1060,
    n912,
    n837,
    n1003
  );


  nor
  g1346
  (
    n1175,
    n1049,
    n1005,
    n1050,
    n878
  );


  or
  g1347
  (
    n1211,
    n1077,
    n840,
    n889,
    n1050
  );


  xor
  g1348
  (
    n1148,
    n906,
    n887,
    n844,
    n1007
  );


  or
  g1349
  (
    n1226,
    n1051,
    n1077,
    n1023,
    n911
  );


  nor
  g1350
  (
    n1206,
    n923,
    n1045,
    n1086,
    n911
  );


  nor
  g1351
  (
    n1482,
    n892,
    n740,
    n925,
    n1035
  );


  and
  g1352
  (
    n1451,
    n1039,
    n1073,
    n902,
    n1083
  );


  xnor
  g1353
  (
    n1370,
    n1011,
    n888,
    n1030,
    n1063
  );


  nand
  g1354
  (
    n1461,
    n851,
    n1002,
    n1075,
    n988
  );


  nand
  g1355
  (
    n1188,
    n1018,
    n893,
    n1054,
    n1076
  );


  nand
  g1356
  (
    n1397,
    n1018,
    n1036,
    n1011,
    n867
  );


  xor
  g1357
  (
    n1421,
    n890,
    n885,
    n928,
    n875
  );


  nor
  g1358
  (
    n1433,
    n898,
    n991,
    n840,
    n1011
  );


  or
  g1359
  (
    n1099,
    n859,
    n1076,
    n874,
    n881
  );


  xor
  g1360
  (
    n1349,
    n834,
    n1084,
    n880,
    n913
  );


  xnor
  g1361
  (
    n1324,
    n1050,
    n1014,
    n920,
    n921
  );


  xor
  g1362
  (
    n1489,
    n1006,
    n888,
    n1010,
    n853
  );


  and
  g1363
  (
    n1469,
    n920,
    n1058,
    n837,
    n1049
  );


  nor
  g1364
  (
    n1350,
    n922,
    n868,
    n908,
    n1004
  );


  or
  g1365
  (
    n1123,
    n877,
    n959,
    n1016,
    n1054
  );


  xor
  g1366
  (
    n1165,
    n1015,
    n867,
    n1017,
    n1009
  );


  xnor
  g1367
  (
    n1234,
    n1019,
    n844,
    n1023,
    n847
  );


  and
  g1368
  (
    n1147,
    n927,
    n992,
    n1017,
    n1051
  );


  nand
  g1369
  (
    n1189,
    n1063,
    n1030,
    n926,
    n849
  );


  xor
  g1370
  (
    n1428,
    n845,
    n905,
    n867,
    n1048
  );


  nand
  g1371
  (
    n1444,
    n1086,
    n908,
    n1088,
    n1042
  );


  or
  g1372
  (
    n1353,
    n854,
    n1020,
    n843,
    n835
  );


  or
  g1373
  (
    n1330,
    n1074,
    n836,
    n911,
    n896
  );


  xor
  g1374
  (
    n1325,
    n1006,
    n904,
    n841,
    n918
  );


  and
  g1375
  (
    n1432,
    n992,
    n842,
    n926,
    n855
  );


  xnor
  g1376
  (
    n1279,
    n910,
    n1014,
    n1069,
    n894
  );


  xnor
  g1377
  (
    n1122,
    n850,
    n857,
    n1087,
    n844
  );


  xor
  g1378
  (
    n1194,
    n894,
    n925,
    n889,
    n850
  );


  xor
  g1379
  (
    n1505,
    n871,
    n839,
    n856,
    n740
  );


  or
  g1380
  (
    n1269,
    n1029,
    n1033,
    n1048,
    n1044
  );


  nor
  g1381
  (
    n1300,
    n917,
    n895,
    n1003,
    n870
  );


  or
  g1382
  (
    n1497,
    n839,
    n874,
    n1032,
    n741
  );


  nor
  g1383
  (
    n1394,
    n1032,
    n990,
    n887,
    n994
  );


  or
  g1384
  (
    n1128,
    n866,
    n1055,
    n860,
    n1029
  );


  nor
  g1385
  (
    n1381,
    n1059,
    n1072,
    n909,
    n1009
  );


  or
  g1386
  (
    n1235,
    n1007,
    n1060,
    n865,
    n999
  );


  or
  g1387
  (
    n1321,
    n1052,
    n997,
    n854,
    n1020
  );


  and
  g1388
  (
    n1264,
    n999,
    n865,
    n876,
    n1032
  );


  or
  g1389
  (
    n1471,
    n1065,
    n890,
    n1089,
    n1036
  );


  and
  g1390
  (
    n1095,
    n1007,
    n1025,
    n907,
    n986
  );


  nand
  g1391
  (
    n1395,
    n1001,
    n1038,
    n988,
    n912
  );


  nand
  g1392
  (
    n1388,
    n997,
    n889,
    n1080,
    n993
  );


  nor
  g1393
  (
    n1155,
    n1042,
    n1023,
    n885,
    n868
  );


  nand
  g1394
  (
    n1392,
    n899,
    n915,
    n872,
    n1030
  );


  nand
  g1395
  (
    n1094,
    n1010,
    n888,
    n1062,
    n862
  );


  xnor
  g1396
  (
    n1110,
    n884,
    n1040,
    n999
  );


  or
  g1397
  (
    n1485,
    n1028,
    n862,
    n874,
    n1045
  );


  and
  g1398
  (
    n1500,
    n886,
    n1039,
    n907,
    n914
  );


  and
  g1399
  (
    n1157,
    n842,
    n843,
    n997,
    n1031
  );


  xor
  g1400
  (
    n1238,
    n1045,
    n1085,
    n856,
    n1034
  );


  nand
  g1401
  (
    n1478,
    n861,
    n890,
    n902,
    n878
  );


  and
  g1402
  (
    n1139,
    n1057,
    n883,
    n873,
    n1022
  );


  nand
  g1403
  (
    n1266,
    n1034,
    n880,
    n1033,
    n1071
  );


  xnor
  g1404
  (
    n1365,
    n900,
    n1000,
    n1019,
    n842
  );


  nor
  g1405
  (
    n1481,
    n1022,
    n1079,
    n1008,
    n1062
  );


  or
  g1406
  (
    n1501,
    n902,
    n987,
    n1020,
    n919
  );


  xor
  g1407
  (
    n1281,
    n1053,
    n1048,
    n895,
    n928
  );


  xor
  g1408
  (
    n1304,
    n1082,
    n905,
    n1021,
    n992
  );


  or
  g1409
  (
    n1495,
    n872,
    n914,
    n853,
    n924
  );


  nand
  g1410
  (
    n1217,
    n926,
    n853,
    n1067,
    n1059
  );


  xnor
  g1411
  (
    n1158,
    n924,
    n886,
    n1066,
    n898
  );


  nand
  g1412
  (
    n1345,
    n900,
    n1002,
    n925,
    n892
  );


  and
  g1413
  (
    n1274,
    n865,
    n1056,
    n1004
  );


  or
  g1414
  (
    n1260,
    n1033,
    n841,
    n1073,
    n856
  );


  nand
  g1415
  (
    n1250,
    n855,
    n894,
    n852,
    n866
  );


  nor
  g1416
  (
    n1092,
    n1043,
    n993,
    n1056,
    n1047
  );


  nand
  g1417
  (
    n1377,
    n851,
    n1021,
    n1049,
    n925
  );


  or
  g1418
  (
    n1484,
    n1073,
    n858,
    n1004,
    n923
  );


  xor
  g1419
  (
    n1403,
    n874,
    n1035,
    n990,
    n864
  );


  xnor
  g1420
  (
    n1467,
    n1007,
    n836,
    n1001,
    n995
  );


  nand
  g1421
  (
    n1236,
    n1038,
    n856,
    n1071,
    n848
  );


  and
  g1422
  (
    n1140,
    n837,
    n988,
    n880,
    n1073
  );


  xnor
  g1423
  (
    n1137,
    n994,
    n858,
    n1068,
    n847
  );


  xor
  g1424
  (
    n1460,
    n986,
    n857,
    n1028,
    n910
  );


  and
  g1425
  (
    n1296,
    n864,
    n988,
    n1063,
    n1028
  );


  nor
  g1426
  (
    n1263,
    n1083,
    n1068,
    n893,
    n1025
  );


  nor
  g1427
  (
    n1373,
    n871,
    n869,
    n860,
    n1057
  );


  xor
  g1428
  (
    n1337,
    n1074,
    n863,
    n917,
    n1055
  );


  or
  g1429
  (
    n1352,
    n1085,
    n1017,
    n1037,
    n917
  );


  nand
  g1430
  (
    n1361,
    n1018,
    n1027,
    n1008,
    n861
  );


  or
  g1431
  (
    n1273,
    n895,
    n912,
    n897,
    n1076
  );


  nor
  g1432
  (
    n1115,
    n928,
    n850,
    n739,
    n897
  );


  xor
  g1433
  (
    n1169,
    n849,
    n1031,
    n1036,
    n959
  );


  nor
  g1434
  (
    n1437,
    n994,
    n875,
    n1081,
    n1038
  );


  nor
  g1435
  (
    n1302,
    n993,
    n989,
    n889
  );


  xnor
  g1436
  (
    n1268,
    n1024,
    n1033,
    n1065,
    n1037
  );


  nand
  g1437
  (
    n1315,
    n987,
    n1066,
    n884,
    n869
  );


  nand
  g1438
  (
    n1271,
    n1022,
    n1016,
    n1072,
    n840
  );


  xnor
  g1439
  (
    n1387,
    n1063,
    n998,
    n1061,
    n1057
  );


  nor
  g1440
  (
    n1176,
    n1017,
    n1078,
    n838,
    n1062
  );


  xnor
  g1441
  (
    n1311,
    n1029,
    n852,
    n906,
    n854
  );


  or
  g1442
  (
    n1298,
    n1076,
    n893,
    n899,
    n1023
  );


  xor
  g1443
  (
    n1118,
    n839,
    n1075,
    n1087,
    n1040
  );


  xor
  g1444
  (
    n1283,
    n998,
    n865,
    n1029,
    n1046
  );


  nand
  g1445
  (
    n1472,
    n1016,
    n860,
    n863,
    n999
  );


  nor
  g1446
  (
    KeyWire_0_8,
    n857,
    n1089,
    n1039,
    n927
  );


  xor
  g1447
  (
    n1420,
    n847,
    n1047,
    n996,
    n836
  );


  and
  g1448
  (
    n1136,
    n899,
    n869,
    n924
  );


  xor
  g1449
  (
    n1205,
    n887,
    n1030,
    n896,
    n877
  );


  nand
  g1450
  (
    n1493,
    n909,
    n1088,
    n919,
    n1064
  );


  xnor
  g1451
  (
    n1504,
    n1006,
    n870,
    n867,
    n891
  );


  xnor
  g1452
  (
    KeyWire_0_27,
    n862,
    n990,
    n887,
    n998
  );


  or
  g1453
  (
    n1177,
    n1050,
    n1024,
    n1021,
    n892
  );


  nor
  g1454
  (
    n1219,
    n886,
    n1060,
    n990,
    n995
  );


  nand
  g1455
  (
    n1168,
    n1010,
    n885,
    n1046,
    n914
  );


  xor
  g1456
  (
    n1376,
    n1064,
    n870,
    n921,
    n846
  );


  xnor
  g1457
  (
    n1470,
    n916,
    n915,
    n995,
    n1054
  );


  xor
  g1458
  (
    n1477,
    n1045,
    n1037,
    n898,
    n859
  );


  and
  g1459
  (
    n1367,
    n1071,
    n833,
    n906,
    n850
  );


  nand
  g1460
  (
    n1310,
    n913,
    n852,
    n854,
    n1025
  );


  nand
  g1461
  (
    n1117,
    n992,
    n797,
    n922,
    n864
  );


  xor
  g1462
  (
    n1276,
    n883,
    n1065,
    n996,
    n907
  );


  and
  g1463
  (
    n1486,
    n910,
    n926,
    n858,
    n846
  );


  or
  g1464
  (
    n1141,
    n871,
    n845,
    n1077,
    n958
  );


  nand
  g1465
  (
    n1224,
    n1014,
    n1048,
    n845,
    n909
  );


  and
  g1466
  (
    n1405,
    n892,
    n1069,
    n1055,
    n904
  );


  xnor
  g1467
  (
    n1195,
    n919,
    n995,
    n907,
    n842
  );


  nor
  g1468
  (
    n1384,
    n848,
    n1027,
    n1058,
    n878
  );


  xor
  g1469
  (
    n1313,
    n855,
    n876,
    n1086,
    n913
  );


  not
  g1470
  (
    n2923,
    n1367
  );


  buf
  g1471
  (
    n2752,
    n1249
  );


  buf
  g1472
  (
    n2199,
    n1371
  );


  buf
  g1473
  (
    n2708,
    n1238
  );


  not
  g1474
  (
    n2699,
    n1236
  );


  buf
  g1475
  (
    n2693,
    n1119
  );


  not
  g1476
  (
    n1844,
    n1290
  );


  not
  g1477
  (
    n2812,
    n1332
  );


  not
  g1478
  (
    n1820,
    n945
  );


  buf
  g1479
  (
    n1858,
    n1296
  );


  buf
  g1480
  (
    n1853,
    n1254
  );


  buf
  g1481
  (
    n2212,
    n1323
  );


  buf
  g1482
  (
    n2616,
    n1131
  );


  buf
  g1483
  (
    n1695,
    n1246
  );


  not
  g1484
  (
    n2328,
    n1261
  );


  not
  g1485
  (
    n1908,
    n1256
  );


  not
  g1486
  (
    n1624,
    n1102
  );


  not
  g1487
  (
    n2494,
    n1410
  );


  not
  g1488
  (
    n2039,
    n1135
  );


  not
  g1489
  (
    n2093,
    n1296
  );


  not
  g1490
  (
    n2889,
    n1102
  );


  not
  g1491
  (
    n2443,
    n1413
  );


  buf
  g1492
  (
    n1718,
    n1106
  );


  not
  g1493
  (
    n2056,
    n1466
  );


  buf
  g1494
  (
    n1726,
    n1126
  );


  not
  g1495
  (
    n2075,
    n1311
  );


  buf
  g1496
  (
    n1637,
    n1125
  );


  not
  g1497
  (
    n2166,
    n1423
  );


  buf
  g1498
  (
    n1724,
    n1255
  );


  buf
  g1499
  (
    n2305,
    n1457
  );


  not
  g1500
  (
    n2054,
    n1419
  );


  not
  g1501
  (
    n1780,
    n1168
  );


  not
  g1502
  (
    n2241,
    n1304
  );


  not
  g1503
  (
    n1770,
    n1194
  );


  buf
  g1504
  (
    n2644,
    n1500
  );


  buf
  g1505
  (
    n1872,
    n1370
  );


  not
  g1506
  (
    n2685,
    n1102
  );


  not
  g1507
  (
    n2163,
    n1411
  );


  buf
  g1508
  (
    n2810,
    n1111
  );


  not
  g1509
  (
    n1921,
    n1143
  );


  buf
  g1510
  (
    n2100,
    n1107
  );


  buf
  g1511
  (
    n1702,
    n1359
  );


  not
  g1512
  (
    n2230,
    n1503
  );


  buf
  g1513
  (
    n2541,
    n1481
  );


  buf
  g1514
  (
    n2769,
    n1161
  );


  buf
  g1515
  (
    n2854,
    n1316
  );


  not
  g1516
  (
    n2485,
    n1153
  );


  buf
  g1517
  (
    n2144,
    n1469
  );


  buf
  g1518
  (
    n2098,
    n1095
  );


  not
  g1519
  (
    n2292,
    n1379
  );


  buf
  g1520
  (
    n2283,
    n1137
  );


  not
  g1521
  (
    n2505,
    n1472
  );


  buf
  g1522
  (
    n2101,
    n1126
  );


  not
  g1523
  (
    n2829,
    n1343
  );


  buf
  g1524
  (
    n2436,
    n1472
  );


  buf
  g1525
  (
    n1936,
    n1216
  );


  buf
  g1526
  (
    n2944,
    n1250
  );


  buf
  g1527
  (
    n1534,
    n758
  );


  not
  g1528
  (
    n2120,
    n1191
  );


  not
  g1529
  (
    n2004,
    n1465
  );


  buf
  g1530
  (
    n2050,
    n1300
  );


  not
  g1531
  (
    KeyWire_0_28,
    n1448
  );


  buf
  g1532
  (
    n2828,
    n1500
  );


  not
  g1533
  (
    n2073,
    n1183
  );


  not
  g1534
  (
    n2891,
    n1229
  );


  not
  g1535
  (
    n2245,
    n1205
  );


  not
  g1536
  (
    n2370,
    n1114
  );


  buf
  g1537
  (
    n2739,
    n1443
  );


  buf
  g1538
  (
    n2216,
    n1369
  );


  not
  g1539
  (
    n1962,
    n1317
  );


  buf
  g1540
  (
    n2387,
    n1342
  );


  buf
  g1541
  (
    n2161,
    n1180
  );


  buf
  g1542
  (
    n2182,
    n1346
  );


  buf
  g1543
  (
    n2574,
    n1226
  );


  not
  g1544
  (
    n2081,
    n1389
  );


  buf
  g1545
  (
    n2643,
    n1493
  );


  buf
  g1546
  (
    n1794,
    n1352
  );


  not
  g1547
  (
    n2326,
    n1436
  );


  not
  g1548
  (
    n1982,
    n1104
  );


  not
  g1549
  (
    n2884,
    n1234
  );


  buf
  g1550
  (
    n2853,
    n1129
  );


  buf
  g1551
  (
    n1738,
    n1294
  );


  not
  g1552
  (
    n2503,
    n1470
  );


  buf
  g1553
  (
    n2400,
    n1150
  );


  buf
  g1554
  (
    n2822,
    n1138
  );


  buf
  g1555
  (
    n2442,
    n1375
  );


  buf
  g1556
  (
    n1697,
    n1345
  );


  not
  g1557
  (
    n1896,
    n1491
  );


  buf
  g1558
  (
    n2607,
    n1217
  );


  buf
  g1559
  (
    n1805,
    n1474
  );


  buf
  g1560
  (
    n2476,
    n1267
  );


  not
  g1561
  (
    n2395,
    n1233
  );


  buf
  g1562
  (
    n2823,
    n1373
  );


  buf
  g1563
  (
    n2730,
    n1141
  );


  not
  g1564
  (
    n1741,
    n1171
  );


  buf
  g1565
  (
    n1958,
    n1470
  );


  buf
  g1566
  (
    n2512,
    n1166
  );


  not
  g1567
  (
    n2169,
    n1502
  );


  not
  g1568
  (
    n1880,
    n1366
  );


  not
  g1569
  (
    n2529,
    n1252
  );


  not
  g1570
  (
    KeyWire_0_12,
    n1092
  );


  buf
  g1571
  (
    n1747,
    n1351
  );


  not
  g1572
  (
    n2521,
    n1103
  );


  buf
  g1573
  (
    n2669,
    n1182
  );


  buf
  g1574
  (
    n2256,
    n1490
  );


  buf
  g1575
  (
    n2229,
    n1282
  );


  buf
  g1576
  (
    n1535,
    n1315
  );


  buf
  g1577
  (
    n1898,
    n1379
  );


  not
  g1578
  (
    n2303,
    n1091
  );


  not
  g1579
  (
    n2630,
    n1091
  );


  not
  g1580
  (
    n2549,
    n1431
  );


  not
  g1581
  (
    n2900,
    n1221
  );


  not
  g1582
  (
    n2536,
    n1450
  );


  buf
  g1583
  (
    n2638,
    n1117
  );


  buf
  g1584
  (
    n2467,
    n1407
  );


  not
  g1585
  (
    n2105,
    n1457
  );


  not
  g1586
  (
    n1745,
    n1220
  );


  not
  g1587
  (
    n2293,
    n1356
  );


  buf
  g1588
  (
    n2573,
    n1187
  );


  buf
  g1589
  (
    n2194,
    n1478
  );


  not
  g1590
  (
    n2817,
    n1142
  );


  buf
  g1591
  (
    n1732,
    n1383
  );


  not
  g1592
  (
    n1949,
    n1321
  );


  not
  g1593
  (
    n2200,
    n1264
  );


  not
  g1594
  (
    n2763,
    n1232
  );


  not
  g1595
  (
    n2294,
    n1178
  );


  buf
  g1596
  (
    n1873,
    n1434
  );


  buf
  g1597
  (
    n2715,
    n1227
  );


  buf
  g1598
  (
    n1801,
    n1495
  );


  buf
  g1599
  (
    n2116,
    n1302
  );


  buf
  g1600
  (
    n2121,
    n1432
  );


  not
  g1601
  (
    n1727,
    n1090
  );


  buf
  g1602
  (
    n2367,
    n1427
  );


  buf
  g1603
  (
    n1803,
    n1208
  );


  not
  g1604
  (
    n1787,
    n1360
  );


  not
  g1605
  (
    n2878,
    n1319
  );


  buf
  g1606
  (
    n2240,
    n1285
  );


  buf
  g1607
  (
    n2402,
    n1492
  );


  not
  g1608
  (
    n2193,
    n1127
  );


  not
  g1609
  (
    n1591,
    n1111
  );


  buf
  g1610
  (
    n2479,
    n1202
  );


  not
  g1611
  (
    n2099,
    n1275
  );


  buf
  g1612
  (
    n1890,
    n1255
  );


  not
  g1613
  (
    n2765,
    n1367
  );


  buf
  g1614
  (
    n2445,
    n1481
  );


  buf
  g1615
  (
    KeyWire_0_15,
    n1274
  );


  buf
  g1616
  (
    n1980,
    n1162
  );


  buf
  g1617
  (
    n1640,
    n1127
  );


  not
  g1618
  (
    n1733,
    n1202
  );


  not
  g1619
  (
    n2041,
    n1365
  );


  not
  g1620
  (
    n2091,
    n1394
  );


  buf
  g1621
  (
    n2185,
    n1349
  );


  buf
  g1622
  (
    n2597,
    n1429
  );


  not
  g1623
  (
    n2351,
    n1373
  );


  not
  g1624
  (
    n2538,
    n1224
  );


  not
  g1625
  (
    n1966,
    n1209
  );


  buf
  g1626
  (
    n1709,
    n1445
  );


  not
  g1627
  (
    n2290,
    n1403
  );


  buf
  g1628
  (
    n1778,
    n1407
  );


  buf
  g1629
  (
    n1541,
    n1251
  );


  not
  g1630
  (
    n2278,
    n1494
  );


  not
  g1631
  (
    n1932,
    n1132
  );


  buf
  g1632
  (
    n2787,
    n1193
  );


  not
  g1633
  (
    n1600,
    n1418
  );


  buf
  g1634
  (
    n1542,
    n1237
  );


  not
  g1635
  (
    n2510,
    n1292
  );


  buf
  g1636
  (
    n1720,
    n1377
  );


  buf
  g1637
  (
    n2309,
    n1422
  );


  buf
  g1638
  (
    n1996,
    n1099
  );


  buf
  g1639
  (
    n2811,
    n1279
  );


  buf
  g1640
  (
    n2352,
    n1274
  );


  buf
  g1641
  (
    n1943,
    n1234
  );


  not
  g1642
  (
    n2393,
    n1187
  );


  not
  g1643
  (
    n2191,
    n1125
  );


  not
  g1644
  (
    n1562,
    n1215
  );


  buf
  g1645
  (
    n2855,
    n1156
  );


  not
  g1646
  (
    n2224,
    n1241
  );


  buf
  g1647
  (
    n2090,
    n1099
  );


  buf
  g1648
  (
    n2672,
    n1323
  );


  not
  g1649
  (
    KeyWire_0_24,
    n1094
  );


  buf
  g1650
  (
    n1598,
    n1156
  );


  not
  g1651
  (
    n1522,
    n1279
  );


  not
  g1652
  (
    n2686,
    n1178
  );


  buf
  g1653
  (
    n1631,
    n1275
  );


  not
  g1654
  (
    n1831,
    n1332
  );


  not
  g1655
  (
    n1836,
    n1378
  );


  buf
  g1656
  (
    n2776,
    n1144
  );


  not
  g1657
  (
    n1776,
    n1354
  );


  not
  g1658
  (
    n2180,
    n1434
  );


  buf
  g1659
  (
    n2474,
    n1484
  );


  buf
  g1660
  (
    n2652,
    n1095
  );


  buf
  g1661
  (
    n2526,
    n1198
  );


  buf
  g1662
  (
    n1626,
    n1100
  );


  buf
  g1663
  (
    n2319,
    n1373
  );


  buf
  g1664
  (
    n1817,
    n1142
  );


  buf
  g1665
  (
    n1603,
    n1158
  );


  not
  g1666
  (
    n1691,
    n1195
  );


  buf
  g1667
  (
    n1516,
    n1486
  );


  buf
  g1668
  (
    n1531,
    n1214
  );


  buf
  g1669
  (
    n2463,
    n1347
  );


  not
  g1670
  (
    n2945,
    n1195
  );


  buf
  g1671
  (
    n2464,
    n1268
  );


  not
  g1672
  (
    n2483,
    n1333
  );


  buf
  g1673
  (
    n2883,
    n1166
  );


  not
  g1674
  (
    n2628,
    n1257
  );


  buf
  g1675
  (
    n2665,
    n1337
  );


  buf
  g1676
  (
    n2846,
    n1343
  );


  buf
  g1677
  (
    n1763,
    n1352
  );


  not
  g1678
  (
    n2710,
    n1476
  );


  not
  g1679
  (
    n1582,
    n1203
  );


  not
  g1680
  (
    n1886,
    n1334
  );


  buf
  g1681
  (
    n2767,
    n1362
  );


  not
  g1682
  (
    n1795,
    n744
  );


  not
  g1683
  (
    n2653,
    n1394
  );


  not
  g1684
  (
    n2800,
    n1201
  );


  not
  g1685
  (
    n2928,
    n1167
  );


  buf
  g1686
  (
    n2189,
    n1276
  );


  not
  g1687
  (
    n2178,
    n1287
  );


  buf
  g1688
  (
    KeyWire_0_21,
    n1417
  );


  buf
  g1689
  (
    n2190,
    n1328
  );


  not
  g1690
  (
    n2488,
    n1195
  );


  buf
  g1691
  (
    n2288,
    n1335
  );


  buf
  g1692
  (
    n1586,
    n1281
  );


  buf
  g1693
  (
    n2655,
    n1204
  );


  not
  g1694
  (
    n2789,
    n1459
  );


  buf
  g1695
  (
    n2729,
    n1105
  );


  not
  g1696
  (
    n2097,
    n1335
  );


  buf
  g1697
  (
    n2297,
    n1262
  );


  buf
  g1698
  (
    n1760,
    n1338
  );


  not
  g1699
  (
    n2219,
    n1322
  );


  not
  g1700
  (
    n2143,
    n1217
  );


  buf
  g1701
  (
    n2357,
    n1154
  );


  not
  g1702
  (
    n2355,
    n1208
  );


  buf
  g1703
  (
    n2439,
    n1299
  );


  not
  g1704
  (
    n1604,
    n1256
  );


  buf
  g1705
  (
    n2542,
    n1165
  );


  not
  g1706
  (
    n2602,
    n1302
  );


  not
  g1707
  (
    n2028,
    n1318
  );


  buf
  g1708
  (
    n2580,
    n1217
  );


  buf
  g1709
  (
    n2816,
    n1397
  );


  buf
  g1710
  (
    n2223,
    n1331
  );


  not
  g1711
  (
    n2210,
    n1315
  );


  buf
  g1712
  (
    n1951,
    n1247
  );


  buf
  g1713
  (
    n2718,
    n1238
  );


  buf
  g1714
  (
    n1781,
    n1172
  );


  buf
  g1715
  (
    n2704,
    n1414
  );


  buf
  g1716
  (
    n1566,
    n1462
  );


  not
  g1717
  (
    n2493,
    n1156
  );


  buf
  g1718
  (
    n1926,
    n1188
  );


  buf
  g1719
  (
    n1986,
    n1500
  );


  buf
  g1720
  (
    n1601,
    n1194
  );


  not
  g1721
  (
    n1707,
    n1184
  );


  buf
  g1722
  (
    n1749,
    n1109
  );


  buf
  g1723
  (
    n2943,
    n1496
  );


  buf
  g1724
  (
    n1569,
    n1327
  );


  not
  g1725
  (
    n1532,
    n1151
  );


  buf
  g1726
  (
    n2057,
    n1193
  );


  buf
  g1727
  (
    n2372,
    n1112
  );


  not
  g1728
  (
    n2936,
    n1295
  );


  not
  g1729
  (
    n1656,
    n1112
  );


  buf
  g1730
  (
    n2598,
    n1414
  );


  not
  g1731
  (
    n1889,
    n1242
  );


  not
  g1732
  (
    n2455,
    n1312
  );


  buf
  g1733
  (
    n2373,
    n743
  );


  not
  g1734
  (
    n2796,
    n1467
  );


  not
  g1735
  (
    n1617,
    n1263
  );


  buf
  g1736
  (
    n1554,
    n1463
  );


  buf
  g1737
  (
    n2660,
    n1497
  );


  buf
  g1738
  (
    n2871,
    n1347
  );


  buf
  g1739
  (
    n1857,
    n1116
  );


  not
  g1740
  (
    n1620,
    n1491
  );


  buf
  g1741
  (
    n2264,
    n1101
  );


  not
  g1742
  (
    n2566,
    n1472
  );


  not
  g1743
  (
    n2209,
    n1104
  );


  not
  g1744
  (
    n2786,
    n1409
  );


  not
  g1745
  (
    n2504,
    n1289
  );


  buf
  g1746
  (
    n2452,
    n1337
  );


  buf
  g1747
  (
    n2024,
    n1321
  );


  not
  g1748
  (
    n2807,
    n1394
  );


  not
  g1749
  (
    n1929,
    n1230
  );


  not
  g1750
  (
    n2938,
    n1391
  );


  buf
  g1751
  (
    n2000,
    n1368
  );


  buf
  g1752
  (
    n2712,
    n1468
  );


  buf
  g1753
  (
    n2226,
    n1126
  );


  buf
  g1754
  (
    n2501,
    n1418
  );


  buf
  g1755
  (
    n2301,
    n1474
  );


  buf
  g1756
  (
    n1708,
    n1246
  );


  not
  g1757
  (
    n2904,
    n755
  );


  not
  g1758
  (
    n2777,
    n1434
  );


  buf
  g1759
  (
    n2155,
    n1272
  );


  not
  g1760
  (
    n1988,
    n1296
  );


  buf
  g1761
  (
    n1648,
    n1299
  );


  not
  g1762
  (
    n1550,
    n1138
  );


  not
  g1763
  (
    n1610,
    n1437
  );


  not
  g1764
  (
    n2696,
    n1107
  );


  buf
  g1765
  (
    n2124,
    n1396
  );


  not
  g1766
  (
    n1662,
    n1331
  );


  buf
  g1767
  (
    n1616,
    n1381
  );


  not
  g1768
  (
    n2341,
    n1240
  );


  buf
  g1769
  (
    n2023,
    n1309
  );


  not
  g1770
  (
    n2629,
    n1432
  );


  buf
  g1771
  (
    n2137,
    n1180
  );


  not
  g1772
  (
    n1901,
    n1162
  );


  not
  g1773
  (
    n2403,
    n1165
  );


  buf
  g1774
  (
    n2614,
    n1180
  );


  not
  g1775
  (
    n2286,
    n1318
  );


  not
  g1776
  (
    n1997,
    n1330
  );


  not
  g1777
  (
    n2595,
    n1471
  );


  buf
  g1778
  (
    n1979,
    n1236
  );


  not
  g1779
  (
    n2415,
    n1357
  );


  not
  g1780
  (
    n2103,
    n1154
  );


  buf
  g1781
  (
    n1536,
    n1181
  );


  buf
  g1782
  (
    n2579,
    n1210
  );


  buf
  g1783
  (
    n2324,
    n1295
  );


  not
  g1784
  (
    n2379,
    n1101
  );


  buf
  g1785
  (
    n2697,
    n1301
  );


  buf
  g1786
  (
    n2077,
    n1131
  );


  not
  g1787
  (
    n2336,
    n1321
  );


  buf
  g1788
  (
    n1928,
    n1260
  );


  not
  g1789
  (
    n1814,
    n1110
  );


  not
  g1790
  (
    n1521,
    n1451
  );


  buf
  g1791
  (
    n2658,
    n1448
  );


  not
  g1792
  (
    n2572,
    n1257
  );


  buf
  g1793
  (
    n1838,
    n1489
  );


  not
  g1794
  (
    n2497,
    n1175
  );


  buf
  g1795
  (
    n2533,
    n1326
  );


  buf
  g1796
  (
    n1694,
    n1269
  );


  buf
  g1797
  (
    n2071,
    n1147
  );


  buf
  g1798
  (
    n1903,
    n1122
  );


  not
  g1799
  (
    n1677,
    n1090
  );


  buf
  g1800
  (
    n2555,
    n1205
  );


  not
  g1801
  (
    n2847,
    n1250
  );


  buf
  g1802
  (
    n1835,
    n1481
  );


  not
  g1803
  (
    n2411,
    n1292
  );


  not
  g1804
  (
    n2620,
    n1093
  );


  buf
  g1805
  (
    n1735,
    n1124
  );


  not
  g1806
  (
    n1692,
    n1160
  );


  buf
  g1807
  (
    n2480,
    n1174
  );


  buf
  g1808
  (
    n1578,
    n1458
  );


  not
  g1809
  (
    n1852,
    n1182
  );


  not
  g1810
  (
    n2437,
    n1327
  );


  not
  g1811
  (
    n2170,
    n1240
  );


  buf
  g1812
  (
    n2779,
    n1315
  );


  buf
  g1813
  (
    n2895,
    n1340
  );


  not
  g1814
  (
    n2306,
    n1278
  );


  not
  g1815
  (
    n2175,
    n1396
  );


  buf
  g1816
  (
    n1555,
    n1265
  );


  buf
  g1817
  (
    n2640,
    n1336
  );


  buf
  g1818
  (
    n2197,
    n1486
  );


  buf
  g1819
  (
    n1827,
    n1321
  );


  buf
  g1820
  (
    n2112,
    n752
  );


  buf
  g1821
  (
    n2903,
    n1103
  );


  buf
  g1822
  (
    n2364,
    n1341
  );


  buf
  g1823
  (
    n2864,
    n1288
  );


  buf
  g1824
  (
    n2618,
    n1255
  );


  not
  g1825
  (
    n2388,
    n1356
  );


  not
  g1826
  (
    n2666,
    n1208
  );


  buf
  g1827
  (
    n1676,
    n1224
  );


  buf
  g1828
  (
    n2405,
    n1479
  );


  not
  g1829
  (
    n1792,
    n1370
  );


  not
  g1830
  (
    n2211,
    n1259
  );


  buf
  g1831
  (
    n1682,
    n1161
  );


  not
  g1832
  (
    n1788,
    n1294
  );


  buf
  g1833
  (
    n1995,
    n1189
  );


  not
  g1834
  (
    n2322,
    n1316
  );


  buf
  g1835
  (
    n2583,
    n1171
  );


  not
  g1836
  (
    n2850,
    n1376
  );


  buf
  g1837
  (
    n2140,
    n1122
  );


  buf
  g1838
  (
    n2570,
    n1388
  );


  not
  g1839
  (
    n2773,
    n1410
  );


  not
  g1840
  (
    n1529,
    n1397
  );


  buf
  g1841
  (
    n1973,
    n1173
  );


  not
  g1842
  (
    n1866,
    n1416
  );


  not
  g1843
  (
    n2361,
    n1311
  );


  buf
  g1844
  (
    n2296,
    n1409
  );


  not
  g1845
  (
    n2065,
    n1279
  );


  not
  g1846
  (
    n2253,
    n1150
  );


  not
  g1847
  (
    n2042,
    n1359
  );


  buf
  g1848
  (
    n2856,
    n1403
  );


  not
  g1849
  (
    n2742,
    n1340
  );


  not
  g1850
  (
    n2375,
    n1358
  );


  buf
  g1851
  (
    n2478,
    n1355
  );


  buf
  g1852
  (
    n1681,
    n1094
  );


  not
  g1853
  (
    n2734,
    n1242
  );


  not
  g1854
  (
    n1574,
    n1258
  );


  buf
  g1855
  (
    n1629,
    n1370
  );


  buf
  g1856
  (
    n2601,
    n1367
  );


  not
  g1857
  (
    n2695,
    n1169
  );


  buf
  g1858
  (
    n1525,
    n1479
  );


  not
  g1859
  (
    n2744,
    n1242
  );


  buf
  g1860
  (
    n1567,
    n1183
  );


  not
  g1861
  (
    n1742,
    n1322
  );


  not
  g1862
  (
    n1905,
    n1101
  );


  not
  g1863
  (
    n2410,
    n1312
  );


  not
  g1864
  (
    n2179,
    n1172
  );


  buf
  g1865
  (
    n2063,
    n1459
  );


  buf
  g1866
  (
    n1875,
    n1351
  );


  not
  g1867
  (
    n2876,
    n1234
  );


  buf
  g1868
  (
    n1751,
    n1488
  );


  not
  g1869
  (
    n2337,
    n1203
  );


  buf
  g1870
  (
    n1800,
    n1460
  );


  not
  g1871
  (
    n2225,
    n1105
  );


  buf
  g1872
  (
    n2756,
    n1278
  );


  buf
  g1873
  (
    n1613,
    n1265
  );


  not
  g1874
  (
    n1714,
    n1117
  );


  buf
  g1875
  (
    n1641,
    n1447
  );


  not
  g1876
  (
    n1878,
    n1271
  );


  buf
  g1877
  (
    n1678,
    n1436
  );


  buf
  g1878
  (
    n2320,
    n1130
  );


  buf
  g1879
  (
    n2758,
    n1272
  );


  buf
  g1880
  (
    n1607,
    n1349
  );


  not
  g1881
  (
    n1548,
    n1265
  );


  not
  g1882
  (
    n2298,
    n1397
  );


  not
  g1883
  (
    n1659,
    n1476
  );


  not
  g1884
  (
    n2381,
    n1369
  );


  not
  g1885
  (
    n2743,
    n1424
  );


  buf
  g1886
  (
    n1867,
    n1420
  );


  buf
  g1887
  (
    KeyWire_0_25,
    n1408
  );


  buf
  g1888
  (
    n2915,
    n1387
  );


  not
  g1889
  (
    n1918,
    n1459
  );


  buf
  g1890
  (
    n2171,
    n1158
  );


  buf
  g1891
  (
    n1605,
    n1221
  );


  not
  g1892
  (
    n1925,
    n1375
  );


  not
  g1893
  (
    n2051,
    n1442
  );


  buf
  g1894
  (
    n1736,
    n1152
  );


  buf
  g1895
  (
    n1762,
    n1231
  );


  buf
  g1896
  (
    n1619,
    n1206
  );


  buf
  g1897
  (
    n1560,
    n1288
  );


  buf
  g1898
  (
    n1618,
    n1416
  );


  not
  g1899
  (
    n1876,
    n1345
  );


  not
  g1900
  (
    n2887,
    n1197
  );


  buf
  g1901
  (
    n2668,
    n1185
  );


  buf
  g1902
  (
    n2899,
    n1349
  );


  not
  g1903
  (
    n1654,
    n1189
  );


  buf
  g1904
  (
    n2490,
    n1250
  );


  buf
  g1905
  (
    KeyWire_0_20,
    n1365
  );


  not
  g1906
  (
    n2236,
    n1432
  );


  buf
  g1907
  (
    n2088,
    n1422
  );


  buf
  g1908
  (
    n2457,
    n1339
  );


  buf
  g1909
  (
    n2867,
    n1310
  );


  buf
  g1910
  (
    n1609,
    n1176
  );


  buf
  g1911
  (
    n2596,
    n1437
  );


  not
  g1912
  (
    n2362,
    n1311
  );


  not
  g1913
  (
    n1859,
    n1333
  );


  buf
  g1914
  (
    n2879,
    n1471
  );


  not
  g1915
  (
    n2425,
    n1467
  );


  buf
  g1916
  (
    n1796,
    n1291
  );


  not
  g1917
  (
    n2208,
    n1477
  );


  not
  g1918
  (
    n2724,
    n1334
  );


  not
  g1919
  (
    n2006,
    n1423
  );


  buf
  g1920
  (
    n2913,
    n1253
  );


  not
  g1921
  (
    n2839,
    n1268
  );


  buf
  g1922
  (
    n2513,
    n1395
  );


  buf
  g1923
  (
    n1954,
    n1172
  );


  buf
  g1924
  (
    n2397,
    n1447
  );


  buf
  g1925
  (
    n2550,
    n1232
  );


  buf
  g1926
  (
    n1759,
    n1451
  );


  buf
  g1927
  (
    n2238,
    n1443
  );


  buf
  g1928
  (
    n2432,
    n1243
  );


  not
  g1929
  (
    n1571,
    n1136
  );


  not
  g1930
  (
    n1734,
    n1164
  );


  not
  g1931
  (
    n1664,
    n1504
  );


  not
  g1932
  (
    n2207,
    n1429
  );


  buf
  g1933
  (
    n1899,
    n1465
  );


  buf
  g1934
  (
    n2295,
    n1384
  );


  buf
  g1935
  (
    n2213,
    n1342
  );


  not
  g1936
  (
    n2183,
    n1353
  );


  not
  g1937
  (
    n2522,
    n1308
  );


  not
  g1938
  (
    n2792,
    n1422
  );


  not
  g1939
  (
    n1930,
    n1456
  );


  not
  g1940
  (
    n2688,
    n1319
  );


  buf
  g1941
  (
    n2637,
    n1501
  );


  not
  g1942
  (
    n2645,
    n1403
  );


  not
  g1943
  (
    n2918,
    n1179
  );


  buf
  g1944
  (
    n2118,
    n1445
  );


  not
  g1945
  (
    n1777,
    n1481
  );


  buf
  g1946
  (
    n2621,
    n1475
  );


  buf
  g1947
  (
    n2263,
    n1114
  );


  not
  g1948
  (
    n2131,
    n1228
  );


  not
  g1949
  (
    n2237,
    n1121
  );


  buf
  g1950
  (
    n2506,
    n1128
  );


  buf
  g1951
  (
    n2473,
    n1109
  );


  buf
  g1952
  (
    n1723,
    n1302
  );


  buf
  g1953
  (
    n1753,
    n1346
  );


  buf
  g1954
  (
    n1790,
    n1207
  );


  not
  g1955
  (
    n2577,
    n1189
  );


  not
  g1956
  (
    n2070,
    n1121
  );


  not
  g1957
  (
    n1960,
    n1316
  );


  not
  g1958
  (
    n2138,
    n1153
  );


  not
  g1959
  (
    n2592,
    n1305
  );


  not
  g1960
  (
    n2673,
    n1360
  );


  buf
  g1961
  (
    n2424,
    n1176
  );


  buf
  g1962
  (
    n1539,
    n1502
  );


  buf
  g1963
  (
    n2611,
    n1245
  );


  buf
  g1964
  (
    n2428,
    n1384
  );


  not
  g1965
  (
    n2429,
    n1258
  );


  buf
  g1966
  (
    n1766,
    n1092
  );


  not
  g1967
  (
    n1863,
    n1436
  );


  buf
  g1968
  (
    n2085,
    n1387
  );


  not
  g1969
  (
    n1684,
    n1493
  );


  not
  g1970
  (
    n2080,
    n1443
  );


  not
  g1971
  (
    n1552,
    n1420
  );


  buf
  g1972
  (
    n1860,
    n1263
  );


  not
  g1973
  (
    n2087,
    n1492
  );


  not
  g1974
  (
    n2126,
    n1407
  );


  not
  g1975
  (
    n1842,
    n1234
  );


  not
  g1976
  (
    n2222,
    n1473
  );


  not
  g1977
  (
    n2196,
    n1423
  );


  buf
  g1978
  (
    n1608,
    n1219
  );


  buf
  g1979
  (
    n2029,
    n1263
  );


  not
  g1980
  (
    n2165,
    n1276
  );


  not
  g1981
  (
    n2654,
    n1128
  );


  not
  g1982
  (
    n2593,
    n1438
  );


  buf
  g1983
  (
    n2881,
    n1501
  );


  not
  g1984
  (
    n2114,
    n1371
  );


  buf
  g1985
  (
    n1511,
    n1301
  );


  buf
  g1986
  (
    n2444,
    n1292
  );


  not
  g1987
  (
    n2349,
    n1330
  );


  buf
  g1988
  (
    n2308,
    n1341
  );


  buf
  g1989
  (
    n2935,
    n1313
  );


  buf
  g1990
  (
    n1666,
    n1104
  );


  not
  g1991
  (
    n2279,
    n1097
  );


  buf
  g1992
  (
    n2865,
    n1218
  );


  buf
  g1993
  (
    n1957,
    n1450
  );


  not
  g1994
  (
    n2287,
    n1291
  );


  buf
  g1995
  (
    n2670,
    n1491
  );


  buf
  g1996
  (
    n1826,
    n1380
  );


  not
  g1997
  (
    n1639,
    n1241
  );


  buf
  g1998
  (
    n1512,
    n1287
  );


  not
  g1999
  (
    n1611,
    n1407
  );


  buf
  g2000
  (
    n2426,
    n1308
  );


  buf
  g2001
  (
    n1865,
    n1303
  );


  not
  g2002
  (
    n1785,
    n1133
  );


  buf
  g2003
  (
    n1965,
    n1203
  );


  not
  g2004
  (
    n2026,
    n1306
  );


  not
  g2005
  (
    n2342,
    n1090
  );


  buf
  g2006
  (
    n2698,
    n1141
  );


  not
  g2007
  (
    n1602,
    n1278
  );


  buf
  g2008
  (
    n2667,
    n1408
  );


  buf
  g2009
  (
    n1775,
    n1499
  );


  buf
  g2010
  (
    n2396,
    n1276
  );


  buf
  g2011
  (
    n1750,
    n1272
  );


  buf
  g2012
  (
    n2391,
    n1162
  );


  not
  g2013
  (
    n2262,
    n1235
  );


  buf
  g2014
  (
    n2774,
    n1490
  );


  buf
  g2015
  (
    n2509,
    n1456
  );


  buf
  g2016
  (
    n2458,
    n1320
  );


  not
  g2017
  (
    n1944,
    n1185
  );


  not
  g2018
  (
    n2824,
    n1108
  );


  buf
  g2019
  (
    n2939,
    n1119
  );


  buf
  g2020
  (
    n2782,
    n1469
  );


  not
  g2021
  (
    n2886,
    n1093
  );


  not
  g2022
  (
    n1769,
    n1427
  );


  not
  g2023
  (
    n2684,
    n1129
  );


  not
  g2024
  (
    n2383,
    n1158
  );


  not
  g2025
  (
    n2151,
    n1361
  );


  buf
  g2026
  (
    n1523,
    n1342
  );


  buf
  g2027
  (
    n2033,
    n1167
  );


  not
  g2028
  (
    n2076,
    n1287
  );


  not
  g2029
  (
    n2427,
    n1433
  );


  not
  g2030
  (
    n2877,
    n1444
  );


  buf
  g2031
  (
    n2221,
    n1350
  );


  buf
  g2032
  (
    n2551,
    n1157
  );


  not
  g2033
  (
    n2117,
    n1289
  );


  not
  g2034
  (
    n2735,
    n1261
  );


  buf
  g2035
  (
    n2567,
    n1413
  );


  not
  g2036
  (
    n2858,
    n1396
  );


  buf
  g2037
  (
    n1513,
    n1094
  );


  buf
  g2038
  (
    n1924,
    n1148
  );


  buf
  g2039
  (
    n2502,
    n1203
  );


  not
  g2040
  (
    n2896,
    n1271
  );


  not
  g2041
  (
    n2079,
    n748
  );


  not
  g2042
  (
    n2150,
    n1372
  );


  not
  g2043
  (
    n2941,
    n1397
  );


  not
  g2044
  (
    n1825,
    n1453
  );


  not
  g2045
  (
    n1894,
    n1120
  );


  not
  g2046
  (
    n2167,
    n1236
  );


  buf
  g2047
  (
    n2046,
    n1222
  );


  not
  g2048
  (
    n1871,
    n1458
  );


  not
  g2049
  (
    n1969,
    n1276
  );


  buf
  g2050
  (
    n1597,
    n1404
  );


  buf
  g2051
  (
    n2047,
    n1412
  );


  buf
  g2052
  (
    n2157,
    n1292
  );


  not
  g2053
  (
    n1856,
    n1475
  );


  not
  g2054
  (
    n2683,
    n1504
  );


  buf
  g2055
  (
    n2930,
    n1307
  );


  not
  g2056
  (
    n1855,
    n1495
  );


  buf
  g2057
  (
    n2032,
    n1212
  );


  buf
  g2058
  (
    n1900,
    n1448
  );


  not
  g2059
  (
    n1565,
    n1291
  );


  not
  g2060
  (
    n1689,
    n1320
  );


  buf
  g2061
  (
    n1704,
    n1199
  );


  not
  g2062
  (
    n2300,
    n1283
  );


  buf
  g2063
  (
    n2450,
    n1176
  );


  buf
  g2064
  (
    n2691,
    n1107
  );


  buf
  g2065
  (
    n1947,
    n1290
  );


  buf
  g2066
  (
    n1757,
    n1425
  );


  buf
  g2067
  (
    n2746,
    n1265
  );


  not
  g2068
  (
    n2713,
    n1361
  );


  not
  g2069
  (
    n2017,
    n1199
  );


  not
  g2070
  (
    n2946,
    n1156
  );


  not
  g2071
  (
    n2560,
    n1213
  );


  buf
  g2072
  (
    n1799,
    n1226
  );


  not
  g2073
  (
    n2492,
    n1229
  );


  not
  g2074
  (
    n1985,
    n1209
  );


  not
  g2075
  (
    n1804,
    n1322
  );


  not
  g2076
  (
    n2408,
    n1248
  );


  buf
  g2077
  (
    n2419,
    n1406
  );


  not
  g2078
  (
    n2423,
    n1285
  );


  not
  g2079
  (
    n2417,
    n1196
  );


  buf
  g2080
  (
    n1927,
    n1152
  );


  buf
  g2081
  (
    n1625,
    n1358
  );


  not
  g2082
  (
    n2109,
    n1454
  );


  not
  g2083
  (
    n2471,
    n1189
  );


  buf
  g2084
  (
    n2347,
    n1115
  );


  not
  g2085
  (
    n2626,
    n1318
  );


  not
  g2086
  (
    n1614,
    n1307
  );


  buf
  g2087
  (
    n2631,
    n1134
  );


  not
  g2088
  (
    n2358,
    n1288
  );


  not
  g2089
  (
    n2612,
    n1098
  );


  not
  g2090
  (
    n1862,
    n1293
  );


  buf
  g2091
  (
    n2385,
    n1162
  );


  not
  g2092
  (
    n2721,
    n1260
  );


  buf
  g2093
  (
    n2244,
    n1173
  );


  buf
  g2094
  (
    n1893,
    n1464
  );


  buf
  g2095
  (
    n2826,
    n1500
  );


  buf
  g2096
  (
    n2663,
    n1124
  );


  buf
  g2097
  (
    n2078,
    n753
  );


  not
  g2098
  (
    n2518,
    n1177
  );


  not
  g2099
  (
    KeyWire_0_0,
    n1229
  );


  not
  g2100
  (
    n1612,
    n1446
  );


  not
  g2101
  (
    n1711,
    n1431
  );


  buf
  g2102
  (
    n2258,
    n1155
  );


  buf
  g2103
  (
    n1514,
    n1411
  );


  buf
  g2104
  (
    n1646,
    n1480
  );


  not
  g2105
  (
    n2246,
    n1425
  );


  not
  g2106
  (
    n1774,
    n1400
  );


  not
  g2107
  (
    n2281,
    n754
  );


  buf
  g2108
  (
    n1716,
    n1489
  );


  not
  g2109
  (
    n2359,
    n1324
  );


  not
  g2110
  (
    n2761,
    n1307
  );


  buf
  g2111
  (
    n2627,
    n1401
  );


  not
  g2112
  (
    n2162,
    n1132
  );


  buf
  g2113
  (
    n2239,
    n1131
  );


  buf
  g2114
  (
    n2345,
    n1283
  );


  not
  g2115
  (
    n2753,
    n1350
  );


  buf
  g2116
  (
    n1885,
    n1426
  );


  buf
  g2117
  (
    n2511,
    n1290
  );


  not
  g2118
  (
    n2872,
    n1479
  );


  buf
  g2119
  (
    n2482,
    n756
  );


  not
  g2120
  (
    n2642,
    n1171
  );


  buf
  g2121
  (
    n2553,
    n1277
  );


  not
  g2122
  (
    n2142,
    n1186
  );


  not
  g2123
  (
    n1561,
    n1275
  );


  not
  g2124
  (
    n1623,
    n1497
  );


  buf
  g2125
  (
    n2354,
    n1406
  );


  not
  g2126
  (
    n2802,
    n1412
  );


  not
  g2127
  (
    n2418,
    n1229
  );


  not
  g2128
  (
    n1789,
    n1391
  );


  buf
  g2129
  (
    n2366,
    n1462
  );


  not
  g2130
  (
    n1904,
    n1184
  );


  buf
  g2131
  (
    n1728,
    n1424
  );


  not
  g2132
  (
    n2153,
    n1482
  );


  not
  g2133
  (
    n2556,
    n1301
  );


  buf
  g2134
  (
    n2885,
    n1226
  );


  buf
  g2135
  (
    n2610,
    n1120
  );


  buf
  g2136
  (
    n2465,
    n1478
  );


  not
  g2137
  (
    n2333,
    n745
  );


  not
  g2138
  (
    n1764,
    n1144
  );


  not
  g2139
  (
    n2716,
    n1194
  );


  not
  g2140
  (
    n2043,
    n1465
  );


  not
  g2141
  (
    n2331,
    n1129
  );


  not
  g2142
  (
    n1994,
    n1293
  );


  not
  g2143
  (
    n1948,
    n1329
  );


  buf
  g2144
  (
    n1978,
    n1105
  );


  not
  g2145
  (
    n1647,
    n1213
  );


  not
  g2146
  (
    n2067,
    n1446
  );


  not
  g2147
  (
    n2624,
    n1357
  );


  not
  g2148
  (
    n1710,
    n1468
  );


  buf
  g2149
  (
    n2745,
    n1096
  );


  not
  g2150
  (
    n2527,
    n1474
  );


  not
  g2151
  (
    n2815,
    n1134
  );


  not
  g2152
  (
    n2737,
    n1379
  );


  not
  g2153
  (
    n1668,
    n1167
  );


  buf
  g2154
  (
    n2532,
    n1355
  );


  not
  g2155
  (
    n2316,
    n1477
  );


  buf
  g2156
  (
    n1848,
    n1369
  );


  not
  g2157
  (
    n1746,
    n1447
  );


  not
  g2158
  (
    n1821,
    n1328
  );


  not
  g2159
  (
    n2948,
    n1257
  );


  buf
  g2160
  (
    n2852,
    n1439
  );


  not
  g2161
  (
    n1690,
    n1149
  );


  buf
  g2162
  (
    n2917,
    n1391
  );


  not
  g2163
  (
    n1808,
    n1428
  );


  buf
  g2164
  (
    n1740,
    n1471
  );


  buf
  g2165
  (
    n1627,
    n1148
  );


  not
  g2166
  (
    n2537,
    n1410
  );


  not
  g2167
  (
    n1705,
    n1411
  );


  not
  g2168
  (
    n2590,
    n1478
  );


  buf
  g2169
  (
    n1851,
    n1264
  );


  not
  g2170
  (
    n1971,
    n1145
  );


  not
  g2171
  (
    n2731,
    n1459
  );


  buf
  g2172
  (
    n2430,
    n1464
  );


  buf
  g2173
  (
    n2035,
    n1489
  );


  not
  g2174
  (
    n2340,
    n1210
  );


  buf
  g2175
  (
    n2055,
    n1169
  );


  not
  g2176
  (
    n2108,
    n1331
  );


  not
  g2177
  (
    n1675,
    n1418
  );


  not
  g2178
  (
    n1665,
    n1490
  );


  buf
  g2179
  (
    n2520,
    n1409
  );


  not
  g2180
  (
    n2656,
    n1165
  );


  buf
  g2181
  (
    n1606,
    n1259
  );


  buf
  g2182
  (
    n2269,
    n1483
  );


  not
  g2183
  (
    n2096,
    n1467
  );


  buf
  g2184
  (
    KeyWire_0_16,
    n1461
  );


  buf
  g2185
  (
    n2875,
    n1289
  );


  not
  g2186
  (
    n2384,
    n1122
  );


  not
  g2187
  (
    n2636,
    n1365
  );


  not
  g2188
  (
    n1595,
    n1117
  );


  not
  g2189
  (
    n2146,
    n1341
  );


  not
  g2190
  (
    n1791,
    n1304
  );


  buf
  g2191
  (
    n1955,
    n1103
  );


  not
  g2192
  (
    n1888,
    n1145
  );


  not
  g2193
  (
    n2282,
    n1303
  );


  not
  g2194
  (
    n1829,
    n1104
  );


  not
  g2195
  (
    n1528,
    n1451
  );


  not
  g2196
  (
    n2129,
    n1103
  );


  not
  g2197
  (
    n1509,
    n1116
  );


  not
  g2198
  (
    n1592,
    n1366
  );


  buf
  g2199
  (
    n2844,
    n1468
  );


  not
  g2200
  (
    n2330,
    n1378
  );


  not
  g2201
  (
    n2931,
    n1306
  );


  buf
  g2202
  (
    n1919,
    n1427
  );


  buf
  g2203
  (
    n2793,
    n1362
  );


  not
  g2204
  (
    n2217,
    n1259
  );


  not
  g2205
  (
    n2940,
    n1175
  );


  buf
  g2206
  (
    n1628,
    n1360
  );


  not
  g2207
  (
    n2818,
    n1320
  );


  not
  g2208
  (
    n2353,
    n949
  );


  buf
  g2209
  (
    n1946,
    n1406
  );


  buf
  g2210
  (
    n2016,
    n1423
  );


  buf
  g2211
  (
    n2898,
    n1452
  );


  not
  g2212
  (
    n1722,
    n1127
  );


  not
  g2213
  (
    n2849,
    n1357
  );


  buf
  g2214
  (
    n2481,
    n1212
  );


  buf
  g2215
  (
    n1583,
    n1128
  );


  buf
  g2216
  (
    n2662,
    n1332
  );


  not
  g2217
  (
    n2307,
    n1483
  );


  buf
  g2218
  (
    n2104,
    n1364
  );


  buf
  g2219
  (
    n1968,
    n1295
  );


  buf
  g2220
  (
    n2186,
    n1501
  );


  not
  g2221
  (
    n2912,
    n1456
  );


  not
  g2222
  (
    n1621,
    n1327
  );


  buf
  g2223
  (
    n2469,
    n1151
  );


  not
  g2224
  (
    n1599,
    n1294
  );


  buf
  g2225
  (
    n1588,
    n1503
  );


  not
  g2226
  (
    n1630,
    n1303
  );


  not
  g2227
  (
    n2472,
    n1192
  );


  buf
  g2228
  (
    n2231,
    n1137
  );


  buf
  g2229
  (
    n2181,
    n1148
  );


  buf
  g2230
  (
    n2534,
    n1415
  );


  buf
  g2231
  (
    n1992,
    n1197
  );


  not
  g2232
  (
    n1941,
    n1338
  );


  buf
  g2233
  (
    n2312,
    n1113
  );


  buf
  g2234
  (
    n2634,
    n1105
  );


  buf
  g2235
  (
    n1655,
    n1186
  );


  not
  g2236
  (
    n2335,
    n1262
  );


  not
  g2237
  (
    n1884,
    n1223
  );


  not
  g2238
  (
    n2271,
    n1190
  );


  not
  g2239
  (
    n2814,
    n1504
  );


  buf
  g2240
  (
    n2382,
    n1446
  );


  buf
  g2241
  (
    n2559,
    n1492
  );


  buf
  g2242
  (
    n2188,
    n1417
  );


  buf
  g2243
  (
    n2926,
    n1215
  );


  not
  g2244
  (
    n1510,
    n1419
  );


  buf
  g2245
  (
    n2438,
    n1280
  );


  not
  g2246
  (
    n1593,
    n1486
  );


  buf
  g2247
  (
    n1622,
    n1159
  );


  not
  g2248
  (
    n2496,
    n1308
  );


  buf
  g2249
  (
    n2072,
    n1390
  );


  not
  g2250
  (
    n1674,
    n1121
  );


  buf
  g2251
  (
    n2001,
    n1251
  );


  not
  g2252
  (
    n1538,
    n1484
  );


  buf
  g2253
  (
    n1897,
    n1138
  );


  buf
  g2254
  (
    n2413,
    n1436
  );


  buf
  g2255
  (
    n2617,
    n1386
  );


  buf
  g2256
  (
    n1843,
    n1108
  );


  not
  g2257
  (
    n1515,
    n1238
  );


  buf
  g2258
  (
    n1633,
    n1288
  );


  not
  g2259
  (
    n1696,
    n1225
  );


  not
  g2260
  (
    n2013,
    n1140
  );


  not
  g2261
  (
    n1549,
    n1416
  );


  not
  g2262
  (
    n2275,
    n1359
  );


  not
  g2263
  (
    n2622,
    n1220
  );


  not
  g2264
  (
    n1524,
    n1226
  );


  buf
  g2265
  (
    n1840,
    n1309
  );


  not
  g2266
  (
    n1570,
    n1477
  );


  buf
  g2267
  (
    n2257,
    n1334
  );


  not
  g2268
  (
    n2819,
    n1193
  );


  not
  g2269
  (
    n1652,
    n1116
  );


  not
  g2270
  (
    n2859,
    n1317
  );


  not
  g2271
  (
    n2920,
    n1404
  );


  buf
  g2272
  (
    n2921,
    n1304
  );


  not
  g2273
  (
    n1573,
    n1277
  );


  buf
  g2274
  (
    n2156,
    n1282
  );


  buf
  g2275
  (
    n2249,
    n1445
  );


  not
  g2276
  (
    n1772,
    n1243
  );


  buf
  g2277
  (
    n2798,
    n1101
  );


  buf
  g2278
  (
    n2933,
    n1413
  );


  buf
  g2279
  (
    n2005,
    n1297
  );


  not
  g2280
  (
    n2768,
    n1206
  );


  not
  g2281
  (
    n1748,
    n1354
  );


  buf
  g2282
  (
    n2568,
    n1179
  );


  buf
  g2283
  (
    n2148,
    n1273
  );


  not
  g2284
  (
    n1956,
    n1193
  );


  buf
  g2285
  (
    n1934,
    n1426
  );


  not
  g2286
  (
    n1877,
    n1327
  );


  not
  g2287
  (
    n2646,
    n1257
  );


  buf
  g2288
  (
    n2632,
    n1244
  );


  buf
  g2289
  (
    n2111,
    n1493
  );


  not
  g2290
  (
    n2299,
    n1463
  );


  buf
  g2291
  (
    n2014,
    n1191
  );


  not
  g2292
  (
    n1998,
    n1424
  );


  buf
  g2293
  (
    n2475,
    n1433
  );


  not
  g2294
  (
    n2044,
    n1314
  );


  not
  g2295
  (
    n2795,
    n1228
  );


  not
  g2296
  (
    n2198,
    n1386
  );


  not
  g2297
  (
    n2897,
    n1116
  );


  buf
  g2298
  (
    n2007,
    n1454
  );


  not
  g2299
  (
    n2414,
    n1441
  );


  not
  g2300
  (
    n2581,
    n1348
  );


  not
  g2301
  (
    n1717,
    n1223
  );


  buf
  g2302
  (
    n2924,
    n1381
  );


  buf
  g2303
  (
    n2563,
    n1114
  );


  not
  g2304
  (
    n2902,
    n1184
  );


  not
  g2305
  (
    n2564,
    n1446
  );


  buf
  g2306
  (
    n1937,
    n1453
  );


  not
  g2307
  (
    n2003,
    n1094
  );


  not
  g2308
  (
    n2441,
    n1106
  );


  not
  g2309
  (
    n2220,
    n1190
  );


  not
  g2310
  (
    n1784,
    n1449
  );


  buf
  g2311
  (
    n1923,
    n1207
  );


  not
  g2312
  (
    n1916,
    n1244
  );


  buf
  g2313
  (
    n2343,
    n1198
  );


  buf
  g2314
  (
    n1911,
    n1222
  );


  buf
  g2315
  (
    n2435,
    n1246
  );


  buf
  g2316
  (
    n1910,
    n1426
  );


  buf
  g2317
  (
    n2242,
    n1341
  );


  not
  g2318
  (
    n2546,
    n1285
  );


  buf
  g2319
  (
    n1822,
    n1233
  );


  not
  g2320
  (
    n1587,
    n1137
  );


  not
  g2321
  (
    n2569,
    n1166
  );


  not
  g2322
  (
    n1797,
    n1262
  );


  buf
  g2323
  (
    n2508,
    n1487
  );


  not
  g2324
  (
    n1712,
    n1419
  );


  buf
  g2325
  (
    n2516,
    n1198
  );


  not
  g2326
  (
    n2113,
    n1099
  );


  buf
  g2327
  (
    n2582,
    n1235
  );


  buf
  g2328
  (
    n2594,
    n1112
  );


  not
  g2329
  (
    n1984,
    n1111
  );


  buf
  g2330
  (
    n2535,
    n1480
  );


  buf
  g2331
  (
    n2325,
    n1221
  );


  not
  g2332
  (
    n2377,
    n1412
  );


  buf
  g2333
  (
    n2722,
    n1470
  );


  buf
  g2334
  (
    n1658,
    n1351
  );


  buf
  g2335
  (
    n2135,
    n1118
  );


  not
  g2336
  (
    n2031,
    n1261
  );


  not
  g2337
  (
    n2647,
    n1387
  );


  buf
  g2338
  (
    n2929,
    n1499
  );


  buf
  g2339
  (
    n2762,
    n1139
  );


  buf
  g2340
  (
    n1981,
    n1177
  );


  not
  g2341
  (
    n2407,
    n1389
  );


  not
  g2342
  (
    n2780,
    n1209
  );


  not
  g2343
  (
    n2368,
    n1488
  );


  not
  g2344
  (
    n2749,
    n1329
  );


  not
  g2345
  (
    n1518,
    n1297
  );


  not
  g2346
  (
    n2030,
    n1421
  );


  not
  g2347
  (
    n1577,
    n1354
  );


  buf
  g2348
  (
    n2804,
    n946
  );


  buf
  g2349
  (
    n1508,
    n1437
  );


  buf
  g2350
  (
    n2952,
    n1335
  );


  not
  g2351
  (
    n2820,
    n1241
  );


  not
  g2352
  (
    n1783,
    n1334
  );


  buf
  g2353
  (
    n1963,
    n1339
  );


  not
  g2354
  (
    n2784,
    n1505
  );


  buf
  g2355
  (
    n2204,
    n749
  );


  buf
  g2356
  (
    n2736,
    n1503
  );


  buf
  g2357
  (
    n2778,
    n1196
  );


  buf
  g2358
  (
    n2565,
    n1482
  );


  buf
  g2359
  (
    n1807,
    n1269
  );


  buf
  g2360
  (
    n1752,
    n1386
  );


  buf
  g2361
  (
    n2813,
    n1473
  );


  buf
  g2362
  (
    n2421,
    n1499
  );


  buf
  g2363
  (
    n2115,
    n1097
  );


  not
  g2364
  (
    n2701,
    n1106
  );


  not
  g2365
  (
    n1959,
    n1393
  );


  not
  g2366
  (
    n1558,
    n1095
  );


  not
  g2367
  (
    n2950,
    n1350
  );


  not
  g2368
  (
    n2932,
    n1204
  );


  not
  g2369
  (
    n2908,
    n1183
  );


  buf
  g2370
  (
    n2619,
    n1375
  );


  buf
  g2371
  (
    n2870,
    n1387
  );


  buf
  g2372
  (
    n2557,
    n1225
  );


  buf
  g2373
  (
    n1729,
    n1421
  );


  buf
  g2374
  (
    n2022,
    n1208
  );


  buf
  g2375
  (
    n2727,
    n750
  );


  not
  g2376
  (
    n1744,
    n1335
  );


  not
  g2377
  (
    n1719,
    n1157
  );


  buf
  g2378
  (
    n2376,
    n1209
  );


  buf
  g2379
  (
    n1557,
    n1382
  );


  buf
  g2380
  (
    n2390,
    n1244
  );


  not
  g2381
  (
    n2747,
    n1173
  );


  buf
  g2382
  (
    n1942,
    n1239
  );


  buf
  g2383
  (
    n2315,
    n1155
  );


  buf
  g2384
  (
    n2801,
    n1123
  );


  buf
  g2385
  (
    n2010,
    n1133
  );


  not
  g2386
  (
    n2661,
    n1159
  );


  buf
  g2387
  (
    n1935,
    n1361
  );


  not
  g2388
  (
    n1667,
    n1132
  );


  buf
  g2389
  (
    n1828,
    n1204
  );


  not
  g2390
  (
    n1615,
    n1278
  );


  not
  g2391
  (
    n2329,
    n1380
  );


  buf
  g2392
  (
    n1809,
    n1460
  );


  buf
  g2393
  (
    n2547,
    n1143
  );


  buf
  g2394
  (
    n2446,
    n1360
  );


  not
  g2395
  (
    n2552,
    n1337
  );


  not
  g2396
  (
    n1931,
    n1470
  );


  buf
  g2397
  (
    n1638,
    n1457
  );


  buf
  g2398
  (
    n2095,
    n1236
  );


  buf
  g2399
  (
    n2754,
    n1270
  );


  buf
  g2400
  (
    n2466,
    n1425
  );


  not
  g2401
  (
    n2291,
    n1476
  );


  buf
  g2402
  (
    n1887,
    n1168
  );


  buf
  g2403
  (
    n2657,
    n1151
  );


  buf
  g2404
  (
    n1643,
    n1143
  );


  not
  g2405
  (
    n2159,
    n1345
  );


  buf
  g2406
  (
    n1756,
    n1164
  );


  buf
  g2407
  (
    n2401,
    n1205
  );


  buf
  g2408
  (
    n1771,
    n1224
  );


  not
  g2409
  (
    n2909,
    n1487
  );


  not
  g2410
  (
    n1861,
    n1149
  );


  not
  g2411
  (
    n2461,
    n1169
  );


  not
  g2412
  (
    n1670,
    n1133
  );


  not
  g2413
  (
    n1779,
    n1496
  );


  not
  g2414
  (
    n1758,
    n1495
  );


  buf
  g2415
  (
    n2680,
    n1431
  );


  buf
  g2416
  (
    n1964,
    n1333
  );


  buf
  g2417
  (
    n2927,
    n1422
  );


  buf
  g2418
  (
    n2470,
    n1128
  );


  buf
  g2419
  (
    n2059,
    n1285
  );


  not
  g2420
  (
    n1649,
    n1259
  );


  buf
  g2421
  (
    n2227,
    n1115
  );


  not
  g2422
  (
    n2600,
    n1126
  );


  not
  g2423
  (
    n2709,
    n1175
  );


  not
  g2424
  (
    n2832,
    n1364
  );


  not
  g2425
  (
    n2498,
    n1372
  );


  not
  g2426
  (
    n2060,
    n1273
  );


  not
  g2427
  (
    n2766,
    n1120
  );


  not
  g2428
  (
    n1642,
    n1290
  );


  buf
  g2429
  (
    n2803,
    n1252
  );


  buf
  g2430
  (
    n2623,
    n1157
  );


  not
  g2431
  (
    n2679,
    n1158
  );


  buf
  g2432
  (
    n2251,
    n1349
  );


  not
  g2433
  (
    n2456,
    n1248
  );


  not
  g2434
  (
    n1879,
    n1402
  );


  buf
  g2435
  (
    n1874,
    n1451
  );


  buf
  g2436
  (
    n2788,
    n1198
  );


  buf
  g2437
  (
    n2528,
    n1399
  );


  buf
  g2438
  (
    n2916,
    n1380
  );


  not
  g2439
  (
    n1739,
    n1326
  );


  buf
  g2440
  (
    n1824,
    n1196
  );


  not
  g2441
  (
    n2515,
    n1249
  );


  not
  g2442
  (
    n2845,
    n1443
  );


  not
  g2443
  (
    n2133,
    n1373
  );


  not
  g2444
  (
    n1895,
    n1232
  );


  not
  g2445
  (
    n1933,
    n1306
  );


  not
  g2446
  (
    n2588,
    n1113
  );


  buf
  g2447
  (
    n1868,
    n1462
  );


  not
  g2448
  (
    n2084,
    n1181
  );


  not
  g2449
  (
    n2525,
    n1475
  );


  buf
  g2450
  (
    n2717,
    n1320
  );


  not
  g2451
  (
    n1909,
    n1096
  );


  not
  g2452
  (
    n2232,
    n1441
  );


  buf
  g2453
  (
    n1519,
    n1450
  );


  buf
  g2454
  (
    n2651,
    n1284
  );


  not
  g2455
  (
    n2173,
    n1164
  );


  not
  g2456
  (
    n2857,
    n1453
  );


  buf
  g2457
  (
    n2489,
    n1331
  );


  buf
  g2458
  (
    n2276,
    n1440
  );


  buf
  g2459
  (
    n2821,
    n1417
  );


  buf
  g2460
  (
    n2523,
    n1228
  );


  buf
  g2461
  (
    n2019,
    n1281
  );


  not
  g2462
  (
    n2422,
    n1140
  );


  not
  g2463
  (
    n1520,
    n1342
  );


  not
  g2464
  (
    n2843,
    n1318
  );


  not
  g2465
  (
    n1833,
    n1227
  );


  buf
  g2466
  (
    n1517,
    n1444
  );


  not
  g2467
  (
    n2514,
    n1129
  );


  buf
  g2468
  (
    n2702,
    n1277
  );


  not
  g2469
  (
    n2720,
    n1188
  );


  not
  g2470
  (
    n2139,
    n1139
  );


  buf
  g2471
  (
    n1699,
    n1454
  );


  not
  g2472
  (
    n2615,
    n1200
  );


  buf
  g2473
  (
    n1673,
    n1371
  );


  buf
  g2474
  (
    n1912,
    n1192
  );


  buf
  g2475
  (
    n1556,
    n1314
  );


  buf
  g2476
  (
    n1703,
    n1132
  );


  not
  g2477
  (
    n2350,
    n1330
  );


  not
  g2478
  (
    n2834,
    n1496
  );


  not
  g2479
  (
    n2248,
    n1237
  );


  buf
  g2480
  (
    n2507,
    n1348
  );


  not
  g2481
  (
    n2554,
    n1398
  );


  buf
  g2482
  (
    n1830,
    n1480
  );


  not
  g2483
  (
    n2284,
    n1472
  );


  buf
  g2484
  (
    n1812,
    n1220
  );


  buf
  g2485
  (
    n2205,
    n1169
  );


  buf
  g2486
  (
    n2741,
    n1431
  );


  not
  g2487
  (
    n2036,
    n1274
  );


  not
  g2488
  (
    n2906,
    n1395
  );


  not
  g2489
  (
    n2433,
    n1145
  );


  buf
  g2490
  (
    n1891,
    n1213
  );


  buf
  g2491
  (
    n2740,
    n1406
  );


  not
  g2492
  (
    n2910,
    n1235
  );


  buf
  g2493
  (
    n2842,
    n1439
  );


  buf
  g2494
  (
    n1553,
    n1283
  );


  buf
  g2495
  (
    n2771,
    n1161
  );


  not
  g2496
  (
    n2015,
    n1264
  );


  buf
  g2497
  (
    n2706,
    n1098
  );


  not
  g2498
  (
    n2321,
    n1346
  );


  not
  g2499
  (
    n2049,
    n1297
  );


  buf
  g2500
  (
    n2833,
    n1252
  );


  not
  g2501
  (
    n1713,
    n1113
  );


  buf
  g2502
  (
    n1914,
    n1190
  );


  not
  g2503
  (
    n2835,
    n1179
  );


  buf
  g2504
  (
    n2705,
    n1147
  );


  buf
  g2505
  (
    n2311,
    n1223
  );


  not
  g2506
  (
    n2202,
    n1400
  );


  buf
  g2507
  (
    n2893,
    n1336
  );


  buf
  g2508
  (
    n1902,
    n1417
  );


  buf
  g2509
  (
    n2711,
    n1420
  );


  not
  g2510
  (
    n1813,
    n1247
  );


  buf
  g2511
  (
    n2589,
    n1386
  );


  buf
  g2512
  (
    n2561,
    n1165
  );


  buf
  g2513
  (
    n2726,
    n1249
  );


  not
  g2514
  (
    n1645,
    n1311
  );


  buf
  g2515
  (
    n1506,
    n1219
  );


  buf
  g2516
  (
    n2434,
    n1286
  );


  buf
  g2517
  (
    n1698,
    n1146
  );


  not
  g2518
  (
    n2677,
    n1494
  );


  not
  g2519
  (
    n1672,
    n1497
  );


  not
  g2520
  (
    n2892,
    n1130
  );


  buf
  g2521
  (
    n1754,
    n1297
  );


  not
  g2522
  (
    n1815,
    n1328
  );


  buf
  g2523
  (
    n2544,
    n1485
  );


  buf
  g2524
  (
    n2136,
    n1442
  );


  not
  g2525
  (
    n1564,
    n1171
  );


  buf
  g2526
  (
    n1802,
    n1204
  );


  not
  g2527
  (
    n2270,
    n1218
  );


  not
  g2528
  (
    n1685,
    n1181
  );


  not
  g2529
  (
    n2045,
    n1214
  );


  buf
  g2530
  (
    n1693,
    n1498
  );


  not
  g2531
  (
    n2951,
    n1433
  );


  buf
  g2532
  (
    n2468,
    n1438
  );


  buf
  g2533
  (
    n2584,
    n1174
  );


  buf
  g2534
  (
    n1584,
    n1307
  );


  not
  g2535
  (
    n2453,
    n1255
  );


  buf
  g2536
  (
    n1989,
    n1281
  );


  not
  g2537
  (
    n1987,
    n1091
  );


  buf
  g2538
  (
    n2603,
    n1227
  );


  buf
  g2539
  (
    n2639,
    n1399
  );


  buf
  g2540
  (
    n2332,
    n1505
  );


  buf
  g2541
  (
    n2243,
    n1385
  );


  buf
  g2542
  (
    n1967,
    n1279
  );


  buf
  g2543
  (
    n2781,
    n1217
  );


  not
  g2544
  (
    n2831,
    n1376
  );


  buf
  g2545
  (
    n2002,
    n1170
  );


  not
  g2546
  (
    n1846,
    n1461
  );


  buf
  g2547
  (
    n1761,
    n1478
  );


  buf
  g2548
  (
    n1687,
    n1402
  );


  buf
  g2549
  (
    n2274,
    n1391
  );


  buf
  g2550
  (
    n2025,
    n1383
  );


  not
  g2551
  (
    n2040,
    n1190
  );


  not
  g2552
  (
    n2323,
    n1445
  );


  buf
  g2553
  (
    n1938,
    n1298
  );


  buf
  g2554
  (
    n2228,
    n1161
  );


  buf
  g2555
  (
    n1773,
    n1177
  );


  buf
  g2556
  (
    n2317,
    n1271
  );


  not
  g2557
  (
    n1547,
    n1237
  );


  not
  g2558
  (
    n2947,
    n1352
  );


  buf
  g2559
  (
    n2123,
    n1108
  );


  not
  g2560
  (
    n2723,
    n1487
  );


  buf
  g2561
  (
    n1533,
    n1344
  );


  buf
  g2562
  (
    n2591,
    n1230
  );


  buf
  g2563
  (
    n2459,
    n1200
  );


  buf
  g2564
  (
    n1585,
    n1140
  );


  not
  g2565
  (
    n2911,
    n1383
  );


  buf
  g2566
  (
    n1743,
    n1344
  );


  not
  g2567
  (
    n2531,
    n1145
  );


  not
  g2568
  (
    n2234,
    n1244
  );


  not
  g2569
  (
    n1635,
    n1358
  );


  buf
  g2570
  (
    n2676,
    n1106
  );


  not
  g2571
  (
    n1819,
    n1293
  );


  buf
  g2572
  (
    n2339,
    n1477
  );


  buf
  g2573
  (
    n2808,
    n1142
  );


  buf
  g2574
  (
    n2690,
    n1170
  );


  not
  g2575
  (
    n1590,
    n1310
  );


  buf
  g2576
  (
    n2371,
    n1399
  );


  buf
  g2577
  (
    n2280,
    n1268
  );


  not
  g2578
  (
    n2641,
    n1139
  );


  buf
  g2579
  (
    n1661,
    n1159
  );


  buf
  g2580
  (
    n2250,
    n1118
  );


  not
  g2581
  (
    n2868,
    n1463
  );


  not
  g2582
  (
    n2083,
    n1310
  );


  buf
  g2583
  (
    n2094,
    n1353
  );


  not
  g2584
  (
    n2692,
    n1253
  );


  buf
  g2585
  (
    n2725,
    n1458
  );


  not
  g2586
  (
    n2119,
    n1207
  );


  buf
  g2587
  (
    n2447,
    n1212
  );


  buf
  g2588
  (
    n1999,
    n1466
  );


  buf
  g2589
  (
    n1977,
    n1404
  );


  buf
  g2590
  (
    n1634,
    n1429
  );


  not
  g2591
  (
    n2477,
    n1480
  );


  buf
  g2592
  (
    n2406,
    n1220
  );


  not
  g2593
  (
    n2548,
    n1225
  );


  not
  g2594
  (
    n2374,
    n1464
  );


  not
  g2595
  (
    n2922,
    n1322
  );


  buf
  g2596
  (
    n2107,
    n1233
  );


  buf
  g2597
  (
    n2703,
    n1254
  );


  not
  g2598
  (
    n2874,
    n1488
  );


  not
  g2599
  (
    n2841,
    n1272
  );


  buf
  g2600
  (
    n2604,
    n1504
  );


  buf
  g2601
  (
    n2034,
    n1450
  );


  buf
  g2602
  (
    n1864,
    n1280
  );


  buf
  g2603
  (
    n2266,
    n1484
  );


  buf
  g2604
  (
    n2235,
    n1214
  );


  not
  g2605
  (
    n1993,
    n1092
  );


  buf
  g2606
  (
    n2174,
    n1130
  );


  buf
  g2607
  (
    n2334,
    n1238
  );


  not
  g2608
  (
    n2764,
    n1280
  );


  not
  g2609
  (
    n1854,
    n1124
  );


  buf
  g2610
  (
    n2195,
    n1231
  );


  not
  g2611
  (
    n2412,
    n1424
  );


  not
  g2612
  (
    n1847,
    n1401
  );


  buf
  g2613
  (
    n2149,
    n1374
  );


  not
  g2614
  (
    n2608,
    n1338
  );


  not
  g2615
  (
    n1688,
    n1258
  );


  not
  g2616
  (
    n2517,
    n1163
  );


  not
  g2617
  (
    n2942,
    n1442
  );


  buf
  g2618
  (
    n2491,
    n1141
  );


  not
  g2619
  (
    n2562,
    n1211
  );


  not
  g2620
  (
    n2086,
    n1395
  );


  buf
  g2621
  (
    n2369,
    n1420
  );


  not
  g2622
  (
    n2318,
    n1235
  );


  not
  g2623
  (
    n2285,
    n1294
  );


  not
  g2624
  (
    n1651,
    n1362
  );


  not
  g2625
  (
    n2187,
    n1332
  );


  buf
  g2626
  (
    n2145,
    n1216
  );


  not
  g2627
  (
    n2011,
    n1384
  );


  buf
  g2628
  (
    n2389,
    n1444
  );


  buf
  g2629
  (
    n2168,
    n1484
  );


  buf
  g2630
  (
    n2649,
    n1108
  );


  not
  g2631
  (
    n2775,
    n1379
  );


  buf
  g2632
  (
    n1544,
    n1385
  );


  not
  g2633
  (
    n1755,
    n759
  );


  not
  g2634
  (
    n2420,
    n1403
  );


  not
  g2635
  (
    n2356,
    n1393
  );


  buf
  g2636
  (
    n2338,
    n1222
  );


  buf
  g2637
  (
    n2484,
    n1394
  );


  not
  g2638
  (
    n1940,
    n1122
  );


  not
  g2639
  (
    n2122,
    n1298
  );


  buf
  g2640
  (
    n2609,
    n1110
  );


  not
  g2641
  (
    n2252,
    n1270
  );


  not
  g2642
  (
    n1632,
    n1141
  );


  buf
  g2643
  (
    n1581,
    n1497
  );


  buf
  g2644
  (
    n2215,
    n1329
  );


  buf
  g2645
  (
    n2650,
    n1125
  );


  not
  g2646
  (
    n2386,
    n1385
  );


  not
  g2647
  (
    n2018,
    n1097
  );


  buf
  g2648
  (
    n2495,
    n1356
  );


  not
  g2649
  (
    n2265,
    n1201
  );


  buf
  g2650
  (
    n1970,
    n1398
  );


  not
  g2651
  (
    n2585,
    n1152
  );


  buf
  g2652
  (
    n1952,
    n1344
  );


  buf
  g2653
  (
    n2048,
    n1348
  );


  not
  g2654
  (
    n2837,
    n1136
  );


  buf
  g2655
  (
    n2134,
    n1491
  );


  not
  g2656
  (
    n1881,
    n757
  );


  buf
  g2657
  (
    n2206,
    n1317
  );


  not
  g2658
  (
    n2606,
    n1306
  );


  not
  g2659
  (
    n2869,
    n1218
  );


  buf
  g2660
  (
    n2327,
    n1392
  );


  not
  g2661
  (
    n2659,
    n1210
  );


  not
  g2662
  (
    KeyWire_0_14,
    n1309
  );


  buf
  g2663
  (
    n1701,
    n1118
  );


  buf
  g2664
  (
    n1976,
    n1323
  );


  buf
  g2665
  (
    n2543,
    n1475
  );


  buf
  g2666
  (
    n2037,
    n1183
  );


  buf
  g2667
  (
    n1540,
    n1233
  );


  buf
  g2668
  (
    n2635,
    n1095
  );


  buf
  g2669
  (
    n2755,
    n1201
  );


  not
  g2670
  (
    n2102,
    n1154
  );


  not
  g2671
  (
    n1636,
    n1345
  );


  buf
  g2672
  (
    n2344,
    n1383
  );


  buf
  g2673
  (
    n2838,
    n1498
  );


  not
  g2674
  (
    n2027,
    n1469
  );


  buf
  g2675
  (
    n2066,
    n1246
  );


  not
  g2676
  (
    n1580,
    n1347
  );


  buf
  g2677
  (
    n1983,
    n1159
  );


  not
  g2678
  (
    n2571,
    n1227
  );


  buf
  g2679
  (
    n1915,
    n1415
  );


  not
  g2680
  (
    n2448,
    n1377
  );


  buf
  g2681
  (
    n2404,
    n1365
  );


  buf
  g2682
  (
    n2880,
    n1201
  );


  not
  g2683
  (
    n2141,
    n1187
  );


  not
  g2684
  (
    n1551,
    n1415
  );


  buf
  g2685
  (
    n2728,
    n1402
  );


  buf
  g2686
  (
    n2068,
    n1325
  );


  buf
  g2687
  (
    n2760,
    n1471
  );


  buf
  g2688
  (
    n2348,
    n1134
  );


  not
  g2689
  (
    n1527,
    n1401
  );


  buf
  g2690
  (
    n1507,
    n1185
  );


  not
  g2691
  (
    n2176,
    n1134
  );


  not
  g2692
  (
    n1782,
    n1142
  );


  not
  g2693
  (
    n2799,
    n1135
  );


  not
  g2694
  (
    n1806,
    n1375
  );


  buf
  g2695
  (
    n1882,
    n1260
  );


  buf
  g2696
  (
    n2530,
    n1400
  );


  not
  g2697
  (
    n2254,
    n1293
  );


  buf
  g2698
  (
    n2578,
    n1115
  );


  not
  g2699
  (
    n2061,
    n1316
  );


  buf
  g2700
  (
    n2794,
    n1414
  );


  not
  g2701
  (
    n2462,
    n1267
  );


  buf
  g2702
  (
    n1870,
    n1372
  );


  not
  g2703
  (
    n2092,
    n1273
  );


  not
  g2704
  (
    n2267,
    n1153
  );


  buf
  g2705
  (
    n2451,
    n1389
  );


  buf
  g2706
  (
    n1793,
    n1219
  );


  not
  g2707
  (
    n2154,
    n1155
  );


  not
  g2708
  (
    n2613,
    n1150
  );


  buf
  g2709
  (
    n2089,
    n1430
  );


  not
  g2710
  (
    n2380,
    n1392
  );


  not
  g2711
  (
    n2790,
    n1485
  );


  buf
  g2712
  (
    n2313,
    n1296
  );


  not
  g2713
  (
    n2689,
    n1207
  );


  not
  g2714
  (
    n2203,
    n1333
  );


  not
  g2715
  (
    n2934,
    n1433
  );


  not
  g2716
  (
    n2247,
    n1200
  );


  not
  g2717
  (
    n1653,
    n1398
  );


  buf
  g2718
  (
    n2772,
    n1300
  );


  not
  g2719
  (
    n1768,
    n1469
  );


  not
  g2720
  (
    n1596,
    n1147
  );


  buf
  g2721
  (
    n2949,
    n1388
  );


  not
  g2722
  (
    n2192,
    n1271
  );


  buf
  g2723
  (
    n1991,
    n1249
  );


  buf
  g2724
  (
    n2860,
    n1168
  );


  not
  g2725
  (
    n2128,
    n1438
  );


  not
  g2726
  (
    n2750,
    n1111
  );


  not
  g2727
  (
    n2805,
    n1239
  );


  buf
  g2728
  (
    n1730,
    n1428
  );


  not
  g2729
  (
    n2147,
    n1231
  );


  buf
  g2730
  (
    n2218,
    n1369
  );


  not
  g2731
  (
    n2836,
    n1269
  );


  not
  g2732
  (
    n2738,
    n1182
  );


  buf
  g2733
  (
    n2009,
    n1427
  );


  not
  g2734
  (
    n2398,
    n1289
  );


  not
  g2735
  (
    n2272,
    n1305
  );


  not
  g2736
  (
    n2863,
    n1123
  );


  not
  g2737
  (
    n1650,
    n1444
  );


  not
  g2738
  (
    n1545,
    n1137
  );


  buf
  g2739
  (
    n1841,
    n1273
  );


  buf
  g2740
  (
    n1765,
    n1270
  );


  not
  g2741
  (
    n2848,
    n1438
  );


  buf
  g2742
  (
    n1660,
    n1460
  );


  not
  g2743
  (
    n1737,
    n1176
  );


  not
  g2744
  (
    n2201,
    n1473
  );


  not
  g2745
  (
    n1945,
    n1160
  );


  not
  g2746
  (
    n1950,
    n1411
  );


  buf
  g2747
  (
    n2392,
    n1237
  );


  buf
  g2748
  (
    n1953,
    n1239
  );


  buf
  g2749
  (
    n1849,
    n1366
  );


  not
  g2750
  (
    n1834,
    n1344
  );


  not
  g2751
  (
    n2082,
    n1266
  );


  buf
  g2752
  (
    n2487,
    n1256
  );


  buf
  g2753
  (
    n2757,
    n1213
  );


  not
  g2754
  (
    n2882,
    n751
  );


  buf
  g2755
  (
    n2233,
    n1184
  );


  buf
  g2756
  (
    n2785,
    n1425
  );


  not
  g2757
  (
    n2255,
    n1185
  );


  not
  g2758
  (
    n1883,
    n1317
  );


  not
  g2759
  (
    n2901,
    n1264
  );


  buf
  g2760
  (
    n2851,
    n1251
  );


  buf
  g2761
  (
    n2012,
    n1354
  );


  buf
  g2762
  (
    n1572,
    n1457
  );


  buf
  g2763
  (
    n2289,
    n1465
  );


  buf
  g2764
  (
    n2440,
    n1347
  );


  not
  g2765
  (
    n2273,
    n1352
  );


  not
  g2766
  (
    n2416,
    n1202
  );


  not
  g2767
  (
    n2925,
    n1143
  );


  buf
  g2768
  (
    n1839,
    n1096
  );


  buf
  g2769
  (
    n2460,
    n1483
  );


  not
  g2770
  (
    n2519,
    n1179
  );


  not
  g2771
  (
    n2346,
    n1300
  );


  buf
  g2772
  (
    n2177,
    n1270
  );


  buf
  g2773
  (
    n2587,
    n1170
  );


  not
  g2774
  (
    n2454,
    n1197
  );


  buf
  g2775
  (
    n2132,
    n1282
  );


  not
  g2776
  (
    n2919,
    n1300
  );


  not
  g2777
  (
    n1706,
    n1100
  );


  buf
  g2778
  (
    n1939,
    n1426
  );


  buf
  g2779
  (
    n2671,
    n1127
  );


  not
  g2780
  (
    n2674,
    n1133
  );


  not
  g2781
  (
    n2558,
    n1340
  );


  not
  g2782
  (
    n2733,
    n747
  );


  buf
  g2783
  (
    n2791,
    n1241
  );


  not
  g2784
  (
    n1669,
    n1371
  );


  buf
  g2785
  (
    n2399,
    n1266
  );


  not
  g2786
  (
    n1644,
    n1363
  );


  buf
  g2787
  (
    n1906,
    n1146
  );


  buf
  g2788
  (
    n2052,
    n1467
  );


  not
  g2789
  (
    n2158,
    n1494
  );


  buf
  g2790
  (
    KeyWire_0_9,
    n1214
  );


  not
  g2791
  (
    n2675,
    n1196
  );


  not
  g2792
  (
    n2605,
    n1440
  );


  buf
  g2793
  (
    n1913,
    n1100
  );


  buf
  g2794
  (
    n2625,
    n1112
  );


  buf
  g2795
  (
    n1683,
    n1195
  );


  not
  g2796
  (
    n2021,
    n1199
  );


  buf
  g2797
  (
    n2540,
    n1151
  );


  not
  g2798
  (
    n2363,
    n1455
  );


  not
  g2799
  (
    n2304,
    n1388
  );


  buf
  g2800
  (
    n1832,
    n1372
  );


  not
  g2801
  (
    n1594,
    n1256
  );


  buf
  g2802
  (
    n1568,
    n1305
  );


  not
  g2803
  (
    n2064,
    n1153
  );


  buf
  g2804
  (
    n2069,
    n1430
  );


  not
  g2805
  (
    n2873,
    n1242
  );


  buf
  g2806
  (
    n2888,
    n1343
  );


  not
  g2807
  (
    n2314,
    n1197
  );


  buf
  g2808
  (
    n1530,
    n1305
  );


  not
  g2809
  (
    n2020,
    n1324
  );


  not
  g2810
  (
    n2214,
    n1148
  );


  buf
  g2811
  (
    n1563,
    n1368
  );


  buf
  g2812
  (
    n2937,
    n1188
  );


  buf
  g2813
  (
    n2310,
    n1295
  );


  buf
  g2814
  (
    n2110,
    n1222
  );


  buf
  g2815
  (
    n2809,
    n1495
  );


  buf
  g2816
  (
    n2861,
    n1174
  );


  buf
  g2817
  (
    n1810,
    n1218
  );


  buf
  g2818
  (
    n2866,
    n1168
  );


  not
  g2819
  (
    n2806,
    n1326
  );


  not
  g2820
  (
    n1837,
    n1366
  );


  buf
  g2821
  (
    n2127,
    n1339
  );


  buf
  g2822
  (
    n2008,
    n1370
  );


  buf
  g2823
  (
    n2074,
    n1206
  );


  buf
  g2824
  (
    n1922,
    n1390
  );


  not
  g2825
  (
    n1700,
    n1224
  );


  not
  g2826
  (
    n1798,
    n1498
  );


  buf
  g2827
  (
    n2714,
    n1415
  );


  buf
  g2828
  (
    n1907,
    n1435
  );


  not
  g2829
  (
    n2694,
    n1359
  );


  not
  g2830
  (
    n1990,
    n1434
  );


  not
  g2831
  (
    n2707,
    n746
  );


  not
  g2832
  (
    n1543,
    n1337
  );


  not
  g2833
  (
    n1657,
    n1125
  );


  buf
  g2834
  (
    n2164,
    n1138
  );


  buf
  g2835
  (
    n2905,
    n1376
  );


  buf
  g2836
  (
    n1823,
    n1319
  );


  xor
  g2837
  (
    n2682,
    n1362,
    n1303,
    n1313
  );


  xor
  g2838
  (
    n1546,
    n1339,
    n1382,
    n1392,
    n1329
  );


  xor
  g2839
  (
    n2748,
    n1374,
    n1413,
    n1378,
    n1325
  );


  nand
  g2840
  (
    n1721,
    n1378,
    n1463,
    n1419,
    n1247
  );


  xnor
  g2841
  (
    n2053,
    n1262,
    n1254,
    n1152,
    n1368
  );


  xnor
  g2842
  (
    n1818,
    n1118,
    n1408,
    n1343,
    n1200
  );


  and
  g2843
  (
    n1917,
    n1286,
    n1430,
    n1228,
    n1231
  );


  nor
  g2844
  (
    n2106,
    n1247,
    n1385,
    n1144,
    n1473
  );


  xor
  g2845
  (
    n2681,
    n1199,
    n1405,
    n1123,
    n1248
  );


  xor
  g2846
  (
    n1845,
    n1187,
    n1091,
    n1455,
    n1485
  );


  xor
  g2847
  (
    n2062,
    n1323,
    n1314,
    n1263,
    n1390
  );


  nand
  g2848
  (
    n2125,
    n1476,
    n1312,
    n1486,
    n1440
  );


  xor
  g2849
  (
    n2524,
    n1251,
    n1319,
    n1099,
    n1166
  );


  xnor
  g2850
  (
    n2261,
    n1429,
    n1435,
    n1358,
    n1266
  );


  and
  g2851
  (
    n2268,
    n1502,
    n1421,
    n1282,
    n1402
  );


  nor
  g2852
  (
    n2797,
    n1330,
    n1191,
    n1215,
    n1211
  );


  or
  g2853
  (
    n1892,
    n1230,
    n1455,
    n1496,
    n1109
  );


  and
  g2854
  (
    n2751,
    n1192,
    n1268,
    n1284,
    n1348
  );


  xor
  g2855
  (
    n1920,
    n1312,
    n1452,
    n1350,
    n1377
  );


  or
  g2856
  (
    n2770,
    n1121,
    n1401,
    n1328,
    n1150
  );


  or
  g2857
  (
    n2783,
    n1167,
    n1474,
    n1325,
    n1163
  );


  nand
  g2858
  (
    n2825,
    n1174,
    n1490,
    n1340,
    n1131
  );


  xor
  g2859
  (
    n2058,
    n1240,
    n1109,
    n1314,
    n1376
  );


  nand
  g2860
  (
    n1575,
    n1186,
    n1449,
    n1170,
    n1405
  );


  xnor
  g2861
  (
    n2365,
    n1277,
    n1194,
    n1499,
    n1448
  );


  xnor
  g2862
  (
    n1680,
    n1435,
    n1177,
    n1102,
    n1501
  );


  and
  g2863
  (
    n2545,
    n1418,
    n1113,
    n1462,
    n1291
  );


  and
  g2864
  (
    n2038,
    n1304,
    n1136,
    n1178,
    n1180
  );


  xor
  g2865
  (
    n1974,
    n1243,
    n1346,
    n1466,
    n1219
  );


  nor
  g2866
  (
    n1537,
    n1093,
    n1147,
    n1313,
    n1100
  );


  nor
  g2867
  (
    n2152,
    n1442,
    n1382,
    n1326,
    n1281
  );


  xnor
  g2868
  (
    n2449,
    n1163,
    n1230,
    n1287,
    n1243
  );


  and
  g2869
  (
    n2648,
    n1206,
    n1136,
    n1299,
    n1155
  );


  xnor
  g2870
  (
    n2830,
    n1483,
    n1405,
    n1191,
    n1096
  );


  xor
  g2871
  (
    n2277,
    n1280,
    n1325,
    n1178,
    n1298
  );


  nor
  g2872
  (
    n1786,
    n1250,
    n1173,
    n1098,
    n1119
  );


  nor
  g2873
  (
    n1576,
    n1149,
    n1149,
    n1267,
    n1223
  );


  nor
  g2874
  (
    n2360,
    n1452,
    n1468,
    n1439,
    n1324
  );


  or
  g2875
  (
    n1975,
    n1202,
    n1252,
    n1458,
    n1374
  );


  xnor
  g2876
  (
    n2719,
    n1410,
    n1245,
    n1388,
    n1363
  );


  xor
  g2877
  (
    n1972,
    n1245,
    n1440,
    n1389,
    n1482
  );


  nor
  g2878
  (
    n2499,
    n1393,
    n1188,
    n1441,
    n1428
  );


  nand
  g2879
  (
    n1686,
    n1211,
    n1461,
    n1090,
    n1239
  );


  and
  g2880
  (
    n1725,
    n1455,
    n1502,
    n1210,
    n1412
  );


  nor
  g2881
  (
    n2184,
    n1093,
    n1301,
    n1464,
    n1146
  );


  nor
  g2882
  (
    n2259,
    n1398,
    n1205,
    n1225,
    n1216
  );


  nand
  g2883
  (
    n2431,
    n1286,
    n1216,
    n1175,
    n1356
  );


  xor
  g2884
  (
    n2732,
    n1120,
    n1253,
    n1416,
    n1098
  );


  and
  g2885
  (
    n2862,
    n1498,
    n1160,
    n1404
  );


  or
  g2886
  (
    n1869,
    n1503,
    n1157,
    n1274,
    n1232
  );


  or
  g2887
  (
    n1589,
    n1164,
    n1107,
    n1135,
    n1357
  );


  nand
  g2888
  (
    n2827,
    n1254,
    n1381,
    n1353,
    n1461
  );


  xor
  g2889
  (
    n1663,
    n1374,
    n1382,
    n1505,
    n1286
  );


  or
  g2890
  (
    n1559,
    n1505,
    n1212,
    n1135,
    n1309
  );


  xor
  g2891
  (
    KeyWire_0_26,
    n1302,
    n1258,
    n1368,
    n1310
  );


  or
  g2892
  (
    n1679,
    n1119,
    n1351,
    n1494,
    n1324
  );


  or
  g2893
  (
    n2260,
    n1110,
    n1454,
    n1353,
    n1240
  );


  nand
  g2894
  (
    n1850,
    n1380,
    n1097,
    n1482,
    n1267
  );


  or
  g2895
  (
    n2409,
    n1181,
    n1432,
    n1449,
    n1260
  );


  and
  g2896
  (
    n2378,
    n1253,
    n1215,
    n1488,
    n1275
  );


  and
  g2897
  (
    n2172,
    n947,
    n1456,
    n1123,
    n1364
  );


  and
  g2898
  (
    n2586,
    n1355,
    n1466,
    n1144,
    n1110
  );


  xnor
  g2899
  (
    n2302,
    n1182,
    n1154,
    n1493,
    n1336
  );


  and
  g2900
  (
    n2160,
    n1338,
    n1315,
    n1487,
    n1363
  );


  xor
  g2901
  (
    n1816,
    n1299,
    n1492,
    n1130,
    n1114
  );


  nand
  g2902
  (
    n1961,
    n1452,
    n1313,
    n1479,
    n1146
  );


  or
  g2903
  (
    n2840,
    n1284,
    n1283,
    n1117,
    n1460
  );


  nor
  g2904
  (
    n2914,
    n1453,
    n1092,
    n1430,
    n1435
  );


  nor
  g2905
  (
    n1526,
    n948,
    n1367,
    n1384,
    n1361
  );


  nand
  g2906
  (
    n2486,
    n1284,
    n1447,
    n1124,
    n1115
  );


  nor
  g2907
  (
    n2394,
    n1248,
    n1390,
    n1485,
    n1409
  );


  nand
  g2908
  (
    n2894,
    n1439,
    n1298,
    n1377,
    n1392
  );


  xor
  g2909
  (
    n2539,
    n1399,
    n1221,
    n1163,
    n1336
  );


  nand
  g2910
  (
    n1811,
    n1393,
    n1364,
    n1396,
    n1139
  );


  xnor
  g2911
  (
    n1579,
    n1363,
    n1449,
    n1414,
    n1381
  );


  xnor
  g2912
  (
    n2907,
    n1245,
    n1441,
    n1405,
    n1395
  );


  nand
  g2913
  (
    n2633,
    n1269,
    n1140,
    n1428,
    n1261
  );


  or
  g2914
  (
    n2664,
    n1308,
    n1355,
    n1400,
    n1172
  );


  and
  g2915
  (
    n1715,
    n1408,
    n1437,
    n1489,
    n1211
  );


  xnor
  g2916
  (
    n1671,
    n1421,
    n1186,
    n1266,
    n1192
  );


  or
  g2917
  (
    n3360,
    n2883,
    n1622,
    n1893,
    n2558
  );


  nor
  g2918
  (
    n3022,
    n2053,
    n2504,
    n711,
    n2404
  );


  nor
  g2919
  (
    n2954,
    n1539,
    n1850,
    n1772,
    n626
  );


  xor
  g2920
  (
    n3066,
    n2187,
    n2903,
    n2274,
    n2878
  );


  xnor
  g2921
  (
    n3061,
    n2792,
    n2608,
    n2767,
    n1723
  );


  xnor
  g2922
  (
    n3337,
    n1562,
    n575,
    n2913,
    n2951
  );


  or
  g2923
  (
    n3382,
    n2252,
    n583,
    n2600,
    n1606
  );


  nor
  g2924
  (
    n3117,
    n2625,
    n2925,
    n2890,
    n2340
  );


  nand
  g2925
  (
    n3326,
    n2921,
    n2943,
    n1820,
    n2935
  );


  nor
  g2926
  (
    n3282,
    n1546,
    n1596,
    n2950,
    n2924
  );


  or
  g2927
  (
    n3251,
    n633,
    n2923,
    n2366,
    n2016
  );


  xor
  g2928
  (
    n3311,
    n1863,
    n2322,
    n1766,
    n2627
  );


  xnor
  g2929
  (
    n2999,
    n617,
    n2932,
    n1920,
    n2083
  );


  and
  g2930
  (
    n2968,
    n588,
    n2925,
    n1524,
    n2045
  );


  nand
  g2931
  (
    n3295,
    n2876,
    n1616,
    n2908,
    n2510
  );


  nand
  g2932
  (
    n3158,
    n2677,
    n2934,
    n1954,
    n2006
  );


  xnor
  g2933
  (
    n3071,
    n2530,
    n1838,
    n2546,
    n1669
  );


  and
  g2934
  (
    n3057,
    n2155,
    n2368,
    n2903,
    n2939
  );


  nor
  g2935
  (
    n3380,
    n2775,
    n2809,
    n714,
    n1819
  );


  and
  g2936
  (
    n3277,
    n1679,
    n1752,
    n2098,
    n1673
  );


  nor
  g2937
  (
    n3019,
    n1608,
    n1515,
    n1578,
    n2536
  );


  or
  g2938
  (
    n3049,
    n2400,
    n2419,
    n2167,
    n1624
  );


  nor
  g2939
  (
    n3146,
    n2685,
    n1613,
    n640,
    n2247
  );


  nor
  g2940
  (
    n3042,
    n2810,
    n2916,
    n2671,
    n562
  );


  nor
  g2941
  (
    n2998,
    n1770,
    n2248,
    n2875,
    n2761
  );


  and
  g2942
  (
    n3123,
    n2454,
    n2657,
    n2391,
    n722
  );


  nand
  g2943
  (
    n3035,
    n2173,
    n2700,
    n2909,
    n2883
  );


  or
  g2944
  (
    n3217,
    n2487,
    n2894,
    n2123,
    n2372
  );


  xnor
  g2945
  (
    n3163,
    n2693,
    n2057,
    n2858,
    n2665
  );


  nor
  g2946
  (
    n3064,
    n577,
    n1744,
    n2441,
    n2676
  );


  xnor
  g2947
  (
    n3044,
    n1833,
    n2952,
    n2418,
    n1949
  );


  and
  g2948
  (
    n3140,
    n2463,
    n2184,
    n2888,
    n673
  );


  nor
  g2949
  (
    n3322,
    n1807,
    n666,
    n2236,
    n2226
  );


  and
  g2950
  (
    n3015,
    n2359,
    n1551,
    n2234,
    n2899
  );


  xnor
  g2951
  (
    n3176,
    n1603,
    n646,
    n2119,
    n2477
  );


  xnor
  g2952
  (
    n2979,
    n1984,
    n1696,
    n2576,
    n2833
  );


  nor
  g2953
  (
    n2958,
    n2938,
    n2787,
    n2312,
    n2695
  );


  nand
  g2954
  (
    n2970,
    n2298,
    n2703,
    n1932,
    n670
  );


  nor
  g2955
  (
    n3271,
    n1909,
    n2357,
    n2724,
    n2506
  );


  nor
  g2956
  (
    n3177,
    n2678,
    n2491,
    n2139,
    n2432
  );


  or
  g2957
  (
    n2975,
    n2829,
    n1549,
    n2717,
    n2675
  );


  nor
  g2958
  (
    n3131,
    n2044,
    n1735,
    n2343,
    n1677
  );


  xor
  g2959
  (
    n2993,
    n2853,
    n2905,
    n1563,
    n2497
  );


  nand
  g2960
  (
    n3240,
    n2503,
    n2559,
    n1915,
    n2811
  );


  xnor
  g2961
  (
    n3028,
    n2143,
    n2822,
    n1591,
    n2295
  );


  nand
  g2962
  (
    n3222,
    n2038,
    n2837,
    n2317,
    n2663
  );


  and
  g2963
  (
    n3167,
    n2952,
    n1733,
    n1611,
    n2233
  );


  nor
  g2964
  (
    n3000,
    n1910,
    n2889,
    n2817,
    n1814
  );


  xnor
  g2965
  (
    n3017,
    n2354,
    n1987,
    n2434,
    n2105
  );


  and
  g2966
  (
    n3185,
    n2462,
    n2318,
    n2112,
    n635
  );


  or
  g2967
  (
    n3070,
    n2358,
    n1957,
    n2094,
    n2423
  );


  or
  g2968
  (
    n3384,
    n2320,
    n2393,
    n2100,
    n1921
  );


  xor
  g2969
  (
    n3020,
    n573,
    n2386,
    n1629,
    n2877
  );


  and
  g2970
  (
    n3119,
    n576,
    n662,
    n686,
    n2407
  );


  and
  g2971
  (
    n3237,
    n1790,
    n2189,
    n2946,
    n1834
  );


  nand
  g2972
  (
    n3196,
    n2892,
    n2421,
    n2319,
    n2762
  );


  xnor
  g2973
  (
    n3234,
    n2556,
    n2931,
    n2895,
    n1940
  );


  xnor
  g2974
  (
    KeyWire_0_31,
    n651,
    n2788,
    n2865,
    n570
  );


  nand
  g2975
  (
    n2973,
    n721,
    n1841,
    n2279,
    n2327
  );


  nand
  g2976
  (
    n3108,
    n1878,
    n2363,
    n1727,
    n2235
  );


  xor
  g2977
  (
    n3142,
    n2913,
    n2022,
    n2834,
    n2653
  );


  or
  g2978
  (
    n2974,
    n2058,
    n1598,
    n591,
    n2798
  );


  or
  g2979
  (
    n3180,
    n1753,
    n2308,
    n2471,
    n2548
  );


  nor
  g2980
  (
    n3219,
    n1988,
    n2581,
    n2553,
    n1991
  );


  xor
  g2981
  (
    n3179,
    n2907,
    n1560,
    n2928,
    n1799
  );


  nand
  g2982
  (
    n3264,
    n2780,
    n1851,
    n2425,
    n687
  );


  nor
  g2983
  (
    n3147,
    n1584,
    n2076,
    n2583,
    n579
  );


  nand
  g2984
  (
    n3168,
    n1939,
    n2460,
    n2686,
    n1929
  );


  and
  g2985
  (
    n2989,
    n2718,
    n2396,
    n1881,
    n2244
  );


  xor
  g2986
  (
    n3150,
    n2178,
    n1512,
    n1809,
    n2486
  );


  xor
  g2987
  (
    n3345,
    n2348,
    n2935,
    n2803,
    n2947
  );


  xnor
  g2988
  (
    n3313,
    n2709,
    n2894,
    n2230,
    n2642
  );


  nand
  g2989
  (
    n3133,
    n2158,
    n2197,
    n2249,
    n2301
  );


  nand
  g2990
  (
    n3113,
    n1715,
    n2203,
    n1989,
    n693
  );


  nor
  g2991
  (
    n3077,
    n2710,
    n2104,
    n2746,
    n2728
  );


  nor
  g2992
  (
    n3141,
    n2440,
    n2914,
    n2596,
    n2101
  );


  xnor
  g2993
  (
    n3050,
    n2776,
    n2195,
    n2283,
    n2069
  );


  xor
  g2994
  (
    n3327,
    n2947,
    n2698,
    n1724,
    n2114
  );


  xnor
  g2995
  (
    n3351,
    n2309,
    n1755,
    n2300,
    n2617
  );


  xor
  g2996
  (
    n3210,
    n2606,
    n1971,
    n568,
    n2727
  );


  xor
  g2997
  (
    n3078,
    n619,
    n2289,
    n2871,
    n1784
  );


  nor
  g2998
  (
    n2965,
    n2880,
    n1847,
    n2914,
    n2797
  );


  nor
  g2999
  (
    n3103,
    n1787,
    n2624,
    n2573,
    n2415
  );


  nand
  g3000
  (
    n3280,
    n2108,
    n1618,
    n1590,
    n2771
  );


  and
  g3001
  (
    n3046,
    n1936,
    n2939,
    n1628,
    n683
  );


  nor
  g3002
  (
    n2984,
    n2140,
    n2915,
    n2242,
    n2498
  );


  nor
  g3003
  (
    n3216,
    n2936,
    n1550,
    n2445,
    n1739
  );


  or
  g3004
  (
    n2956,
    n1734,
    n2644,
    n2074,
    n1913
  );


  and
  g3005
  (
    n3181,
    n1545,
    n1623,
    n2681,
    n1721
  );


  or
  g3006
  (
    n3304,
    n2755,
    n2807,
    n2565,
    n2930
  );


  xnor
  g3007
  (
    n3156,
    n699,
    n1544,
    n2569,
    n2383
  );


  or
  g3008
  (
    n2957,
    n2647,
    n2949,
    n2900,
    n1740
  );


  xnor
  g3009
  (
    n3093,
    n1840,
    n2145,
    n1977,
    n2782
  );


  xor
  g3010
  (
    n3135,
    n679,
    n1869,
    n2759,
    n1898
  );


  nand
  g3011
  (
    n3032,
    n1975,
    n655,
    n2349,
    n580
  );


  nor
  g3012
  (
    n3288,
    n2211,
    n2660,
    n1760,
    n2870
  );


  and
  g3013
  (
    n3213,
    n1973,
    n1633,
    n1938,
    n2666
  );


  xor
  g3014
  (
    n3248,
    n1762,
    n1757,
    n2007,
    n1996
  );


  nor
  g3015
  (
    n3162,
    n1896,
    n2153,
    n2455,
    n1901
  );


  xnor
  g3016
  (
    n3225,
    n2088,
    n1575,
    n1717,
    n1506
  );


  nand
  g3017
  (
    n3214,
    n2165,
    n2092,
    n1690,
    n2585
  );


  xnor
  g3018
  (
    n3058,
    n1888,
    n2381,
    n2206,
    n2941
  );


  nand
  g3019
  (
    n3383,
    n2588,
    n678,
    n2918,
    n2004
  );


  xnor
  g3020
  (
    n2982,
    n2943,
    n1535,
    n681,
    n2934
  );


  nand
  g3021
  (
    n3296,
    n2023,
    n2448,
    n571,
    n2652
  );


  or
  g3022
  (
    n3347,
    n1555,
    n1547,
    n1997,
    n2539
  );


  and
  g3023
  (
    n3328,
    n1951,
    n1759,
    n2944,
    n2511
  );


  xor
  g3024
  (
    n3247,
    n2429,
    n2192,
    n1780,
    n2458
  );


  and
  g3025
  (
    n3004,
    n2093,
    n1526,
    n644,
    n1768
  );


  nor
  g3026
  (
    n3395,
    n2011,
    n2476,
    n1805,
    n1602
  );


  nand
  g3027
  (
    n2990,
    n2055,
    n2082,
    n2035,
    n1754
  );


  xnor
  g3028
  (
    n3208,
    n1588,
    n2378,
    n1699,
    n2172
  );


  and
  g3029
  (
    n3105,
    n2879,
    n2648,
    n1680,
    n1976
  );


  or
  g3030
  (
    n3275,
    n1565,
    n2929,
    n2224,
    n2919
  );


  nor
  g3031
  (
    n3193,
    n2018,
    n2282,
    n1706,
    n2439
  );


  xnor
  g3032
  (
    n3012,
    n2870,
    n2063,
    n567,
    n2408
  );


  nor
  g3033
  (
    n3291,
    n2124,
    n1533,
    n2324,
    n2111
  );


  xnor
  g3034
  (
    n3294,
    n1540,
    n1758,
    n2910,
    n2701
  );


  xnor
  g3035
  (
    n3085,
    n2405,
    n2869,
    n658,
    n2937
  );


  xor
  g3036
  (
    n3349,
    n2555,
    n2705,
    n2857,
    n1626
  );


  xor
  g3037
  (
    n3355,
    n2185,
    n1918,
    n1892,
    n1519
  );


  and
  g3038
  (
    n3018,
    n2896,
    n2134,
    n707,
    n2078
  );


  xnor
  g3039
  (
    n3281,
    n1636,
    n2861,
    n709,
    n1845
  );


  nand
  g3040
  (
    n3372,
    n1592,
    n2936,
    n1917,
    n2945
  );


  nand
  g3041
  (
    n3386,
    n2799,
    n2682,
    n2297,
    n2332
  );


  nand
  g3042
  (
    n3377,
    n2468,
    n2730,
    n2937,
    n2863
  );


  xnor
  g3043
  (
    n3243,
    n1955,
    n2737,
    n1937,
    n659
  );


  nand
  g3044
  (
    n3241,
    n2250,
    n2729,
    n1556,
    n663
  );


  and
  g3045
  (
    n3292,
    n2047,
    n618,
    n1671,
    n1781
  );


  xor
  g3046
  (
    n3084,
    n1665,
    n1952,
    n2890,
    n1640
  );


  xnor
  g3047
  (
    n3041,
    n2904,
    n2840,
    n598,
    n2271
  );


  nand
  g3048
  (
    n2986,
    n2561,
    n566,
    n2286,
    n1538
  );


  and
  g3049
  (
    n3220,
    n1998,
    n1612,
    n1972,
    n1944
  );


  or
  g3050
  (
    n3400,
    n1674,
    n1818,
    n2523,
    n1763
  );


  xnor
  g3051
  (
    n3023,
    n2901,
    n2795,
    n1963,
    n2613
  );


  and
  g3052
  (
    n3335,
    n2150,
    n1978,
    n1528,
    n2949
  );


  nor
  g3053
  (
    n3246,
    n2591,
    n2107,
    n2070,
    n2268
  );


  xnor
  g3054
  (
    n3052,
    n2778,
    n2394,
    n2937,
    n2770
  );


  or
  g3055
  (
    n2983,
    n1521,
    n2290,
    n2221,
    n1594
  );


  nor
  g3056
  (
    n2997,
    n1967,
    n1846,
    n2904,
    n2933
  );


  and
  g3057
  (
    n3130,
    n2163,
    n2321,
    n2594,
    n2891
  );


  nand
  g3058
  (
    n3056,
    n1974,
    n2779,
    n1827,
    n2075
  );


  or
  g3059
  (
    n3171,
    n2897,
    n587,
    n2305,
    n2667
  );


  nand
  g3060
  (
    n3283,
    n2010,
    n2768,
    n1558,
    n1965
  );


  xnor
  g3061
  (
    n3266,
    n2912,
    n2944,
    n2072,
    n2512
  );


  xor
  g3062
  (
    n3054,
    n1631,
    n2804,
    n1876,
    n1788
  );


  nor
  g3063
  (
    n3359,
    n2773,
    n2814,
    n2905,
    n569
  );


  and
  g3064
  (
    n3194,
    n2948,
    n1691,
    n2551,
    n1886
  );


  and
  g3065
  (
    n3074,
    n2220,
    n2601,
    n2845,
    n2331
  );


  xnor
  g3066
  (
    n3276,
    n2891,
    n1769,
    n2467,
    n2926
  );


  nand
  g3067
  (
    n3175,
    n1514,
    n2924,
    n2604,
    n2540
  );


  and
  g3068
  (
    n3305,
    n2879,
    n2169,
    n2929,
    n2410
  );


  and
  g3069
  (
    n3317,
    n2839,
    n2641,
    n1871,
    n1999
  );


  xor
  g3070
  (
    n3390,
    n2887,
    n2884,
    n2473,
    n2917
  );


  nand
  g3071
  (
    n3170,
    n2632,
    n2061,
    n1852,
    n2866
  );


  and
  g3072
  (
    n3299,
    n2051,
    n2927,
    n2543,
    n1647
  );


  and
  g3073
  (
    n3010,
    n2831,
    n1595,
    n2599,
    n2572
  );


  xnor
  g3074
  (
    n3204,
    n2882,
    n2699,
    n2219,
    n1570
  );


  nand
  g3075
  (
    n3040,
    n2260,
    n1711,
    n2893,
    n2377
  );


  nand
  g3076
  (
    n3055,
    n1648,
    n2411,
    n669,
    n1803
  );


  xnor
  g3077
  (
    n3006,
    n2501,
    n1899,
    n2735,
    n2259
  );


  nor
  g3078
  (
    n3387,
    n2469,
    n2931,
    n1905,
    n2360
  );


  or
  g3079
  (
    n3375,
    n2616,
    n1554,
    n2213,
    n2524
  );


  xnor
  g3080
  (
    n3086,
    n2106,
    n2888,
    n1773,
    n1522
  );


  xor
  g3081
  (
    n3048,
    n1689,
    n1811,
    n2037,
    n1559
  );


  nor
  g3082
  (
    n3244,
    n1649,
    n2019,
    n2293,
    n1703
  );


  nand
  g3083
  (
    n3357,
    n1738,
    n1935,
    n648,
    n2292
  );


  xor
  g3084
  (
    n3242,
    n2649,
    n2945,
    n620,
    n2352
  );


  and
  g3085
  (
    n3206,
    n2442,
    n1789,
    n2723,
    n2936
  );


  and
  g3086
  (
    n3278,
    n2580,
    n2089,
    n1541,
    n637
  );


  xor
  g3087
  (
    n2962,
    n2680,
    n607,
    n1761,
    n2872
  );


  or
  g3088
  (
    n3106,
    n2951,
    n1927,
    n2867,
    n2071
  );


  or
  g3089
  (
    n3187,
    n2871,
    n2026,
    n2889,
    n1862
  );


  xor
  g3090
  (
    n3339,
    n2866,
    n1891,
    n2520,
    n1904
  );


  and
  g3091
  (
    n3329,
    n2527,
    n2631,
    n1610,
    n2910
  );


  xor
  g3092
  (
    n2981,
    n584,
    n2855,
    n2144,
    n1832
  );


  and
  g3093
  (
    n3104,
    n695,
    n1748,
    n1660,
    n2355
  );


  nand
  g3094
  (
    n3002,
    n1816,
    n2137,
    n1694,
    n2754
  );


  nor
  g3095
  (
    n3399,
    n2908,
    n2567,
    n1826,
    n2873
  );


  nor
  g3096
  (
    n2992,
    n2459,
    n2864,
    n2450,
    n2951
  );


  xnor
  g3097
  (
    n3080,
    n650,
    n1943,
    n1946,
    n2870
  );


  or
  g3098
  (
    n3373,
    n589,
    n2842,
    n1746,
    n2732
  );


  nor
  g3099
  (
    n3095,
    n2127,
    n2480,
    n636,
    n634
  );


  xor
  g3100
  (
    n3063,
    n2948,
    n2256,
    n2210,
    n2182
  );


  nor
  g3101
  (
    n2991,
    n1794,
    n1894,
    n2064,
    n2479
  );


  nor
  g3102
  (
    n3352,
    n585,
    n1849,
    n2838,
    n2854
  );


  or
  g3103
  (
    n3370,
    n2238,
    n1885,
    n1824,
    n2748
  );


  and
  g3104
  (
    n3218,
    n2828,
    n2879,
    n2742,
    n2085
  );


  nor
  g3105
  (
    n3098,
    n1877,
    n1517,
    n2193,
    n2760
  );


  and
  g3106
  (
    n3192,
    n2619,
    n642,
    n2528,
    n1767
  );


  xnor
  g3107
  (
    n3236,
    n2162,
    n2825,
    n2942,
    n1830
  );


  and
  g3108
  (
    n3114,
    n1684,
    n2447,
    n665,
    n1854
  );


  xor
  g3109
  (
    n3051,
    n1880,
    n2841,
    n1749,
    n2427
  );


  and
  g3110
  (
    n3008,
    n2867,
    n2734,
    n2534,
    n1627
  );


  nor
  g3111
  (
    n3231,
    n2231,
    n2346,
    n2886,
    n2827
  );


  or
  g3112
  (
    n3178,
    n613,
    n1645,
    n2118,
    n2593
  );


  xor
  g3113
  (
    n2961,
    n2401,
    n2005,
    n2280,
    n2208
  );


  or
  g3114
  (
    n3200,
    n1751,
    n2382,
    n2066,
    n1798
  );


  nand
  g3115
  (
    n3129,
    n1969,
    n1609,
    n1945,
    n2897
  );


  xnor
  g3116
  (
    n3346,
    n2856,
    n2883,
    n2715,
    n1635
  );


  nand
  g3117
  (
    n3016,
    n2928,
    n557,
    n2952,
    n1527
  );


  or
  g3118
  (
    KeyWire_0_4,
    n2222,
    n671,
    n1779,
    n2518
  );


  xor
  g3119
  (
    n3021,
    n2621,
    n624,
    n2362,
    n2135
  );


  nor
  g3120
  (
    n3274,
    n561,
    n2090,
    n2079,
    n2128
  );


  nor
  g3121
  (
    n3203,
    n627,
    n2753,
    n2711,
    n2704
  );


  or
  g3122
  (
    n3239,
    n2217,
    n2874,
    n2562,
    n1534
  );


  nor
  g3123
  (
    n3396,
    n2579,
    n2232,
    n2867,
    n2042
  );


  xor
  g3124
  (
    n3232,
    n694,
    n2826,
    n2373,
    n2669
  );


  nor
  g3125
  (
    n2959,
    n2397,
    n2876,
    n1750,
    n700
  );


  or
  g3126
  (
    n3120,
    n1776,
    n1567,
    n1870,
    n2942
  );


  and
  g3127
  (
    n3223,
    n1848,
    n1621,
    n2056,
    n1792
  );


  or
  g3128
  (
    n3286,
    n2875,
    n2302,
    n2342,
    n1931
  );


  nand
  g3129
  (
    n3238,
    n628,
    n1693,
    n2261,
    n2882
  );


  nor
  g3130
  (
    n3394,
    n2266,
    n652,
    n2131,
    n2277
  );


  xnor
  g3131
  (
    n2980,
    n2928,
    n2895,
    n1516,
    n682
  );


  xor
  g3132
  (
    n3205,
    n1962,
    n611,
    n1785,
    n2917
  );


  xnor
  g3133
  (
    n3303,
    n2916,
    n2821,
    n1942,
    n632
  );


  and
  g3134
  (
    n3075,
    n2110,
    n2239,
    n2869,
    n1707
  );


  xnor
  g3135
  (
    n3197,
    n2716,
    n2656,
    n2243,
    n2659
  );


  or
  g3136
  (
    n3127,
    n660,
    n1836,
    n2892,
    n1777
  );


  xnor
  g3137
  (
    n3227,
    n2949,
    n2898,
    n1681,
    n2921
  );


  or
  g3138
  (
    n3073,
    n1655,
    n2246,
    n616,
    n2692
  );


  and
  g3139
  (
    n3090,
    n710,
    n647,
    n2612,
    n2938
  );


  nand
  g3140
  (
    n3371,
    n2229,
    n2923,
    n1651,
    n622
  );


  and
  g3141
  (
    n2987,
    n1736,
    n2919,
    n2033,
    n2338
  );


  and
  g3142
  (
    n3233,
    n2915,
    n2347,
    n1685,
    n1662
  );


  and
  g3143
  (
    n2955,
    n685,
    n2253,
    n2021,
    n2607
  );


  or
  g3144
  (
    n3001,
    n2008,
    n2713,
    n1743,
    n2050
  );


  and
  g3145
  (
    n3285,
    n2578,
    n1889,
    n1634,
    n1985
  );


  or
  g3146
  (
    n3081,
    n2147,
    n1796,
    n656,
    n1964
  );


  xnor
  g3147
  (
    n3254,
    n2940,
    n2328,
    n2191,
    n2877
  );


  nor
  g3148
  (
    n3159,
    n2747,
    n1656,
    n2750,
    n1804
  );


  and
  g3149
  (
    n3186,
    n2499,
    n2885,
    n2426,
    n2181
  );


  xnor
  g3150
  (
    n3121,
    n1716,
    n2915,
    n698,
    n1536
  );


  or
  g3151
  (
    n3252,
    n2160,
    n2350,
    n2102,
    n2129
  );


  or
  g3152
  (
    n3398,
    n2899,
    n2818,
    n2781,
    n2255
  );


  and
  g3153
  (
    n3367,
    n2334,
    n1857,
    n1605,
    n2036
  );


  nor
  g3154
  (
    n3045,
    n1902,
    n1686,
    n2679,
    n1577
  );


  xor
  g3155
  (
    n3368,
    n2918,
    n2740,
    n1639,
    n2690
  );


  and
  g3156
  (
    n3191,
    n1934,
    n2031,
    n2096,
    n2764
  );


  or
  g3157
  (
    n3038,
    n2892,
    n2482,
    n2899,
    n2922
  );


  xnor
  g3158
  (
    n3290,
    n2529,
    n2950,
    n2387,
    n2307
  );


  nand
  g3159
  (
    n3101,
    n1713,
    n586,
    n1718,
    n2796
  );


  xor
  g3160
  (
    n3312,
    n2945,
    n2634,
    n2582,
    n1919
  );


  or
  g3161
  (
    n3388,
    n2847,
    n2691,
    n1531,
    n2336
  );


  nor
  g3162
  (
    n3364,
    n2603,
    n2605,
    n2012,
    n2938
  );


  and
  g3163
  (
    n3007,
    n2942,
    n2874,
    n2263,
    n2344
  );


  xor
  g3164
  (
    n3257,
    n2436,
    n2784,
    n1589,
    n2880
  );


  xor
  g3165
  (
    n3230,
    n1861,
    n2823,
    n2330,
    n2457
  );


  nand
  g3166
  (
    n3309,
    n2708,
    n2227,
    n2884,
    n2039
  );


  and
  g3167
  (
    n3102,
    n2736,
    n1702,
    n2947,
    n2566
  );


  or
  g3168
  (
    n3195,
    n1960,
    n2375,
    n2223,
    n1714
  );


  xnor
  g3169
  (
    n3182,
    n2757,
    n2122,
    n2353,
    n703
  );


  xnor
  g3170
  (
    n3209,
    n2950,
    n1771,
    n2059,
    n2661
  );


  xnor
  g3171
  (
    n3065,
    n2557,
    n2141,
    n2595,
    n582
  );


  and
  g3172
  (
    n3132,
    n2866,
    n2303,
    n1922,
    n606
  );


  and
  g3173
  (
    KeyWire_0_23,
    n2571,
    n1599,
    n2901,
    n674
  );


  or
  g3174
  (
    n3320,
    n2900,
    n1572,
    n2099,
    n2917
  );


  xnor
  g3175
  (
    n3314,
    n2739,
    n2430,
    n2674,
    n1726
  );


  nand
  g3176
  (
    n3047,
    n2109,
    n2484,
    n2264,
    n2881
  );


  xor
  g3177
  (
    KeyWire_0_1,
    n2517,
    n1529,
    n1672,
    n690
  );


  and
  g3178
  (
    n3107,
    n2926,
    n1676,
    n1641,
    n2485
  );


  nand
  g3179
  (
    n3011,
    n2901,
    n2918,
    n2843,
    n2574
  );


  and
  g3180
  (
    n3224,
    n2862,
    n2877,
    n2509,
    n2041
  );


  xnor
  g3181
  (
    n3343,
    n2889,
    n1644,
    n1981,
    n2869
  );


  or
  g3182
  (
    n3143,
    n639,
    n2687,
    n1858,
    n2902
  );


  xnor
  g3183
  (
    n3165,
    n675,
    n2635,
    n2908,
    n2662
  );


  xor
  g3184
  (
    n3030,
    n2288,
    n1582,
    n2294,
    n1874
  );


  or
  g3185
  (
    n3361,
    n1800,
    n2801,
    n2905,
    n2909
  );


  and
  g3186
  (
    n3344,
    n1741,
    n615,
    n2844,
    n630
  );


  and
  g3187
  (
    n3083,
    n2228,
    n1756,
    n2130,
    n2910
  );


  or
  g3188
  (
    n3258,
    n1842,
    n2577,
    n1813,
    n1709
  );


  and
  g3189
  (
    n3112,
    n2152,
    n1666,
    n2950,
    n1925
  );


  nor
  g3190
  (
    n3211,
    n2549,
    n2944,
    n2508,
    n2202
  );


  xnor
  g3191
  (
    n3226,
    n1638,
    n2592,
    n629,
    n2630
  );


  or
  g3192
  (
    n3365,
    n2417,
    n2726,
    n2437,
    n2376
  );


  nor
  g3193
  (
    n3145,
    n2205,
    n1687,
    n2744,
    n661
  );


  and
  g3194
  (
    n3184,
    n1879,
    n2488,
    n2694,
    n2590
  );


  or
  g3195
  (
    n3354,
    n2552,
    n2951,
    n2281,
    n1810
  );


  nor
  g3196
  (
    n3092,
    n2878,
    n1630,
    n1958,
    n2783
  );


  or
  g3197
  (
    n3279,
    n2623,
    n1865,
    n2424,
    n2752
  );


  xor
  g3198
  (
    KeyWire_0_17,
    n716,
    n2873,
    n2628,
    n2765
  );


  xor
  g3199
  (
    n3273,
    n621,
    n581,
    n2860,
    n1895
  );


  and
  g3200
  (
    n2996,
    n2464,
    n2493,
    n1507,
    n2859
  );


  xor
  g3201
  (
    n3255,
    n1525,
    n2422,
    n1720,
    n2478
  );


  xnor
  g3202
  (
    n3245,
    n1617,
    n2832,
    n1774,
    n2474
  );


  xnor
  g3203
  (
    n3358,
    n2816,
    n1737,
    n1663,
    n2313
  );


  nand
  g3204
  (
    n3316,
    n2526,
    n2584,
    n2174,
    n1574
  );


  and
  g3205
  (
    n3172,
    n1872,
    n1775,
    n2490,
    n2672
  );


  xnor
  g3206
  (
    n3148,
    n2533,
    n2802,
    n1986,
    n676
  );


  xnor
  g3207
  (
    n3341,
    n2766,
    n2461,
    n2179,
    n2030
  );


  or
  g3208
  (
    n3272,
    n2712,
    n2003,
    n2149,
    n1828
  );


  or
  g3209
  (
    n3053,
    n1532,
    n597,
    n654,
    n1923
  );


  nand
  g3210
  (
    n3268,
    n1646,
    n2900,
    n2615,
    n2519
  );


  xor
  g3211
  (
    n3153,
    n2941,
    n2367,
    n1791,
    n2329
  );


  or
  g3212
  (
    n3139,
    n2749,
    n1586,
    n2240,
    n1571
  );


  nor
  g3213
  (
    n3137,
    n1583,
    n1990,
    n2284,
    n2345
  );


  nand
  g3214
  (
    n2978,
    n2560,
    n2000,
    n2609,
    n2946
  );


  nor
  g3215
  (
    n3087,
    n2180,
    n2341,
    n1508,
    n1597
  );


  nor
  g3216
  (
    n2960,
    n1601,
    n2875,
    n2385,
    n1860
  );


  nand
  g3217
  (
    n3253,
    n1956,
    n2412,
    n2873,
    n2444
  );


  and
  g3218
  (
    n3198,
    n643,
    n1897,
    n645,
    n2815
  );


  xnor
  g3219
  (
    n3166,
    n2587,
    n2638,
    n2670,
    n1619
  );


  and
  g3220
  (
    n3363,
    n2646,
    n2893,
    n2920,
    n2291
  );


  nor
  g3221
  (
    n3321,
    n2911,
    n697,
    n2380,
    n2922
  );


  or
  g3222
  (
    n3289,
    n2171,
    n2121,
    n2920,
    n1947
  );


  nand
  g3223
  (
    n3332,
    n2323,
    n1822,
    n2333,
    n564
  );


  nand
  g3224
  (
    KeyWire_0_2,
    n1786,
    n1668,
    n704,
    n1692
  );


  xor
  g3225
  (
    n3300,
    n1579,
    n1625,
    n1853,
    n2199
  );


  xnor
  g3226
  (
    n3310,
    n2156,
    n2743,
    n2697,
    n2550
  );


  nor
  g3227
  (
    n3385,
    n688,
    n2673,
    n2287,
    n2084
  );


  or
  g3228
  (
    n3259,
    n1831,
    n2916,
    n2888,
    n2922
  );


  xor
  g3229
  (
    n3207,
    n1793,
    n1953,
    n2032,
    n2927
  );


  and
  g3230
  (
    n3319,
    n1698,
    n1513,
    n1906,
    n1548
  );


  nand
  g3231
  (
    n3183,
    n2785,
    n2115,
    n2392,
    n2898
  );


  nand
  g3232
  (
    n3079,
    n2138,
    n2772,
    n2505,
    n2852
  );


  and
  g3233
  (
    n3138,
    n1764,
    n1585,
    n2914,
    n719
  );


  and
  g3234
  (
    n2969,
    n2414,
    n1725,
    n1979,
    n2390
  );


  xor
  g3235
  (
    n3014,
    n2745,
    n2887,
    n2446,
    n2065
  );


  nand
  g3236
  (
    n3342,
    n1837,
    n631,
    n2911,
    n2909
  );


  nor
  g3237
  (
    n3025,
    n2148,
    n2542,
    n2315,
    n625
  );


  and
  g3238
  (
    n3069,
    n1884,
    n2514,
    n2258,
    n2696
  );


  nand
  g3239
  (
    n3128,
    n1632,
    n1950,
    n2403,
    n2048
  );


  nand
  g3240
  (
    n3161,
    n2871,
    n2758,
    n2515,
    n2884
  );


  nor
  g3241
  (
    n2964,
    n2120,
    n2610,
    n2894,
    n692
  );


  or
  g3242
  (
    n3350,
    n2880,
    n2570,
    n2146,
    n2465
  );


  nor
  g3243
  (
    n3089,
    n1587,
    n2351,
    n1557,
    n2453
  );


  xor
  g3244
  (
    n3270,
    n2849,
    n641,
    n1712,
    n677
  );


  nor
  g3245
  (
    n3284,
    n723,
    n2554,
    n2731,
    n1867
  );


  xnor
  g3246
  (
    n3379,
    n2416,
    n2819,
    n2650,
    n2080
  );


  nor
  g3247
  (
    n2966,
    n2126,
    n2891,
    n1523,
    n1835
  );


  nor
  g3248
  (
    n3067,
    n2371,
    n2428,
    n2060,
    n717
  );


  xnor
  g3249
  (
    n3099,
    n1882,
    n590,
    n696,
    n705
  );


  xnor
  g3250
  (
    n3323,
    n2933,
    n1537,
    n1914,
    n715
  );


  or
  g3251
  (
    n3397,
    n2456,
    n1637,
    n1722,
    n2939
  );


  xnor
  g3252
  (
    n3091,
    n2002,
    n2212,
    n2903,
    n2769
  );


  xnor
  g3253
  (
    n3338,
    n2887,
    n1568,
    n2275,
    n2733
  );


  xnor
  g3254
  (
    n3189,
    n1778,
    n2200,
    n2640,
    n1900
  );


  xnor
  g3255
  (
    n3155,
    n2923,
    n1747,
    n1855,
    n1866
  );


  xor
  g3256
  (
    n3260,
    n2886,
    n2159,
    n1765,
    n2738
  );


  xor
  g3257
  (
    n3324,
    n2902,
    n2311,
    n2046,
    n2316
  );


  nand
  g3258
  (
    n3235,
    n593,
    n1657,
    n2117,
    n2335
  );


  or
  g3259
  (
    n2967,
    n1710,
    n2168,
    n2943,
    n605
  );


  nand
  g3260
  (
    n3331,
    n2846,
    n2756,
    n2241,
    n1675
  );


  nor
  g3261
  (
    n3212,
    n2502,
    n604,
    n2932,
    n1994
  );


  nor
  g3262
  (
    n3293,
    n2751,
    n1983,
    n2113,
    n2489
  );


  nand
  g3263
  (
    n3115,
    n2741,
    n2904,
    n574,
    n2614
  );


  xnor
  g3264
  (
    n3076,
    n1658,
    n2722,
    n2949,
    n2216
  );


  or
  g3265
  (
    n3391,
    n565,
    n2885,
    n2568,
    n1890
  );


  and
  g3266
  (
    n2977,
    n2029,
    n2668,
    n603,
    n2805
  );


  and
  g3267
  (
    n3059,
    n2872,
    n664,
    n1817,
    n2285
  );


  or
  g3268
  (
    n3308,
    n2516,
    n600,
    n1815,
    n1806
  );


  and
  g3269
  (
    n3125,
    n2868,
    n2452,
    n2091,
    n2254
  );


  xor
  g3270
  (
    n3122,
    n2525,
    n2868,
    n2812,
    n2443
  );


  xnor
  g3271
  (
    n3124,
    n2014,
    n2545,
    n2885,
    n2830
  );


  and
  g3272
  (
    n3221,
    n2874,
    n2194,
    n2878,
    n1670
  );


  and
  g3273
  (
    n3333,
    n2081,
    n2125,
    n2306,
    n1511
  );


  nor
  g3274
  (
    n3381,
    n1652,
    n1552,
    n2020,
    n2299
  );


  or
  g3275
  (
    n3348,
    n2824,
    n2496,
    n2714,
    n2622
  );


  or
  g3276
  (
    n3190,
    n1966,
    n2218,
    n1614,
    n2720
  );


  xor
  g3277
  (
    n3301,
    n2643,
    n578,
    n2409,
    n609
  );


  and
  g3278
  (
    n3249,
    n2925,
    n1650,
    n2684,
    n1961
  );


  nor
  g3279
  (
    n3157,
    n1530,
    n2073,
    n2370,
    n2806
  );


  xnor
  g3280
  (
    n3039,
    n2547,
    n1859,
    n2902,
    n2924
  );


  nand
  g3281
  (
    n3013,
    n2310,
    n2532,
    n1843,
    n2188
  );


  and
  g3282
  (
    n3340,
    n1941,
    n1821,
    n1992,
    n1982
  );


  xnor
  g3283
  (
    n3027,
    n2043,
    n2136,
    n2872,
    n2896
  );


  nor
  g3284
  (
    n3353,
    n667,
    n559,
    n1580,
    n2406
  );


  nor
  g3285
  (
    n3250,
    n2470,
    n2237,
    n2379,
    n653
  );


  and
  g3286
  (
    n3376,
    n1607,
    n1566,
    n2906,
    n2215
  );


  xor
  g3287
  (
    n3062,
    n1948,
    n1561,
    n1700,
    n1520
  );


  and
  g3288
  (
    n2971,
    n1732,
    n680,
    n1701,
    n2719
  );


  and
  g3289
  (
    n3009,
    n708,
    n1730,
    n1542,
    n2209
  );


  xnor
  g3290
  (
    n3096,
    n1728,
    n1697,
    n1553,
    n2929
  );


  xor
  g3291
  (
    n3389,
    n1678,
    n2025,
    n712,
    n1664
  );


  xor
  g3292
  (
    n3261,
    n2868,
    n2541,
    n2267,
    n2633
  );


  xnor
  g3293
  (
    n2963,
    n2337,
    n2702,
    n2395,
    n2688
  );


  nor
  g3294
  (
    n3068,
    n2881,
    n706,
    n2774,
    n2017
  );


  xor
  g3295
  (
    n2994,
    n2164,
    n1968,
    n1729,
    n649
  );


  nand
  g3296
  (
    n3306,
    n1661,
    n1916,
    n2794,
    n2040
  );


  xnor
  g3297
  (
    KeyWire_0_6,
    n2214,
    n1604,
    n2521,
    n1783
  );


  xnor
  g3298
  (
    n3318,
    n595,
    n2494,
    n1908,
    n1995
  );


  and
  g3299
  (
    n3154,
    n2940,
    n2538,
    n1970,
    n1695
  );


  xnor
  g3300
  (
    KeyWire_0_3,
    n2522,
    n1569,
    n2791,
    n2907
  );


  xor
  g3301
  (
    n3188,
    n2890,
    n2848,
    n1683,
    n2201
  );


  and
  g3302
  (
    n3201,
    n718,
    n2157,
    n2177,
    n2586
  );


  and
  g3303
  (
    n3031,
    n1745,
    n2198,
    n2912,
    n713
  );


  nor
  g3304
  (
    n3136,
    n2251,
    n1868,
    n1839,
    n2449
  );


  nor
  g3305
  (
    n3082,
    n2431,
    n1654,
    n2898,
    n2658
  );


  and
  g3306
  (
    n2972,
    n2369,
    n2433,
    n2912,
    n1719
  );


  or
  g3307
  (
    n2985,
    n2133,
    n2151,
    n2262,
    n1659
  );


  or
  g3308
  (
    n3199,
    n1812,
    n2930,
    n2361,
    n2027
  );


  and
  g3309
  (
    n3356,
    n2068,
    n2850,
    n2637,
    n2820
  );


  xnor
  g3310
  (
    n3126,
    n2276,
    n2836,
    n560,
    n2273
  );


  or
  g3311
  (
    n3325,
    n2906,
    n2813,
    n2257,
    n2933
  );


  or
  g3312
  (
    KeyWire_0_29,
    n2095,
    n1510,
    n1705,
    n1742
  );


  nor
  g3313
  (
    n3037,
    n614,
    n2906,
    n2103,
    n2655
  );


  nor
  g3314
  (
    n3374,
    n689,
    n623,
    n2196,
    n2513
  );


  or
  g3315
  (
    n2995,
    n2654,
    n2611,
    n2927,
    n2265
  );


  or
  g3316
  (
    n3116,
    n2049,
    n1615,
    n1907,
    n2175
  );


  or
  g3317
  (
    n3362,
    n2921,
    n2620,
    n2777,
    n2013
  );


  nand
  g3318
  (
    n3033,
    n2941,
    n2725,
    n2399,
    n1873
  );


  nor
  g3319
  (
    n3298,
    n668,
    n2270,
    n672,
    n1509
  );


  nor
  g3320
  (
    n3366,
    n599,
    n1704,
    n2931,
    n2897
  );


  xor
  g3321
  (
    n3169,
    n2024,
    n2438,
    n2015,
    n2911
  );


  nor
  g3322
  (
    n3174,
    n2154,
    n2808,
    n1797,
    n684
  );


  nand
  g3323
  (
    n3315,
    n1829,
    n2790,
    n2535,
    n1823
  );


  and
  g3324
  (
    n3072,
    n2389,
    n610,
    n2054,
    n1620
  );


  xor
  g3325
  (
    n3302,
    n2451,
    n2161,
    n2296,
    n1912
  );


  xnor
  g3326
  (
    n3111,
    n1825,
    n1795,
    n2314,
    n2278
  );


  and
  g3327
  (
    n3024,
    n2086,
    n2882,
    n2388,
    n2001
  );


  xnor
  g3328
  (
    n3267,
    n2721,
    n2398,
    n2475,
    n1864
  );


  nor
  g3329
  (
    n3265,
    n691,
    n2402,
    n2786,
    n2598
  );


  or
  g3330
  (
    n3392,
    n2876,
    n2664,
    n2935,
    n1924
  );


  nand
  g3331
  (
    n3307,
    n2930,
    n2507,
    n1593,
    n1573
  );


  and
  g3332
  (
    n3151,
    n2618,
    n2835,
    n2435,
    n2531
  );


  nor
  g3333
  (
    n3269,
    n1708,
    n2028,
    n2763,
    n2920
  );


  nand
  g3334
  (
    n3334,
    n2062,
    n2683,
    n2946,
    n2034
  );


  nand
  g3335
  (
    n3149,
    n2940,
    n2204,
    n1643,
    n1801
  );


  xor
  g3336
  (
    n3256,
    n657,
    n612,
    n2420,
    n2097
  );


  nand
  g3337
  (
    n3036,
    n602,
    n2926,
    n2142,
    n1581
  );


  or
  g3338
  (
    n3097,
    n2597,
    n2183,
    n2800,
    n2537
  );


  or
  g3339
  (
    n3215,
    n2374,
    n2689,
    n638,
    n1933
  );


  xor
  g3340
  (
    n3109,
    n2563,
    n2645,
    n596,
    n2907
  );


  nand
  g3341
  (
    n3152,
    n2483,
    n1903,
    n2575,
    n1911
  );


  xnor
  g3342
  (
    n3336,
    n1930,
    n2052,
    n2170,
    n2919
  );


  nor
  g3343
  (
    n3378,
    n2225,
    n2895,
    n2564,
    n1875
  );


  nand
  g3344
  (
    n3263,
    n2384,
    n2364,
    n2851,
    n2881
  );


  xnor
  g3345
  (
    n2953,
    n2365,
    n2626,
    n2706,
    n2492
  );


  nand
  g3346
  (
    n3088,
    n720,
    n1883,
    n2495,
    n2481
  );


  or
  g3347
  (
    n2976,
    n2304,
    n2186,
    n2602,
    n2116
  );


  and
  g3348
  (
    n3297,
    n1808,
    n1802,
    n594,
    n2245
  );


  or
  g3349
  (
    n3160,
    n1844,
    n2207,
    n2886,
    n608
  );


  xnor
  g3350
  (
    n3164,
    n1667,
    n1564,
    n1600,
    n2067
  );


  and
  g3351
  (
    n3026,
    n2793,
    n2166,
    n2589,
    n2639
  );


  or
  g3352
  (
    n3262,
    n2707,
    n2789,
    n558,
    n2472
  );


  xor
  g3353
  (
    n3228,
    n1576,
    n1782,
    n2077,
    n1887
  );


  nand
  g3354
  (
    n3287,
    n2948,
    n2629,
    n2190,
    n601
  );


  and
  g3355
  (
    n3369,
    n2356,
    n2325,
    n563,
    n702
  );


  and
  g3356
  (
    n3202,
    n2544,
    n2913,
    n1856,
    n2413
  );


  or
  g3357
  (
    n3118,
    n1993,
    n2896,
    n2952,
    n1959
  );


  nor
  g3358
  (
    n3100,
    n1518,
    n2932,
    n1928,
    n2132
  );


  nand
  g3359
  (
    n3134,
    n2500,
    n1642,
    n2176,
    n1682
  );


  nand
  g3360
  (
    n3094,
    n2651,
    n2934,
    n1731,
    n2009
  );


  and
  g3361
  (
    n3173,
    n2339,
    n592,
    n2326,
    n2466
  );


  and
  g3362
  (
    n3110,
    n2269,
    n2087,
    n1926,
    n1653
  );


  and
  g3363
  (
    n3144,
    n572,
    n1543,
    n2636,
    n701
  );


  and
  g3364
  (
    n3060,
    n1980,
    n1688,
    n2893,
    n2272
  );


  nand
  g3365
  (
    n3408,
    n3068,
    n3230,
    n3087,
    n3203
  );


  nand
  g3366
  (
    n3448,
    n3222,
    n3323,
    n3310,
    n2993
  );


  or
  g3367
  (
    n3410,
    n3034,
    n3114,
    n3062,
    n3107
  );


  nor
  g3368
  (
    n3466,
    n3022,
    n3132,
    n2990,
    n3357
  );


  or
  g3369
  (
    n3441,
    n3227,
    n3264,
    n3290,
    n3151
  );


  and
  g3370
  (
    n3403,
    n3375,
    n3024,
    n3214,
    n3134
  );


  or
  g3371
  (
    n3501,
    n3250,
    n3188,
    n3113,
    n3279
  );


  and
  g3372
  (
    n3415,
    n2956,
    n3398,
    n3352,
    n3268
  );


  nor
  g3373
  (
    n3507,
    n3328,
    n3297,
    n3054,
    n2968
  );


  xor
  g3374
  (
    n3449,
    n3187,
    n3213,
    n3365,
    n3347
  );


  xnor
  g3375
  (
    n3499,
    n2964,
    n3399,
    n3017,
    n3000
  );


  or
  g3376
  (
    n3480,
    n3393,
    n2982,
    n3362,
    n3021
  );


  nand
  g3377
  (
    n3496,
    n3124,
    n3023,
    n2997,
    n3197
  );


  and
  g3378
  (
    n3454,
    n3096,
    n2991,
    n3207,
    n3129
  );


  xnor
  g3379
  (
    n3478,
    n3205,
    n3261,
    n3329,
    n3358
  );


  xor
  g3380
  (
    n3412,
    n3144,
    n3141,
    n3184,
    n2959
  );


  or
  g3381
  (
    n3430,
    n3066,
    n3104,
    n3039,
    n3179
  );


  nor
  g3382
  (
    n3492,
    n2963,
    n3135,
    n3170,
    n3217
  );


  xor
  g3383
  (
    n3498,
    n2977,
    n3225,
    n3138,
    n2966
  );


  xor
  g3384
  (
    n3468,
    n3314,
    n3367,
    n3341,
    n3288
  );


  and
  g3385
  (
    n3455,
    n3254,
    n3089,
    n3007,
    n3074
  );


  xor
  g3386
  (
    n3413,
    n3048,
    n3332,
    n3152,
    n3313
  );


  nor
  g3387
  (
    n3424,
    n3277,
    n3094,
    n3031,
    n3337
  );


  xor
  g3388
  (
    n3457,
    n2979,
    n3292,
    n3164,
    n3052
  );


  xnor
  g3389
  (
    n3489,
    n3079,
    n3145,
    n2976,
    n3005
  );


  xor
  g3390
  (
    n3476,
    n3208,
    n3331,
    n3065,
    n3162
  );


  xnor
  g3391
  (
    n3479,
    n3231,
    n2996,
    n2969,
    n3339
  );


  nor
  g3392
  (
    n3422,
    n3157,
    n3333,
    n2992,
    n3026
  );


  xor
  g3393
  (
    n3405,
    n3287,
    n3259,
    n3055,
    n3371
  );


  or
  g3394
  (
    n3429,
    n3088,
    n3059,
    n3140,
    n3042
  );


  xor
  g3395
  (
    n3426,
    n3016,
    n3040,
    n3274,
    n3117
  );


  nand
  g3396
  (
    n3447,
    n3190,
    n3136,
    n3298,
    n3169
  );


  xor
  g3397
  (
    n3481,
    n3180,
    n3330,
    n3355,
    n3194
  );


  xnor
  g3398
  (
    n3484,
    n3370,
    n3378,
    n3100,
    n3098
  );


  nand
  g3399
  (
    n3470,
    n3221,
    n3252,
    n3216,
    n2962
  );


  xor
  g3400
  (
    n3474,
    n3201,
    n3251,
    n3368,
    n3106
  );


  and
  g3401
  (
    n3488,
    n3206,
    n3155,
    n3245,
    n3163
  );


  xnor
  g3402
  (
    n3450,
    n3272,
    n2961,
    n3032,
    n3383
  );


  xnor
  g3403
  (
    n3465,
    n3168,
    n3395,
    n3043,
    n3236
  );


  nor
  g3404
  (
    n3458,
    n3020,
    n3220,
    n3004,
    n3072
  );


  xor
  g3405
  (
    n3434,
    n3076,
    n3182,
    n3394,
    n3030
  );


  and
  g3406
  (
    n3491,
    n3340,
    n3263,
    n3183,
    n3189
  );


  nand
  g3407
  (
    n3443,
    n2989,
    n3050,
    n3233,
    n3051
  );


  xor
  g3408
  (
    n3437,
    n3064,
    n3359,
    n3239,
    n3391
  );


  nand
  g3409
  (
    n3475,
    n2978,
    n3271,
    n3353,
    n3160
  );


  nor
  g3410
  (
    n3417,
    n3255,
    n3033,
    n3177,
    n3266
  );


  nor
  g3411
  (
    n3510,
    n3047,
    n3241,
    n3092,
    n3118
  );


  or
  g3412
  (
    n3504,
    n3396,
    n3384,
    n3120,
    n3376
  );


  nor
  g3413
  (
    n3414,
    n3278,
    n3166,
    n3283,
    n3161
  );


  nor
  g3414
  (
    KeyWire_0_22,
    n3348,
    n3081,
    n3270,
    n2988
  );


  xnor
  g3415
  (
    n3461,
    n3006,
    n3149,
    n3176,
    n3392
  );


  and
  g3416
  (
    n3446,
    n3008,
    n3351,
    n3281,
    n3148
  );


  xor
  g3417
  (
    n3485,
    n3125,
    n3354,
    n3010,
    n3025
  );


  nor
  g3418
  (
    n3432,
    n3364,
    n3105,
    n3244,
    n3069
  );


  xnor
  g3419
  (
    n3503,
    n3049,
    n3301,
    n3192,
    n3285
  );


  nor
  g3420
  (
    n3460,
    n3058,
    n3037,
    n3318,
    n3174
  );


  nor
  g3421
  (
    n3471,
    n3173,
    n3334,
    n3369,
    n3193
  );


  xnor
  g3422
  (
    n3469,
    n3265,
    n3284,
    n3103,
    n3159
  );


  xnor
  g3423
  (
    n3512,
    n3224,
    n3002,
    n2999,
    n3322
  );


  nand
  g3424
  (
    n3459,
    n3046,
    n3146,
    n3232,
    n3204
  );


  or
  g3425
  (
    n3483,
    n3085,
    n3108,
    n3299,
    n3181
  );


  nand
  g3426
  (
    n3444,
    n3360,
    n3015,
    n3202,
    n3260
  );


  nor
  g3427
  (
    n3473,
    n3209,
    n3242,
    n3372,
    n3253
  );


  xor
  g3428
  (
    n3464,
    n2957,
    n3400,
    n3112,
    n3029
  );


  or
  g3429
  (
    n3453,
    n2985,
    n3133,
    n2974,
    n3056
  );


  or
  g3430
  (
    n3467,
    n3321,
    n3045,
    n3116,
    n3027
  );


  xor
  g3431
  (
    n3497,
    n3178,
    n3342,
    n3309,
    n3256
  );


  nor
  g3432
  (
    n3442,
    n3061,
    n2995,
    n3381,
    n3044
  );


  or
  g3433
  (
    n3490,
    n3228,
    n3386,
    n3142,
    n3316
  );


  or
  g3434
  (
    n3416,
    n3198,
    n3101,
    n3057,
    n2984
  );


  xor
  g3435
  (
    n3486,
    n3327,
    n3326,
    n3280,
    n3397
  );


  nor
  g3436
  (
    n3508,
    n3093,
    n3035,
    n3175,
    n3003
  );


  xnor
  g3437
  (
    n3477,
    n3078,
    n3382,
    n3165,
    n3041
  );


  xnor
  g3438
  (
    n3511,
    n3257,
    n3122,
    n3086,
    n3235
  );


  or
  g3439
  (
    n3433,
    n3223,
    n3338,
    n3186,
    n2986
  );


  nand
  g3440
  (
    n3463,
    n3071,
    n2994,
    n2987,
    n3014
  );


  xor
  g3441
  (
    n3419,
    n3325,
    n2955,
    n3345,
    n3293
  );


  xnor
  g3442
  (
    n3494,
    n3147,
    n3324,
    n3269,
    n3246
  );


  or
  g3443
  (
    n3482,
    n2980,
    n3077,
    n3247,
    n3082
  );


  or
  g3444
  (
    n3456,
    n3387,
    n3249,
    n3097,
    n3080
  );


  nor
  g3445
  (
    n3425,
    n3215,
    n3300,
    n3028,
    n3315
  );


  nor
  g3446
  (
    n3505,
    n2971,
    n3248,
    n2983,
    n3361
  );


  xnor
  g3447
  (
    n3401,
    n3126,
    n3294,
    n3139,
    n3090
  );


  or
  g3448
  (
    n3502,
    n3350,
    n3200,
    n3356,
    n3019
  );


  nand
  g3449
  (
    n3495,
    n3154,
    n3291,
    n3060,
    n3335
  );


  xor
  g3450
  (
    n3452,
    n3067,
    n2970,
    n3267,
    n3380
  );


  or
  g3451
  (
    n3509,
    n3238,
    n3296,
    n3091,
    n3343
  );


  and
  g3452
  (
    n3440,
    n3075,
    n3128,
    n3303,
    n3185
  );


  nor
  g3453
  (
    n3500,
    n3011,
    n3336,
    n3258,
    n3262
  );


  or
  g3454
  (
    n3418,
    n3095,
    n3363,
    n3304,
    n3115
  );


  nand
  g3455
  (
    n3402,
    n3346,
    n3084,
    n3317,
    n3312
  );


  xor
  g3456
  (
    n3406,
    n3289,
    n3385,
    n3012,
    n3374
  );


  and
  g3457
  (
    n3439,
    n3110,
    n3295,
    n3156,
    n3311
  );


  or
  g3458
  (
    n3451,
    n3109,
    n3275,
    n2972,
    n3036
  );


  xnor
  g3459
  (
    KeyWire_0_13,
    n3349,
    n3237,
    n3276,
    n3171
  );


  nand
  g3460
  (
    n3472,
    n3111,
    n3196,
    n3273,
    n3282
  );


  nand
  g3461
  (
    n3428,
    n3240,
    n3308,
    n3320,
    n3377
  );


  nand
  g3462
  (
    n3427,
    n2998,
    n3307,
    n2958,
    n3199
  );


  xor
  g3463
  (
    n3506,
    n3153,
    n3243,
    n3131,
    n3195
  );


  xor
  g3464
  (
    n3421,
    n3305,
    n2981,
    n3212,
    n3302
  );


  nor
  g3465
  (
    n3420,
    n3390,
    n3226,
    n3319,
    n3123
  );


  nand
  g3466
  (
    n3435,
    n2960,
    n3211,
    n3013,
    n3083
  );


  and
  g3467
  (
    n3438,
    n3172,
    n3001,
    n3070,
    n2973
  );


  or
  g3468
  (
    n3436,
    n3102,
    n3018,
    n3379,
    n3210
  );


  or
  g3469
  (
    n3445,
    n3127,
    n3219,
    n3167,
    n3137
  );


  or
  g3470
  (
    n3407,
    n3099,
    n3234,
    n3150,
    n2975
  );


  xnor
  g3471
  (
    n3411,
    n3130,
    n3389,
    n2954,
    n2965
  );


  nand
  g3472
  (
    n3431,
    n3053,
    n3366,
    n3143,
    n3344
  );


  xor
  g3473
  (
    n3404,
    n3073,
    n3229,
    n3038,
    n3121
  );


  nand
  g3474
  (
    n3487,
    n2967,
    n3388,
    n3286,
    n3218
  );


  nand
  g3475
  (
    n3423,
    n2953,
    n3158,
    n3063,
    n3009
  );


  nand
  g3476
  (
    n3462,
    n3119,
    n3191,
    n3373,
    n3306
  );


  and
  g3477
  (
    n3520,
    n3450,
    n3468,
    n3405,
    n3414
  );


  nor
  g3478
  (
    n3515,
    n3466,
    n3461,
    n3483,
    n3492
  );


  nor
  g3479
  (
    n3516,
    n3420,
    n3409,
    n3509,
    n3458
  );


  or
  g3480
  (
    n3532,
    n3453,
    n3472,
    n3448,
    n3449
  );


  xnor
  g3481
  (
    n3538,
    n3498,
    n3417,
    n3457,
    n3416
  );


  nor
  g3482
  (
    n3537,
    n3402,
    n3452,
    n3506,
    n3488
  );


  xor
  g3483
  (
    n3536,
    n3493,
    n3428,
    n3437,
    n3475
  );


  or
  g3484
  (
    n3523,
    n3412,
    n3486,
    n3438,
    n3499
  );


  nor
  g3485
  (
    n3521,
    n3446,
    n3403,
    n3445,
    n3463
  );


  xor
  g3486
  (
    n3514,
    n3429,
    n3441,
    n3422,
    n3454
  );


  xnor
  g3487
  (
    n3525,
    n3508,
    n3465,
    n3479,
    n3431
  );


  xnor
  g3488
  (
    n3513,
    n3502,
    n3482,
    n3473,
    n3469
  );


  nor
  g3489
  (
    n3526,
    n3408,
    n3467,
    n3497,
    n3470
  );


  nor
  g3490
  (
    n3534,
    n3451,
    n3415,
    n3474,
    n3510
  );


  xor
  g3491
  (
    n3528,
    n3495,
    n3496,
    n3478,
    n3512
  );


  xnor
  g3492
  (
    n3540,
    n3443,
    n3411,
    n3435,
    n3494
  );


  xor
  g3493
  (
    n3524,
    n3421,
    n3442,
    n3434,
    n3455
  );


  and
  g3494
  (
    n3519,
    n3410,
    n3406,
    n3501,
    n3476
  );


  xor
  g3495
  (
    n3539,
    n3511,
    n3419,
    n3464,
    n3433
  );


  xor
  g3496
  (
    n3527,
    n3423,
    n3430,
    n3503,
    n3490
  );


  xor
  g3497
  (
    n3533,
    n3500,
    n3484,
    n3407,
    n3481
  );


  nand
  g3498
  (
    n3530,
    n3427,
    n3480,
    n3491,
    n3444
  );


  nor
  g3499
  (
    n3522,
    n3447,
    n3505,
    n3485,
    n3418
  );


  xnor
  g3500
  (
    n3529,
    n3425,
    n3507,
    n3440,
    n3487
  );


  xnor
  g3501
  (
    n3517,
    n3504,
    n3456,
    n3459,
    n3462
  );


  nor
  g3502
  (
    n3531,
    n3436,
    n3477,
    n3424,
    n3439
  );


  and
  g3503
  (
    n3518,
    n3401,
    n3489,
    n3404,
    n3432
  );


  or
  g3504
  (
    n3535,
    n3460,
    n3426,
    n3471,
    n3413
  );


  nand
  g3505
  (
    n3546,
    n3522,
    n3531,
    n3538,
    n3514
  );


  nand
  g3506
  (
    n3543,
    n3526,
    n3516,
    n3535,
    n3521
  );


  nor
  g3507
  (
    n3541,
    n3513,
    n3519,
    n3515,
    n3528
  );


  nand
  g3508
  (
    n3542,
    n3540,
    n3537,
    n3517,
    n3536
  );


  and
  g3509
  (
    n3544,
    n3518,
    n3523,
    n3539,
    n3525
  );


  nor
  g3510
  (
    n3545,
    n3527,
    n3524,
    n3532,
    n3530
  );


  or
  g3511
  (
    n3547,
    n3534,
    n3533,
    n3520,
    n3529
  );


  xnor
  KeyGate_0_0
  (
    n1767,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n3034,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n3003,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n3393,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n3229,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n1385,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n3005,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n860,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1322,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n2759,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n544,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1440,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n2575,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n3409,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n2687,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n2678,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n2700,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n3029,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n907,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n350,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n2599,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1731,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n3493,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n2988,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n2130,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n2576,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n2890,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1153,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n2500,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n3043,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n996,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n3330,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

