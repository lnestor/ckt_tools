// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1368_61_7 written by SynthGen on 2021/05/24 19:42:18
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1368_61_7 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20,
 n1085, n1156, n1190, n1183, n1187, n1186, n1184, n1181,
 n1182, n1207, n1379, n1374, n1384, n1376, n1383, n1387,
 n1381, n1385, n1382, n1377, n1378, n1373, n1380, n1388,
 n1375, n1386);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20;

output n1085, n1156, n1190, n1183, n1187, n1186, n1184, n1181,
 n1182, n1207, n1379, n1374, n1384, n1376, n1383, n1387,
 n1381, n1385, n1382, n1377, n1378, n1373, n1380, n1388,
 n1375, n1386;

wire n21, n22, n23, n24, n25, n26, n27, n28,
 n29, n30, n31, n32, n33, n34, n35, n36,
 n37, n38, n39, n40, n41, n42, n43, n44,
 n45, n46, n47, n48, n49, n50, n51, n52,
 n53, n54, n55, n56, n57, n58, n59, n60,
 n61, n62, n63, n64, n65, n66, n67, n68,
 n69, n70, n71, n72, n73, n74, n75, n76,
 n77, n78, n79, n80, n81, n82, n83, n84,
 n85, n86, n87, n88, n89, n90, n91, n92,
 n93, n94, n95, n96, n97, n98, n99, n100,
 n101, n102, n103, n104, n105, n106, n107, n108,
 n109, n110, n111, n112, n113, n114, n115, n116,
 n117, n118, n119, n120, n121, n122, n123, n124,
 n125, n126, n127, n128, n129, n130, n131, n132,
 n133, n134, n135, n136, n137, n138, n139, n140,
 n141, n142, n143, n144, n145, n146, n147, n148,
 n149, n150, n151, n152, n153, n154, n155, n156,
 n157, n158, n159, n160, n161, n162, n163, n164,
 n165, n166, n167, n168, n169, n170, n171, n172,
 n173, n174, n175, n176, n177, n178, n179, n180,
 n181, n182, n183, n184, n185, n186, n187, n188,
 n189, n190, n191, n192, n193, n194, n195, n196,
 n197, n198, n199, n200, n201, n202, n203, n204,
 n205, n206, n207, n208, n209, n210, n211, n212,
 n213, n214, n215, n216, n217, n218, n219, n220,
 n221, n222, n223, n224, n225, n226, n227, n228,
 n229, n230, n231, n232, n233, n234, n235, n236,
 n237, n238, n239, n240, n241, n242, n243, n244,
 n245, n246, n247, n248, n249, n250, n251, n252,
 n253, n254, n255, n256, n257, n258, n259, n260,
 n261, n262, n263, n264, n265, n266, n267, n268,
 n269, n270, n271, n272, n273, n274, n275, n276,
 n277, n278, n279, n280, n281, n282, n283, n284,
 n285, n286, n287, n288, n289, n290, n291, n292,
 n293, n294, n295, n296, n297, n298, n299, n300,
 n301, n302, n303, n304, n305, n306, n307, n308,
 n309, n310, n311, n312, n313, n314, n315, n316,
 n317, n318, n319, n320, n321, n322, n323, n324,
 n325, n326, n327, n328, n329, n330, n331, n332,
 n333, n334, n335, n336, n337, n338, n339, n340,
 n341, n342, n343, n344, n345, n346, n347, n348,
 n349, n350, n351, n352, n353, n354, n355, n356,
 n357, n358, n359, n360, n361, n362, n363, n364,
 n365, n366, n367, n368, n369, n370, n371, n372,
 n373, n374, n375, n376, n377, n378, n379, n380,
 n381, n382, n383, n384, n385, n386, n387, n388,
 n389, n390, n391, n392, n393, n394, n395, n396,
 n397, n398, n399, n400, n401, n402, n403, n404,
 n405, n406, n407, n408, n409, n410, n411, n412,
 n413, n414, n415, n416, n417, n418, n419, n420,
 n421, n422, n423, n424, n425, n426, n427, n428,
 n429, n430, n431, n432, n433, n434, n435, n436,
 n437, n438, n439, n440, n441, n442, n443, n444,
 n445, n446, n447, n448, n449, n450, n451, n452,
 n453, n454, n455, n456, n457, n458, n459, n460,
 n461, n462, n463, n464, n465, n466, n467, n468,
 n469, n470, n471, n472, n473, n474, n475, n476,
 n477, n478, n479, n480, n481, n482, n483, n484,
 n485, n486, n487, n488, n489, n490, n491, n492,
 n493, n494, n495, n496, n497, n498, n499, n500,
 n501, n502, n503, n504, n505, n506, n507, n508,
 n509, n510, n511, n512, n513, n514, n515, n516,
 n517, n518, n519, n520, n521, n522, n523, n524,
 n525, n526, n527, n528, n529, n530, n531, n532,
 n533, n534, n535, n536, n537, n538, n539, n540,
 n541, n542, n543, n544, n545, n546, n547, n548,
 n549, n550, n551, n552, n553, n554, n555, n556,
 n557, n558, n559, n560, n561, n562, n563, n564,
 n565, n566, n567, n568, n569, n570, n571, n572,
 n573, n574, n575, n576, n577, n578, n579, n580,
 n581, n582, n583, n584, n585, n586, n587, n588,
 n589, n590, n591, n592, n593, n594, n595, n596,
 n597, n598, n599, n600, n601, n602, n603, n604,
 n605, n606, n607, n608, n609, n610, n611, n612,
 n613, n614, n615, n616, n617, n618, n619, n620,
 n621, n622, n623, n624, n625, n626, n627, n628,
 n629, n630, n631, n632, n633, n634, n635, n636,
 n637, n638, n639, n640, n641, n642, n643, n644,
 n645, n646, n647, n648, n649, n650, n651, n652,
 n653, n654, n655, n656, n657, n658, n659, n660,
 n661, n662, n663, n664, n665, n666, n667, n668,
 n669, n670, n671, n672, n673, n674, n675, n676,
 n677, n678, n679, n680, n681, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n758, n759, n760, n761, n762, n763, n764,
 n765, n766, n767, n768, n769, n770, n771, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n840, n841, n842, n843, n844,
 n845, n846, n847, n848, n849, n850, n851, n852,
 n853, n854, n855, n856, n857, n858, n859, n860,
 n861, n862, n863, n864, n865, n866, n867, n868,
 n869, n870, n871, n872, n873, n874, n875, n876,
 n877, n878, n879, n880, n881, n882, n883, n884,
 n885, n886, n887, n888, n889, n890, n891, n892,
 n893, n894, n895, n896, n897, n898, n899, n900,
 n901, n902, n903, n904, n905, n906, n907, n908,
 n909, n910, n911, n912, n913, n914, n915, n916,
 n917, n918, n919, n920, n921, n922, n923, n924,
 n925, n926, n927, n928, n929, n930, n931, n932,
 n933, n934, n935, n936, n937, n938, n939, n940,
 n941, n942, n943, n944, n945, n946, n947, n948,
 n949, n950, n951, n952, n953, n954, n955, n956,
 n957, n958, n959, n960, n961, n962, n963, n964,
 n965, n966, n967, n968, n969, n970, n971, n972,
 n973, n974, n975, n976, n977, n978, n979, n980,
 n981, n982, n983, n984, n985, n986, n987, n988,
 n989, n990, n991, n992, n993, n994, n995, n996,
 n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
 n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
 n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
 n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
 n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
 n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
 n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
 n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
 n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
 n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
 n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
 n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
 n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
 n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
 n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
 n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
 n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
 n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
 n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
 n1150, n1151, n1152, n1153, n1154, n1155, n1157, n1158,
 n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
 n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
 n1175, n1176, n1177, n1178, n1179, n1180, n1185, n1188,
 n1189, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
 n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
 n1206, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
 n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
 n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
 n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
 n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
 n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
 n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
 n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
 n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
 n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
 n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
 n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
 n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
 n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
 n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
 n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
 n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
 n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
 n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
 n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
 n1367, n1368, n1369, n1370, n1371, n1372;

buf  g0 (n50, n7);
buf  g1 (n36, n13);
buf  g2 (n22, n10);
not  g3 (n64, n3);
not  g4 (n31, n8);
buf  g5 (n63, n4);
not  g6 (n52, n10);
not  g7 (n54, n2);
not  g8 (n60, n3);
buf  g9 (n53, n8);
not  g10 (n41, n9);
buf  g11 (n33, n6);
not  g12 (n25, n2);
buf  g13 (n48, n3);
not  g14 (n40, n4);
buf  g15 (n62, n1);
buf  g16 (n42, n5);
not  g17 (n29, n10);
not  g18 (n47, n9);
buf  g19 (n57, n13);
buf  g20 (n55, n8);
not  g21 (n38, n4);
not  g22 (n69, n7);
buf  g23 (n49, n11);
not  g24 (n61, n1);
buf  g25 (n70, n9);
not  g26 (n56, n9);
not  g27 (n45, n7);
buf  g28 (n34, n7);
not  g29 (n46, n12);
not  g30 (n23, n6);
not  g31 (n68, n12);
not  g32 (n43, n6);
not  g33 (n26, n5);
buf  g34 (n44, n4);
buf  g35 (n72, n13);
buf  g36 (n28, n5);
not  g37 (n24, n2);
not  g38 (n21, n1);
not  g39 (n67, n11);
not  g40 (n39, n11);
not  g41 (n32, n10);
not  g42 (n35, n6);
not  g43 (n37, n3);
not  g44 (n59, n13);
buf  g45 (n65, n11);
not  g46 (n27, n12);
not  g47 (n51, n1);
buf  g48 (n71, n8);
not  g49 (n58, n5);
buf  g50 (n66, n2);
not  g51 (n30, n12);
buf  g52 (n77, n23);
buf  g53 (n74, n21);
buf  g54 (n81, n23);
buf  g55 (n85, n22);
not  g56 (n80, n22);
buf  g57 (n88, n21);
buf  g58 (n79, n23);
buf  g59 (n82, n24);
buf  g60 (n76, n21);
not  g61 (n78, n22);
buf  g62 (n73, n22);
buf  g63 (n75, n24);
not  g64 (n87, n21);
buf  g65 (n83, n24);
buf  g66 (n84, n24);
not  g67 (n86, n23);
not  g68 (n121, n88);
buf  g69 (n111, n75);
not  g70 (n118, n86);
not  g71 (n95, n75);
not  g72 (n136, n84);
not  g73 (n130, n79);
buf  g74 (n92, n88);
buf  g75 (n116, n84);
buf  g76 (n123, n82);
not  g77 (n151, n79);
not  g78 (n102, n87);
buf  g79 (n140, n83);
buf  g80 (n104, n81);
buf  g81 (n97, n76);
not  g82 (n139, n77);
buf  g83 (n101, n80);
not  g84 (n109, n81);
buf  g85 (n126, n73);
not  g86 (n93, n75);
not  g87 (n100, n80);
not  g88 (n146, n86);
not  g89 (n94, n87);
not  g90 (n113, n87);
buf  g91 (n132, n73);
not  g92 (n149, n78);
not  g93 (n137, n86);
not  g94 (n135, n84);
not  g95 (n127, n77);
not  g96 (n133, n80);
buf  g97 (n124, n78);
not  g98 (n131, n75);
buf  g99 (n115, n85);
not  g100 (n99, n87);
buf  g101 (n129, n74);
not  g102 (n107, n81);
buf  g103 (n114, n85);
buf  g104 (n110, n88);
not  g105 (n119, n74);
not  g106 (n98, n82);
buf  g107 (n108, n86);
not  g108 (n103, n79);
buf  g109 (n144, n88);
buf  g110 (n89, n80);
buf  g111 (n122, n82);
not  g112 (n125, n79);
buf  g113 (n143, n77);
not  g114 (n142, n83);
buf  g115 (n128, n74);
buf  g116 (n105, n81);
not  g117 (n120, n83);
not  g118 (n145, n77);
buf  g119 (n152, n73);
not  g120 (n134, n76);
buf  g121 (n90, n76);
buf  g122 (n106, n85);
buf  g123 (n141, n73);
buf  g124 (n112, n82);
not  g125 (n91, n85);
buf  g126 (n147, n74);
buf  g127 (n117, n78);
buf  g128 (n150, n78);
not  g129 (n96, n76);
not  g130 (n138, n83);
not  g131 (n148, n84);
buf  g132 (n363, n107);
not  g133 (n378, n106);
buf  g134 (n293, n133);
not  g135 (n219, n124);
not  g136 (n391, n100);
not  g137 (n181, n105);
not  g138 (n257, n103);
not  g139 (n227, n90);
not  g140 (n262, n146);
buf  g141 (n407, n98);
buf  g142 (n312, n127);
not  g143 (n264, n129);
not  g144 (n287, n117);
not  g145 (n197, n142);
buf  g146 (n153, n137);
not  g147 (n232, n103);
buf  g148 (n292, n113);
buf  g149 (n225, n133);
not  g150 (n216, n95);
buf  g151 (n268, n111);
buf  g152 (n375, n95);
not  g153 (n280, n98);
not  g154 (n234, n89);
not  g155 (n291, n95);
buf  g156 (n275, n98);
buf  g157 (n206, n114);
not  g158 (n175, n139);
not  g159 (n230, n125);
buf  g160 (n200, n101);
not  g161 (n254, n133);
buf  g162 (n303, n90);
buf  g163 (n408, n126);
buf  g164 (n324, n129);
buf  g165 (n172, n131);
buf  g166 (n241, n115);
not  g167 (n349, n151);
not  g168 (n272, n131);
buf  g169 (n315, n109);
not  g170 (n191, n109);
not  g171 (n156, n145);
buf  g172 (n309, n107);
buf  g173 (n158, n121);
not  g174 (n278, n130);
buf  g175 (n339, n102);
buf  g176 (n320, n93);
not  g177 (n251, n147);
not  g178 (n194, n100);
buf  g179 (n282, n107);
not  g180 (n304, n152);
not  g181 (n405, n108);
buf  g182 (n226, n119);
not  g183 (n166, n112);
buf  g184 (n169, n123);
not  g185 (n396, n106);
not  g186 (n160, n99);
not  g187 (n331, n101);
buf  g188 (n285, n135);
not  g189 (n178, n104);
buf  g190 (n371, n133);
buf  g191 (n299, n101);
buf  g192 (n192, n113);
not  g193 (n188, n94);
buf  g194 (n372, n93);
not  g195 (n177, n126);
buf  g196 (n246, n151);
not  g197 (n301, n148);
not  g198 (n247, n104);
buf  g199 (n328, n138);
not  g200 (n354, n150);
buf  g201 (n353, n97);
not  g202 (n267, n113);
buf  g203 (n343, n89);
not  g204 (n389, n121);
buf  g205 (n394, n139);
buf  g206 (n259, n114);
not  g207 (n332, n140);
buf  g208 (n316, n108);
buf  g209 (n388, n99);
buf  g210 (n215, n140);
buf  g211 (n159, n108);
not  g212 (n229, n96);
buf  g213 (n295, n110);
not  g214 (n239, n123);
not  g215 (n252, n103);
buf  g216 (n333, n114);
not  g217 (n163, n146);
buf  g218 (n189, n140);
not  g219 (n345, n146);
buf  g220 (n243, n122);
buf  g221 (n351, n110);
not  g222 (n390, n117);
not  g223 (n233, n104);
buf  g224 (n167, n142);
buf  g225 (n171, n149);
not  g226 (n196, n119);
not  g227 (n381, n89);
not  g228 (n360, n149);
not  g229 (n401, n103);
not  g230 (n183, n129);
buf  g231 (n176, n151);
buf  g232 (n179, n120);
not  g233 (n223, n110);
not  g234 (n366, n116);
buf  g235 (n224, n143);
not  g236 (n329, n111);
not  g237 (n297, n95);
not  g238 (n323, n117);
buf  g239 (n248, n97);
not  g240 (n350, n147);
not  g241 (n319, n147);
not  g242 (n213, n130);
not  g243 (n256, n131);
not  g244 (n348, n109);
buf  g245 (n164, n128);
not  g246 (n393, n116);
buf  g247 (n231, n115);
not  g248 (n209, n102);
buf  g249 (n325, n115);
buf  g250 (n255, n130);
not  g251 (n313, n126);
not  g252 (n369, n146);
buf  g253 (n168, n144);
buf  g254 (n218, n99);
not  g255 (n242, n152);
buf  g256 (n337, n144);
buf  g257 (n249, n137);
not  g258 (n161, n119);
not  g259 (n207, n105);
buf  g260 (n258, n118);
buf  g261 (n380, n91);
buf  g262 (n211, n134);
not  g263 (n279, n112);
buf  g264 (n187, n145);
buf  g265 (n203, n114);
buf  g266 (n346, n118);
not  g267 (n352, n92);
buf  g268 (n221, n121);
buf  g269 (n308, n93);
buf  g270 (n162, n132);
not  g271 (n347, n97);
not  g272 (n374, n94);
not  g273 (n261, n141);
not  g274 (n253, n125);
buf  g275 (n386, n134);
buf  g276 (n359, n130);
not  g277 (n170, n124);
buf  g278 (n190, n93);
not  g279 (n377, n126);
not  g280 (n318, n148);
buf  g281 (n327, n96);
buf  g282 (n289, n136);
buf  g283 (n344, n123);
buf  g284 (n382, n148);
not  g285 (n288, n92);
buf  g286 (n199, n96);
not  g287 (n306, n141);
buf  g288 (n311, n118);
buf  g289 (n155, n128);
not  g290 (n214, n92);
not  g291 (n245, n109);
buf  g292 (n269, n144);
buf  g293 (n307, n116);
buf  g294 (n404, n91);
not  g295 (n220, n134);
not  g296 (n342, n100);
buf  g297 (n367, n102);
buf  g298 (n321, n102);
buf  g299 (n370, n138);
not  g300 (n387, n125);
not  g301 (n173, n108);
buf  g302 (n357, n107);
buf  g303 (n198, n138);
buf  g304 (n195, n144);
buf  g305 (n338, n134);
buf  g306 (n202, n92);
not  g307 (n298, n111);
not  g308 (n368, n136);
not  g309 (n286, n121);
not  g310 (n326, n136);
not  g311 (n193, n101);
not  g312 (n385, n141);
buf  g313 (n228, n151);
buf  g314 (n277, n94);
buf  g315 (n317, n110);
not  g316 (n365, n116);
buf  g317 (n373, n127);
not  g318 (n263, n105);
buf  g319 (n398, n135);
not  g320 (n154, n131);
buf  g321 (n157, n137);
buf  g322 (n266, n90);
buf  g323 (n336, n124);
buf  g324 (n235, n142);
buf  g325 (n182, n120);
not  g326 (n204, n132);
buf  g327 (n201, n143);
not  g328 (n237, n119);
buf  g329 (n205, n135);
not  g330 (n395, n100);
buf  g331 (n270, n143);
not  g332 (n364, n140);
buf  g333 (n384, n122);
not  g334 (n184, n115);
buf  g335 (n244, n150);
not  g336 (n217, n128);
not  g337 (n302, n112);
buf  g338 (n402, n94);
buf  g339 (n208, n99);
buf  g340 (n362, n148);
not  g341 (n273, n139);
not  g342 (n334, n136);
buf  g343 (n281, n147);
buf  g344 (n271, n143);
not  g345 (n305, n90);
buf  g346 (n238, n111);
not  g347 (n403, n104);
not  g348 (n300, n129);
buf  g349 (n212, n113);
not  g350 (n356, n118);
buf  g351 (n180, n124);
not  g352 (n400, n135);
not  g353 (n361, n106);
not  g354 (n210, n106);
not  g355 (n379, n128);
buf  g356 (n296, n96);
not  g357 (n335, n145);
buf  g358 (n274, n105);
buf  g359 (n236, n132);
not  g360 (n406, n120);
buf  g361 (n165, n137);
buf  g362 (n376, n91);
buf  g363 (n283, n120);
buf  g364 (n222, n97);
buf  g365 (n186, n149);
not  g366 (n265, n145);
buf  g367 (n310, n149);
buf  g368 (n250, n150);
buf  g369 (n341, n139);
buf  g370 (n314, n150);
buf  g371 (n399, n141);
not  g372 (n294, n112);
not  g373 (n397, n142);
not  g374 (n174, n152);
buf  g375 (n355, n91);
not  g376 (n290, n98);
not  g377 (n383, n122);
buf  g378 (n392, n138);
buf  g379 (n260, n125);
buf  g380 (n240, n117);
not  g381 (n185, n127);
buf  g382 (n358, n89);
buf  g383 (n276, n132);
not  g384 (n340, n123);
not  g385 (n330, n122);
not  g386 (n284, n127);
not  g387 (n322, n152);
buf  g388 (n525, n303);
not  g389 (n608, n158);
buf  g390 (n645, n298);
buf  g391 (n764, n258);
not  g392 (n524, n296);
buf  g393 (n651, n301);
not  g394 (n708, n344);
buf  g395 (n478, n321);
not  g396 (n567, n382);
buf  g397 (n595, n209);
not  g398 (n670, n181);
not  g399 (n769, n155);
buf  g400 (n863, n272);
buf  g401 (n600, n325);
buf  g402 (n606, n335);
buf  g403 (n793, n332);
not  g404 (n804, n201);
buf  g405 (n466, n224);
not  g406 (n726, n209);
buf  g407 (n579, n153);
not  g408 (n449, n358);
not  g409 (n687, n371);
buf  g410 (n720, n198);
buf  g411 (n429, n265);
buf  g412 (n508, n305);
buf  g413 (n551, n312);
buf  g414 (n701, n220);
buf  g415 (n689, n159);
buf  g416 (n656, n183);
not  g417 (n775, n215);
not  g418 (n534, n325);
buf  g419 (n628, n333);
not  g420 (n712, n261);
buf  g421 (n597, n298);
not  g422 (n441, n246);
buf  g423 (n660, n168);
not  g424 (n735, n369);
not  g425 (n667, n165);
buf  g426 (n554, n224);
buf  g427 (n640, n311);
not  g428 (n682, n295);
buf  g429 (n706, n160);
not  g430 (n635, n197);
buf  g431 (n768, n247);
buf  g432 (n621, n178);
not  g433 (n455, n185);
buf  g434 (n728, n191);
buf  g435 (n851, n196);
buf  g436 (n632, n254);
buf  g437 (n605, n274);
not  g438 (n853, n369);
not  g439 (n770, n377);
buf  g440 (n634, n324);
not  g441 (n734, n328);
not  g442 (n432, n321);
not  g443 (n812, n335);
buf  g444 (n574, n219);
buf  g445 (n655, n203);
not  g446 (n420, n206);
buf  g447 (n710, n308);
buf  g448 (n813, n258);
not  g449 (n631, n281);
not  g450 (n531, n270);
buf  g451 (n564, n291);
not  g452 (n657, n277);
buf  g453 (n841, n169);
not  g454 (n518, n356);
not  g455 (n474, n242);
buf  g456 (n443, n255);
buf  g457 (n861, n189);
buf  g458 (n497, n296);
buf  g459 (n529, n208);
not  g460 (n457, n341);
not  g461 (n566, n292);
buf  g462 (n596, n230);
not  g463 (n544, n161);
buf  g464 (n521, n282);
not  g465 (n583, n311);
buf  g466 (n830, n235);
not  g467 (n479, n176);
not  g468 (n470, n319);
not  g469 (n649, n313);
buf  g470 (n550, n317);
buf  g471 (n724, n381);
buf  g472 (n498, n320);
buf  g473 (n753, n286);
not  g474 (n797, n189);
buf  g475 (n654, n238);
buf  g476 (n584, n183);
not  g477 (n523, n257);
not  g478 (n811, n293);
not  g479 (n481, n226);
not  g480 (n762, n249);
buf  g481 (n836, n188);
not  g482 (n504, n348);
buf  g483 (n425, n300);
buf  g484 (n555, n193);
not  g485 (n718, n323);
buf  g486 (n743, n320);
buf  g487 (n448, n285);
not  g488 (n843, n161);
not  g489 (n738, n230);
buf  g490 (n615, n277);
not  g491 (n527, n267);
not  g492 (n757, n207);
not  g493 (n549, n228);
not  g494 (n677, n364);
not  g495 (n451, n297);
not  g496 (n696, n275);
not  g497 (n717, n238);
buf  g498 (n761, n302);
not  g499 (n664, n200);
buf  g500 (n759, n171);
not  g501 (n548, n276);
buf  g502 (n642, n186);
not  g503 (n599, n169);
buf  g504 (n417, n165);
buf  g505 (n580, n309);
not  g506 (n705, n376);
not  g507 (n781, n156);
not  g508 (n590, n359);
not  g509 (n674, n246);
buf  g510 (n601, n207);
not  g511 (n739, n237);
not  g512 (n730, n319);
buf  g513 (n460, n170);
not  g514 (n570, n175);
buf  g515 (n581, n383);
buf  g516 (n828, n194);
not  g517 (n777, n231);
not  g518 (n623, n281);
not  g519 (n754, n361);
not  g520 (n752, n247);
not  g521 (n442, n366);
not  g522 (n607, n287);
buf  g523 (n446, n281);
buf  g524 (n681, n316);
buf  g525 (n780, n238);
not  g526 (n428, n195);
not  g527 (n507, n251);
buf  g528 (n736, n371);
buf  g529 (n435, n300);
buf  g530 (n644, n177);
not  g531 (n773, n214);
buf  g532 (n639, n383);
buf  g533 (n465, n180);
not  g534 (n411, n261);
buf  g535 (n447, n190);
not  g536 (n509, n299);
buf  g537 (n473, n193);
not  g538 (n622, n290);
not  g539 (n445, n322);
not  g540 (n800, n367);
not  g541 (n790, n337);
not  g542 (n782, n320);
buf  g543 (n665, n189);
buf  g544 (n758, n353);
buf  g545 (n823, n355);
buf  g546 (n543, n285);
buf  g547 (n522, n259);
buf  g548 (n412, n269);
not  g549 (n589, n185);
buf  g550 (n496, n296);
buf  g551 (n568, n341);
buf  g552 (n732, n376);
buf  g553 (n819, n374);
not  g554 (n515, n351);
buf  g555 (n467, n271);
buf  g556 (n462, n252);
not  g557 (n704, n275);
not  g558 (n697, n381);
buf  g559 (n791, n239);
buf  g560 (n535, n204);
not  g561 (n629, n198);
not  g562 (n666, n182);
not  g563 (n808, n249);
buf  g564 (n532, n232);
not  g565 (n715, n377);
not  g566 (n783, n329);
not  g567 (n627, n338);
not  g568 (n516, n166);
not  g569 (n835, n360);
not  g570 (n845, n382);
not  g571 (n494, n299);
buf  g572 (n848, n349);
buf  g573 (n713, n305);
not  g574 (n691, n328);
buf  g575 (n868, n256);
not  g576 (n472, n208);
buf  g577 (n703, n311);
not  g578 (n831, n182);
not  g579 (n611, n249);
not  g580 (n821, n218);
not  g581 (n740, n350);
buf  g582 (n533, n365);
buf  g583 (n434, n302);
buf  g584 (n476, n349);
buf  g585 (n513, n369);
not  g586 (n727, n341);
not  g587 (n433, n211);
buf  g588 (n716, n321);
buf  g589 (n413, n175);
buf  g590 (n771, n375);
not  g591 (n569, n253);
not  g592 (n636, n314);
buf  g593 (n785, n355);
buf  g594 (n858, n352);
buf  g595 (n490, n242);
not  g596 (n698, n346);
not  g597 (n850, n164);
not  g598 (n721, n327);
buf  g599 (n860, n285);
buf  g600 (n461, n217);
not  g601 (n862, n237);
not  g602 (n495, n350);
not  g603 (n440, n241);
not  g604 (n719, n322);
buf  g605 (n668, n186);
buf  g606 (n854, n370);
not  g607 (n573, n234);
buf  g608 (n816, n178);
not  g609 (n849, n207);
not  g610 (n626, n337);
buf  g611 (n675, n174);
buf  g612 (n801, n373);
buf  g613 (n633, n339);
not  g614 (n475, n353);
not  g615 (n514, n168);
not  g616 (n709, n378);
buf  g617 (n690, n267);
not  g618 (n563, n223);
buf  g619 (n603, n343);
buf  g620 (n744, n286);
not  g621 (n653, n305);
buf  g622 (n419, n339);
buf  g623 (n766, n272);
buf  g624 (n820, n354);
not  g625 (n686, n329);
buf  g626 (n788, n216);
buf  g627 (n410, n181);
buf  g628 (n829, n255);
buf  g629 (n598, n357);
buf  g630 (n827, n351);
not  g631 (n431, n222);
buf  g632 (n520, n211);
buf  g633 (n663, n336);
buf  g634 (n612, n273);
not  g635 (n439, n273);
not  g636 (n810, n227);
not  g637 (n814, n321);
not  g638 (n505, n170);
buf  g639 (n729, n266);
buf  g640 (n484, n163);
buf  g641 (n616, n293);
buf  g642 (n685, n342);
buf  g643 (n444, n196);
not  g644 (n426, n325);
not  g645 (n561, n158);
not  g646 (n693, n232);
buf  g647 (n585, n280);
buf  g648 (n414, n217);
buf  g649 (n671, n240);
not  g650 (n463, n352);
not  g651 (n625, n222);
not  g652 (n702, n252);
buf  g653 (n844, n179);
not  g654 (n486, n181);
not  g655 (n593, n198);
buf  g656 (n565, n226);
buf  g657 (n415, n192);
not  g658 (n792, n234);
buf  g659 (n855, n251);
not  g660 (n669, n214);
not  g661 (n409, n245);
not  g662 (n838, n301);
not  g663 (n760, n194);
buf  g664 (n511, n286);
buf  g665 (n604, n371);
not  g666 (n798, n342);
not  g667 (n436, n261);
not  g668 (n711, n304);
not  g669 (n803, n268);
buf  g670 (n547, n195);
buf  g671 (n765, n318);
buf  g672 (n650, n357);
buf  g673 (n648, n255);
buf  g674 (n748, n378);
not  g675 (n834, n292);
buf  g676 (n530, n265);
buf  g677 (n679, n288);
not  g678 (n491, n285);
not  g679 (n742, n164);
buf  g680 (n528, n220);
buf  g681 (n503, n233);
not  g682 (n613, n313);
buf  g683 (n556, n367);
buf  g684 (n506, n249);
not  g685 (n469, n326);
buf  g686 (n501, n312);
not  g687 (n763, n348);
buf  g688 (n587, n372);
buf  g689 (n733, n209);
not  g690 (n707, n329);
nand g691 (n847, n192, n173, n299, n252);
xor  g692 (n746, n305, n259, n287, n334);
xnor g693 (n624, n209, n232, n334, n205);
nor  g694 (n438, n365, n361, n366, n295);
xor  g695 (n856, n203, n268, n309, n343);
or   g696 (n416, n326, n256, n289, n294);
nand g697 (n558, n253, n212, n258, n363);
and  g698 (n794, n172, n205, n163, n347);
and  g699 (n807, n366, n203, n303, n352);
nand g700 (n646, n373, n368, n220, n173);
xnor g701 (n576, n166, n158, n309, n159);
and  g702 (n714, n244, n184, n383, n247);
nor  g703 (n582, n360, n171, n371);
xor  g704 (n480, n243, n154, n190, n341);
xor  g705 (n661, n179, n161, n172, n257);
and  g706 (n817, n317, n155, n260, n225);
or   g707 (n865, n282, n372, n344, n363);
xor  g708 (n609, n354, n235, n368, n231);
xnor g709 (n619, n274, n345, n180, n292);
or   g710 (n591, n293, n375, n304, n263);
nand g711 (n500, n337, n230, n236, n192);
nor  g712 (n471, n244, n376, n368, n197);
xnor g713 (n418, n180, n270, n343, n306);
nor  g714 (n539, n166, n190, n294, n282);
nand g715 (n699, n298, n284, n178, n233);
or   g716 (n552, n307, n284, n289, n260);
xor  g717 (n477, n252, n342, n333, n177);
xnor g718 (n557, n378, n161, n353, n291);
nand g719 (n560, n329, n277, n229, n362);
nand g720 (n731, n279, n162, n345, n336);
or   g721 (n617, n200, n159, n273, n356);
xor  g722 (n741, n376, n303, n202, n193);
and  g723 (n837, n266, n214, n301, n176);
xnor g724 (n662, n322, n157, n362, n280);
nand g725 (n786, n298, n345, n170, n168);
nor  g726 (n450, n157, n340, n175, n262);
xnor g727 (n423, n241, n380, n246, n236);
nand g728 (n519, n202, n204, n175, n372);
and  g729 (n795, n160, n304, n224, n356);
and  g730 (n747, n334, n251, n220, n309);
nor  g731 (n852, n153, n297, n348, n234);
or   g732 (n859, n255, n296, n294, n283);
nor  g733 (n542, n312, n273, n269, n370);
or   g734 (n620, n184, n278, n239, n287);
xor  g735 (n592, n362, n236, n187, n323);
xor  g736 (n774, n333, n336, n358, n271);
nor  g737 (n421, n370, n275, n384, n172);
xor  g738 (n424, n262, n183, n380, n228);
and  g739 (n572, n356, n340, n155, n283);
xnor g740 (n637, n354, n327, n316, n266);
nor  g741 (n453, n225, n233, n218, n240);
nand g742 (n846, n384, n187, n267, n237);
nor  g743 (n692, n269, n314, n217, n228);
and  g744 (n614, n287, n290, n211, n174);
and  g745 (n430, n317, n300, n274, n257);
and  g746 (n652, n154, n295, n203, n223);
xor  g747 (n559, n325, n335, n385, n239);
and  g748 (n586, n346, n163, n208, n326);
or   g749 (n772, n205, n330, n372, n263);
or   g750 (n594, n167, n171, n250, n254);
xor  g751 (n684, n377, n331, n153, n158);
nand g752 (n799, n253, n210, n242, n165);
and  g753 (n749, n313, n290, n324, n253);
nor  g754 (n575, n170, n278, n324, n229);
nor  g755 (n537, n188, n278, n165, n202);
xnor g756 (n683, n355, n206, n385, n369);
and  g757 (n482, n227, n258, n174, n320);
nand g758 (n456, n272, n382, n340, n364);
nor  g759 (n641, n223, n350, n221, n367);
nor  g760 (n737, n315, n283, n306, n223);
xnor g761 (n695, n266, n229, n308, n339);
nor  g762 (n458, n373, n207, n187, n182);
xnor g763 (n751, n184, n169, n172, n347);
xnor g764 (n673, n381, n196, n359, n338);
or   g765 (n776, n206, n244, n297, n199);
xor  g766 (n643, n202, n316, n283, n242);
and  g767 (n745, n195, n234, n355, n357);
xor  g768 (n755, n327, n289, n354, n264);
nor  g769 (n545, n270, n201, n328, n237);
and  g770 (n540, n167, n183, n228, n240);
nor  g771 (n756, n310, n156, n385, n339);
xnor g772 (n502, n315, n199, n162, n224);
nor  g773 (n825, n210, n335, n180, n154);
xnor g774 (n802, n238, n312, n222, n247);
or   g775 (n489, n254, n204, n348, n259);
xor  g776 (n767, n260, n375, n221, n251);
nand g777 (n676, n212, n338, n384, n310);
and  g778 (n842, n248, n248, n278, n179);
nand g779 (n678, n324, n381, n166, n290);
nand g780 (n680, n153, n213, n186, n212);
xnor g781 (n840, n215, n188, n182, n241);
nor  g782 (n536, n245, n360, n367, n232);
and  g783 (n658, n276, n306, n268, n257);
xnor g784 (n546, n289, n268, n322, n357);
nor  g785 (n722, n306, n365, n340, n279);
or   g786 (n778, n307, n245, n374, n155);
nor  g787 (n672, n297, n331, n374, n186);
xnor g788 (n541, n157, n215, n177, n213);
or   g789 (n725, n157, n279, n292, n344);
nand g790 (n839, n334, n383, n250, n302);
or   g791 (n796, n318, n200, n256, n194);
or   g792 (n610, n314, n353, n248, n291);
nand g793 (n805, n198, n256, n303, n264);
xor  g794 (n789, n184, n178, n230, n374);
and  g795 (n809, n222, n227, n188, n214);
or   g796 (n468, n279, n363, n194, n302);
xnor g797 (n452, n187, n219, n338, n301);
xnor g798 (n487, n179, n288, n167, n262);
nor  g799 (n857, n375, n264, n177, n208);
or   g800 (n806, n277, n346, n216, n250);
and  g801 (n824, n377, n201, n337, n364);
xor  g802 (n826, n358, n307, n164, n216);
xnor g803 (n577, n318, n293, n196, n362);
nor  g804 (n499, n210, n271, n254, n310);
and  g805 (n818, n211, n352, n244, n344);
nor  g806 (n517, n330, n239, n304, n332);
nand g807 (n700, n311, n176, n317, n160);
and  g808 (n833, n260, n243, n176, n313);
and  g809 (n694, n332, n380, n314, n229);
and  g810 (n485, n225, n379, n360, n274);
xnor g811 (n483, n235, n212, n272, n199);
xnor g812 (n459, n349, n181, n307, n330);
nand g813 (n867, n225, n327, n219, n351);
xnor g814 (n630, n378, n323, n231, n347);
nor  g815 (n815, n246, n382, n333, n288);
nand g816 (n562, n261, n156, n345, n219);
or   g817 (n538, n169, n190, n363, n245);
and  g818 (n659, n280, n384, n213, n275);
or   g819 (n427, n280, n379, n351, n276);
or   g820 (n864, n271, n295, n217, n343);
xor  g821 (n750, n191, n213, n288, n195);
xor  g822 (n784, n159, n226, n233, n264);
and  g823 (n464, n262, n365, n250, n197);
nor  g824 (n638, n294, n284, n197, n160);
xnor g825 (n787, n361, n221, n346, n248);
nor  g826 (n422, n206, n358, n240, n270);
xnor g827 (n454, n379, n235, n241, n173);
xnor g828 (n588, n336, n163, n259, n319);
xor  g829 (n618, n276, n359, n286, n221);
xnor g830 (n822, n349, n193, n189, n373);
and  g831 (n493, n215, n263, n174, n330);
and  g832 (n553, n361, n300, n366, n204);
nand g833 (n510, n218, n318, n299, n319);
or   g834 (n647, n162, n359, n173, n205);
or   g835 (n866, n370, n192, n281, n231);
and  g836 (n832, n380, n331, n326, n284);
nor  g837 (n492, n315, n342, n243);
xor  g838 (n779, n368, n210, n328, n263);
xnor g839 (n512, n364, n350, n218, n282);
nand g840 (n578, n310, n185, n267, n226);
xnor g841 (n488, n308, n236, n162, n227);
xor  g842 (n526, n316, n379, n216, n199);
or   g843 (n571, n191, n168, n265, n315);
xnor g844 (n688, n265, n332, n185, n164);
or   g845 (n602, n191, n154, n323, n156);
and  g846 (n723, n200, n201, n347, n308);
and  g847 (n437, n291, n167, n269, n331);
buf  g848 (n874, n409);
buf  g849 (n870, n427);
xor  g850 (n877, n416, n432, n419, n437);
nand g851 (n872, n412, n413, n429, n424);
xor  g852 (n875, n417, n431, n425, n414);
nand g853 (n869, n435, n438, n428, n420);
xor  g854 (n873, n433, n418, n430, n423);
or   g855 (n871, n426, n434, n410, n411);
xor  g856 (n876, n422, n421, n415, n436);
xnor g857 (n883, n869, n459, n467, n458);
and  g858 (n884, n870, n461, n455, n439);
nand g859 (n885, n460, n877, n444, n448);
nor  g860 (n879, n876, n466, n446, n443);
and  g861 (n878, n440, n449, n871, n451);
nor  g862 (n880, n872, n874, n877, n457);
nor  g863 (n882, n450, n442, n456, n462);
and  g864 (n886, n875, n873, n463, n454);
and  g865 (n881, n464, n445, n452, n447);
and  g866 (n887, n465, n441, n468, n453);
not  g867 (n888, n879);
buf  g868 (n893, n469);
buf  g869 (n889, n470);
buf  g870 (n890, n878);
nand g871 (n891, n472, n878);
and  g872 (n892, n471, n879, n878);
not  g873 (n895, n888);
buf  g874 (n897, n888);
buf  g875 (n894, n888);
not  g876 (n896, n888);
not  g877 (n898, n889);
nor  g878 (n900, n474, n895, n894);
xnor g879 (n899, n475, n476, n473);
or   g880 (n902, n880, n882, n900, n477);
and  g881 (n905, n879, n881, n880);
or   g882 (n904, n879, n900, n882, n899);
or   g883 (n903, n882, n880, n881, n900);
xnor g884 (n901, n900, n881, n882);
not  g885 (n908, n903);
buf  g886 (n909, n901);
not  g887 (n906, n903);
buf  g888 (n912, n901);
not  g889 (n907, n901);
buf  g890 (n911, n902);
not  g891 (n913, n902);
not  g892 (n910, n902);
not  g893 (n917, n908);
not  g894 (n916, n909);
buf  g895 (n914, n907);
buf  g896 (n915, n906);
buf  g897 (n918, n917);
buf  g898 (n930, n478);
not  g899 (n919, n914);
not  g900 (n929, n914);
not  g901 (n923, n896);
buf  g902 (n927, n897);
not  g903 (n920, n917);
buf  g904 (n921, n480);
not  g905 (n928, n916);
buf  g906 (n926, n915);
not  g907 (n925, n916);
not  g908 (n931, n914);
xor  g909 (n932, n481, n479);
xnor g910 (n924, n915, n914, n482, n917);
or   g911 (n922, n915, n916);
not  g912 (n941, n408);
buf  g913 (n946, n391);
buf  g914 (n974, n399);
not  g915 (n964, n393);
not  g916 (n991, n395);
not  g917 (n981, n928);
buf  g918 (n960, n927);
not  g919 (n953, n926);
buf  g920 (n985, n396);
buf  g921 (n956, n406);
not  g922 (n984, n921);
buf  g923 (n943, n406);
buf  g924 (n967, n400);
not  g925 (n935, n394);
not  g926 (n954, n408);
not  g927 (n972, n395);
not  g928 (n979, n925);
buf  g929 (n950, n932);
buf  g930 (n934, n407);
buf  g931 (n947, n920);
buf  g932 (n978, n386);
not  g933 (n949, n929);
nor  g934 (n970, n393, n391);
xor  g935 (n973, n387, n406, n403, n407);
xor  g936 (n977, n925, n931, n919, n390);
xor  g937 (n989, n388, n921, n399, n394);
xnor g938 (n976, n390, n923, n925, n396);
nand g939 (n966, n407, n930, n386, n408);
xor  g940 (n962, n386, n403, n398, n922);
xnor g941 (n942, n404, n485, n918, n923);
xnor g942 (n968, n405, n911, n926, n391);
xor  g943 (n990, n483, n407, n922, n931);
nand g944 (n965, n929, n402, n927, n398);
xnor g945 (n982, n932, n921, n924, n926);
and  g946 (n948, n395, n390, n401, n392);
and  g947 (n959, n400, n905, n904, n388);
and  g948 (n958, n389, n389, n928, n405);
or   g949 (n961, n904, n918, n392, n927);
nand g950 (n980, n917, n486, n388, n393);
and  g951 (n971, n488, n919, n397, n399);
or   g952 (n986, n930, n388, n387, n401);
and  g953 (n936, n397, n402, n398, n924);
nor  g954 (n944, n920, n904, n385, n924);
nor  g955 (n957, n389, n903, n919, n931);
or   g956 (n983, n930, n404, n932, n400);
xnor g957 (n939, n905, n387, n928, n912);
xor  g958 (n938, n921, n394, n392);
xnor g959 (n992, n404, n390, n401, n930);
xor  g960 (n945, n905, n403, n918, n922);
nor  g961 (n937, n927, n402, n931, n405);
or   g962 (n933, n925, n398, n402, n920);
xnor g963 (n963, n923, n386, n397, n919);
and  g964 (n969, n401, n397, n389, n920);
nand g965 (n952, n924, n406, n484, n913);
xor  g966 (n955, n387, n400, n923, n393);
nor  g967 (n987, n396, n926, n487, n922);
xnor g968 (n951, n918, n928, n932, n391);
xor  g969 (n988, n404, n408, n910, n405);
xor  g970 (n975, n905, n396, n392, n403);
nor  g971 (n940, n399, n395, n929);
buf  g972 (n997, n935);
not  g973 (n1001, n938);
not  g974 (n1002, n942);
not  g975 (n995, n934);
not  g976 (n993, n493);
buf  g977 (n996, n936);
buf  g978 (n998, n489);
buf  g979 (n999, n940);
nand g980 (n1000, n937, n490, n939);
xor  g981 (n994, n492, n941, n491, n933);
xor  g982 (n1016, n1001, n1002, n993);
nor  g983 (n1011, n962, n948, n946, n950);
nand g984 (n1007, n949, n973, n961, n965);
nand g985 (n1003, n978, n495, n1000, n975);
xnor g986 (n1013, n959, n971, n947, n997);
xnor g987 (n1015, n945, n952, n994, n951);
nor  g988 (n1010, n975, n963, n943, n976);
xnor g989 (n1004, n966, n977, n964, n974);
nor  g990 (n1005, n958, n494, n976, n999);
nand g991 (n1012, n977, n970, n998, n954);
nand g992 (n1018, n976, n978, n974);
xnor g993 (n1006, n956, n955, n972, n957);
xnor g994 (n1017, n996, n953, n1000, n1001);
or   g995 (n1014, n969, n968, n1001, n974);
nand g996 (n1009, n995, n944, n967, n1002);
nand g997 (n1008, n1000, n975, n960, n977);
nand g998 (n1019, n498, n980, n501, n883);
xnor g999 (n1025, n979, n1006, n883, n884);
or   g1000 (n1020, n980, n979, n496);
nor  g1001 (n1024, n1003, n980, n1004, n503);
nor  g1002 (n1026, n981, n1009);
nand g1003 (n1021, n1005, n1007, n883, n884);
nand g1004 (n1022, n500, n1008, n499, n883);
and  g1005 (n1023, n497, n981, n502, n504);
buf  g1006 (n1032, n1022);
buf  g1007 (n1027, n1020);
buf  g1008 (n1033, n1021);
buf  g1009 (n1031, n505);
buf  g1010 (n1029, n1024);
buf  g1011 (n1028, n1019);
xnor g1012 (n1030, n1023, n1025);
and  g1013 (n1035, n1027, n511, n508, n506);
xor  g1014 (n1034, n1027, n509, n507, n510);
buf  g1015 (n1040, n1035);
not  g1016 (n1038, n1035);
buf  g1017 (n1039, n1034);
not  g1018 (n1036, n1035);
buf  g1019 (n1037, n1034);
not  g1020 (n1043, n1037);
buf  g1021 (n1044, n1036);
buf  g1022 (n1041, n512);
or   g1023 (n1042, n1039, n1038);
not  g1024 (n1047, n1042);
buf  g1025 (n1048, n1044);
not  g1026 (n1049, n1044);
buf  g1027 (n1045, n1043);
buf  g1028 (n1046, n1041);
not  g1029 (n1063, n531);
not  g1030 (n1050, n521);
not  g1031 (n1060, n1047);
buf  g1032 (n1065, n530);
not  g1033 (n1056, n1049);
buf  g1034 (n1068, n1048);
not  g1035 (n1062, n528);
buf  g1036 (n1064, n520);
buf  g1037 (n1059, n1046);
buf  g1038 (n1058, n519);
not  g1039 (n1052, n1048);
buf  g1040 (n1057, n514);
or   g1041 (n1061, n1046, n1045);
or   g1042 (n1054, n516, n517, n1047, n1048);
xnor g1043 (n1067, n518, n1045, n1049);
nor  g1044 (n1066, n522, n515, n525, n529);
xor  g1045 (n1053, n1045, n1049, n524, n513);
nand g1046 (n1055, n527, n1046, n1047, n526);
or   g1047 (n1051, n523, n1046, n1048, n1047);
not  g1048 (n1072, n1053);
not  g1049 (n1074, n1054);
buf  g1050 (n1073, n1056);
not  g1051 (n1075, n1055);
not  g1052 (n1069, n1050);
buf  g1053 (n1070, n1052);
buf  g1054 (n1071, n1051);
not  g1055 (n1077, n1069);
buf  g1056 (n1076, n1070);
xor  g1057 (n1081, n532, n535, n537, n539);
nor  g1058 (n1080, n541, n1077, n542, n534);
and  g1059 (n1079, n538, n1076, n540, n533);
xor  g1060 (n1078, n536, n1077, n543);
not  g1061 (n1083, n1061);
or   g1062 (n1082, n1059, n1057, n1060, n1061);
or   g1063 (n1084, n1079, n1078, n1080, n1058);
xor  g1064 (n1086, n1063, n1062);
or   g1065 (n1085, n1082, n884, n1083);
xor  g1066 (n1087, n546, n545, n544, n1086);
or   g1067 (n1089, n898, n897);
xnor g1068 (n1088, n1087, n898);
nand g1069 (n1091, n548, n1010, n1081, n547);
or   g1070 (n1090, n1009, n1089, n1010, n1088);
not  g1071 (n1092, n1090);
not  g1072 (n1093, n890);
or   g1073 (n1096, n1091, n889, n983);
nand g1074 (n1097, n1090, n982, n1084);
nand g1075 (n1095, n1091, n1044, n889);
or   g1076 (n1094, n982, n1010, n889, n1091);
nand g1077 (n1098, n1091, n1087, n982, n1090);
xor  g1078 (n1106, n985, n989, n988, n987);
nor  g1079 (n1099, n984, n983, n1095, n1093);
nand g1080 (n1101, n990, n986, n987);
xnor g1081 (n1103, n1097, n990, n985, n988);
and  g1082 (n1104, n1097, n984, n1094, n985);
nand g1083 (n1100, n984, n987, n990, n983);
and  g1084 (n1105, n989, n991, n986, n1096);
or   g1085 (n1102, n989, n1097, n1092, n988);
xnor g1086 (n1107, n1103, n1065, n991);
xor  g1087 (n1109, n1063, n1067, n1102, n992);
xnor g1088 (n1110, n1099, n1104, n1066, n1067);
or   g1089 (n1111, n992, n1064, n1101, n1100);
nor  g1090 (n1113, n992, n1067, n1064);
xor  g1091 (n1112, n1066, n1066, n1065, n1063);
or   g1092 (n1108, n1066, n991, n1067, n1105);
xnor g1093 (n1117, n1012, n1013, n1040, n1109);
nand g1094 (n1118, n1072, n1110, n1071, n1012);
xnor g1095 (n1115, n1108, n1012, n1014, n1013);
and  g1096 (n1116, n1013, n1014, n1011);
xor  g1097 (n1114, n1107, n1111, n1011);
nand g1098 (n1119, n549, n558, n554, n556);
or   g1099 (n1121, n1115, n553, n555, n560);
nor  g1100 (n1120, n551, n1116, n1114, n1117);
or   g1101 (n1122, n550, n559, n557, n552);
buf  g1102 (n1123, n1068);
or   g1103 (n1125, n1113, n1112, n1106, n1122);
nor  g1104 (n1124, n1098, n1121, n1119, n1118);
nand g1105 (n1126, n1098, n1098, n1049, n1120);
buf  g1106 (n1129, n1123);
not  g1107 (n1127, n1123);
buf  g1108 (n1128, n1123);
nor  g1109 (n1132, n575, n571, n1129, n570);
nor  g1110 (n1133, n561, n1129, n569, n562);
xor  g1111 (n1131, n563, n572, n573, n568);
nand g1112 (n1134, n1128, n567, n1127, n1129);
and  g1113 (n1130, n574, n566, n565, n564);
buf  g1114 (n1136, n1124);
not  g1115 (n1135, n1131);
not  g1116 (n1139, n1130);
not  g1117 (n1137, n1133);
xnor g1118 (n1138, n1132, n1134);
and  g1119 (n1141, n1124, n1125);
nand g1120 (n1140, n1124, n1136, n1135, n1125);
not  g1121 (n1142, n1141);
not  g1122 (n1143, n1140);
not  g1123 (n1145, n1142);
buf  g1124 (n1149, n1143);
not  g1125 (n1148, n578);
buf  g1126 (n1147, n1143);
not  g1127 (n1150, n577);
not  g1128 (n1144, n1142);
and  g1129 (n1146, n576, n1142, n1143);
xor  g1130 (n1151, n586, n580, n589, n587);
and  g1131 (n1154, n591, n582, n595, n1144);
xnor g1132 (n1153, n585, n596, n1145, n579);
xor  g1133 (n1152, n1145, n1144, n590);
or   g1134 (n1155, n588, n583, n581, n592);
xor  g1135 (n1156, n584, n593, n1144, n594);
buf  g1136 (n1159, n597);
not  g1137 (n1157, n1153);
buf  g1138 (n1158, n1154);
nand g1139 (n1160, n1152, n1155);
xnor g1140 (n1162, n886, n887, n885);
nand g1141 (n1163, n886, n887, n885, n1157);
nor  g1142 (n1161, n1160, n885, n1158);
xnor g1143 (n1164, n887, n1159, n886);
nor  g1144 (n1175, n611, n604, n1147, n612);
xor  g1145 (n1169, n1147, n1161, n891, n605);
xor  g1146 (n1178, n1162, n892, n1147, n1148);
and  g1147 (n1165, n890, n890, n1146, n615);
and  g1148 (n1171, n613, n891, n1164);
xnor g1149 (n1170, n606, n609, n890, n610);
xor  g1150 (n1180, n599, n607, n614, n1161);
xnor g1151 (n1168, n1164, n1146, n1163);
and  g1152 (n1173, n1162, n608, n603, n1149);
or   g1153 (n1177, n892, n1164, n1162, n1148);
xor  g1154 (n1174, n892, n1148, n1161, n1147);
xnor g1155 (n1166, n1164, n1163, n1145);
xnor g1156 (n1179, n601, n1145, n891, n1148);
and  g1157 (n1176, n598, n1161, n602, n892);
or   g1158 (n1172, n600, n1162, n893);
xnor g1159 (n1167, n1146, n893, n1163);
nor  g1160 (n1181, n1172, n630, n637, n1149);
nand g1161 (n1184, n632, n1173, n1149, n633);
and  g1162 (n1182, n1165, n1168, n620, n1170);
xnor g1163 (n1189, n629, n619, n617, n1169);
xnor g1164 (n1190, n641, n638, n640, n642);
xnor g1165 (n1183, n1175, n1149, n1174, n626);
xnor g1166 (n1191, n623, n639, n644, n635);
and  g1167 (n1186, n628, n1167, n634, n1150);
nand g1168 (n1188, n621, n622, n643, n616);
or   g1169 (n1187, n625, n627, n1171, n636);
and  g1170 (n1185, n618, n631, n624, n1166);
nand g1171 (n1193, n1178, n1179, n1156, n1176);
xor  g1172 (n1195, n1177, n1075, n1180);
or   g1173 (n1194, n1188, n1074, n1189, n1191);
or   g1174 (n1192, n1190, n1180, n1073);
buf  g1175 (n1196, n1193);
buf  g1176 (n1197, n1192);
xnor g1177 (n1200, n651, n654, n646, n647);
xnor g1178 (n1198, n649, n650, n1193, n1196);
nor  g1179 (n1199, n1138, n652, n656, n1196);
and  g1180 (n1203, n1196, n1138, n655);
or   g1181 (n1201, n1139, n1139, n653, n1196);
xor  g1182 (n1205, n648, n645, n1197);
or   g1183 (n1204, n1139, n1139, n1137, n1194);
xor  g1184 (n1202, n1197, n1137);
nor  g1185 (n1206, n1198, n657, n1126, n658);
nor  g1186 (n1208, n1199, n1195, n1206);
xnor g1187 (n1207, n1194, n1194, n1195, n1206);
not  g1188 (n1209, n1208);
not  g1189 (n1211, n1209);
buf  g1190 (n1210, n1209);
nor  g1191 (n1214, n1204, n1017, n1015);
nand g1192 (n1216, n1203, n1016, n1210);
or   g1193 (n1213, n1018, n1211, n1017);
nand g1194 (n1215, n1201, n1200, n1018, n1016);
and  g1195 (n1218, n1211, n1016, n1205, n1015);
nor  g1196 (n1212, n1211, n1202, n1210, n1018);
nor  g1197 (n1217, n1211, n1018, n1015, n1016);
nand g1198 (n1235, n726, n668, n684, n660);
nand g1199 (n1230, n678, n733, n719, n718);
nor  g1200 (n1219, n725, n723, n679, n662);
nor  g1201 (n1233, n691, n1216, n710, n698);
xor  g1202 (n1239, n674, n1214, n1215, n671);
nand g1203 (n1223, n666, n721, n664, n1212);
or   g1204 (n1245, n659, n1216, n1213, n734);
xor  g1205 (n1238, n672, n1218, n735);
and  g1206 (n1220, n703, n675, n1214, n1217);
or   g1207 (n1234, n1218, n1217, n730, n699);
xnor g1208 (n1227, n676, n737, n692, n717);
xor  g1209 (n1240, n724, n727, n1215, n704);
and  g1210 (n1244, n686, n1215, n701, n689);
xor  g1211 (n1243, n702, n696, n706, n1212);
or   g1212 (n1237, n1214, n673, n708, n716);
or   g1213 (n1232, n1026, n731, n663, n728);
nor  g1214 (n1242, n736, n681, n688, n732);
nor  g1215 (n1225, n682, n693, n695, n713);
nand g1216 (n1231, n1216, n1214, n714, n1212);
xor  g1217 (n1224, n669, n715, n700, n1217);
xor  g1218 (n1221, n665, n722, n1126, n707);
and  g1219 (n1222, n683, n705, n1213, n1217);
nand g1220 (n1246, n711, n1215, n685, n1212);
nand g1221 (n1226, n1218, n661, n720, n709);
xnor g1222 (n1229, n670, n697, n687, n1126);
xor  g1223 (n1236, n1216, n1213, n680);
nor  g1224 (n1228, n667, n729, n738, n690);
nand g1225 (n1241, n694, n1126, n677, n712);
or   g1226 (n1277, n795, n1244, n864, n787);
xor  g1227 (n1265, n1031, n803, n791, n757);
and  g1228 (n1248, n20, n745, n838, n1233);
nand g1229 (n1250, n17, n827, n1228, n774);
and  g1230 (n1279, n1028, n1224, n1239, n775);
nor  g1231 (n1286, n742, n790, n1240, n842);
nand g1232 (n1258, n15, n17, n14, n1229);
xnor g1233 (n1303, n756, n847, n1032, n862);
and  g1234 (n1301, n763, n853, n1243, n1028);
nor  g1235 (n1257, n754, n840, n1032, n753);
nor  g1236 (n1291, n1030, n1230, n1245, n819);
nand g1237 (n1304, n750, n761, n15, n1239);
and  g1238 (n1247, n867, n1243, n764, n849);
and  g1239 (n1263, n1238, n826, n814, n794);
and  g1240 (n1283, n848, n868, n1231, n1033);
xor  g1241 (n1260, n1246, n1221, n743, n866);
xor  g1242 (n1298, n845, n856, n779, n1241);
or   g1243 (n1288, n804, n1225, n1234, n813);
and  g1244 (n1280, n18, n1238, n1246, n1231);
xnor g1245 (n1282, n18, n839, n837, n1033);
nand g1246 (n1281, n786, n14, n19, n796);
or   g1247 (n1274, n824, n785, n802, n18);
or   g1248 (n1256, n800, n805, n1227, n860);
or   g1249 (n1297, n828, n799, n1241, n1237);
nor  g1250 (n1259, n863, n815, n1236, n841);
nand g1251 (n1289, n823, n780, n1239, n766);
nand g1252 (n1271, n788, n859, n835, n1235);
nor  g1253 (n1264, n1029, n830, n850, n1236);
xor  g1254 (n1262, n772, n1233, n1238, n744);
nand g1255 (n1273, n752, n20, n822, n1028);
nand g1256 (n1290, n749, n19, n861, n1235);
nor  g1257 (n1296, n793, n739, n769, n817);
or   g1258 (n1295, n1234, n1234, n1031, n16);
nand g1259 (n1307, n851, n810, n1246, n16);
nor  g1260 (n1272, n852, n773, n1032, n1033);
xnor g1261 (n1308, n1241, n17, n1150, n759);
or   g1262 (n1253, n15, n1031, n801, n1242);
xor  g1263 (n1267, n834, n833, n748, n747);
nor  g1264 (n1270, n1226, n843, n1030, n776);
and  g1265 (n1300, n829, n818, n846, n865);
nand g1266 (n1268, n858, n760, n1220, n1232);
xor  g1267 (n1305, n1242, n782, n1245, n1244);
or   g1268 (n1285, n820, n832, n1032, n778);
xor  g1269 (n1306, n811, n1236, n771, n1029);
nand g1270 (n1293, n831, n1027, n784, n751);
xnor g1271 (n1287, n812, n777, n770, n1219);
xnor g1272 (n1254, n781, n1150, n807, n16);
nor  g1273 (n1269, n1223, n857, n14, n19);
nor  g1274 (n1251, n20, n1244, n1242, n768);
or   g1275 (n1249, n855, n1028, n18, n1230);
nor  g1276 (n1302, n1030, n1243, n1033, n1029);
nor  g1277 (n1294, n1231, n1240, n1029, n1237);
xor  g1278 (n1275, n767, n740, n806, n16);
xor  g1279 (n1292, n1030, n765, n1233, n1245);
nand g1280 (n1276, n854, n1232, n1237, n783);
and  g1281 (n1266, n825, n1150, n836, n758);
xor  g1282 (n1261, n1232, n1222, n1240, n821);
xor  g1283 (n1284, n19, n792, n1031, n844);
xnor g1284 (n1255, n1230, n798, n17, n816);
or   g1285 (n1278, n1235, n741, n14, n762);
or   g1286 (n1252, n808, n789, n809, n797);
nor  g1287 (n1299, n755, n20, n746, n15);
or   g1288 (n1313, n28, n25, n41, n1305);
nand g1289 (n1369, n52, n60, n32, n71);
and  g1290 (n1318, n28, n55, n65, n27);
and  g1291 (n1349, n26, n1284, n35, n55);
nor  g1292 (n1332, n38, n1251, n57, n29);
and  g1293 (n1337, n46, n1272, n65, n1308);
nor  g1294 (n1359, n43, n27, n1253, n1261);
or   g1295 (n1366, n1296, n1293, n72);
and  g1296 (n1362, n48, n1275, n39, n58);
xnor g1297 (n1314, n62, n43, n42, n52);
nand g1298 (n1339, n1249, n1289, n1297, n35);
xor  g1299 (n1317, n48, n62, n31, n45);
nand g1300 (n1324, n60, n1264, n1255, n47);
and  g1301 (n1320, n1270, n1282, n42, n1304);
and  g1302 (n1331, n32, n37, n1248, n51);
nor  g1303 (n1370, n52, n1263, n26, n66);
nand g1304 (n1354, n1280, n1266, n70, n60);
or   g1305 (n1351, n30, n47, n56, n59);
nor  g1306 (n1371, n25, n1301, n46, n1285);
and  g1307 (n1311, n36, n67, n1256, n43);
or   g1308 (n1346, n53, n68, n36, n64);
or   g1309 (n1322, n72, n41, n44, n46);
or   g1310 (n1355, n1295, n1278, n51, n42);
nand g1311 (n1343, n31, n1271, n61, n54);
or   g1312 (n1364, n1307, n33, n1258, n56);
xor  g1313 (n1334, n34, n56, n57, n45);
and  g1314 (n1360, n40, n48, n50, n1268);
and  g1315 (n1353, n49, n38, n28, n25);
nor  g1316 (n1336, n58, n41, n35, n68);
nand g1317 (n1372, n40, n52, n50, n35);
xor  g1318 (n1357, n69, n44, n61, n68);
nor  g1319 (n1309, n30, n38, n50, n69);
nor  g1320 (n1358, n49, n31, n62, n58);
nor  g1321 (n1352, n61, n65, n1303, n66);
or   g1322 (n1325, n1302, n59, n1250, n57);
xor  g1323 (n1330, n30, n26, n68, n45);
nor  g1324 (n1328, n51, n60, n1292, n44);
and  g1325 (n1335, n53, n1277, n63, n37);
xnor g1326 (n1368, n1287, n46, n1291, n63);
xnor g1327 (n1327, n70, n1269, n33, n47);
and  g1328 (n1341, n31, n34, n1267, n45);
nand g1329 (n1333, n28, n26, n55, n1283);
and  g1330 (n1350, n27, n64, n32, n69);
nor  g1331 (n1363, n58, n71, n29, n50);
nand g1332 (n1338, n63, n34, n61, n54);
nand g1333 (n1321, n1276, n1308, n71, n62);
and  g1334 (n1367, n29, n1288, n34, n1294);
or   g1335 (n1315, n59, n39, n33, n1286);
xor  g1336 (n1342, n70, n54, n1274, n63);
xor  g1337 (n1348, n1265, n1299, n37, n69);
or   g1338 (n1365, n1281, n36, n51, n47);
xor  g1339 (n1323, n65, n37, n38, n27);
and  g1340 (n1361, n55, n72, n48, n64);
xor  g1341 (n1310, n49, n70, n56, n32);
nand g1342 (n1344, n1300, n41, n71, n53);
nor  g1343 (n1345, n1247, n1259, n49, n64);
xnor g1344 (n1340, n54, n25, n42, n1260);
nor  g1345 (n1319, n1257, n57, n1298, n1308);
nor  g1346 (n1347, n67, n67, n30, n1252);
nor  g1347 (n1356, n1273, n44, n59, n36);
xor  g1348 (n1312, n66, n1290, n67, n40);
xor  g1349 (n1316, n1254, n1262, n39, n40);
xor  g1350 (n1329, n53, n29, n33, n39);
xnor g1351 (n1326, n1279, n1306, n66, n43);
xor  g1352 (n1383, n1322, n1348, n1372, n1344);
nand g1353 (n1378, n1337, n1342, n1316, n1362);
nand g1354 (n1385, n1351, n1371, n1336, n1310);
nand g1355 (n1380, n1357, n1321, n1320, n1364);
and  g1356 (n1373, n1361, n1353, n1358, n1341);
nor  g1357 (n1388, n1328, n1329, n1331, n1347);
or   g1358 (n1377, n1365, n1313, n1309, n1324);
xnor g1359 (n1384, n1355, n1367, n1345, n1354);
or   g1360 (n1375, n1360, n1340, n1366, n1334);
nor  g1361 (n1382, n1350, n1325, n1359, n1327);
xor  g1362 (n1387, n1318, n1323, n1335, n1332);
nor  g1363 (n1376, n1346, n1369, n1339, n1338);
nor  g1364 (n1386, n1311, n1356, n1333, n1312);
xor  g1365 (n1381, n1326, n1314, n1368, n1363);
xnor g1366 (n1374, n1349, n1317, n1343, n1352);
nor  g1367 (n1379, n1315, n1330, n1319, n1370);
endmodule
