// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_201 written by SynthGen on 2021/04/05 11:23:24
module Stat_2000_201( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1069, n1036, n1901, n2024, n2031, n2020, n2030, n2009,
 n2023, n2026, n2018, n2022, n2019, n2011, n2021, n2012,
 n2005, n2017, n2007, n2016, n2013, n2004, n2032, n2014,
 n2025, n2010, n2028, n2015, n2027, n2006, n2029, n2008);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1069, n1036, n1901, n2024, n2031, n2020, n2030, n2009,
 n2023, n2026, n2018, n2022, n2019, n2011, n2021, n2012,
 n2005, n2017, n2007, n2016, n2013, n2004, n2032, n2014,
 n2025, n2010, n2028, n2015, n2027, n2006, n2029, n2008;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1902, n1903, n1904, n1905, n1906, n1907,
 n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
 n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
 n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
 n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
 n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
 n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
 n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
 n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
 n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
 n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
 n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
 n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003;

not  g0 (n145, n32);
buf  g1 (n116, n2);
buf  g2 (n130, n24);
buf  g3 (n141, n6);
buf  g4 (n67, n13);
not  g5 (n126, n2);
not  g6 (n46, n21);
buf  g7 (n79, n18);
not  g8 (n53, n31);
not  g9 (n151, n27);
buf  g10 (n146, n8);
not  g11 (n107, n21);
buf  g12 (n57, n17);
buf  g13 (n62, n30);
not  g14 (n66, n32);
buf  g15 (n132, n6);
buf  g16 (n148, n18);
buf  g17 (n85, n20);
not  g18 (n56, n5);
not  g19 (n54, n11);
not  g20 (n104, n4);
buf  g21 (n92, n23);
not  g22 (n33, n7);
not  g23 (n105, n19);
buf  g24 (n68, n28);
buf  g25 (n50, n16);
not  g26 (n38, n23);
buf  g27 (n39, n3);
not  g28 (n119, n26);
buf  g29 (n65, n7);
not  g30 (n125, n17);
buf  g31 (n81, n11);
not  g32 (n60, n31);
buf  g33 (n43, n29);
buf  g34 (n99, n21);
buf  g35 (n111, n1);
not  g36 (n110, n1);
buf  g37 (n159, n17);
buf  g38 (n51, n26);
not  g39 (n106, n4);
buf  g40 (n91, n10);
buf  g41 (n143, n20);
not  g42 (n147, n29);
not  g43 (n109, n26);
not  g44 (n112, n17);
not  g45 (n113, n28);
buf  g46 (n101, n15);
not  g47 (n97, n14);
buf  g48 (n88, n7);
not  g49 (n78, n29);
buf  g50 (n140, n11);
not  g51 (n74, n14);
buf  g52 (n156, n3);
buf  g53 (n87, n1);
not  g54 (n135, n8);
buf  g55 (n73, n30);
buf  g56 (n63, n18);
buf  g57 (n34, n16);
not  g58 (n58, n11);
not  g59 (n86, n20);
buf  g60 (n83, n27);
buf  g61 (n100, n25);
buf  g62 (n52, n5);
not  g63 (n42, n16);
buf  g64 (n36, n13);
buf  g65 (n123, n22);
buf  g66 (n98, n1);
not  g67 (n72, n23);
buf  g68 (n82, n26);
buf  g69 (n155, n15);
not  g70 (n121, n23);
buf  g71 (n136, n18);
buf  g72 (n102, n8);
not  g73 (n71, n9);
not  g74 (n127, n2);
buf  g75 (n61, n27);
buf  g76 (n158, n6);
not  g77 (n84, n22);
not  g78 (n55, n9);
not  g79 (n49, n19);
buf  g80 (n118, n15);
not  g81 (n144, n22);
buf  g82 (n69, n24);
buf  g83 (n59, n2);
not  g84 (n77, n28);
not  g85 (n120, n24);
buf  g86 (n142, n19);
buf  g87 (n133, n9);
buf  g88 (n95, n28);
not  g89 (n80, n13);
not  g90 (n89, n5);
not  g91 (n35, n7);
buf  g92 (n138, n24);
buf  g93 (n137, n31);
not  g94 (n40, n16);
not  g95 (n48, n10);
buf  g96 (n124, n29);
buf  g97 (n70, n30);
not  g98 (n157, n32);
buf  g99 (n108, n31);
not  g100 (n64, n8);
not  g101 (n115, n19);
buf  g102 (n117, n3);
buf  g103 (n150, n9);
not  g104 (n96, n5);
buf  g105 (n131, n25);
not  g106 (n37, n13);
buf  g107 (n114, n10);
buf  g108 (n41, n14);
buf  g109 (n154, n3);
buf  g110 (n103, n4);
buf  g111 (n122, n21);
not  g112 (n134, n27);
buf  g113 (n139, n12);
not  g114 (n153, n4);
not  g115 (n93, n12);
not  g116 (n149, n12);
not  g117 (n152, n12);
not  g118 (n129, n15);
buf  g119 (n44, n25);
not  g120 (n47, n20);
buf  g121 (n75, n14);
not  g122 (n76, n10);
buf  g123 (n90, n6);
buf  g124 (n128, n30);
buf  g125 (n45, n22);
not  g126 (n94, n25);
not  g127 (n399, n91);
buf  g128 (n175, n51);
not  g129 (n662, n40);
not  g130 (n514, n37);
not  g131 (n663, n156);
not  g132 (n340, n66);
buf  g133 (n327, n152);
not  g134 (n550, n62);
not  g135 (n497, n78);
not  g136 (n513, n146);
not  g137 (n600, n156);
not  g138 (n469, n46);
buf  g139 (n527, n143);
buf  g140 (n632, n104);
not  g141 (n197, n69);
buf  g142 (n230, n138);
not  g143 (n451, n124);
not  g144 (n416, n108);
buf  g145 (n471, n49);
not  g146 (n552, n69);
buf  g147 (n348, n50);
not  g148 (n524, n74);
buf  g149 (n459, n33);
not  g150 (n634, n122);
not  g151 (n216, n92);
buf  g152 (n371, n76);
not  g153 (n617, n38);
not  g154 (n402, n37);
buf  g155 (n473, n33);
buf  g156 (n183, n58);
buf  g157 (n211, n106);
buf  g158 (n379, n154);
buf  g159 (n453, n113);
buf  g160 (n384, n54);
buf  g161 (n176, n84);
buf  g162 (n648, n39);
buf  g163 (n330, n68);
buf  g164 (n201, n100);
not  g165 (n179, n130);
buf  g166 (n406, n108);
not  g167 (n498, n102);
not  g168 (n202, n66);
buf  g169 (n626, n99);
not  g170 (n364, n135);
buf  g171 (n658, n76);
not  g172 (n217, n154);
buf  g173 (n564, n59);
not  g174 (n533, n61);
not  g175 (n590, n117);
not  g176 (n253, n76);
not  g177 (n544, n84);
buf  g178 (n562, n78);
buf  g179 (n418, n148);
not  g180 (n549, n94);
not  g181 (n643, n155);
not  g182 (n357, n146);
not  g183 (n646, n33);
not  g184 (n267, n98);
buf  g185 (n488, n124);
not  g186 (n342, n36);
buf  g187 (n667, n101);
not  g188 (n186, n118);
buf  g189 (n571, n88);
buf  g190 (n581, n124);
buf  g191 (n325, n128);
not  g192 (n242, n108);
not  g193 (n509, n87);
buf  g194 (n535, n145);
not  g195 (n236, n139);
not  g196 (n422, n68);
buf  g197 (n461, n55);
buf  g198 (n203, n130);
buf  g199 (n583, n105);
not  g200 (n466, n132);
buf  g201 (n537, n47);
buf  g202 (n538, n46);
buf  g203 (n647, n111);
not  g204 (n353, n79);
not  g205 (n413, n91);
buf  g206 (n446, n125);
buf  g207 (n394, n92);
not  g208 (n610, n78);
buf  g209 (n561, n85);
buf  g210 (n246, n119);
not  g211 (n243, n158);
buf  g212 (n226, n54);
not  g213 (n288, n65);
not  g214 (n219, n111);
not  g215 (n569, n96);
not  g216 (n547, n94);
buf  g217 (n664, n143);
buf  g218 (n511, n76);
not  g219 (n304, n39);
not  g220 (n350, n144);
buf  g221 (n287, n148);
buf  g222 (n409, n138);
not  g223 (n380, n102);
not  g224 (n387, n149);
not  g225 (n199, n81);
not  g226 (n339, n99);
not  g227 (n563, n81);
buf  g228 (n265, n107);
not  g229 (n574, n60);
not  g230 (n444, n114);
buf  g231 (n652, n94);
buf  g232 (n361, n68);
not  g233 (n629, n92);
buf  g234 (n595, n93);
not  g235 (n349, n133);
not  g236 (n536, n73);
not  g237 (n255, n52);
buf  g238 (n337, n146);
not  g239 (n531, n38);
not  g240 (n518, n135);
buf  g241 (n496, n132);
not  g242 (n290, n112);
not  g243 (n316, n150);
buf  g244 (n597, n113);
buf  g245 (n633, n103);
not  g246 (n294, n52);
not  g247 (n654, n60);
buf  g248 (n485, n93);
not  g249 (n463, n92);
not  g250 (n400, n132);
not  g251 (n307, n34);
not  g252 (n336, n33);
buf  g253 (n480, n106);
not  g254 (n167, n49);
not  g255 (n378, n112);
buf  g256 (n502, n87);
not  g257 (n188, n109);
not  g258 (n492, n157);
buf  g259 (n331, n96);
buf  g260 (n576, n57);
not  g261 (n543, n109);
not  g262 (n508, n139);
buf  g263 (n411, n121);
not  g264 (n171, n86);
buf  g265 (n495, n103);
buf  g266 (n209, n113);
buf  g267 (n443, n152);
not  g268 (n232, n85);
not  g269 (n620, n96);
not  g270 (n630, n115);
not  g271 (n441, n136);
buf  g272 (n185, n65);
not  g273 (n315, n116);
buf  g274 (n439, n73);
buf  g275 (n368, n151);
buf  g276 (n417, n40);
buf  g277 (n631, n149);
not  g278 (n475, n115);
not  g279 (n570, n159);
buf  g280 (n427, n134);
buf  g281 (n559, n71);
not  g282 (n401, n69);
buf  g283 (n546, n128);
not  g284 (n656, n85);
buf  g285 (n636, n135);
buf  g286 (n362, n104);
not  g287 (n397, n42);
buf  g288 (n189, n102);
not  g289 (n404, n81);
buf  g290 (n582, n47);
not  g291 (n604, n47);
not  g292 (n333, n36);
not  g293 (n472, n127);
not  g294 (n248, n126);
not  g295 (n528, n89);
not  g296 (n258, n143);
buf  g297 (n395, n97);
not  g298 (n355, n90);
not  g299 (n205, n58);
not  g300 (n273, n86);
not  g301 (n251, n70);
buf  g302 (n231, n139);
not  g303 (n212, n42);
buf  g304 (n244, n77);
buf  g305 (n615, n95);
not  g306 (n187, n120);
not  g307 (n602, n141);
buf  g308 (n424, n144);
buf  g309 (n181, n88);
not  g310 (n366, n63);
not  g311 (n506, n43);
buf  g312 (n593, n86);
buf  g313 (n296, n123);
buf  g314 (n426, n37);
buf  g315 (n510, n51);
buf  g316 (n437, n131);
buf  g317 (n291, n59);
not  g318 (n207, n145);
not  g319 (n445, n113);
not  g320 (n623, n115);
buf  g321 (n341, n73);
buf  g322 (n609, n34);
not  g323 (n343, n139);
not  g324 (n430, n64);
buf  g325 (n180, n72);
buf  g326 (n660, n153);
not  g327 (n650, n149);
buf  g328 (n190, n118);
not  g329 (n486, n123);
buf  g330 (n539, n45);
buf  g331 (n173, n125);
not  g332 (n584, n117);
not  g333 (n522, n54);
not  g334 (n436, n82);
not  g335 (n354, n151);
not  g336 (n503, n142);
not  g337 (n454, n62);
not  g338 (n312, n72);
buf  g339 (n655, n140);
buf  g340 (n318, n58);
buf  g341 (n194, n116);
buf  g342 (n228, n89);
not  g343 (n249, n157);
buf  g344 (n612, n138);
not  g345 (n618, n151);
buf  g346 (n271, n73);
buf  g347 (n237, n60);
buf  g348 (n160, n130);
not  g349 (n196, n41);
not  g350 (n640, n44);
not  g351 (n580, n137);
buf  g352 (n616, n84);
buf  g353 (n286, n141);
buf  g354 (n462, n107);
not  g355 (n554, n140);
buf  g356 (n499, n89);
buf  g357 (n585, n152);
not  g358 (n365, n41);
buf  g359 (n659, n61);
not  g360 (n545, n110);
not  g361 (n260, n120);
buf  g362 (n392, n147);
not  g363 (n182, n34);
not  g364 (n346, n64);
buf  g365 (n532, n112);
buf  g366 (n234, n119);
buf  g367 (n611, n137);
buf  g368 (n603, n146);
not  g369 (n192, n118);
not  g370 (n589, n158);
buf  g371 (n405, n157);
not  g372 (n592, n68);
buf  g373 (n359, n74);
not  g374 (n165, n90);
not  g375 (n245, n57);
buf  g376 (n625, n93);
buf  g377 (n627, n36);
not  g378 (n521, n66);
buf  g379 (n279, n151);
not  g380 (n484, n70);
buf  g381 (n568, n74);
not  g382 (n391, n77);
not  g383 (n526, n106);
not  g384 (n601, n93);
not  g385 (n651, n48);
not  g386 (n573, n42);
buf  g387 (n322, n62);
buf  g388 (n588, n134);
buf  g389 (n283, n152);
not  g390 (n374, n138);
not  g391 (n222, n148);
buf  g392 (n501, n83);
buf  g393 (n320, n64);
not  g394 (n324, n63);
not  g395 (n308, n147);
buf  g396 (n272, n35);
not  g397 (n591, n79);
buf  g398 (n345, n91);
buf  g399 (n375, n79);
buf  g400 (n565, n136);
buf  g401 (n386, n72);
not  g402 (n504, n35);
not  g403 (n238, n87);
buf  g404 (n619, n140);
buf  g405 (n530, n89);
buf  g406 (n500, n98);
not  g407 (n420, n105);
not  g408 (n206, n38);
not  g409 (n373, n35);
not  g410 (n390, n80);
not  g411 (n607, n67);
buf  g412 (n332, n53);
not  g413 (n363, n121);
buf  g414 (n464, n48);
buf  g415 (n520, n129);
not  g416 (n313, n34);
not  g417 (n487, n71);
not  g418 (n637, n144);
buf  g419 (n447, n136);
buf  g420 (n195, n65);
buf  g421 (n452, n45);
buf  g422 (n319, n125);
buf  g423 (n227, n121);
buf  g424 (n270, n147);
buf  g425 (n263, n70);
not  g426 (n164, n112);
not  g427 (n557, n107);
buf  g428 (n661, n115);
buf  g429 (n281, n55);
not  g430 (n275, n114);
not  g431 (n352, n55);
buf  g432 (n264, n124);
not  g433 (n598, n52);
buf  g434 (n382, n129);
buf  g435 (n262, n50);
not  g436 (n621, n155);
buf  g437 (n274, n129);
buf  g438 (n577, n100);
not  g439 (n635, n158);
not  g440 (n624, n88);
buf  g441 (n414, n117);
buf  g442 (n323, n153);
buf  g443 (n385, n79);
not  g444 (n177, n41);
not  g445 (n478, n140);
not  g446 (n204, n119);
buf  g447 (n622, n136);
not  g448 (n259, n109);
buf  g449 (n280, n131);
buf  g450 (n241, n83);
buf  g451 (n200, n103);
buf  g452 (n169, n144);
not  g453 (n435, n155);
buf  g454 (n299, n56);
not  g455 (n567, n119);
buf  g456 (n184, n127);
not  g457 (n172, n43);
buf  g458 (n221, n75);
not  g459 (n542, n46);
not  g460 (n377, n127);
buf  g461 (n408, n142);
buf  g462 (n208, n154);
not  g463 (n193, n59);
not  g464 (n335, n98);
buf  g465 (n317, n153);
not  g466 (n305, n63);
buf  g467 (n376, n49);
not  g468 (n470, n110);
not  g469 (n419, n122);
buf  g470 (n481, n126);
not  g471 (n489, n125);
not  g472 (n170, n104);
buf  g473 (n289, n56);
buf  g474 (n523, n67);
not  g475 (n415, n40);
not  g476 (n553, n106);
not  g477 (n638, n116);
buf  g478 (n358, n109);
buf  g479 (n605, n53);
buf  g480 (n455, n47);
buf  g481 (n163, n100);
not  g482 (n220, n56);
buf  g483 (n556, n101);
buf  g484 (n393, n129);
not  g485 (n301, n137);
not  g486 (n293, n128);
buf  g487 (n644, n130);
buf  g488 (n256, n137);
buf  g489 (n225, n99);
not  g490 (n210, n102);
buf  g491 (n449, n71);
buf  g492 (n328, n131);
not  g493 (n347, n75);
not  g494 (n282, n50);
not  g495 (n174, n97);
buf  g496 (n512, n159);
not  g497 (n433, n111);
not  g498 (n295, n77);
not  g499 (n587, n58);
not  g500 (n423, n80);
buf  g501 (n292, n43);
buf  g502 (n560, n120);
buf  g503 (n344, n110);
not  g504 (n596, n87);
buf  g505 (n572, n105);
buf  g506 (n429, n45);
not  g507 (n474, n114);
buf  g508 (n410, n135);
buf  g509 (n306, n155);
not  g510 (n303, n128);
not  g511 (n614, n52);
not  g512 (n389, n150);
not  g513 (n613, n45);
not  g514 (n541, n84);
buf  g515 (n440, n83);
buf  g516 (n298, n150);
buf  g517 (n431, n65);
not  g518 (n442, n95);
not  g519 (n278, n41);
not  g520 (n398, n134);
not  g521 (n266, n145);
buf  g522 (n608, n150);
not  g523 (n356, n156);
not  g524 (n642, n158);
not  g525 (n493, n120);
buf  g526 (n240, n56);
not  g527 (n168, n37);
buf  g528 (n428, n69);
not  g529 (n314, n108);
not  g530 (n606, n74);
not  g531 (n224, n127);
not  g532 (n566, n148);
buf  g533 (n425, n114);
buf  g534 (n178, n63);
not  g535 (n465, n141);
buf  g536 (n250, n70);
not  g537 (n233, n62);
not  g538 (n482, n156);
not  g539 (n310, n133);
not  g540 (n551, n101);
not  g541 (n548, n116);
buf  g542 (n434, n48);
not  g543 (n653, n80);
not  g544 (n507, n42);
not  g545 (n457, n36);
buf  g546 (n456, n55);
not  g547 (n494, n82);
buf  g548 (n468, n122);
not  g549 (n338, n49);
buf  g550 (n460, n57);
buf  g551 (n639, n133);
buf  g552 (n257, n153);
buf  g553 (n284, n97);
buf  g554 (n599, n77);
not  g555 (n421, n100);
not  g556 (n229, n39);
buf  g557 (n311, n64);
not  g558 (n476, n78);
not  g559 (n477, n61);
not  g560 (n351, n59);
not  g561 (n370, n82);
not  g562 (n525, n117);
buf  g563 (n329, n94);
buf  g564 (n448, n159);
buf  g565 (n369, n71);
buf  g566 (n223, n51);
not  g567 (n277, n81);
buf  g568 (n309, n97);
not  g569 (n285, n142);
not  g570 (n388, n35);
buf  g571 (n235, n61);
not  g572 (n360, n96);
not  g573 (n594, n75);
buf  g574 (n529, n154);
buf  g575 (n555, n85);
not  g576 (n252, n39);
buf  g577 (n458, n90);
buf  g578 (n450, n66);
not  g579 (n166, n44);
buf  g580 (n641, n134);
buf  g581 (n628, n101);
buf  g582 (n491, n57);
buf  g583 (n579, n82);
buf  g584 (n645, n54);
not  g585 (n432, n159);
buf  g586 (n540, n131);
buf  g587 (n517, n111);
buf  g588 (n586, n95);
buf  g589 (n516, n123);
buf  g590 (n575, n118);
buf  g591 (n534, n60);
buf  g592 (n578, n132);
not  g593 (n297, n145);
buf  g594 (n490, n51);
not  g595 (n326, n126);
buf  g596 (n479, n90);
buf  g597 (n247, n147);
not  g598 (n334, n107);
not  g599 (n218, n104);
not  g600 (n383, n122);
not  g601 (n261, n123);
not  g602 (n396, n126);
buf  g603 (n649, n105);
not  g604 (n269, n38);
buf  g605 (n438, n143);
buf  g606 (n483, n110);
buf  g607 (n302, n44);
not  g608 (n321, n86);
not  g609 (n214, n53);
buf  g610 (n558, n80);
not  g611 (n191, n43);
not  g612 (n239, n46);
not  g613 (n162, n67);
not  g614 (n215, n141);
not  g615 (n381, n44);
buf  g616 (n467, n99);
not  g617 (n657, n95);
not  g618 (n412, n103);
buf  g619 (n407, n88);
not  g620 (n665, n72);
not  g621 (n403, n83);
not  g622 (n505, n149);
buf  g623 (n161, n53);
buf  g624 (n519, n157);
buf  g625 (n367, n133);
buf  g626 (n213, n48);
not  g627 (n268, n50);
not  g628 (n300, n75);
not  g629 (n666, n121);
not  g630 (n276, n91);
not  g631 (n515, n40);
buf  g632 (n372, n98);
not  g633 (n254, n142);
buf  g634 (n198, n67);
buf  g635 (n784, n308);
not  g636 (n879, n427);
buf  g637 (n677, n377);
not  g638 (n811, n447);
not  g639 (n858, n358);
not  g640 (n672, n468);
not  g641 (n913, n369);
not  g642 (n698, n316);
not  g643 (n793, n206);
buf  g644 (n730, n380);
buf  g645 (n739, n553);
buf  g646 (n794, n565);
not  g647 (n919, n549);
not  g648 (n866, n276);
not  g649 (n831, n490);
buf  g650 (n916, n559);
buf  g651 (n914, n265);
not  g652 (n843, n554);
buf  g653 (n851, n224);
buf  g654 (n818, n504);
not  g655 (n878, n323);
not  g656 (n817, n240);
buf  g657 (n892, n246);
buf  g658 (n734, n214);
buf  g659 (n829, n357);
buf  g660 (n671, n275);
buf  g661 (n722, n235);
not  g662 (n751, n328);
buf  g663 (n714, n415);
buf  g664 (n876, n486);
buf  g665 (n826, n500);
not  g666 (n754, n386);
buf  g667 (n915, n300);
buf  g668 (n740, n229);
buf  g669 (n798, n330);
buf  g670 (n732, n250);
buf  g671 (n788, n351);
buf  g672 (n676, n399);
not  g673 (n761, n267);
not  g674 (n670, n301);
buf  g675 (n787, n459);
not  g676 (n762, n186);
not  g677 (n716, n251);
buf  g678 (n924, n527);
buf  g679 (n709, n493);
not  g680 (n796, n187);
not  g681 (n713, n203);
not  g682 (n891, n462);
not  g683 (n790, n383);
not  g684 (n691, n370);
not  g685 (n907, n464);
not  g686 (n680, n482);
buf  g687 (n721, n537);
buf  g688 (n723, n457);
not  g689 (n932, n506);
not  g690 (n888, n329);
buf  g691 (n899, n238);
not  g692 (n773, n181);
not  g693 (n690, n485);
not  g694 (n717, n465);
buf  g695 (n792, n172);
not  g696 (n872, n405);
buf  g697 (n682, n349);
not  g698 (n725, n228);
buf  g699 (n750, n350);
buf  g700 (n674, n322);
buf  g701 (n705, n563);
buf  g702 (n711, n178);
buf  g703 (n745, n575);
not  g704 (n812, n197);
buf  g705 (n718, n389);
not  g706 (n724, n494);
buf  g707 (n930, n560);
not  g708 (n673, n419);
not  g709 (n805, n217);
not  g710 (n766, n492);
not  g711 (n862, n470);
not  g712 (n871, n367);
not  g713 (n869, n288);
not  g714 (n885, n564);
not  g715 (n854, n574);
not  g716 (n845, n518);
buf  g717 (n702, n422);
buf  g718 (n810, n437);
not  g719 (n696, n339);
buf  g720 (n837, n579);
buf  g721 (n802, n283);
not  g722 (n777, n438);
buf  g723 (n883, n365);
buf  g724 (n921, n484);
not  g725 (n875, n539);
buf  g726 (n808, n223);
not  g727 (n688, n523);
not  g728 (n853, n298);
not  g729 (n731, n261);
buf  g730 (n873, n208);
buf  g731 (n737, n222);
buf  g732 (n746, n215);
buf  g733 (n807, n184);
not  g734 (n785, n216);
not  g735 (n749, n403);
not  g736 (n701, n234);
not  g737 (n779, n268);
not  g738 (n848, n277);
buf  g739 (n694, n175);
buf  g740 (n755, n204);
not  g741 (n896, n176);
buf  g742 (n855, n376);
not  g743 (n706, n513);
buf  g744 (n840, n286);
not  g745 (n909, n347);
not  g746 (n923, n372);
not  g747 (n703, n243);
not  g748 (n804, n356);
not  g749 (n776, n368);
buf  g750 (n849, n558);
buf  g751 (n870, n211);
not  g752 (n668, n289);
not  g753 (n936, n318);
not  g754 (n799, n555);
not  g755 (n859, n269);
and  g756 (n738, n543, n279);
or   g757 (n775, n291, n418);
xor  g758 (n707, n408, n515);
xor  g759 (n882, n202, n331);
xnor g760 (n757, n168, n429);
xnor g761 (n693, n471, n233);
xor  g762 (n772, n432, n454);
xor  g763 (n823, n430, n189);
xor  g764 (n748, n311, n535);
xor  g765 (n720, n232, n502);
xor  g766 (n685, n461, n236);
and  g767 (n774, n538, n337);
nand g768 (n860, n325, n548);
nand g769 (n928, n312, n340);
nand g770 (n767, n381, n508);
or   g771 (n874, n402, n561);
nand g772 (n763, n573, n534);
xnor g773 (n678, n266, n442);
or   g774 (n898, n584, n374);
or   g775 (n783, n314, n580);
xor  g776 (n911, n517, n570);
nand g777 (n927, n556, n388);
nor  g778 (n768, n509, n213);
xor  g779 (n736, n507, n257);
or   g780 (n704, n373, n263);
and  g781 (n926, n307, n285);
nor  g782 (n675, n274, n396);
xor  g783 (n841, n505, n463);
or   g784 (n764, n533, n446);
nand g785 (n850, n362, n487);
xnor g786 (n758, n363, n452);
nand g787 (n903, n218, n551);
xnor g788 (n809, n467, n207);
xnor g789 (n814, n503, n581);
xor  g790 (n938, n491, n434);
or   g791 (n828, n576, n210);
xor  g792 (n669, n520, n393);
xor  g793 (n712, n273, n571);
xnor g794 (n827, n302, n443);
or   g795 (n931, n309, n237);
or   g796 (n729, n253, n526);
xnor g797 (n897, n220, n466);
xor  g798 (n819, n425, n310);
and  g799 (n834, n428, n477);
xnor g800 (n789, n209, n315);
nor  g801 (n863, n359, n201);
or   g802 (n697, n530, n199);
xor  g803 (n781, n426, n242);
nand g804 (n902, n449, n212);
xor  g805 (n686, n542, n583);
and  g806 (n679, n258, n395);
nand g807 (n733, n541, n497);
and  g808 (n816, n510, n255);
nand g809 (n906, n336, n180);
xor  g810 (n735, n287, n448);
or   g811 (n846, n424, n173);
nand g812 (n795, n163, n499);
xnor g813 (n778, n247, n552);
and  g814 (n681, n196, n192);
and  g815 (n825, n327, n294);
nor  g816 (n824, n413, n456);
nor  g817 (n822, n566, n171);
nor  g818 (n838, n183, n352);
xor  g819 (n884, n512, n572);
nor  g820 (n877, n444, n441);
nand g821 (n868, n519, n296);
nand g822 (n900, n264, n185);
nand g823 (n727, n451, n227);
and  g824 (n861, n360, n525);
xnor g825 (n743, n390, n321);
xnor g826 (n925, n416, n343);
and  g827 (n760, n225, n378);
nand g828 (n832, n406, n511);
and  g829 (n803, n332, n320);
xnor g830 (n801, n557, n342);
nor  g831 (n769, n221, n411);
and  g832 (n857, n480, n407);
xnor g833 (n747, n398, n475);
nor  g834 (n889, n160, n167);
nand g835 (n800, n540, n170);
xnor g836 (n700, n293, n546);
xor  g837 (n695, n384, n578);
and  g838 (n833, n479, n272);
xor  g839 (n821, n324, n420);
xnor g840 (n842, n544, n524);
and  g841 (n893, n241, n379);
or   g842 (n847, n483, n182);
xor  g843 (n922, n385, n319);
nand g844 (n920, n495, n231);
and  g845 (n744, n259, n194);
nor  g846 (n905, n473, n521);
nand g847 (n683, n165, n387);
xor  g848 (n856, n476, n421);
xnor g849 (n782, n412, n547);
and  g850 (n904, n278, n562);
nor  g851 (n689, n290, n392);
xnor g852 (n917, n353, n219);
nor  g853 (n687, n179, n436);
nor  g854 (n940, n439, n472);
xor  g855 (n895, n453, n254);
and  g856 (n867, n305, n409);
nor  g857 (n937, n306, n582);
and  g858 (n881, n177, n366);
nand g859 (n933, n361, n433);
and  g860 (n699, n334, n166);
nand g861 (n806, n488, n417);
and  g862 (n852, n256, n391);
nor  g863 (n728, n280, n371);
nand g864 (n742, n404, n193);
xnor g865 (n886, n317, n198);
or   g866 (n929, n262, n364);
nand g867 (n887, n445, n478);
nor  g868 (n934, n252, n354);
and  g869 (n813, n498, n355);
nand g870 (n835, n460, n410);
or   g871 (n692, n375, n496);
or   g872 (n839, n397, n458);
or   g873 (n890, n346, n239);
or   g874 (n765, n516, n401);
xor  g875 (n791, n394, n450);
nand g876 (n710, n169, n501);
nand g877 (n880, n423, n313);
nand g878 (n759, n270, n297);
or   g879 (n726, n435, n474);
nor  g880 (n830, n248, n304);
and  g881 (n752, n226, n205);
or   g882 (n797, n284, n200);
nor  g883 (n708, n333, n244);
and  g884 (n780, n348, n469);
nand g885 (n939, n536, n245);
nand g886 (n901, n271, n545);
and  g887 (n836, n522, n550);
nor  g888 (n844, n514, n338);
or   g889 (n918, n303, n299);
or   g890 (n715, n260, n195);
xnor g891 (n894, n341, n230);
nor  g892 (n865, n292, n191);
xnor g893 (n815, n345, n455);
xnor g894 (n770, n568, n295);
nor  g895 (n910, n489, n382);
xnor g896 (n935, n281, n161);
xnor g897 (n771, n431, n528);
and  g898 (n864, n249, n440);
or   g899 (n753, n174, n567);
xnor g900 (n684, n164, n532);
nand g901 (n756, n400, n531);
nand g902 (n741, n282, n529);
xnor g903 (n912, n190, n481);
and  g904 (n820, n569, n326);
xnor g905 (n786, n414, n344);
nor  g906 (n908, n162, n188);
nand g907 (n719, n577, n335);
buf  g908 (n955, n683);
buf  g909 (n957, n672);
buf  g910 (n943, n693);
not  g911 (n953, n676);
buf  g912 (n956, n686);
not  g913 (n958, n692);
not  g914 (n949, n689);
not  g915 (n948, n694);
not  g916 (n951, n677);
not  g917 (n942, n681);
not  g918 (n959, n679);
buf  g919 (n960, n671);
not  g920 (n950, n695);
not  g921 (n952, n670);
and  g922 (n961, n674, n691);
or   g923 (n947, n685, n682);
or   g924 (n945, n675, n680);
nor  g925 (n946, n688, n687);
nand g926 (n944, n696, n684);
and  g927 (n954, n669, n673);
nor  g928 (n941, n678, n690);
not  g929 (n969, n714);
buf  g930 (n971, n953);
buf  g931 (n981, n945);
not  g932 (n977, n961);
buf  g933 (n978, n698);
buf  g934 (n982, n713);
buf  g935 (n962, n700);
not  g936 (n980, n956);
buf  g937 (n979, n958);
not  g938 (n974, n702);
not  g939 (n965, n722);
buf  g940 (n963, n721);
buf  g941 (n966, n952);
or   g942 (n975, n705, n955, n943);
nor  g943 (n964, n716, n697, n708, n941);
or   g944 (n968, n719, n951, n717, n706);
and  g945 (n967, n709, n954, n960, n701);
and  g946 (n983, n703, n944, n710, n949);
nand g947 (n970, n942, n948, n699, n950);
and  g948 (n973, n704, n946, n718, n957);
and  g949 (n972, n707, n715, n720, n961);
or   g950 (n976, n712, n947, n711, n959);
buf  g951 (n1030, n734);
buf  g952 (n985, n737);
not  g953 (n994, n970);
buf  g954 (n1016, n755);
buf  g955 (n1029, n736);
buf  g956 (n992, n733);
buf  g957 (n996, n972);
not  g958 (n1003, n962);
buf  g959 (n1024, n962);
not  g960 (n1012, n730);
not  g961 (n986, n749);
buf  g962 (n993, n963);
not  g963 (n1026, n735);
buf  g964 (n1027, n771);
not  g965 (n989, n723);
buf  g966 (n997, n728);
buf  g967 (n1023, n751);
buf  g968 (n1013, n759);
buf  g969 (n1014, n964);
not  g970 (n1006, n761);
not  g971 (n1005, n732);
not  g972 (n1009, n750);
buf  g973 (n1001, n969);
buf  g974 (n1010, n738);
buf  g975 (n1008, n770);
buf  g976 (n999, n970);
not  g977 (n1025, n968);
not  g978 (n995, n739);
not  g979 (n990, n967);
not  g980 (n1017, n724);
buf  g981 (n1000, n966);
not  g982 (n987, n760);
or   g983 (n1002, n731, n974);
xor  g984 (n1020, n963, n966, n970, n962);
xnor g985 (n1018, n965, n774, n773, n973);
xnor g986 (n1022, n971, n965, n968, n772);
or   g987 (n1019, n968, n972, n971, n766);
xor  g988 (n1021, n725, n746, n971, n963);
or   g989 (n998, n964, n740, n963, n741);
nand g990 (n984, n742, n745, n969, n754);
xor  g991 (n1015, n752, n763, n748, n973);
or   g992 (n991, n972, n970, n964, n756);
or   g993 (n1004, n962, n767, n968, n744);
or   g994 (n1031, n747, n753, n973, n727);
and  g995 (n988, n967, n973, n765, n764);
nand g996 (n1028, n769, n743, n972, n967);
and  g997 (n1033, n974, n965, n969);
xnor g998 (n1007, n757, n966, n726);
nor  g999 (n1032, n964, n729, n967, n762);
or   g1000 (n1011, n768, n758, n965, n971);
and  g1001 (n1051, n1002, n1006, n1000, n1014);
xor  g1002 (n1062, n1008, n1010, n981, n1001);
nor  g1003 (n1048, n986, n989, n978, n999);
and  g1004 (n1074, n988, n988, n997, n993);
nand g1005 (n1038, n982, n974, n978, n590);
xnor g1006 (n1043, n1006, n992, n991, n1008);
xnor g1007 (n1068, n994, n1007, n980, n1012);
and  g1008 (n1058, n1001, n979, n1013, n977);
nand g1009 (n1035, n588, n997, n1004, n1014);
or   g1010 (n1041, n998, n989, n975, n985);
and  g1011 (n1073, n1001, n589, n1005, n992);
and  g1012 (n1066, n1007, n1010, n974);
or   g1013 (n1075, n591, n1011, n987, n998);
or   g1014 (n1047, n1006, n996, n993, n1012);
and  g1015 (n1036, n775, n1002, n1009, n995);
xnor g1016 (n1069, n978, n995, n986, n1009);
and  g1017 (n1053, n1004, n985, n979);
xnor g1018 (n1061, n975, n994, n1011, n988);
or   g1019 (n1040, n981, n986, n980, n976);
xor  g1020 (n1072, n982, n1001, n992, n1000);
xnor g1021 (n1070, n1015, n987, n998, n995);
and  g1022 (n1037, n1013, n976, n990);
and  g1023 (n1055, n977, n1003, n975, n979);
xnor g1024 (n1059, n586, n992, n1003, n585);
and  g1025 (n1042, n983, n991, n1014, n977);
nand g1026 (n1063, n987, n1012, n1011, n980);
xor  g1027 (n1045, n978, n983, n1006, n1011);
xnor g1028 (n1049, n989, n1003, n991, n1005);
nor  g1029 (n1067, n1005, n985, n1010, n988);
xor  g1030 (n1034, n1007, n1014, n995, n990);
xnor g1031 (n1044, n1003, n996, n983, n998);
nand g1032 (n1064, n1008, n986, n981, n999);
xor  g1033 (n1060, n975, n982, n976, n1002);
xor  g1034 (n1057, n996, n987, n1000, n1005);
xor  g1035 (n1071, n982, n976, n1012, n1013);
xnor g1036 (n1054, n1002, n997, n1004, n1009);
nand g1037 (n1065, n999, n994, n587, n979);
and  g1038 (n1052, n994, n991, n977, n1004);
or   g1039 (n1039, n1009, n983, n997, n990);
xnor g1040 (n1046, n989, n993, n981, n1000);
or   g1041 (n1050, n1007, n980, n984, n993);
or   g1042 (n1056, n996, n1013, n999, n1008);
buf  g1043 (n1078, n1036);
not  g1044 (n1076, n778);
xor  g1045 (n1079, n1038, n779, n781, n777);
xnor g1046 (n1077, n780, n776, n1037, n1039);
buf  g1047 (n1088, n1016);
xor  g1048 (n1091, n790, n1079);
or   g1049 (n1089, n1078, n1076, n1077, n784);
and  g1050 (n1090, n788, n787, n1019, n1020);
or   g1051 (n1084, n1015, n1020, n783, n782);
nor  g1052 (n1083, n1018, n1079, n789, n1021);
or   g1053 (n1085, n797, n1040, n1021, n1016);
nor  g1054 (n1081, n1016, n1076, n1015, n1041);
nand g1055 (n1095, n1019, n1020, n793, n1079);
nor  g1056 (n1093, n796, n1018, n1017, n1077);
or   g1057 (n1094, n785, n1019, n1042, n1018);
xnor g1058 (n1086, n1078, n1078, n786, n794);
nand g1059 (n1087, n1077, n1019, n1017);
or   g1060 (n1092, n1017, n792, n1076, n1079);
xnor g1061 (n1080, n795, n1078, n1076, n1018);
nor  g1062 (n1082, n1020, n1015, n791, n1077);
buf  g1063 (n1099, n1080);
not  g1064 (n1097, n1082);
buf  g1065 (n1096, n1081);
not  g1066 (n1098, n1083);
not  g1067 (n1108, n1099);
buf  g1068 (n1109, n1098);
not  g1069 (n1105, n1097);
not  g1070 (n1107, n1099);
not  g1071 (n1110, n1098);
buf  g1072 (n1106, n1096);
not  g1073 (n1100, n1097);
not  g1074 (n1103, n1099);
not  g1075 (n1113, n1099);
buf  g1076 (n1111, n1097);
buf  g1077 (n1112, n1097);
buf  g1078 (n1101, n1096);
buf  g1079 (n1114, n1096);
buf  g1080 (n1115, n1098);
not  g1081 (n1104, n1096);
not  g1082 (n1102, n1098);
buf  g1083 (n1163, n1109);
buf  g1084 (n1161, n1066);
not  g1085 (n1154, n1059);
not  g1086 (n1176, n1108);
not  g1087 (n1178, n1111);
buf  g1088 (n1172, n1107);
not  g1089 (n1121, n802);
buf  g1090 (n1117, n808);
not  g1091 (n1139, n1061);
buf  g1092 (n1122, n1107);
buf  g1093 (n1137, n1101);
not  g1094 (n1157, n1055);
buf  g1095 (n1124, n1060);
not  g1096 (n1156, n1074);
not  g1097 (n1149, n799);
buf  g1098 (n1119, n1069);
not  g1099 (n1158, n1106);
not  g1100 (n1164, n1075);
buf  g1101 (n1116, n1109);
buf  g1102 (n1162, n1114);
not  g1103 (n1135, n1053);
buf  g1104 (n1118, n1073);
buf  g1105 (n1127, n811);
not  g1106 (n1142, n1113);
not  g1107 (n1171, n1113);
not  g1108 (n1175, n1114);
buf  g1109 (n1131, n1070);
not  g1110 (n1152, n1100);
not  g1111 (n1159, n1115);
not  g1112 (n1165, n1045);
not  g1113 (n1179, n1050);
not  g1114 (n1173, n804);
not  g1115 (n1169, n1108);
not  g1116 (n1170, n1047);
not  g1117 (n1174, n1115);
buf  g1118 (n1151, n1107);
buf  g1119 (n1148, n1101);
buf  g1120 (n1140, n809);
buf  g1121 (n1129, n1071);
not  g1122 (n1125, n1049);
buf  g1123 (n1130, n801);
buf  g1124 (n1155, n1057);
not  g1125 (n1143, n1063);
buf  g1126 (n1128, n1106);
not  g1127 (n1138, n1107);
not  g1128 (n1177, n810);
xor  g1129 (n1150, n1052, n1056, n816);
xor  g1130 (n1147, n1111, n1110, n1062, n813);
xor  g1131 (n1145, n1112, n1106, n1108, n1105);
nor  g1132 (n1153, n1072, n1113, n1104, n1048);
nor  g1133 (n1136, n1104, n1102, n815, n1100);
xor  g1134 (n1134, n1102, n1110, n1105, n1043);
xor  g1135 (n1141, n1067, n1111, n1064, n1100);
nand g1136 (n1126, n1108, n1112, n1109, n1101);
nand g1137 (n1120, n1044, n1113, n1101, n803);
or   g1138 (n1133, n1103, n1104, n1068, n1115);
xor  g1139 (n1166, n1103, n1110, n806, n1051);
or   g1140 (n1144, n798, n1103, n807, n1106);
or   g1141 (n1167, n1109, n1112, n812, n1114);
and  g1142 (n1168, n1105, n1046, n1054, n814);
nand g1143 (n1146, n1065, n1102, n805, n800);
nor  g1144 (n1132, n1115, n1103, n1111, n1105);
xnor g1145 (n1160, n1114, n1104, n1102, n1110);
or   g1146 (n1123, n817, n1100, n1112, n1058);
buf  g1147 (n1190, n1025);
buf  g1148 (n1227, n824);
buf  g1149 (n1246, n1128);
not  g1150 (n1216, n1175);
not  g1151 (n1245, n1170);
not  g1152 (n1192, n1169);
buf  g1153 (n1218, n1169);
not  g1154 (n1234, n822);
not  g1155 (n1211, n1174);
buf  g1156 (n1244, n1168);
buf  g1157 (n1237, n1029);
buf  g1158 (n1254, n1151);
buf  g1159 (n1180, n1119);
not  g1160 (n1213, n1024);
buf  g1161 (n1191, n1137);
not  g1162 (n1240, n1123);
buf  g1163 (n1224, n1126);
not  g1164 (n1184, n1025);
not  g1165 (n1195, n1023);
buf  g1166 (n1201, n821);
not  g1167 (n1206, n1134);
buf  g1168 (n1188, n1133);
not  g1169 (n1247, n1164);
buf  g1170 (n1231, n1027);
buf  g1171 (n1209, n1132);
buf  g1172 (n1223, n1136);
buf  g1173 (n1243, n1026);
buf  g1174 (n1225, n1140);
buf  g1175 (n1251, n1030);
not  g1176 (n1226, n1177);
not  g1177 (n1181, n1174);
buf  g1178 (n1239, n1120);
buf  g1179 (n1249, n1127);
not  g1180 (n1199, n1176);
not  g1181 (n1235, n1029);
buf  g1182 (n1241, n1118);
not  g1183 (n1242, n1149);
buf  g1184 (n1222, n1117);
buf  g1185 (n1250, n1028);
buf  g1186 (n1238, n1142);
not  g1187 (n1220, n1138);
buf  g1188 (n1210, n1158);
not  g1189 (n1230, n1139);
buf  g1190 (n1207, n1172);
buf  g1191 (n1186, n1178);
not  g1192 (n1200, n825);
not  g1193 (n1183, n1024);
not  g1194 (n1229, n1116);
buf  g1195 (n1204, n1165);
buf  g1196 (n1196, n1026);
buf  g1197 (n1233, n1173);
not  g1198 (n1185, n1179);
not  g1199 (n1253, n1026);
not  g1200 (n1208, n1157);
and  g1201 (n1217, n1159, n1161, n1153);
nor  g1202 (n1203, n1171, n1124, n1177);
xnor g1203 (n1212, n1024, n1028, n1027);
nor  g1204 (n1197, n1144, n1141, n1146);
or   g1205 (n1189, n1154, n818, n1022);
xor  g1206 (n1193, n819, n1122, n1025);
or   g1207 (n1255, n1029, n1028, n1022);
or   g1208 (n1205, n1030, n1029, n1145);
and  g1209 (n1214, n1030, n1170, n1176);
or   g1210 (n1232, n1130, n1023, n1152);
nor  g1211 (n1194, n1163, n1131, n1171);
xnor g1212 (n1182, n1155, n1026, n1028);
nand g1213 (n1256, n1166, n1156, n1021);
and  g1214 (n1198, n1023, n1135, n1178);
or   g1215 (n1202, n1160, n1121, n1025);
nand g1216 (n1215, n823, n1030, n1024);
nand g1217 (n1236, n820, n1027, n1168);
xnor g1218 (n1219, n1175, n1027, n1021);
or   g1219 (n1248, n1148, n1023, n1167);
nand g1220 (n1187, n1022, n1172, n1129);
nor  g1221 (n1228, n1173, n1022, n1125);
xor  g1222 (n1252, n1150, n1179, n1162);
and  g1223 (n1221, n1147, n1143, n1167);
not  g1224 (n1351, n1184);
buf  g1225 (n1265, n1243);
not  g1226 (n1347, n1091);
not  g1227 (n1417, n1215);
buf  g1228 (n1534, n1227);
buf  g1229 (n1546, n1205);
not  g1230 (n1562, n1092);
not  g1231 (n1276, n1187);
buf  g1232 (n1560, n1221);
buf  g1233 (n1271, n1216);
buf  g1234 (n1537, n1182);
not  g1235 (n1517, n1093);
buf  g1236 (n1559, n1182);
not  g1237 (n1521, n1203);
not  g1238 (n1413, n1202);
not  g1239 (n1399, n1217);
buf  g1240 (n1329, n1031);
not  g1241 (n1535, n1256);
not  g1242 (n1371, n1195);
buf  g1243 (n1311, n1214);
buf  g1244 (n1488, n1246);
not  g1245 (n1526, n1213);
not  g1246 (n1424, n1212);
buf  g1247 (n1389, n1252);
buf  g1248 (n1414, n1245);
not  g1249 (n1304, n1183);
not  g1250 (n1278, n1224);
buf  g1251 (n1490, n1223);
not  g1252 (n1392, n1092);
not  g1253 (n1268, n1089);
not  g1254 (n1477, n1239);
not  g1255 (n1492, n1189);
buf  g1256 (n1259, n1244);
buf  g1257 (n1307, n1231);
buf  g1258 (n1367, n1246);
buf  g1259 (n1461, n1199);
buf  g1260 (n1445, n1216);
buf  g1261 (n1544, n1090);
not  g1262 (n1495, n1252);
not  g1263 (n1470, n1201);
buf  g1264 (n1390, n1200);
not  g1265 (n1522, n1219);
not  g1266 (n1302, n1212);
not  g1267 (n1485, n1185);
not  g1268 (n1398, n1184);
buf  g1269 (n1527, n1186);
not  g1270 (n1549, n1212);
buf  g1271 (n1502, n1233);
not  g1272 (n1442, n1253);
buf  g1273 (n1403, n1199);
not  g1274 (n1496, n1240);
buf  g1275 (n1383, n1229);
not  g1276 (n1400, n1033);
buf  g1277 (n1558, n1194);
not  g1278 (n1459, n1192);
buf  g1279 (n1482, n1236);
not  g1280 (n1260, n1245);
not  g1281 (n1419, n1089);
not  g1282 (n1292, n1228);
not  g1283 (n1531, n1241);
buf  g1284 (n1375, n1206);
not  g1285 (n1282, n1252);
buf  g1286 (n1530, n1237);
buf  g1287 (n1323, n1213);
not  g1288 (n1291, n1227);
buf  g1289 (n1491, n1189);
buf  g1290 (n1473, n1238);
buf  g1291 (n1415, n1210);
not  g1292 (n1339, n1186);
not  g1293 (n1324, n1212);
buf  g1294 (n1368, n1185);
not  g1295 (n1464, n1196);
not  g1296 (n1303, n1092);
buf  g1297 (n1543, n1250);
not  g1298 (n1499, n1090);
not  g1299 (n1360, n1180);
not  g1300 (n1258, n1234);
not  g1301 (n1377, n1226);
not  g1302 (n1466, n1094);
not  g1303 (n1447, n1187);
buf  g1304 (n1452, n1254);
not  g1305 (n1538, n1088);
buf  g1306 (n1474, n1253);
buf  g1307 (n1518, n1238);
buf  g1308 (n1336, n1086);
not  g1309 (n1362, n1243);
not  g1310 (n1536, n1219);
not  g1311 (n1489, n1202);
not  g1312 (n1355, n1085);
not  g1313 (n1410, n1237);
not  g1314 (n1366, n1229);
buf  g1315 (n1273, n1181);
not  g1316 (n1457, n1197);
buf  g1317 (n1342, n1198);
not  g1318 (n1372, n1195);
buf  g1319 (n1272, n1095);
buf  g1320 (n1553, n826);
buf  g1321 (n1333, n1240);
not  g1322 (n1402, n1204);
buf  g1323 (n1523, n1244);
buf  g1324 (n1280, n1191);
buf  g1325 (n1545, n1204);
not  g1326 (n1467, n1207);
buf  g1327 (n1564, n1221);
buf  g1328 (n1369, n1254);
not  g1329 (n1483, n1247);
not  g1330 (n1263, n1032);
buf  g1331 (n1386, n1213);
buf  g1332 (n1438, n1090);
buf  g1333 (n1328, n1191);
buf  g1334 (n1327, n1256);
not  g1335 (n1346, n1249);
not  g1336 (n1556, n1213);
buf  g1337 (n1266, n1200);
buf  g1338 (n1451, n1214);
buf  g1339 (n1388, n1188);
not  g1340 (n1465, n1206);
buf  g1341 (n1541, n1182);
not  g1342 (n1349, n1229);
buf  g1343 (n1500, n1191);
buf  g1344 (n1335, n1248);
buf  g1345 (n1296, n1221);
not  g1346 (n1270, n1245);
not  g1347 (n1279, n1185);
buf  g1348 (n1503, n1189);
buf  g1349 (n1281, n1232);
not  g1350 (n1441, n1226);
buf  g1351 (n1365, n1201);
buf  g1352 (n1345, n1199);
not  g1353 (n1520, n1180);
not  g1354 (n1338, n1187);
not  g1355 (n1401, n1241);
not  g1356 (n1509, n1207);
not  g1357 (n1421, n1232);
not  g1358 (n1325, n1237);
not  g1359 (n1449, n1248);
buf  g1360 (n1439, n1215);
buf  g1361 (n1533, n1215);
not  g1362 (n1540, n1233);
not  g1363 (n1411, n1235);
not  g1364 (n1408, n1234);
buf  g1365 (n1486, n1206);
not  g1366 (n1370, n1222);
not  g1367 (n1440, n1244);
not  g1368 (n1397, n1235);
not  g1369 (n1340, n1246);
buf  g1370 (n1454, n1253);
not  g1371 (n1288, n1190);
buf  g1372 (n1548, n1230);
buf  g1373 (n1469, n1095);
not  g1374 (n1409, n1215);
not  g1375 (n1284, n1245);
not  g1376 (n1275, n1190);
buf  g1377 (n1498, n1218);
buf  g1378 (n1379, n1242);
not  g1379 (n1404, n1190);
not  g1380 (n1354, n1225);
not  g1381 (n1396, n1255);
buf  g1382 (n1374, n1187);
not  g1383 (n1310, n828);
buf  g1384 (n1315, n1249);
not  g1385 (n1317, n1209);
buf  g1386 (n1332, n1236);
buf  g1387 (n1460, n1234);
buf  g1388 (n1269, n1198);
buf  g1389 (n1446, n1239);
buf  g1390 (n1437, n1197);
not  g1391 (n1394, n1033);
not  g1392 (n1391, n1192);
not  g1393 (n1519, n1247);
not  g1394 (n1289, n1220);
buf  g1395 (n1429, n1207);
buf  g1396 (n1384, n1254);
buf  g1397 (n1287, n1180);
buf  g1398 (n1352, n1188);
buf  g1399 (n1475, n1224);
buf  g1400 (n1443, n1094);
buf  g1401 (n1395, n1249);
not  g1402 (n1453, n1203);
not  g1403 (n1416, n1220);
buf  g1404 (n1381, n1227);
buf  g1405 (n1434, n1250);
buf  g1406 (n1293, n1225);
buf  g1407 (n1277, n1243);
not  g1408 (n1331, n1214);
buf  g1409 (n1285, n1235);
buf  g1410 (n1380, n1194);
not  g1411 (n1484, n1194);
buf  g1412 (n1343, n1236);
not  g1413 (n1539, n1183);
buf  g1414 (n1450, n1197);
not  g1415 (n1322, n1095);
not  g1416 (n1330, n1093);
buf  g1417 (n1478, n1211);
not  g1418 (n1510, n1188);
not  g1419 (n1418, n1031);
not  g1420 (n1507, n1205);
buf  g1421 (n1525, n1216);
buf  g1422 (n1373, n1197);
not  g1423 (n1427, n1180);
buf  g1424 (n1309, n1196);
not  g1425 (n1480, n1238);
buf  g1426 (n1295, n1252);
not  g1427 (n1358, n1204);
not  g1428 (n1514, n1089);
buf  g1429 (n1341, n1235);
buf  g1430 (n1456, n1193);
buf  g1431 (n1513, n1200);
buf  g1432 (n1363, n1087);
not  g1433 (n1528, n1230);
buf  g1434 (n1353, n1241);
buf  g1435 (n1298, n1203);
not  g1436 (n1504, n829);
not  g1437 (n1356, n1243);
not  g1438 (n1542, n1251);
buf  g1439 (n1448, n1211);
not  g1440 (n1344, n1226);
buf  g1441 (n1359, n1223);
not  g1442 (n1364, n1227);
buf  g1443 (n1497, n1218);
buf  g1444 (n1547, n1242);
buf  g1445 (n1301, n1208);
not  g1446 (n1436, n1199);
not  g1447 (n1426, n1233);
buf  g1448 (n1493, n1203);
buf  g1449 (n1382, n1186);
not  g1450 (n1348, n1225);
not  g1451 (n1501, n1196);
not  g1452 (n1506, n1201);
buf  g1453 (n1290, n1189);
buf  g1454 (n1468, n1247);
not  g1455 (n1378, n1248);
not  g1456 (n1308, n1210);
buf  g1457 (n1387, n1186);
not  g1458 (n1274, n1208);
not  g1459 (n1350, n1088);
not  g1460 (n1508, n1032);
not  g1461 (n1334, n1250);
buf  g1462 (n1283, n1207);
not  g1463 (n1524, n1225);
buf  g1464 (n1420, n1087);
not  g1465 (n1430, n1089);
not  g1466 (n1405, n1032);
buf  g1467 (n1512, n1239);
not  g1468 (n1425, n1248);
not  g1469 (n1312, n1200);
not  g1470 (n1264, n1239);
buf  g1471 (n1479, n1234);
not  g1472 (n1433, n1088);
not  g1473 (n1494, n1221);
buf  g1474 (n1529, n1211);
not  g1475 (n1423, n1206);
not  g1476 (n1516, n1210);
buf  g1477 (n1376, n1222);
not  g1478 (n1505, n1222);
buf  g1479 (n1257, n1233);
not  g1480 (n1294, n1208);
not  g1481 (n1435, n1184);
buf  g1482 (n1431, n1093);
buf  g1483 (n1321, n1181);
not  g1484 (n1472, n1244);
buf  g1485 (n1550, n1214);
buf  g1486 (n1552, n1241);
buf  g1487 (n1305, n827);
not  g1488 (n1455, n1185);
not  g1489 (n1297, n1224);
buf  g1490 (n1393, n1217);
not  g1491 (n1481, n1217);
buf  g1492 (n1511, n1188);
not  g1493 (n1563, n1198);
not  g1494 (n1267, n1222);
buf  g1495 (n1412, n1230);
not  g1496 (n1561, n1183);
buf  g1497 (n1471, n1231);
buf  g1498 (n1361, n1251);
buf  g1499 (n1314, n1211);
not  g1500 (n1337, n1255);
buf  g1501 (n1326, n1093);
not  g1502 (n1318, n1192);
not  g1503 (n1428, n1181);
buf  g1504 (n1407, n1190);
not  g1505 (n1406, n1193);
not  g1506 (n1313, n1242);
not  g1507 (n1532, n1095);
not  g1508 (n1487, n1192);
not  g1509 (n1320, n1228);
not  g1510 (n1444, n1209);
not  g1511 (n1385, n1228);
buf  g1512 (n1463, n1087);
and  g1513 (n1299, n1208, n1092);
or   g1514 (n1300, n1033, n1255, n1205, n1236);
or   g1515 (n1261, n1250, n1196, n1084, n1224);
xor  g1516 (n1422, n1094, n1219, n1242);
nand g1517 (n1554, n1232, n1246, n1091, n1240);
or   g1518 (n1316, n1229, n1220, n1210, n1183);
nand g1519 (n1306, n1088, n1247, n1216, n1094);
nor  g1520 (n1319, n1220, n1031, n1255, n1209);
nor  g1521 (n1555, n1240, n1218, n1228, n1195);
or   g1522 (n1551, n1201, n1249, n1091, n1223);
nand g1523 (n1286, n1256, n1031, n1209, n1230);
and  g1524 (n1476, n1198, n1087, n1204, n1251);
nor  g1525 (n1557, n1194, n1205, n1202, n1253);
nand g1526 (n1462, n1217, n1193, n1091, n1251);
xor  g1527 (n1262, n1090, n1237, n1182, n1032);
xor  g1528 (n1357, n1223, n1256, n1184, n1033);
xnor g1529 (n1432, n1181, n1193, n1254, n1226);
and  g1530 (n1515, n1218, n1238, n1231);
and  g1531 (n1458, n1195, n1191, n1202, n1232);
not  g1532 (n1645, n1472);
not  g1533 (n1737, n1507);
not  g1534 (n1649, n1312);
not  g1535 (n1621, n1259);
buf  g1536 (n1816, n1485);
not  g1537 (n1594, n1307);
not  g1538 (n1579, n1509);
buf  g1539 (n1712, n1355);
buf  g1540 (n1730, n1359);
buf  g1541 (n1828, n1379);
buf  g1542 (n1731, n1477);
not  g1543 (n1820, n1428);
buf  g1544 (n1804, n1384);
not  g1545 (n1679, n1419);
buf  g1546 (n1698, n1516);
not  g1547 (n1700, n1383);
not  g1548 (n1636, n1293);
not  g1549 (n1702, n1394);
buf  g1550 (n1654, n1513);
not  g1551 (n1843, n1290);
not  g1552 (n1623, n1381);
buf  g1553 (n1622, n1413);
not  g1554 (n1755, n1340);
not  g1555 (n1761, n1382);
not  g1556 (n1681, n1471);
buf  g1557 (n1682, n1469);
not  g1558 (n1817, n1323);
not  g1559 (n1687, n1498);
not  g1560 (n1769, n1511);
buf  g1561 (n1609, n1508);
not  g1562 (n1600, n1273);
not  g1563 (n1741, n1346);
buf  g1564 (n1632, n839);
not  g1565 (n1604, n1459);
not  g1566 (n1775, n1352);
buf  g1567 (n1661, n1350);
not  g1568 (n1836, n1351);
not  g1569 (n1619, n1427);
not  g1570 (n1629, n1455);
buf  g1571 (n1767, n1305);
not  g1572 (n1710, n1389);
not  g1573 (n1568, n1461);
buf  g1574 (n1720, n838);
buf  g1575 (n1806, n1429);
not  g1576 (n1764, n831);
not  g1577 (n1652, n1300);
not  g1578 (n1567, n1466);
buf  g1579 (n1813, n1411);
not  g1580 (n1736, n833);
buf  g1581 (n1718, n1424);
buf  g1582 (n1824, n1500);
not  g1583 (n1822, n1366);
not  g1584 (n1840, n1354);
not  g1585 (n1848, n1341);
not  g1586 (n1653, n1514);
not  g1587 (n1626, n1304);
buf  g1588 (n1795, n1326);
not  g1589 (n1798, n1270);
buf  g1590 (n1808, n1422);
not  g1591 (n1605, n1322);
not  g1592 (n1655, n1298);
not  g1593 (n1639, n1264);
not  g1594 (n1677, n1439);
not  g1595 (n1777, n1452);
not  g1596 (n1608, n1515);
not  g1597 (n1762, n1473);
not  g1598 (n1722, n1414);
buf  g1599 (n1650, n1514);
not  g1600 (n1829, n1296);
buf  g1601 (n1792, n1283);
not  g1602 (n1750, n1506);
not  g1603 (n1791, n1479);
buf  g1604 (n1754, n1368);
buf  g1605 (n1625, n1504);
not  g1606 (n1749, n1316);
not  g1607 (n1664, n1332);
not  g1608 (n1672, n1313);
buf  g1609 (n1656, n1391);
not  g1610 (n1815, n1501);
buf  g1611 (n1714, n1276);
not  g1612 (n1756, n1513);
buf  g1613 (n1760, n1421);
buf  g1614 (n1703, n1328);
buf  g1615 (n1646, n1345);
buf  g1616 (n1685, n1361);
not  g1617 (n1582, n1438);
buf  g1618 (n1739, n1436);
not  g1619 (n1787, n1426);
buf  g1620 (n1577, n1433);
not  g1621 (n1724, n1430);
buf  g1622 (n1591, n1462);
buf  g1623 (n1837, n1321);
not  g1624 (n1690, n1288);
not  g1625 (n1835, n1501);
not  g1626 (n1606, n1364);
buf  g1627 (n1706, n1498);
not  g1628 (n1805, n1263);
buf  g1629 (n1595, n1510);
not  g1630 (n1638, n1487);
not  g1631 (n1721, n1517);
not  g1632 (n1707, n1417);
buf  g1633 (n1733, n1301);
buf  g1634 (n1847, n1286);
not  g1635 (n1734, n1339);
buf  g1636 (n1744, n1490);
buf  g1637 (n1635, n1274);
buf  g1638 (n1607, n1310);
not  g1639 (n1785, n1465);
not  g1640 (n1746, n1376);
buf  g1641 (n1779, n1437);
not  g1642 (n1716, n1358);
buf  g1643 (n1642, n1517);
buf  g1644 (n1678, n1292);
not  g1645 (n1797, n1375);
not  g1646 (n1573, n1458);
not  g1647 (n1788, n1509);
not  g1648 (n1599, n836);
buf  g1649 (n1647, n1484);
not  g1650 (n1615, n1454);
buf  g1651 (n1659, n1453);
not  g1652 (n1651, n1299);
not  g1653 (n1711, n1447);
not  g1654 (n1570, n1360);
buf  g1655 (n1832, n1343);
not  g1656 (n1772, n1491);
not  g1657 (n1657, n1499);
buf  g1658 (n1589, n1262);
not  g1659 (n1633, n1496);
buf  g1660 (n1793, n1518);
buf  g1661 (n1598, n1444);
not  g1662 (n1807, n1372);
not  g1663 (n1794, n1367);
buf  g1664 (n1644, n1400);
buf  g1665 (n1827, n1327);
buf  g1666 (n1770, n1395);
not  g1667 (n1766, n1333);
buf  g1668 (n1705, n1277);
not  g1669 (n1812, n835);
not  g1670 (n1694, n1309);
not  g1671 (n1727, n1502);
buf  g1672 (n1819, n1441);
buf  g1673 (n1774, n1324);
not  g1674 (n1715, n1377);
buf  g1675 (n1743, n832);
buf  g1676 (n1838, n1482);
not  g1677 (n1631, n1331);
not  g1678 (n1686, n1335);
buf  g1679 (n1809, n1480);
buf  g1680 (n1680, n1319);
not  g1681 (n1637, n1435);
buf  g1682 (n1616, n1289);
not  g1683 (n1666, n1317);
buf  g1684 (n1611, n1415);
not  g1685 (n1839, n1378);
not  g1686 (n1610, n1420);
buf  g1687 (n1796, n1409);
not  g1688 (n1596, n1334);
buf  g1689 (n1811, n1291);
buf  g1690 (n1784, n837);
not  g1691 (n1586, n1260);
not  g1692 (n1576, n1418);
not  g1693 (n1778, n1311);
not  g1694 (n1726, n1468);
buf  g1695 (n1783, n1503);
not  g1696 (n1683, n1392);
not  g1697 (n1768, n1515);
buf  g1698 (n1660, n1497);
buf  g1699 (n1574, n1365);
buf  g1700 (n1663, n1385);
buf  g1701 (n1738, n1257);
not  g1702 (n1713, n1295);
buf  g1703 (n1575, n1464);
not  g1704 (n1691, n1388);
buf  g1705 (n1693, n1369);
buf  g1706 (n1701, n1280);
not  g1707 (n1799, n1315);
not  g1708 (n1845, n1393);
buf  g1709 (n1849, n1373);
not  g1710 (n1790, n1338);
not  g1711 (n1640, n1267);
not  g1712 (n1833, n1460);
buf  g1713 (n1617, n1488);
buf  g1714 (n1588, n1478);
not  g1715 (n1803, n1470);
not  g1716 (n1627, n1272);
buf  g1717 (n1800, n1399);
not  g1718 (n1723, n1398);
not  g1719 (n1593, n1320);
buf  g1720 (n1628, n1318);
buf  g1721 (n1821, n1329);
not  g1722 (n1587, n1505);
buf  g1723 (n1745, n1261);
not  g1724 (n1771, n1281);
buf  g1725 (n1844, n1390);
buf  g1726 (n1668, n1440);
buf  g1727 (n1748, n1463);
buf  g1728 (n1758, n1476);
buf  g1729 (n1602, n1407);
not  g1730 (n1665, n1431);
not  g1731 (n1842, n1297);
buf  g1732 (n1565, n1287);
not  g1733 (n1620, n1496);
buf  g1734 (n1671, n1505);
buf  g1735 (n1614, n1502);
not  g1736 (n1584, n1475);
buf  g1737 (n1825, n1412);
buf  g1738 (n1773, n1467);
not  g1739 (n1566, n1405);
not  g1740 (n1592, n830);
not  g1741 (n1572, n1337);
buf  g1742 (n1674, n1284);
not  g1743 (n1676, n1474);
not  g1744 (n1728, n1493);
buf  g1745 (n1673, n1344);
not  g1746 (n1846, n1396);
buf  g1747 (n1675, n1483);
buf  g1748 (n1747, n1265);
not  g1749 (n1776, n1397);
buf  g1750 (n1752, n1269);
buf  g1751 (n1603, n1357);
buf  g1752 (n1740, n1353);
buf  g1753 (n1782, n1499);
buf  g1754 (n1709, n834);
not  g1755 (n1597, n1374);
not  g1756 (n1802, n1503);
buf  g1757 (n1688, n1275);
buf  g1758 (n1830, n1268);
not  g1759 (n1814, n1348);
not  g1760 (n1634, n1278);
not  g1761 (n1630, n1282);
buf  g1762 (n1669, n1442);
buf  g1763 (n1751, n1512);
not  g1764 (n1753, n1303);
buf  g1765 (n1667, n1402);
buf  g1766 (n1571, n1443);
not  g1767 (n1658, n1495);
not  g1768 (n1581, n1342);
not  g1769 (n1708, n1457);
buf  g1770 (n1624, n1266);
buf  g1771 (n1696, n1271);
not  g1772 (n1834, n1404);
not  g1773 (n1725, n1449);
not  g1774 (n1735, n1508);
buf  g1775 (n1670, n1371);
not  g1776 (n1612, n1362);
not  g1777 (n1601, n1425);
buf  g1778 (n1643, n1294);
buf  g1779 (n1826, n1349);
buf  g1780 (n1692, n1279);
buf  g1781 (n1590, n1451);
buf  g1782 (n1719, n1347);
buf  g1783 (n1662, n1423);
buf  g1784 (n1818, n1336);
buf  g1785 (n1569, n1387);
buf  g1786 (n1580, n1356);
buf  g1787 (n1763, n1330);
buf  g1788 (n1583, n1306);
not  g1789 (n1789, n1386);
not  g1790 (n1695, n1445);
not  g1791 (n1831, n1302);
buf  g1792 (n1841, n1308);
buf  g1793 (n1648, n1504);
not  g1794 (n1717, n1506);
buf  g1795 (n1585, n1456);
buf  g1796 (n1618, n1408);
buf  g1797 (n1613, n1450);
not  g1798 (n1729, n1494);
not  g1799 (n1732, n1416);
not  g1800 (n1786, n1448);
buf  g1801 (n1697, n1511);
not  g1802 (n1757, n1370);
not  g1803 (n1781, n1481);
buf  g1804 (n1742, n1486);
buf  g1805 (n1801, n1363);
buf  g1806 (n1689, n1518);
buf  g1807 (n1578, n1325);
buf  g1808 (n1810, n1446);
buf  g1809 (n1765, n1403);
buf  g1810 (n1759, n1410);
not  g1811 (n1704, n1500);
buf  g1812 (n1641, n1258);
nor  g1813 (n1699, n1497, n1314);
or   g1814 (n1823, n1401, n1432, n1492, n1516);
xor  g1815 (n1684, n1434, n1512, n1285, n1380);
nor  g1816 (n1780, n1489, n1406, n1507, n1510);
nand g1817 (n1868, n1565, n1546, n1531, n1556);
and  g1818 (n1867, n1555, n1545, n1527, n1534);
and  g1819 (n1859, n1563, n1527, n1529, n1562);
and  g1820 (n1862, n1544, n1601, n1547, n1572);
nor  g1821 (n1871, n1576, n1549, n1519, n1534);
or   g1822 (n1882, n1598, n1540, n1589, n1561);
nor  g1823 (n1850, n1525, n1522, n1564, n1550);
or   g1824 (n1866, n1548, n1526, n1539, n1558);
and  g1825 (n1851, n1543, n1536, n1551, n1559);
or   g1826 (n1881, n1520, n1550, n1557, n1600);
or   g1827 (n1865, n1569, n841, n1563, n1523);
and  g1828 (n1880, n1592, n1547, n1566, n1539);
and  g1829 (n1876, n1593, n1586, n1528, n1555);
xor  g1830 (n1852, n1519, n1524, n1560, n1591);
xor  g1831 (n1853, n1583, n1523, n1554, n1521);
or   g1832 (n1856, n1579, n1532, n1548, n1526);
nor  g1833 (n1858, n1538, n1549, n1567, n1546);
or   g1834 (n1874, n1522, n1573, n1562, n1528);
and  g1835 (n1857, n1584, n1552, n1544, n1560);
xor  g1836 (n1863, n1541, n1533, n1596, n1531);
xnor g1837 (n1878, n1538, n1568, n1578, n1597);
nand g1838 (n1870, n1552, n1558, n1540, n1542);
xor  g1839 (n1854, n1587, n1577, n1532, n1554);
nor  g1840 (n1864, n1556, n1525, n1542, n1588);
xnor g1841 (n1872, n1571, n1543, n1529, n1585);
xnor g1842 (n1869, n1530, n1590, n1581, n1524);
xnor g1843 (n1873, n1553, n1533, n1530, n1574);
nor  g1844 (n1855, n1535, n1521, n1561, n1564);
or   g1845 (n1879, n1551, n1545, n1570, n1537);
xor  g1846 (n1861, n1537, n1541, n842, n1520);
and  g1847 (n1860, n1559, n1594, n1535, n840);
and  g1848 (n1877, n1575, n1582, n1536, n1557);
nor  g1849 (n1875, n1595, n1599, n1580, n1553);
xor  g1850 (n1899, n856, n1636, n848, n1668);
or   g1851 (n1903, n844, n1618, n1651, n1670);
nand g1852 (n1914, n1684, n1851, n1661, n1641);
nand g1853 (n1883, n1624, n852, n1676, n1867);
xor  g1854 (n1904, n1626, n1650, n1666, n1652);
and  g1855 (n1888, n1631, n1629, n1603, n1663);
and  g1856 (n1894, n1667, n1678, n1665, n1680);
nor  g1857 (n1887, n1644, n1672, n1604, n1874);
xor  g1858 (n1892, n1632, n1669, n857, n1860);
and  g1859 (n1905, n1648, n1616, n1662, n1862);
and  g1860 (n1900, n1611, n1628, n1683, n1637);
or   g1861 (n1910, n1674, n1645, n1621, n1612);
or   g1862 (n1913, n846, n1659, n1646, n1614);
and  g1863 (n1891, n1878, n1877, n853, n1639);
or   g1864 (n1897, n1864, n1605, n1620, n1615);
and  g1865 (n1884, n1607, n1859, n1857, n1660);
or   g1866 (n1890, n1868, n1664, n1872, n1633);
nand g1867 (n1885, n1619, n1634, n847, n1870);
nand g1868 (n1909, n1609, n1643, n1630, n1653);
or   g1869 (n1886, n1871, n1649, n1856, n1855);
or   g1870 (n1893, n1606, n1866, n850, n1865);
or   g1871 (n1911, n1854, n849, n851, n1640);
xnor g1872 (n1915, n1617, n1681, n1602, n1858);
nor  g1873 (n1896, n1677, n1682, n1608, n1873);
or   g1874 (n1907, n1625, n1679, n1879, n1623);
or   g1875 (n1895, n1655, n1622, n1673, n858);
nor  g1876 (n1898, n843, n1642, n1853, n1613);
xor  g1877 (n1901, n1657, n1880, n1869, n854);
nor  g1878 (n1912, n1658, n1861, n1863, n1876);
and  g1879 (n1902, n1627, n1647, n1850, n1881);
or   g1880 (n1908, n1675, n1671, n1875, n1654);
or   g1881 (n1889, n1610, n845, n1638, n1635);
xor  g1882 (n1906, n1852, n1656, n855, n1882);
xor  g1883 (n1962, n1815, n1733, n1801, n1914);
or   g1884 (n1922, n1808, n1911, n1766, n1915);
xnor g1885 (n1970, n1763, n1845, n1883, n1848);
nor  g1886 (n1943, n1823, n1755, n1915, n1890);
nor  g1887 (n1959, n1903, n1703, n1701, n1782);
or   g1888 (n1949, n1836, n1906, n1786, n1696);
nor  g1889 (n1920, n1728, n1826, n1803, n1912);
xor  g1890 (n1960, n1788, n1685, n1746, n1888);
xor  g1891 (n1952, n1821, n1840, n1694, n1708);
nand g1892 (n1946, n1912, n1812, n1764, n1749);
nor  g1893 (n1929, n1712, n1887, n1898, n1839);
nor  g1894 (n1945, n1720, n1910, n1734, n1715);
and  g1895 (n1917, n1834, n1906, n1779, n1907);
nand g1896 (n1936, n1692, n1790, n1783, n1741);
xnor g1897 (n1916, n1902, n1742, n1835, n1752);
nand g1898 (n1925, n1698, n1817, n1841, n1705);
nor  g1899 (n1933, n1737, n1828, n1898, n1699);
and  g1900 (n1935, n1904, n1736, n1909, n1702);
or   g1901 (n1944, n1690, n1789, n1796, n1908);
xnor g1902 (n1967, n1889, n1785, n1787, n1884);
and  g1903 (n1931, n1740, n1802, n1748, n1793);
or   g1904 (n1941, n1822, n1791, n1739, n1724);
or   g1905 (n1924, n1804, n1846, n1833, n1885);
xnor g1906 (n1923, n1757, n1732, n1907, n1908);
xor  g1907 (n1955, n1813, n1723, n1894, n1776);
and  g1908 (n1937, n1896, n1816, n1899, n1838);
or   g1909 (n1953, n1716, n1767, n1847, n1758);
or   g1910 (n1940, n1792, n1735, n1901, n1807);
xor  g1911 (n1948, n1704, n1795, n1814, n1777);
nor  g1912 (n1966, n1778, n1827, n1711, n1831);
xnor g1913 (n1954, n1905, n1754, n1902, n1909);
and  g1914 (n1932, n1904, n1900, n1718, n1818);
xor  g1915 (n1942, n1829, n1709, n1892, n1805);
nand g1916 (n1958, n1913, n1900, n1714, n1775);
or   g1917 (n1934, n1780, n1731, n1768, n1842);
nor  g1918 (n1918, n1717, n1891, n1726, n1799);
or   g1919 (n1930, n1914, n1781, n1722, n1738);
or   g1920 (n1961, n1769, n1830, n1751, n1825);
nand g1921 (n1947, n1761, n1773, n1695, n1800);
and  g1922 (n1938, n1913, n1798, n1905, n1771);
and  g1923 (n1957, n1914, n1697, n1837, n1910);
xor  g1924 (n1964, n1725, n1730, n1819, n1901);
xnor g1925 (n1939, n1688, n1832, n1843, n1750);
xnor g1926 (n1956, n1721, n1765, n1753, n1747);
nor  g1927 (n1968, n1756, n1707, n1744, n1810);
nor  g1928 (n1965, n1844, n1691, n1745, n1686);
and  g1929 (n1963, n1762, n1719, n1784, n1759);
xor  g1930 (n1921, n1897, n1820, n1774, n1915);
nor  g1931 (n1919, n1914, n1794, n1700, n1809);
and  g1932 (n1928, n1729, n1743, n1903, n1893);
xor  g1933 (n1927, n1689, n1899, n1797, n1886);
xnor g1934 (n1950, n1710, n1895, n1706, n1760);
nand g1935 (n1926, n1911, n1806, n1687, n1770);
or   g1936 (n1951, n1824, n1693, n1727, n1772);
and  g1937 (n1969, n1713, n1811, n1915, n1849);
xor  g1938 (n1999, n619, n1950, n1952, n610);
and  g1939 (n1996, n1958, n1967, n609, n594);
nor  g1940 (n1989, n1919, n607, n1924, n614);
nand g1941 (n1997, n600, n1933, n645, n1941);
and  g1942 (n1982, n625, n629, n1943, n664);
xnor g1943 (n1976, n1963, n627, n1937, n1938);
and  g1944 (n1995, n640, n646, n1931, n633);
nor  g1945 (n2000, n1921, n595, n1929, n1939);
xor  g1946 (n1974, n620, n636, n606, n653);
xor  g1947 (n1985, n616, n1957, n654, n596);
nand g1948 (n1987, n1944, n32, n662, n650);
or   g1949 (n1980, n1970, n651, n644, n1923);
and  g1950 (n1984, n624, n1916, n603, n1936);
xnor g1951 (n1994, n643, n638, n1966, n660);
xnor g1952 (n2002, n1918, n648, n1925, n1965);
xor  g1953 (n1977, n647, n666, n604, n1951);
xnor g1954 (n1990, n621, n626, n659, n1917);
nand g1955 (n2003, n658, n599, n1947, n1945);
xor  g1956 (n1972, n1964, n1935, n593, n1946);
xor  g1957 (n1998, n613, n641, n1959, n649);
xor  g1958 (n1971, n635, n661, n1920, n657);
xor  g1959 (n1979, n1961, n622, n612, n615);
nor  g1960 (n1993, n665, n628, n1940, n1922);
nor  g1961 (n1986, n598, n597, n637, n1969);
and  g1962 (n1983, n631, n634, n642, n1934);
or   g1963 (n1988, n1955, n611, n617, n592);
xnor g1964 (n1973, n1928, n656, n667, n1932);
nor  g1965 (n1992, n1968, n602, n1953, n1948);
and  g1966 (n1981, n655, n1956, n1930, n623);
xor  g1967 (n1975, n608, n605, n618, n601);
nand g1968 (n1991, n1942, n652, n630, n639);
nor  g1969 (n1978, n1954, n663, n1949, n632);
or   g1970 (n2001, n1962, n1960, n1926, n1927);
xnor g1971 (n2031, n1975, n907, n1992, n865);
nor  g1972 (n2032, n1997, n872, n881, n890);
xor  g1973 (n2030, n935, n884, n936, n912);
or   g1974 (n2017, n877, n930, n913, n2000);
nand g1975 (n2005, n908, n901, n1974, n889);
or   g1976 (n2029, n900, n1993, n1988, n920);
xor  g1977 (n2007, n906, n923, n904, n905);
and  g1978 (n2015, n1979, n1973, n859, n1972);
and  g1979 (n2016, n863, n934, n917, n1978);
nand g1980 (n2014, n869, n880, n927, n887);
xnor g1981 (n2028, n2001, n914, n916, n878);
or   g1982 (n2006, n883, n2003, n860, n1991);
xnor g1983 (n2023, n866, n938, n895, n2002);
and  g1984 (n2004, n888, n915, n903, n876);
xnor g1985 (n2010, n911, n861, n862, n1986);
xnor g1986 (n2025, n932, n931, n870, n886);
or   g1987 (n2026, n873, n924, n897, n1984);
or   g1988 (n2008, n885, n871, n1995, n882);
or   g1989 (n2012, n1999, n933, n902, n1983);
xnor g1990 (n2009, n898, n925, n1971, n910);
or   g1991 (n2018, n893, n896, n939, n1976);
xor  g1992 (n2011, n918, n879, n891, n1990);
nor  g1993 (n2027, n868, n1994, n937, n921);
xnor g1994 (n2013, n1985, n864, n875, n922);
and  g1995 (n2024, n892, n1982, n909, n940);
xnor g1996 (n2021, n1998, n919, n899, n928);
xnor g1997 (n2022, n1980, n940, n867, n1981);
and  g1998 (n2019, n926, n894, n1987, n1996);
xor  g1999 (n2020, n929, n874, n1977, n1989);
endmodule
