

module Stat_100_63
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n43,
  n115,
  n88,
  n103,
  n96,
  n97,
  n80,
  n100,
  n66,
  n77,
  n102,
  n75,
  n65,
  n111,
  n78,
  n95,
  n82,
  n106,
  n129,
  n123,
  n121,
  n119,
  n124,
  n125,
  n120,
  n122,
  n127,
  n126,
  n128,
  n132,
  n131,
  n130,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n43;output n115;output n88;output n103;output n96;output n97;output n80;output n100;output n66;output n77;output n102;output n75;output n65;output n111;output n78;output n95;output n82;output n106;output n129;output n123;output n121;output n119;output n124;output n125;output n120;output n122;output n127;output n126;output n128;output n132;output n131;output n130;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n76;wire n79;wire n81;wire n83;wire n84;wire n85;wire n86;wire n87;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n98;wire n99;wire n101;wire n104;wire n105;wire n107;wire n108;wire n109;wire n110;wire n112;wire n113;wire n114;wire n116;wire n117;wire n118;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  not
  g0
  (
    n35,
    n1
  );


  buf
  g1
  (
    n36,
    n2
  );


  buf
  g2
  (
    KeyWire_0_7,
    n1
  );


  not
  g3
  (
    n37,
    n1
  );


  buf
  g4
  (
    n38,
    n1
  );


  not
  g5
  (
    n34,
    n2
  );


  not
  g6
  (
    n40,
    n37
  );


  not
  g7
  (
    n41,
    n37
  );


  buf
  g8
  (
    KeyWire_0_14,
    n2
  );


  buf
  g9
  (
    KeyWire_0_27,
    n3
  );


  nand
  g10
  (
    n39,
    n2,
    n36
  );


  not
  g11
  (
    KeyWire_0_16,
    n43
  );


  buf
  g12
  (
    n46,
    n40
  );


  buf
  g13
  (
    n47,
    n41
  );


  not
  g14
  (
    KeyWire_0_3,
    n42
  );


  buf
  g15
  (
    KeyWire_0_19,
    n44
  );


  buf
  g16
  (
    n58,
    n44
  );


  buf
  g17
  (
    n59,
    n4
  );


  not
  g18
  (
    KeyWire_0_22,
    n5
  );


  buf
  g19
  (
    n56,
    n47
  );


  buf
  g20
  (
    KeyWire_0_8,
    n45
  );


  buf
  g21
  (
    n49,
    n4
  );


  buf
  g22
  (
    n63,
    n46
  );


  buf
  g23
  (
    KeyWire_0_20,
    n6
  );


  buf
  g24
  (
    n62,
    n3
  );


  buf
  g25
  (
    KeyWire_0_26,
    n46
  );


  buf
  g26
  (
    n53,
    n46
  );


  nor
  g27
  (
    n60,
    n45,
    n4,
    n5,
    n46
  );


  nor
  g28
  (
    n57,
    n45,
    n47,
    n44
  );


  xnor
  g29
  (
    n48,
    n44,
    n5,
    n3,
    n4
  );


  or
  g30
  (
    n51,
    n47,
    n45,
    n5,
    n3
  );


  not
  g31
  (
    n110,
    n9
  );


  buf
  g32
  (
    n100,
    n7
  );


  buf
  g33
  (
    n80,
    n59
  );


  buf
  g34
  (
    n108,
    n52
  );


  not
  g35
  (
    KeyWire_0_6,
    n26
  );


  not
  g36
  (
    KeyWire_0_24,
    n23
  );


  buf
  g37
  (
    KeyWire_0_21,
    n19
  );


  not
  g38
  (
    n86,
    n50
  );


  buf
  g39
  (
    n75,
    n38
  );


  not
  g40
  (
    KeyWire_0_9,
    n20
  );


  not
  g41
  (
    n107,
    n60
  );


  not
  g42
  (
    n72,
    n6
  );


  not
  g43
  (
    n68,
    n9
  );


  buf
  g44
  (
    n115,
    n8
  );


  not
  g45
  (
    n81,
    n28
  );


  xor
  g46
  (
    KeyWire_0_10,
    n20,
    n61,
    n10
  );


  xnor
  g47
  (
    KeyWire_0_12,
    n8,
    n14,
    n18,
    n28
  );


  nor
  g48
  (
    KeyWire_0_17,
    n57,
    n56,
    n58,
    n31
  );


  xnor
  g49
  (
    n67,
    n51,
    n56,
    n11,
    n13
  );


  xnor
  g50
  (
    n84,
    n18,
    n61,
    n27,
    n60
  );


  nand
  g51
  (
    n103,
    n53,
    n18,
    n62
  );


  and
  g52
  (
    n79,
    n14,
    n48,
    n31,
    n7
  );


  xor
  g53
  (
    KeyWire_0_23,
    n28,
    n57,
    n60,
    n49
  );


  nor
  g54
  (
    n95,
    n16,
    n32,
    n15,
    n57
  );


  nor
  g55
  (
    KeyWire_0_2,
    n26,
    n12,
    n31,
    n27
  );


  xnor
  g56
  (
    n109,
    n21,
    n12,
    n49,
    n32
  );


  nor
  g57
  (
    n102,
    n28,
    n30,
    n14,
    n16
  );


  xnor
  g58
  (
    n78,
    n32,
    n11,
    n15,
    n54
  );


  or
  g59
  (
    n71,
    n16,
    n63,
    n18,
    n25
  );


  nor
  g60
  (
    n96,
    n53,
    n14,
    n51,
    n57
  );


  nand
  g61
  (
    n93,
    n22,
    n30,
    n63,
    n58
  );


  xor
  g62
  (
    KeyWire_0_5,
    n23,
    n10,
    n37,
    n27
  );


  xor
  g63
  (
    KeyWire_0_13,
    n60,
    n29,
    n6,
    n27
  );


  xor
  g64
  (
    KeyWire_0_30,
    n55,
    n53,
    n12,
    n13
  );


  xnor
  g65
  (
    KeyWire_0_15,
    n52,
    n52,
    n21,
    n16
  );


  and
  g66
  (
    n106,
    n25,
    n19,
    n23,
    n55
  );


  or
  g67
  (
    KeyWire_0_29,
    n26,
    n55,
    n63,
    n29
  );


  xnor
  g68
  (
    KeyWire_0_0,
    n59,
    n52,
    n50,
    n13
  );


  or
  g69
  (
    n91,
    n53,
    n15,
    n19,
    n24
  );


  or
  g70
  (
    n116,
    n58,
    n29,
    n56,
    n62
  );


  and
  g71
  (
    n104,
    n21,
    n38,
    n22,
    n17
  );


  nand
  g72
  (
    n82,
    n23,
    n10,
    n48,
    n51
  );


  xnor
  g73
  (
    n65,
    n20,
    n48,
    n9,
    n13
  );


  and
  g74
  (
    n76,
    n6,
    n63,
    n49,
    n10
  );


  and
  g75
  (
    n113,
    n24,
    n50,
    n7,
    n59
  );


  nor
  g76
  (
    n83,
    n21,
    n24,
    n30
  );


  nand
  g77
  (
    n112,
    n51,
    n54,
    n8,
    n56
  );


  xnor
  g78
  (
    n98,
    n8,
    n22,
    n9,
    n26
  );


  nand
  g79
  (
    n101,
    n20,
    n59,
    n54,
    n17
  );


  nand
  g80
  (
    n77,
    n49,
    n25,
    n29,
    n61
  );


  nor
  g81
  (
    n111,
    n15,
    n31,
    n19,
    n12
  );


  and
  g82
  (
    n90,
    n38,
    n58,
    n22,
    n11
  );


  and
  g83
  (
    n92,
    n55,
    n32,
    n62,
    n48
  );


  nand
  g84
  (
    n114,
    n7,
    n50,
    n25,
    n54
  );


  or
  g85
  (
    n70,
    n11,
    n30,
    n17
  );


  xnor
  g86
  (
    KeyWire_0_1,
    n118,
    n101,
    n107,
    n115
  );


  xnor
  g87
  (
    KeyWire_0_18,
    n95,
    n110,
    n113,
    n103
  );


  xor
  g88
  (
    KeyWire_0_11,
    n115,
    n111,
    n116,
    n118
  );


  xnor
  g89
  (
    n119,
    n86,
    n106,
    n100,
    n84
  );


  nor
  g90
  (
    n132,
    n112,
    n99,
    n94,
    n82
  );


  xnor
  g91
  (
    KeyWire_0_4,
    n80,
    n77,
    n117,
    n93
  );


  and
  g92
  (
    n124,
    n117,
    n97,
    n116,
    n115
  );


  or
  g93
  (
    n128,
    n117,
    n89,
    n104,
    n98
  );


  and
  g94
  (
    KeyWire_0_25,
    n114,
    n116,
    n88,
    n87
  );


  nand
  g95
  (
    n125,
    n105,
    n113,
    n96,
    n92
  );


  nor
  g96
  (
    KeyWire_0_31,
    n85,
    n109,
    n102,
    n78
  );


  nand
  g97
  (
    n129,
    n112,
    n114,
    n90,
    n113
  );


  and
  g98
  (
    KeyWire_0_28,
    n79,
    n108,
    n114,
    n112
  );


  and
  g99
  (
    n121,
    n83,
    n118,
    n81,
    n91
  );


  xor
  KeyGate_0_0
  (
    n87,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n130,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n118,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n45,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n120,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n74,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n117,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n33,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n54,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n97,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n66,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n131,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n105,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n85,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n42,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n99,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n44,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n88,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n122,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n61,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n55,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n94,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n50,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n89,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n73,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n126,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n52,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n43,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n123,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n64,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n69,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n127,
    KeyNOTWire_0_31
  );


endmodule

