

module Stat_714_926
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n737,
  n723,
  n732,
  n729,
  n730,
  n736,
  n725,
  n728,
  n738,
  n726,
  n722,
  n727,
  n719,
  n724,
  n734,
  n731,
  n720,
  n733,
  n735,
  n721,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n737;
  output n723;
  output n732;
  output n729;
  output n730;
  output n736;
  output n725;
  output n728;
  output n738;
  output n726;
  output n722;
  output n727;
  output n719;
  output n724;
  output n734;
  output n731;
  output n720;
  output n733;
  output n735;
  output n721;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n70,
    n6
  );


  not
  g1
  (
    n77,
    n7
  );


  not
  g2
  (
    n29,
    n21
  );


  not
  g3
  (
    n75,
    n13
  );


  not
  g4
  (
    n74,
    n15
  );


  not
  g5
  (
    n67,
    n20
  );


  not
  g6
  (
    n81,
    n17
  );


  buf
  g7
  (
    n97,
    n2
  );


  not
  g8
  (
    n108,
    n23
  );


  not
  g9
  (
    n36,
    n13
  );


  buf
  g10
  (
    n31,
    n15
  );


  buf
  g11
  (
    n58,
    n1
  );


  buf
  g12
  (
    n27,
    n24
  );


  buf
  g13
  (
    n51,
    n4
  );


  buf
  g14
  (
    n88,
    n16
  );


  buf
  g15
  (
    n47,
    n11
  );


  not
  g16
  (
    n102,
    n23
  );


  not
  g17
  (
    n53,
    n8
  );


  buf
  g18
  (
    n99,
    n8
  );


  buf
  g19
  (
    KeyWire_0_1,
    n12
  );


  buf
  g20
  (
    n32,
    n24
  );


  not
  g21
  (
    n64,
    n12
  );


  not
  g22
  (
    n57,
    n12
  );


  not
  g23
  (
    KeyWire_0_6,
    n19
  );


  buf
  g24
  (
    n37,
    n5
  );


  not
  g25
  (
    n69,
    n8
  );


  not
  g26
  (
    n43,
    n22
  );


  not
  g27
  (
    n95,
    n15
  );


  buf
  g28
  (
    KeyWire_0_25,
    n9
  );


  not
  g29
  (
    n33,
    n17
  );


  buf
  g30
  (
    n120,
    n5
  );


  buf
  g31
  (
    n52,
    n6
  );


  not
  g32
  (
    n54,
    n24
  );


  not
  g33
  (
    KeyWire_0_50,
    n18
  );


  not
  g34
  (
    KeyWire_0_22,
    n6
  );


  not
  g35
  (
    KeyWire_0_15,
    n23
  );


  not
  g36
  (
    n79,
    n17
  );


  not
  g37
  (
    n44,
    n24
  );


  not
  g38
  (
    n96,
    n21
  );


  not
  g39
  (
    n65,
    n9
  );


  buf
  g40
  (
    n61,
    n18
  );


  buf
  g41
  (
    n90,
    n2
  );


  not
  g42
  (
    n60,
    n12
  );


  not
  g43
  (
    KeyWire_0_24,
    n8
  );


  buf
  g44
  (
    n100,
    n9
  );


  buf
  g45
  (
    n35,
    n16
  );


  buf
  g46
  (
    n91,
    n20
  );


  buf
  g47
  (
    n101,
    n2
  );


  not
  g48
  (
    n113,
    n3
  );


  buf
  g49
  (
    n116,
    n22
  );


  buf
  g50
  (
    n98,
    n14
  );


  buf
  g51
  (
    KeyWire_0_13,
    n14
  );


  buf
  g52
  (
    n111,
    n10
  );


  not
  g53
  (
    n112,
    n19
  );


  not
  g54
  (
    n45,
    n14
  );


  buf
  g55
  (
    n56,
    n20
  );


  buf
  g56
  (
    n87,
    n4
  );


  not
  g57
  (
    n26,
    n11
  );


  not
  g58
  (
    n83,
    n17
  );


  not
  g59
  (
    n59,
    n18
  );


  not
  g60
  (
    n86,
    n16
  );


  buf
  g61
  (
    n109,
    n7
  );


  buf
  g62
  (
    n39,
    n1
  );


  buf
  g63
  (
    n62,
    n16
  );


  not
  g64
  (
    n42,
    n20
  );


  not
  g65
  (
    n55,
    n11
  );


  not
  g66
  (
    n71,
    n4
  );


  not
  g67
  (
    KeyWire_0_17,
    n1
  );


  not
  g68
  (
    n80,
    n4
  );


  not
  g69
  (
    n103,
    n9
  );


  not
  g70
  (
    n119,
    n14
  );


  buf
  g71
  (
    n50,
    n22
  );


  not
  g72
  (
    n104,
    n19
  );


  buf
  g73
  (
    n34,
    n21
  );


  not
  g74
  (
    n28,
    n3
  );


  buf
  g75
  (
    n41,
    n10
  );


  buf
  g76
  (
    n106,
    n2
  );


  buf
  g77
  (
    n76,
    n10
  );


  not
  g78
  (
    n117,
    n5
  );


  buf
  g79
  (
    n82,
    n6
  );


  not
  g80
  (
    KeyWire_0_47,
    n18
  );


  not
  g81
  (
    n30,
    n1
  );


  not
  g82
  (
    n38,
    n15
  );


  not
  g83
  (
    n89,
    n22
  );


  not
  g84
  (
    n107,
    n19
  );


  not
  g85
  (
    n78,
    n23
  );


  not
  g86
  (
    n105,
    n7
  );


  buf
  g87
  (
    n40,
    n13
  );


  buf
  g88
  (
    n73,
    n7
  );


  not
  g89
  (
    n110,
    n3
  );


  buf
  g90
  (
    n49,
    n21
  );


  buf
  g91
  (
    n94,
    n10
  );


  buf
  g92
  (
    n48,
    n3
  );


  buf
  g93
  (
    n115,
    n11
  );


  buf
  g94
  (
    n85,
    n13
  );


  buf
  g95
  (
    n114,
    n5
  );


  not
  g96
  (
    n277,
    n25
  );


  not
  g97
  (
    n162,
    n29
  );


  buf
  g98
  (
    n266,
    n32
  );


  buf
  g99
  (
    n335,
    n82
  );


  not
  g100
  (
    n329,
    n82
  );


  not
  g101
  (
    n275,
    n84
  );


  not
  g102
  (
    KeyWire_0_32,
    n32
  );


  not
  g103
  (
    n200,
    n66
  );


  buf
  g104
  (
    n150,
    n88
  );


  buf
  g105
  (
    n336,
    n55
  );


  not
  g106
  (
    n367,
    n44
  );


  buf
  g107
  (
    n261,
    n70
  );


  buf
  g108
  (
    n310,
    n64
  );


  not
  g109
  (
    n282,
    n48
  );


  not
  g110
  (
    n229,
    n84
  );


  buf
  g111
  (
    KeyWire_0_12,
    n70
  );


  not
  g112
  (
    n377,
    n67
  );


  buf
  g113
  (
    n273,
    n91
  );


  not
  g114
  (
    n147,
    n51
  );


  not
  g115
  (
    n173,
    n52
  );


  not
  g116
  (
    n340,
    n73
  );


  buf
  g117
  (
    n136,
    n45
  );


  not
  g118
  (
    n214,
    n25
  );


  not
  g119
  (
    n215,
    n39
  );


  buf
  g120
  (
    n308,
    n30
  );


  buf
  g121
  (
    n125,
    n84
  );


  not
  g122
  (
    n148,
    n44
  );


  buf
  g123
  (
    n267,
    n47
  );


  buf
  g124
  (
    n381,
    n60
  );


  buf
  g125
  (
    n145,
    n44
  );


  not
  g126
  (
    n351,
    n82
  );


  not
  g127
  (
    n204,
    n90
  );


  buf
  g128
  (
    n184,
    n89
  );


  not
  g129
  (
    n300,
    n79
  );


  not
  g130
  (
    n211,
    n86
  );


  not
  g131
  (
    n166,
    n57
  );


  not
  g132
  (
    n255,
    n79
  );


  buf
  g133
  (
    n197,
    n55
  );


  buf
  g134
  (
    n155,
    n28
  );


  buf
  g135
  (
    n302,
    n26
  );


  not
  g136
  (
    KeyWire_0_51,
    n77
  );


  not
  g137
  (
    n356,
    n55
  );


  buf
  g138
  (
    n143,
    n37
  );


  not
  g139
  (
    n347,
    n52
  );


  not
  g140
  (
    n203,
    n25
  );


  not
  g141
  (
    n238,
    n73
  );


  buf
  g142
  (
    n318,
    n32
  );


  buf
  g143
  (
    KeyWire_0_20,
    n75
  );


  buf
  g144
  (
    KeyWire_0_60,
    n54
  );


  buf
  g145
  (
    n354,
    n73
  );


  buf
  g146
  (
    n328,
    n62
  );


  not
  g147
  (
    n359,
    n69
  );


  not
  g148
  (
    n361,
    n67
  );


  buf
  g149
  (
    n137,
    n41
  );


  buf
  g150
  (
    n209,
    n75
  );


  buf
  g151
  (
    n231,
    n85
  );


  buf
  g152
  (
    n168,
    n68
  );


  not
  g153
  (
    KeyWire_0_62,
    n77
  );


  buf
  g154
  (
    KeyWire_0_46,
    n31
  );


  not
  g155
  (
    n224,
    n72
  );


  buf
  g156
  (
    n139,
    n58
  );


  buf
  g157
  (
    n126,
    n38
  );


  buf
  g158
  (
    n257,
    n60
  );


  buf
  g159
  (
    n260,
    n67
  );


  buf
  g160
  (
    n364,
    n87
  );


  buf
  g161
  (
    n258,
    n81
  );


  buf
  g162
  (
    n218,
    n78
  );


  not
  g163
  (
    n183,
    n65
  );


  not
  g164
  (
    n297,
    n85
  );


  buf
  g165
  (
    n368,
    n58
  );


  buf
  g166
  (
    n309,
    n61
  );


  not
  g167
  (
    n380,
    n50
  );


  not
  g168
  (
    n191,
    n82
  );


  buf
  g169
  (
    n227,
    n30
  );


  buf
  g170
  (
    n181,
    n45
  );


  not
  g171
  (
    n252,
    n68
  );


  buf
  g172
  (
    n262,
    n48
  );


  not
  g173
  (
    n271,
    n43
  );


  not
  g174
  (
    n212,
    n41
  );


  buf
  g175
  (
    n159,
    n49
  );


  not
  g176
  (
    n226,
    n35
  );


  buf
  g177
  (
    n130,
    n34
  );


  buf
  g178
  (
    n341,
    n76
  );


  buf
  g179
  (
    KeyWire_0_35,
    n83
  );


  buf
  g180
  (
    n121,
    n38
  );


  not
  g181
  (
    n350,
    n36
  );


  not
  g182
  (
    n192,
    n43
  );


  buf
  g183
  (
    n317,
    n80
  );


  not
  g184
  (
    n369,
    n88
  );


  not
  g185
  (
    n259,
    n62
  );


  not
  g186
  (
    n312,
    n49
  );


  not
  g187
  (
    n299,
    n47
  );


  buf
  g188
  (
    n217,
    n51
  );


  not
  g189
  (
    n272,
    n58
  );


  not
  g190
  (
    n342,
    n85
  );


  not
  g191
  (
    n264,
    n43
  );


  buf
  g192
  (
    n338,
    n59
  );


  not
  g193
  (
    n301,
    n31
  );


  buf
  g194
  (
    n248,
    n50
  );


  not
  g195
  (
    n175,
    n61
  );


  buf
  g196
  (
    n287,
    n83
  );


  buf
  g197
  (
    n314,
    n25
  );


  not
  g198
  (
    n236,
    n54
  );


  not
  g199
  (
    KeyWire_0_11,
    n91
  );


  not
  g200
  (
    n144,
    n39
  );


  not
  g201
  (
    n346,
    n27
  );


  buf
  g202
  (
    n169,
    n57
  );


  buf
  g203
  (
    n378,
    n48
  );


  buf
  g204
  (
    n213,
    n26
  );


  buf
  g205
  (
    n131,
    n30
  );


  buf
  g206
  (
    n208,
    n55
  );


  buf
  g207
  (
    KeyWire_0_39,
    n56
  );


  buf
  g208
  (
    n194,
    n86
  );


  not
  g209
  (
    n138,
    n81
  );


  buf
  g210
  (
    n122,
    n69
  );


  buf
  g211
  (
    n298,
    n61
  );


  not
  g212
  (
    n244,
    n89
  );


  buf
  g213
  (
    n253,
    n66
  );


  buf
  g214
  (
    n289,
    n50
  );


  buf
  g215
  (
    n305,
    n65
  );


  buf
  g216
  (
    n296,
    n67
  );


  buf
  g217
  (
    n134,
    n78
  );


  not
  g218
  (
    n201,
    n46
  );


  not
  g219
  (
    n124,
    n77
  );


  not
  g220
  (
    n280,
    n31
  );


  not
  g221
  (
    n243,
    n63
  );


  buf
  g222
  (
    n307,
    n27
  );


  not
  g223
  (
    n156,
    n45
  );


  not
  g224
  (
    n132,
    n42
  );


  not
  g225
  (
    n177,
    n46
  );


  not
  g226
  (
    n355,
    n75
  );


  buf
  g227
  (
    n286,
    n51
  );


  not
  g228
  (
    n372,
    n29
  );


  buf
  g229
  (
    n185,
    n53
  );


  not
  g230
  (
    n163,
    n77
  );


  buf
  g231
  (
    n241,
    n59
  );


  not
  g232
  (
    KeyWire_0_54,
    n60
  );


  buf
  g233
  (
    n327,
    n41
  );


  buf
  g234
  (
    n311,
    n80
  );


  not
  g235
  (
    n158,
    n74
  );


  not
  g236
  (
    n189,
    n49
  );


  buf
  g237
  (
    n193,
    n38
  );


  not
  g238
  (
    n283,
    n40
  );


  not
  g239
  (
    n278,
    n32
  );


  buf
  g240
  (
    n199,
    n26
  );


  buf
  g241
  (
    n270,
    n29
  );


  buf
  g242
  (
    n288,
    n76
  );


  not
  g243
  (
    n379,
    n69
  );


  buf
  g244
  (
    n357,
    n85
  );


  buf
  g245
  (
    n216,
    n56
  );


  not
  g246
  (
    n178,
    n45
  );


  buf
  g247
  (
    n190,
    n48
  );


  buf
  g248
  (
    KeyWire_0_44,
    n68
  );


  buf
  g249
  (
    n157,
    n72
  );


  not
  g250
  (
    n313,
    n36
  );


  buf
  g251
  (
    n320,
    n33
  );


  buf
  g252
  (
    n250,
    n63
  );


  not
  g253
  (
    n172,
    n71
  );


  buf
  g254
  (
    n316,
    n35
  );


  buf
  g255
  (
    n146,
    n56
  );


  buf
  g256
  (
    n123,
    n74
  );


  not
  g257
  (
    n222,
    n78
  );


  not
  g258
  (
    n337,
    n79
  );


  not
  g259
  (
    n174,
    n71
  );


  buf
  g260
  (
    n263,
    n49
  );


  not
  g261
  (
    n234,
    n71
  );


  buf
  g262
  (
    n374,
    n76
  );


  not
  g263
  (
    n149,
    n61
  );


  not
  g264
  (
    n291,
    n28
  );


  not
  g265
  (
    n319,
    n76
  );


  buf
  g266
  (
    n386,
    n75
  );


  not
  g267
  (
    n165,
    n27
  );


  buf
  g268
  (
    n202,
    n78
  );


  buf
  g269
  (
    n240,
    n63
  );


  buf
  g270
  (
    n339,
    n52
  );


  not
  g271
  (
    n304,
    n74
  );


  buf
  g272
  (
    n256,
    n80
  );


  buf
  g273
  (
    KeyWire_0_49,
    n40
  );


  not
  g274
  (
    n269,
    n70
  );


  buf
  g275
  (
    n323,
    n34
  );


  buf
  g276
  (
    n153,
    n74
  );


  buf
  g277
  (
    n207,
    n81
  );


  buf
  g278
  (
    n161,
    n81
  );


  buf
  g279
  (
    n206,
    n43
  );


  not
  g280
  (
    n167,
    n90
  );


  not
  g281
  (
    n141,
    n83
  );


  buf
  g282
  (
    n294,
    n71
  );


  not
  g283
  (
    n362,
    n90
  );


  not
  g284
  (
    n330,
    n46
  );


  buf
  g285
  (
    KeyWire_0_21,
    n34
  );


  buf
  g286
  (
    KeyWire_0_2,
    n83
  );


  not
  g287
  (
    n179,
    n89
  );


  not
  g288
  (
    n268,
    n86
  );


  not
  g289
  (
    n365,
    n31
  );


  buf
  g290
  (
    n233,
    n58
  );


  not
  g291
  (
    n247,
    n91
  );


  buf
  g292
  (
    n290,
    n53
  );


  not
  g293
  (
    KeyWire_0_30,
    n57
  );


  not
  g294
  (
    KeyWire_0_45,
    n59
  );


  not
  g295
  (
    n135,
    n72
  );


  buf
  g296
  (
    n315,
    n53
  );


  buf
  g297
  (
    KeyWire_0_27,
    n62
  );


  not
  g298
  (
    KeyWire_0_38,
    n26
  );


  not
  g299
  (
    n128,
    n65
  );


  buf
  g300
  (
    n344,
    n66
  );


  not
  g301
  (
    n363,
    n84
  );


  buf
  g302
  (
    n187,
    n33
  );


  not
  g303
  (
    n348,
    n88
  );


  not
  g304
  (
    n205,
    n64
  );


  not
  g305
  (
    n343,
    n42
  );


  buf
  g306
  (
    n221,
    n47
  );


  buf
  g307
  (
    n151,
    n80
  );


  not
  g308
  (
    n182,
    n44
  );


  buf
  g309
  (
    n293,
    n62
  );


  buf
  g310
  (
    n322,
    n35
  );


  not
  g311
  (
    n360,
    n68
  );


  not
  g312
  (
    n326,
    n34
  );


  not
  g313
  (
    n152,
    n72
  );


  buf
  g314
  (
    n385,
    n41
  );


  buf
  g315
  (
    n285,
    n69
  );


  buf
  g316
  (
    n129,
    n91
  );


  not
  g317
  (
    n160,
    n36
  );


  not
  g318
  (
    KeyWire_0_31,
    n90
  );


  not
  g319
  (
    n180,
    n29
  );


  buf
  g320
  (
    KeyWire_0_14,
    n86
  );


  buf
  g321
  (
    n333,
    n40
  );


  not
  g322
  (
    n358,
    n46
  );


  not
  g323
  (
    n388,
    n39
  );


  buf
  g324
  (
    n210,
    n87
  );


  not
  g325
  (
    n334,
    n37
  );


  not
  g326
  (
    n375,
    n50
  );


  buf
  g327
  (
    n198,
    n42
  );


  buf
  g328
  (
    n265,
    n87
  );


  buf
  g329
  (
    n292,
    n38
  );


  buf
  g330
  (
    n371,
    n39
  );


  buf
  g331
  (
    n154,
    n65
  );


  buf
  g332
  (
    KeyWire_0_63,
    n40
  );


  not
  g333
  (
    n140,
    n89
  );


  not
  g334
  (
    n171,
    n63
  );


  not
  g335
  (
    n237,
    n64
  );


  not
  g336
  (
    n246,
    n30
  );


  buf
  g337
  (
    n276,
    n52
  );


  not
  g338
  (
    n332,
    n54
  );


  not
  g339
  (
    n254,
    n60
  );


  not
  g340
  (
    n321,
    n79
  );


  buf
  g341
  (
    n232,
    n37
  );


  buf
  g342
  (
    n345,
    n57
  );


  buf
  g343
  (
    n133,
    n47
  );


  buf
  g344
  (
    n303,
    n27
  );


  buf
  g345
  (
    n353,
    n70
  );


  not
  g346
  (
    n225,
    n28
  );


  buf
  g347
  (
    n235,
    n36
  );


  buf
  g348
  (
    n195,
    n73
  );


  buf
  g349
  (
    n164,
    n37
  );


  not
  g350
  (
    n228,
    n53
  );


  buf
  g351
  (
    n370,
    n87
  );


  not
  g352
  (
    n383,
    n56
  );


  buf
  g353
  (
    n306,
    n33
  );


  not
  g354
  (
    n295,
    n51
  );


  buf
  g355
  (
    n279,
    n35
  );


  buf
  g356
  (
    n366,
    n28
  );


  not
  g357
  (
    n384,
    n64
  );


  buf
  g358
  (
    n373,
    n59
  );


  not
  g359
  (
    n219,
    n42
  );


  buf
  g360
  (
    n239,
    n33
  );


  buf
  g361
  (
    n349,
    n54
  );


  buf
  g362
  (
    n376,
    n66
  );


  buf
  g363
  (
    n186,
    n88
  );


  buf
  g364
  (
    n417,
    n139
  );


  buf
  g365
  (
    n420,
    n123
  );


  buf
  g366
  (
    n407,
    n147
  );


  not
  g367
  (
    n390,
    n144
  );


  not
  g368
  (
    n410,
    n142
  );


  not
  g369
  (
    n396,
    n143
  );


  buf
  g370
  (
    n404,
    n127
  );


  buf
  g371
  (
    n403,
    n152
  );


  not
  g372
  (
    n415,
    n121
  );


  not
  g373
  (
    n394,
    n135
  );


  buf
  g374
  (
    n401,
    n122
  );


  buf
  g375
  (
    n414,
    n137
  );


  not
  g376
  (
    n397,
    n140
  );


  not
  g377
  (
    n406,
    n132
  );


  not
  g378
  (
    n411,
    n148
  );


  not
  g379
  (
    n391,
    n128
  );


  buf
  g380
  (
    n413,
    n130
  );


  buf
  g381
  (
    n416,
    n145
  );


  buf
  g382
  (
    n399,
    n141
  );


  not
  g383
  (
    n408,
    n146
  );


  buf
  g384
  (
    n419,
    n125
  );


  not
  g385
  (
    n395,
    n138
  );


  buf
  g386
  (
    n393,
    n149
  );


  not
  g387
  (
    n412,
    n124
  );


  not
  g388
  (
    n409,
    n134
  );


  buf
  g389
  (
    n405,
    n129
  );


  buf
  g390
  (
    n392,
    n133
  );


  not
  g391
  (
    n400,
    n150
  );


  not
  g392
  (
    n389,
    n136
  );


  not
  g393
  (
    KeyWire_0_41,
    n126
  );


  not
  g394
  (
    n418,
    n151
  );


  buf
  g395
  (
    n402,
    n131
  );


  buf
  g396
  (
    KeyWire_0_48,
    n284
  );


  buf
  g397
  (
    KeyWire_0_0,
    n192
  );


  not
  g398
  (
    n445,
    n227
  );


  buf
  g399
  (
    n535,
    n396
  );


  buf
  g400
  (
    n424,
    n406
  );


  buf
  g401
  (
    n509,
    n93
  );


  buf
  g402
  (
    n469,
    n116
  );


  buf
  g403
  (
    n435,
    n222
  );


  not
  g404
  (
    n439,
    n259
  );


  not
  g405
  (
    n493,
    n212
  );


  buf
  g406
  (
    n461,
    n399
  );


  not
  g407
  (
    KeyWire_0_59,
    n113
  );


  buf
  g408
  (
    n454,
    n93
  );


  buf
  g409
  (
    n475,
    n402
  );


  not
  g410
  (
    n449,
    n394
  );


  buf
  g411
  (
    n527,
    n117
  );


  buf
  g412
  (
    KeyWire_0_28,
    n397
  );


  not
  g413
  (
    n426,
    n220
  );


  not
  g414
  (
    n513,
    n92
  );


  buf
  g415
  (
    n458,
    n413
  );


  not
  g416
  (
    KeyWire_0_43,
    n110
  );


  buf
  g417
  (
    n536,
    n406
  );


  not
  g418
  (
    n511,
    n238
  );


  not
  g419
  (
    n456,
    n109
  );


  buf
  g420
  (
    n546,
    n168
  );


  buf
  g421
  (
    n421,
    n92
  );


  buf
  g422
  (
    n491,
    n191
  );


  not
  g423
  (
    n514,
    n162
  );


  buf
  g424
  (
    n450,
    n391
  );


  not
  g425
  (
    n451,
    n165
  );


  buf
  g426
  (
    n470,
    n236
  );


  buf
  g427
  (
    n533,
    n265
  );


  buf
  g428
  (
    n504,
    n184
  );


  not
  g429
  (
    KeyWire_0_9,
    n407
  );


  buf
  g430
  (
    n505,
    n393
  );


  not
  g431
  (
    n486,
    n281
  );


  buf
  g432
  (
    n464,
    n116
  );


  buf
  g433
  (
    n429,
    n100
  );


  buf
  g434
  (
    n482,
    n250
  );


  buf
  g435
  (
    n436,
    n411
  );


  not
  g436
  (
    n489,
    n392
  );


  not
  g437
  (
    n540,
    n418
  );


  not
  g438
  (
    n453,
    n190
  );


  buf
  g439
  (
    n518,
    n104
  );


  xor
  g440
  (
    n471,
    n182,
    n97,
    n411
  );


  and
  g441
  (
    n532,
    n230,
    n408,
    n411,
    n400
  );


  xnor
  g442
  (
    n547,
    n201,
    n105,
    n419,
    n402
  );


  xor
  g443
  (
    n487,
    n99,
    n101,
    n119,
    n414
  );


  xnor
  g444
  (
    n481,
    n416,
    n206,
    n101,
    n392
  );


  or
  g445
  (
    n444,
    n414,
    n117,
    n226,
    n118
  );


  xnor
  g446
  (
    n506,
    n171,
    n110,
    n217,
    n398
  );


  xor
  g447
  (
    n526,
    n163,
    n211,
    n403,
    n274
  );


  xor
  g448
  (
    n483,
    n237,
    n391,
    n241,
    n266
  );


  xor
  g449
  (
    n522,
    n399,
    n228,
    n221,
    n110
  );


  xor
  g450
  (
    n485,
    n405,
    n115,
    n116,
    n395
  );


  and
  g451
  (
    n432,
    n102,
    n160,
    n94,
    n208
  );


  xnor
  g452
  (
    n497,
    n158,
    n98,
    n117,
    n108
  );


  and
  g453
  (
    n541,
    n391,
    n389,
    n108,
    n99
  );


  nor
  g454
  (
    KeyWire_0_58,
    n234,
    n251,
    n155,
    n120
  );


  xnor
  g455
  (
    n447,
    n105,
    n197,
    n412,
    n176
  );


  nor
  g456
  (
    n437,
    n100,
    n94,
    n404,
    n398
  );


  xor
  g457
  (
    n442,
    n413,
    n396,
    n412,
    n416
  );


  and
  g458
  (
    n534,
    n103,
    n119,
    n416,
    n404
  );


  xor
  g459
  (
    n457,
    n235,
    n106,
    n407,
    n260
  );


  or
  g460
  (
    n543,
    n100,
    n103,
    n209,
    n398
  );


  nand
  g461
  (
    KeyWire_0_34,
    n409,
    n252,
    n106,
    n95
  );


  or
  g462
  (
    n434,
    n389,
    n181,
    n413,
    n204
  );


  and
  g463
  (
    n528,
    n223,
    n248,
    n396,
    n103
  );


  nand
  g464
  (
    n519,
    n189,
    n393,
    n117,
    n112
  );


  and
  g465
  (
    n499,
    n268,
    n406,
    n202,
    n396
  );


  nor
  g466
  (
    n517,
    n409,
    n267,
    n405,
    n408
  );


  or
  g467
  (
    n467,
    n93,
    n105,
    n417,
    n264
  );


  xnor
  g468
  (
    n423,
    n98,
    n118,
    n229,
    n103
  );


  and
  g469
  (
    n529,
    n409,
    n115,
    n401,
    n224
  );


  or
  g470
  (
    n459,
    n119,
    n390,
    n169,
    n394
  );


  and
  g471
  (
    n428,
    n95,
    n397,
    n233,
    n177
  );


  xor
  g472
  (
    n476,
    n232,
    n94,
    n419,
    n392
  );


  nor
  g473
  (
    n478,
    n105,
    n401,
    n390,
    n116
  );


  and
  g474
  (
    n498,
    n93,
    n94,
    n178,
    n166
  );


  or
  g475
  (
    n488,
    n108,
    n420,
    n111,
    n271
  );


  or
  g476
  (
    KeyWire_0_36,
    n218,
    n278,
    n243,
    n401
  );


  nand
  g477
  (
    n508,
    n96,
    n399,
    n415,
    n416
  );


  nand
  g478
  (
    n422,
    n404,
    n110,
    n400,
    n156
  );


  or
  g479
  (
    n468,
    n187,
    n113,
    n203,
    n97
  );


  xnor
  g480
  (
    n542,
    n407,
    n282,
    n389,
    n390
  );


  or
  g481
  (
    n495,
    n261,
    n219,
    n215,
    n397
  );


  xnor
  g482
  (
    n544,
    n115,
    n186,
    n258,
    n389
  );


  and
  g483
  (
    KeyWire_0_42,
    n411,
    n198,
    n199,
    n104
  );


  xnor
  g484
  (
    n441,
    n118,
    n253,
    n119,
    n242
  );


  nor
  g485
  (
    n538,
    n288,
    n214,
    n412,
    n112
  );


  or
  g486
  (
    n512,
    n111,
    n417,
    n114,
    n179
  );


  and
  g487
  (
    n500,
    n418,
    n109,
    n415,
    n394
  );


  nand
  g488
  (
    n425,
    n272,
    n244,
    n164,
    n400
  );


  xnor
  g489
  (
    n433,
    n255,
    n101,
    n231,
    n104
  );


  and
  g490
  (
    n452,
    n403,
    n407,
    n269,
    n249
  );


  nand
  g491
  (
    n466,
    n106,
    n405,
    n210,
    n194
  );


  nand
  g492
  (
    n502,
    n414,
    n395,
    n263,
    n409
  );


  nor
  g493
  (
    n438,
    n183,
    n277,
    n96,
    n418
  );


  nand
  g494
  (
    n531,
    n154,
    n205,
    n188,
    n415
  );


  xnor
  g495
  (
    n430,
    n216,
    n98,
    n95,
    n107
  );


  nand
  g496
  (
    n490,
    n403,
    n410,
    n109,
    n280
  );


  and
  g497
  (
    n516,
    n195,
    n245,
    n111,
    n410
  );


  nor
  g498
  (
    n472,
    n403,
    n419,
    n96,
    n417
  );


  and
  g499
  (
    n477,
    n415,
    n412,
    n270,
    n102
  );


  and
  g500
  (
    KeyWire_0_53,
    n262,
    n254,
    n401,
    n400
  );


  and
  g501
  (
    n465,
    n112,
    n390,
    n193,
    n99
  );


  xor
  g502
  (
    n474,
    n239,
    n114,
    n414,
    n112
  );


  xor
  g503
  (
    n507,
    n114,
    n395,
    n170,
    n283
  );


  xnor
  g504
  (
    KeyWire_0_26,
    n405,
    n393,
    n157,
    n102
  );


  xnor
  g505
  (
    n446,
    n257,
    n420,
    n410,
    n106
  );


  nand
  g506
  (
    n473,
    n159,
    n107,
    n101,
    n393
  );


  and
  g507
  (
    n520,
    n419,
    n256,
    n402,
    n97
  );


  or
  g508
  (
    n427,
    n225,
    n96,
    n290,
    n92
  );


  and
  g509
  (
    n503,
    n398,
    n111,
    n402,
    n207
  );


  and
  g510
  (
    n539,
    n95,
    n394,
    n114,
    n418
  );


  xor
  g511
  (
    n463,
    n107,
    n286,
    n406,
    n279
  );


  nor
  g512
  (
    n440,
    n408,
    n395,
    n102,
    n246
  );


  nand
  g513
  (
    n484,
    n185,
    n213,
    n287,
    n275
  );


  nand
  g514
  (
    n501,
    n399,
    n200,
    n285,
    n397
  );


  nand
  g515
  (
    n515,
    n97,
    n108,
    n420,
    n113
  );


  or
  g516
  (
    n530,
    n173,
    n413,
    n417,
    n92
  );


  and
  g517
  (
    n510,
    n410,
    n115,
    n273,
    n100
  );


  nor
  g518
  (
    n431,
    n161,
    n276,
    n247,
    n118
  );


  and
  g519
  (
    n462,
    n240,
    n99,
    n175,
    n174
  );


  and
  g520
  (
    n455,
    n289,
    n113,
    n109,
    n107
  );


  nor
  g521
  (
    n523,
    n391,
    n167,
    n408,
    n98
  );


  nand
  g522
  (
    n480,
    n392,
    n153,
    n404,
    n180
  );


  xnor
  g523
  (
    n537,
    n420,
    n104,
    n196,
    n172
  );


  not
  g524
  (
    n555,
    n424
  );


  not
  g525
  (
    n557,
    n429
  );


  not
  g526
  (
    n553,
    n423
  );


  not
  g527
  (
    n552,
    n426
  );


  not
  g528
  (
    n550,
    n422
  );


  not
  g529
  (
    n551,
    n421
  );


  buf
  g530
  (
    n556,
    n430
  );


  not
  g531
  (
    n549,
    n428
  );


  not
  g532
  (
    n554,
    n425
  );


  buf
  g533
  (
    n558,
    n427
  );


  xnor
  g534
  (
    n563,
    n293,
    n305,
    n300
  );


  xnor
  g535
  (
    n569,
    n326,
    n299,
    n558,
    n302
  );


  nor
  g536
  (
    n560,
    n329,
    n331,
    n330,
    n310
  );


  nor
  g537
  (
    n565,
    n550,
    n334,
    n552,
    n304
  );


  nand
  g538
  (
    KeyWire_0_52,
    n315,
    n322,
    n327,
    n333
  );


  nor
  g539
  (
    n572,
    n312,
    n306,
    n553,
    n308
  );


  xor
  g540
  (
    KeyWire_0_37,
    n556,
    n323,
    n558
  );


  nand
  g541
  (
    n564,
    n551,
    n311,
    n294,
    n324
  );


  xnor
  g542
  (
    n573,
    n321,
    n555,
    n296,
    n557
  );


  xor
  g543
  (
    n570,
    n332,
    n317,
    n335,
    n309
  );


  xnor
  g544
  (
    KeyWire_0_56,
    n295,
    n307,
    n557,
    n554
  );


  nand
  g545
  (
    n568,
    n432,
    n320,
    n557,
    n558
  );


  or
  g546
  (
    n571,
    n325,
    n291,
    n298,
    n557
  );


  or
  g547
  (
    n559,
    n297,
    n292,
    n319,
    n313
  );


  xnor
  g548
  (
    n561,
    n431,
    n318,
    n314,
    n303
  );


  xnor
  g549
  (
    n562,
    n316,
    n301,
    n328,
    n549
  );


  xnor
  g550
  (
    n597,
    n479,
    n339,
    n366,
    n483
  );


  nor
  g551
  (
    n586,
    n477,
    n562,
    n494,
    n485
  );


  xnor
  g552
  (
    n606,
    n356,
    n565,
    n488,
    n492
  );


  and
  g553
  (
    n599,
    n492,
    n570,
    n489,
    n572
  );


  or
  g554
  (
    KeyWire_0_7,
    n449,
    n484,
    n436
  );


  xnor
  g555
  (
    n590,
    n367,
    n489,
    n491,
    n561
  );


  nor
  g556
  (
    n630,
    n482,
    n496,
    n490,
    n434
  );


  nand
  g557
  (
    n602,
    n487,
    n447,
    n441,
    n457
  );


  nand
  g558
  (
    n598,
    n357,
    n440,
    n451,
    n485
  );


  and
  g559
  (
    n631,
    n344,
    n350,
    n493,
    n567
  );


  nor
  g560
  (
    n587,
    n384,
    n358,
    n488,
    n495
  );


  or
  g561
  (
    n625,
    n355,
    n483,
    n573,
    n559
  );


  nor
  g562
  (
    n635,
    n571,
    n480,
    n380,
    n385
  );


  xor
  g563
  (
    KeyWire_0_61,
    n349,
    n453,
    n559,
    n384
  );


  xnor
  g564
  (
    n634,
    n570,
    n572,
    n473,
    n476
  );


  or
  g565
  (
    n575,
    n450,
    n464,
    n572,
    n477
  );


  xnor
  g566
  (
    n591,
    n563,
    n471,
    n378,
    n495
  );


  nor
  g567
  (
    n604,
    n444,
    n571,
    n562,
    n567
  );


  nand
  g568
  (
    KeyWire_0_10,
    n346,
    n478,
    n351,
    n574
  );


  nand
  g569
  (
    n622,
    n560,
    n488,
    n561,
    n490
  );


  xnor
  g570
  (
    n579,
    n562,
    n564,
    n570,
    n495
  );


  or
  g571
  (
    KeyWire_0_40,
    n475,
    n480,
    n568,
    n463
  );


  or
  g572
  (
    n610,
    n479,
    n560,
    n377,
    n488
  );


  nor
  g573
  (
    n637,
    n570,
    n120,
    n470,
    n480
  );


  xnor
  g574
  (
    n624,
    n475,
    n561,
    n486,
    n383
  );


  nor
  g575
  (
    n612,
    n485,
    n559,
    n363,
    n572
  );


  xnor
  g576
  (
    n607,
    n364,
    n448,
    n567,
    n385
  );


  and
  g577
  (
    n617,
    n382,
    n368,
    n491,
    n459
  );


  and
  g578
  (
    n615,
    n492,
    n574,
    n566,
    n342
  );


  or
  g579
  (
    n588,
    n462,
    n569,
    n490,
    n493
  );


  xor
  g580
  (
    n577,
    n566,
    n567,
    n438,
    n472
  );


  and
  g581
  (
    n638,
    n484,
    n481,
    n371,
    n569
  );


  nor
  g582
  (
    KeyWire_0_18,
    n466,
    n484,
    n370,
    n372
  );


  xor
  g583
  (
    n608,
    n347,
    n348,
    n569,
    n475
  );


  xor
  g584
  (
    n583,
    n456,
    n341,
    n383,
    n483
  );


  nand
  g585
  (
    n580,
    n566,
    n560,
    n433,
    n493
  );


  nand
  g586
  (
    n629,
    n487,
    n465,
    n337,
    n446
  );


  or
  g587
  (
    n595,
    n494,
    n375,
    n573,
    n477
  );


  nor
  g588
  (
    n619,
    n478,
    n476,
    n452,
    n361
  );


  xnor
  g589
  (
    n601,
    n385,
    n481,
    n353,
    n574
  );


  nand
  g590
  (
    n589,
    n485,
    n365,
    n491,
    n474
  );


  xnor
  g591
  (
    n584,
    n486,
    n384,
    n482,
    n474
  );


  or
  g592
  (
    n613,
    n571,
    n455,
    n486
  );


  nor
  g593
  (
    n616,
    n566,
    n120,
    n474,
    n483
  );


  xnor
  g594
  (
    n585,
    n482,
    n383,
    n564,
    n569
  );


  or
  g595
  (
    n581,
    n571,
    n564,
    n381,
    n445
  );


  xnor
  g596
  (
    n614,
    n376,
    n383,
    n494,
    n565
  );


  nor
  g597
  (
    KeyWire_0_55,
    n565,
    n336,
    n489,
    n373
  );


  xnor
  g598
  (
    n611,
    n563,
    n481,
    n478,
    n493
  );


  or
  g599
  (
    n596,
    n460,
    n360,
    n382,
    n362
  );


  xor
  g600
  (
    n620,
    n487,
    n561,
    n468,
    n479
  );


  and
  g601
  (
    n582,
    n482,
    n492,
    n479,
    n474
  );


  nor
  g602
  (
    n626,
    n568,
    n568,
    n345,
    n354
  );


  nor
  g603
  (
    n623,
    n487,
    n491,
    n477,
    n559
  );


  xnor
  g604
  (
    n628,
    n469,
    n338,
    n563,
    n476
  );


  nor
  g605
  (
    n605,
    n120,
    n475,
    n480,
    n562
  );


  nor
  g606
  (
    n633,
    n442,
    n458,
    n384,
    n573
  );


  nor
  g607
  (
    n603,
    n443,
    n461,
    n489,
    n478
  );


  nand
  g608
  (
    n632,
    n340,
    n490,
    n481,
    n359
  );


  nor
  g609
  (
    n600,
    n369,
    n564,
    n439,
    n573
  );


  xnor
  g610
  (
    n576,
    n568,
    n435,
    n467,
    n454
  );


  nor
  g611
  (
    n593,
    n476,
    n379,
    n343,
    n495
  );


  and
  g612
  (
    n618,
    n565,
    n574,
    n437,
    n374
  );


  and
  g613
  (
    KeyWire_0_8,
    n352,
    n563,
    n494,
    n560
  );


  xor
  g614
  (
    KeyWire_0_57,
    n621,
    n633,
    n542
  );


  and
  g615
  (
    KeyWire_0_16,
    n537,
    n516,
    n631,
    n499
  );


  xor
  g616
  (
    n666,
    n638,
    n531,
    n504,
    n511
  );


  xor
  g617
  (
    n647,
    n519,
    n511,
    n530,
    n527
  );


  and
  g618
  (
    n655,
    n498,
    n529,
    n525,
    n499
  );


  xor
  g619
  (
    n639,
    n527,
    n530,
    n584,
    n388
  );


  nand
  g620
  (
    n677,
    n517,
    n531,
    n619,
    n519
  );


  xnor
  g621
  (
    n669,
    n541,
    n512,
    n548,
    n540
  );


  xnor
  g622
  (
    n683,
    n542,
    n635,
    n497,
    n540
  );


  nand
  g623
  (
    n694,
    n523,
    n507,
    n385,
    n513
  );


  xor
  g624
  (
    KeyWire_0_29,
    n525,
    n501,
    n537,
    n504
  );


  xnor
  g625
  (
    n697,
    n505,
    n631,
    n538,
    n544
  );


  and
  g626
  (
    n654,
    n634,
    n628,
    n521,
    n510
  );


  nor
  g627
  (
    n675,
    n630,
    n612,
    n544,
    n506
  );


  xor
  g628
  (
    n678,
    n387,
    n526,
    n545,
    n578
  );


  nand
  g629
  (
    n709,
    n507,
    n625,
    n526,
    n590
  );


  nand
  g630
  (
    n688,
    n507,
    n536,
    n520,
    n636
  );


  nor
  g631
  (
    n708,
    n522,
    n496,
    n633,
    n535
  );


  or
  g632
  (
    n679,
    n530,
    n509,
    n536,
    n635
  );


  or
  g633
  (
    n652,
    n513,
    n534,
    n538,
    n501
  );


  or
  g634
  (
    n700,
    n515,
    n501,
    n508,
    n614
  );


  xor
  g635
  (
    n644,
    n615,
    n534,
    n528,
    n637
  );


  and
  g636
  (
    n714,
    n623,
    n602,
    n502,
    n513
  );


  xor
  g637
  (
    n650,
    n535,
    n581,
    n499,
    n526
  );


  xor
  g638
  (
    n640,
    n511,
    n534,
    n503,
    n527
  );


  nor
  g639
  (
    n712,
    n512,
    n636,
    n500,
    n632
  );


  xnor
  g640
  (
    n692,
    n630,
    n616,
    n547,
    n512
  );


  nor
  g641
  (
    n641,
    n386,
    n536,
    n591,
    n496
  );


  nor
  g642
  (
    n667,
    n502,
    n524,
    n533
  );


  or
  g643
  (
    n687,
    n548,
    n523,
    n601,
    n630
  );


  nand
  g644
  (
    KeyWire_0_3,
    n508,
    n522,
    n521,
    n520
  );


  or
  g645
  (
    n686,
    n543,
    n527,
    n537,
    n498
  );


  xor
  g646
  (
    n681,
    n596,
    n524,
    n546,
    n637
  );


  nor
  g647
  (
    n702,
    n617,
    n636,
    n387,
    n522
  );


  xor
  g648
  (
    n704,
    n543,
    n541,
    n577,
    n538
  );


  xor
  g649
  (
    n685,
    n635,
    n629,
    n502,
    n519
  );


  and
  g650
  (
    n718,
    n626,
    n519,
    n634,
    n605
  );


  nor
  g651
  (
    n707,
    n498,
    n628,
    n585,
    n580
  );


  nand
  g652
  (
    n656,
    n515,
    n637,
    n387,
    n636
  );


  xnor
  g653
  (
    KeyWire_0_4,
    n542,
    n386,
    n515,
    n518
  );


  nor
  g654
  (
    n711,
    n620,
    n516,
    n505,
    n544
  );


  xnor
  g655
  (
    n664,
    n627,
    n624,
    n508,
    n517
  );


  nand
  g656
  (
    n663,
    n388,
    n510,
    n517,
    n496
  );


  and
  g657
  (
    n649,
    n539,
    n388,
    n632,
    n528
  );


  or
  g658
  (
    n705,
    n515,
    n511,
    n545,
    n629
  );


  xor
  g659
  (
    n710,
    n509,
    n540,
    n530,
    n630
  );


  xnor
  g660
  (
    n651,
    n631,
    n535,
    n547,
    n506
  );


  or
  g661
  (
    n716,
    n528,
    n547,
    n512,
    n506
  );


  xor
  g662
  (
    n715,
    n388,
    n387,
    n516,
    n503
  );


  nand
  g663
  (
    KeyWire_0_23,
    n522,
    n606,
    n542,
    n539
  );


  xnor
  g664
  (
    n642,
    n541,
    n546,
    n521,
    n507
  );


  xnor
  g665
  (
    n690,
    n505,
    n607,
    n587,
    n531
  );


  nor
  g666
  (
    n698,
    n532,
    n638,
    n548,
    n597
  );


  and
  g667
  (
    n674,
    n618,
    n535,
    n503,
    n613
  );


  and
  g668
  (
    n701,
    n510,
    n622,
    n505,
    n545
  );


  nand
  g669
  (
    n661,
    n548,
    n599,
    n540,
    n603
  );


  xor
  g670
  (
    n646,
    n631,
    n637,
    n506,
    n529
  );


  xnor
  g671
  (
    n676,
    n531,
    n529,
    n386,
    n532
  );


  nand
  g672
  (
    n684,
    n594,
    n576,
    n582,
    n520
  );


  nor
  g673
  (
    n657,
    n510,
    n501,
    n517,
    n588
  );


  and
  g674
  (
    n682,
    n503,
    n497,
    n523,
    n524
  );


  nor
  g675
  (
    n643,
    n529,
    n539,
    n523,
    n600
  );


  and
  g676
  (
    n717,
    n537,
    n514,
    n532,
    n525
  );


  nor
  g677
  (
    n659,
    n498,
    n518,
    n521,
    n538
  );


  xnor
  g678
  (
    n703,
    n545,
    n509,
    n539,
    n638
  );


  or
  g679
  (
    n680,
    n513,
    n575,
    n497,
    n546
  );


  or
  g680
  (
    KeyWire_0_33,
    n546,
    n518,
    n543,
    n533
  );


  nor
  g681
  (
    n673,
    n518,
    n632,
    n533,
    n586
  );


  xnor
  g682
  (
    n706,
    n635,
    n528,
    n604,
    n516
  );


  nand
  g683
  (
    n689,
    n543,
    n633,
    n611,
    n589
  );


  or
  g684
  (
    n653,
    n638,
    n499,
    n627,
    n526
  );


  nand
  g685
  (
    n648,
    n532,
    n508,
    n609,
    n610
  );


  and
  g686
  (
    n693,
    n579,
    n500,
    n541,
    n634
  );


  and
  g687
  (
    n668,
    n598,
    n592,
    n544,
    n608
  );


  or
  g688
  (
    n645,
    n504,
    n502,
    n595,
    n634
  );


  nand
  g689
  (
    n658,
    n536,
    n629,
    n583,
    n386
  );


  and
  g690
  (
    KeyWire_0_19,
    n509,
    n534,
    n629,
    n593
  );


  nand
  g691
  (
    n672,
    n520,
    n504,
    n547,
    n525
  );


  nor
  g692
  (
    n671,
    n500,
    n497,
    n514,
    n533
  );


  xor
  g693
  (
    n695,
    n632,
    n500,
    n514
  );


  nor
  g694
  (
    n731,
    n674,
    n664,
    n680,
    n708
  );


  xor
  g695
  (
    n734,
    n703,
    n685,
    n695,
    n655
  );


  and
  g696
  (
    n732,
    n704,
    n656,
    n699,
    n642
  );


  nand
  g697
  (
    n724,
    n661,
    n673,
    n714,
    n707
  );


  nor
  g698
  (
    n726,
    n698,
    n696,
    n665,
    n706
  );


  nor
  g699
  (
    n737,
    n718,
    n660,
    n640,
    n670
  );


  nor
  g700
  (
    n730,
    n666,
    n643,
    n667,
    n713
  );


  nor
  g701
  (
    n733,
    n689,
    n645,
    n668,
    n697
  );


  nor
  g702
  (
    n722,
    n694,
    n710,
    n717,
    n715
  );


  or
  g703
  (
    n738,
    n671,
    n663,
    n678,
    n675
  );


  or
  g704
  (
    n735,
    n650,
    n676,
    n691,
    n652
  );


  or
  g705
  (
    n728,
    n639,
    n709,
    n690,
    n651
  );


  or
  g706
  (
    n723,
    n688,
    n711,
    n684,
    n692
  );


  nor
  g707
  (
    n719,
    n644,
    n647,
    n679,
    n712
  );


  and
  g708
  (
    n720,
    n669,
    n705,
    n682,
    n657
  );


  or
  g709
  (
    n736,
    n641,
    n654,
    n672,
    n653
  );


  and
  g710
  (
    n725,
    n677,
    n683,
    n693,
    n687
  );


  or
  g711
  (
    n727,
    n686,
    n648,
    n649,
    n700
  );


  and
  g712
  (
    KeyWire_0_5,
    n646,
    n681,
    n702,
    n701
  );


  nand
  g713
  (
    n729,
    n662,
    n716,
    n659,
    n658
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n494,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n25,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n284,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n660,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n662,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n721,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n68,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n594,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n621,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n545,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n636,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n245,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n274,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n63,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n249,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n46,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n665,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n118,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n627,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n699,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n176,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n230,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n84,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n691,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n93,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n72,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n525,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n142,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n524,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n670,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n324,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n220,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n281,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n713,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n448,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n251,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n492,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n574,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n170,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n325,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n578,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n398,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n479,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n496,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n382,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n127,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n196,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n66,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n460,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n242,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n92,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n223,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n567,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n548,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n188,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n609,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n566,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n696,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n521,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n443,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n387,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n592,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n331,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n352,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

