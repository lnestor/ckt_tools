

module Stat_100_59
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n90,
  n113,
  n105,
  n89,
  n92,
  n114,
  n94,
  n118,
  n82,
  n88,
  n111,
  n102,
  n95,
  n119,
  n110,
  n93,
  n101,
  n87,
  n91,
  n97,
  n86,
  n98,
  n107,
  n106,
  n112,
  n117,
  n123,
  n130,
  n132,
  n128,
  n131,
  n129,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n90;
  output n113;
  output n105;
  output n89;
  output n92;
  output n114;
  output n94;
  output n118;
  output n82;
  output n88;
  output n111;
  output n102;
  output n95;
  output n119;
  output n110;
  output n93;
  output n101;
  output n87;
  output n91;
  output n97;
  output n86;
  output n98;
  output n107;
  output n106;
  output n112;
  output n117;
  output n123;
  output n130;
  output n132;
  output n128;
  output n131;
  output n129;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n83;
  wire n84;
  wire n85;
  wire n96;
  wire n99;
  wire n100;
  wire n103;
  wire n104;
  wire n108;
  wire n109;
  wire n115;
  wire n116;
  wire n120;
  wire n121;
  wire n122;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n68,
    n17
  );


  buf
  g1
  (
    KeyWire_0_48,
    n30
  );


  buf
  g2
  (
    KeyWire_0_54,
    n30
  );


  buf
  g3
  (
    n34,
    n6
  );


  not
  g4
  (
    KeyWire_0_20,
    n31
  );


  not
  g5
  (
    n64,
    n14
  );


  buf
  g6
  (
    KeyWire_0_38,
    n11
  );


  not
  g7
  (
    KeyWire_0_33,
    n26
  );


  buf
  g8
  (
    KeyWire_0_9,
    n31
  );


  buf
  g9
  (
    KeyWire_0_34,
    n5
  );


  not
  g10
  (
    KeyWire_0_13,
    n24
  );


  buf
  g11
  (
    n61,
    n23
  );


  buf
  g12
  (
    KeyWire_0_2,
    n32
  );


  not
  g13
  (
    n54,
    n9
  );


  not
  g14
  (
    KeyWire_0_12,
    n18
  );


  buf
  g15
  (
    n71,
    n8
  );


  buf
  g16
  (
    KeyWire_0_58,
    n21
  );


  buf
  g17
  (
    n65,
    n7
  );


  buf
  g18
  (
    n40,
    n20
  );


  not
  g19
  (
    n56,
    n31
  );


  not
  g20
  (
    KeyWire_0_16,
    n15
  );


  not
  g21
  (
    KeyWire_0_24,
    n32
  );


  buf
  g22
  (
    KeyWire_0_11,
    n28
  );


  buf
  g23
  (
    KeyWire_0_1,
    n10
  );


  not
  g24
  (
    KeyWire_0_46,
    n13
  );


  buf
  g25
  (
    n52,
    n12
  );


  not
  g26
  (
    KeyWire_0_43,
    n4
  );


  not
  g27
  (
    KeyWire_0_6,
    n22
  );


  buf
  g28
  (
    n67,
    n2
  );


  buf
  g29
  (
    n59,
    n19
  );


  not
  g30
  (
    n41,
    n29
  );


  buf
  g31
  (
    KeyWire_0_52,
    n25
  );


  not
  g32
  (
    n46,
    n30
  );


  not
  g33
  (
    n60,
    n3
  );


  not
  g34
  (
    n39,
    n1
  );


  buf
  g35
  (
    KeyWire_0_21,
    n27
  );


  buf
  g36
  (
    KeyWire_0_35,
    n31
  );


  buf
  g37
  (
    KeyWire_0_63,
    n32
  );


  buf
  g38
  (
    KeyWire_0_60,
    n16
  );


  not
  g39
  (
    n73,
    n35
  );


  not
  g40
  (
    n76,
    n37
  );


  not
  g41
  (
    n75,
    n37
  );


  not
  g42
  (
    n80,
    n34
  );


  not
  g43
  (
    KeyWire_0_44,
    n36
  );


  not
  g44
  (
    KeyWire_0_17,
    n37
  );


  not
  g45
  (
    KeyWire_0_19,
    n33
  );


  not
  g46
  (
    KeyWire_0_26,
    n36
  );


  buf
  g47
  (
    n72,
    n38
  );


  not
  g48
  (
    KeyWire_0_22,
    n36
  );


  or
  g49
  (
    KeyWire_0_27,
    n76,
    n60,
    n72,
    n59
  );


  xor
  g50
  (
    KeyWire_0_18,
    n60,
    n75,
    n80,
    n48
  );


  or
  g51
  (
    n106,
    n57,
    n56,
    n42,
    n74
  );


  and
  g52
  (
    KeyWire_0_36,
    n57,
    n74,
    n65,
    n44
  );


  nand
  g53
  (
    KeyWire_0_28,
    n43,
    n47,
    n41,
    n46
  );


  or
  g54
  (
    KeyWire_0_47,
    n57,
    n79,
    n80,
    n58
  );


  xor
  g55
  (
    KeyWire_0_4,
    n66,
    n73,
    n46,
    n40
  );


  nand
  g56
  (
    KeyWire_0_23,
    n39,
    n58,
    n55,
    n78
  );


  xnor
  g57
  (
    KeyWire_0_25,
    n63,
    n54,
    n56,
    n46
  );


  xor
  g58
  (
    KeyWire_0_59,
    n66,
    n42,
    n62,
    n77
  );


  nand
  g59
  (
    KeyWire_0_42,
    n50,
    n47,
    n40,
    n79
  );


  xnor
  g60
  (
    KeyWire_0_0,
    n44,
    n47,
    n56,
    n49
  );


  nor
  g61
  (
    n114,
    n78,
    n81,
    n48,
    n40
  );


  or
  g62
  (
    KeyWire_0_50,
    n51,
    n43,
    n48,
    n64
  );


  or
  g63
  (
    KeyWire_0_10,
    n43,
    n66,
    n77,
    n42
  );


  xor
  g64
  (
    KeyWire_0_55,
    n55,
    n57,
    n74,
    n47
  );


  nand
  g65
  (
    n97,
    n58,
    n63,
    n53,
    n51
  );


  nand
  g66
  (
    KeyWire_0_49,
    n56,
    n52,
    n45,
    n75
  );


  nor
  g67
  (
    KeyWire_0_5,
    n61,
    n53,
    n39,
    n54
  );


  or
  g68
  (
    KeyWire_0_29,
    n50,
    n78,
    n41,
    n73
  );


  nor
  g69
  (
    n83,
    n46,
    n80,
    n58,
    n49
  );


  nor
  g70
  (
    KeyWire_0_3,
    n67,
    n78,
    n81,
    n49
  );


  xor
  g71
  (
    n104,
    n48,
    n53,
    n67
  );


  xor
  g72
  (
    KeyWire_0_7,
    n77,
    n60,
    n76,
    n44
  );


  xor
  g73
  (
    KeyWire_0_62,
    n63,
    n50,
    n64,
    n39
  );


  and
  g74
  (
    KeyWire_0_41,
    n79,
    n79,
    n40,
    n72
  );


  xor
  g75
  (
    KeyWire_0_14,
    n44,
    n39,
    n67,
    n66
  );


  or
  g76
  (
    n107,
    n49,
    n73,
    n54,
    n77
  );


  or
  g77
  (
    KeyWire_0_51,
    n61,
    n81,
    n72
  );


  nand
  g78
  (
    n116,
    n74,
    n42,
    n45,
    n38
  );


  xor
  g79
  (
    KeyWire_0_53,
    n55,
    n52,
    n68,
    n75
  );


  or
  g80
  (
    KeyWire_0_32,
    n67,
    n50,
    n55,
    n72
  );


  and
  g81
  (
    KeyWire_0_15,
    n65,
    n52,
    n45,
    n38
  );


  xnor
  g82
  (
    KeyWire_0_8,
    n80,
    n59,
    n64,
    n75
  );


  or
  g83
  (
    n109,
    n76,
    n61,
    n63,
    n38
  );


  and
  g84
  (
    KeyWire_0_57,
    n76,
    n65,
    n59,
    n41
  );


  nor
  g85
  (
    n102,
    n65,
    n61,
    n62,
    n59
  );


  xor
  g86
  (
    KeyWire_0_37,
    n51,
    n43,
    n64,
    n54
  );


  nor
  g87
  (
    KeyWire_0_45,
    n62,
    n62,
    n73,
    n51
  );


  nand
  g88
  (
    n85,
    n60,
    n41,
    n45,
    n52
  );


  not
  g89
  (
    KeyWire_0_56,
    n116
  );


  not
  g90
  (
    KeyWire_0_40,
    n120
  );


  not
  g91
  (
    KeyWire_0_39,
    n118
  );


  nand
  g92
  (
    n124,
    n117,
    n32,
    n119,
    n110
  );


  and
  g93
  (
    KeyWire_0_30,
    n113,
    n109,
    n121,
    n115
  );


  nor
  g94
  (
    n127,
    n112,
    n114,
    n111,
    n108
  );


  nand
  g95
  (
    KeyWire_0_61,
    n69,
    n71,
    n126,
    n125
  );


  or
  g96
  (
    KeyWire_0_31,
    n71,
    n69
  );


  or
  g97
  (
    n128,
    n68,
    n70,
    n123,
    n69
  );


  xor
  g98
  (
    n132,
    n71,
    n68,
    n70
  );


  and
  g99
  (
    n129,
    n124,
    n70,
    n68,
    n127
  );


  xor
  KeyGate_0_0
  (
    n87,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n62,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n51,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n119,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n82,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n112,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n70,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n110,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n89,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n42,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n108,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n50,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n38,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n36,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n121,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n111,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n66,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n77,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n92,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n81,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n53,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n57,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n79,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n86,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n49,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n115,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n74,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n91,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n88,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n90,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n125,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n131,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n100,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n35,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n37,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n45,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n84,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n118,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n63,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n126,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n123,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n94,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n120,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n43,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n78,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n101,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n33,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n103,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n58,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n113,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n95,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n98,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n47,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n93,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n55,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n117,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n122,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n96,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n44,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n105,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n69,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n130,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n99,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n48,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

