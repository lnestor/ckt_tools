

module Stat_2000_202
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n659,
  n657,
  n632,
  n660,
  n627,
  n654,
  n644,
  n628,
  n634,
  n635,
  n646,
  n641,
  n648,
  n661,
  n652,
  n624,
  n906,
  n900,
  n896,
  n910,
  n983,
  n958,
  n1006,
  n973,
  n1017,
  n999,
  n976,
  n1011,
  n967,
  n1943,
  n2031,
  n2032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n659;
  output n657;
  output n632;
  output n660;
  output n627;
  output n654;
  output n644;
  output n628;
  output n634;
  output n635;
  output n646;
  output n641;
  output n648;
  output n661;
  output n652;
  output n624;
  output n906;
  output n900;
  output n896;
  output n910;
  output n983;
  output n958;
  output n1006;
  output n973;
  output n1017;
  output n999;
  output n976;
  output n1011;
  output n967;
  output n1943;
  output n2031;
  output n2032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n625;
  wire n626;
  wire n629;
  wire n630;
  wire n631;
  wire n633;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n642;
  wire n643;
  wire n645;
  wire n647;
  wire n649;
  wire n650;
  wire n651;
  wire n653;
  wire n655;
  wire n656;
  wire n658;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n897;
  wire n898;
  wire n899;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n907;
  wire n908;
  wire n909;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n974;
  wire n975;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n53,
    n26
  );


  buf
  g1
  (
    n125,
    n9
  );


  not
  g2
  (
    n127,
    n4
  );


  not
  g3
  (
    n132,
    n6
  );


  not
  g4
  (
    n99,
    n2
  );


  not
  g5
  (
    n155,
    n14
  );


  not
  g6
  (
    n74,
    n12
  );


  not
  g7
  (
    n76,
    n13
  );


  not
  g8
  (
    n55,
    n20
  );


  buf
  g9
  (
    n157,
    n18
  );


  not
  g10
  (
    n34,
    n11
  );


  buf
  g11
  (
    n87,
    n21
  );


  buf
  g12
  (
    n41,
    n10
  );


  not
  g13
  (
    n129,
    n28
  );


  buf
  g14
  (
    n50,
    n26
  );


  buf
  g15
  (
    n150,
    n25
  );


  buf
  g16
  (
    n82,
    n5
  );


  buf
  g17
  (
    n63,
    n6
  );


  not
  g18
  (
    n124,
    n6
  );


  buf
  g19
  (
    n65,
    n18
  );


  buf
  g20
  (
    n66,
    n15
  );


  buf
  g21
  (
    n100,
    n4
  );


  buf
  g22
  (
    n151,
    n24
  );


  not
  g23
  (
    n89,
    n28
  );


  not
  g24
  (
    n137,
    n25
  );


  buf
  g25
  (
    n154,
    n1
  );


  not
  g26
  (
    n88,
    n7
  );


  not
  g27
  (
    n78,
    n30
  );


  buf
  g28
  (
    n85,
    n25
  );


  buf
  g29
  (
    n111,
    n32
  );


  buf
  g30
  (
    n112,
    n3
  );


  not
  g31
  (
    n62,
    n3
  );


  buf
  g32
  (
    n57,
    n11
  );


  buf
  g33
  (
    n49,
    n16
  );


  not
  g34
  (
    n70,
    n32
  );


  not
  g35
  (
    n114,
    n32
  );


  buf
  g36
  (
    n119,
    n29
  );


  buf
  g37
  (
    n71,
    n29
  );


  not
  g38
  (
    n102,
    n18
  );


  buf
  g39
  (
    n98,
    n32
  );


  not
  g40
  (
    n68,
    n17
  );


  not
  g41
  (
    n54,
    n19
  );


  buf
  g42
  (
    n156,
    n25
  );


  buf
  g43
  (
    n90,
    n21
  );


  buf
  g44
  (
    n46,
    n23
  );


  not
  g45
  (
    n149,
    n26
  );


  buf
  g46
  (
    n110,
    n1
  );


  not
  g47
  (
    n118,
    n27
  );


  not
  g48
  (
    n38,
    n5
  );


  not
  g49
  (
    n69,
    n22
  );


  not
  g50
  (
    n103,
    n29
  );


  not
  g51
  (
    n126,
    n14
  );


  buf
  g52
  (
    n133,
    n8
  );


  buf
  g53
  (
    n160,
    n29
  );


  buf
  g54
  (
    n59,
    n31
  );


  not
  g55
  (
    n152,
    n17
  );


  not
  g56
  (
    n141,
    n6
  );


  not
  g57
  (
    n113,
    n14
  );


  buf
  g58
  (
    n44,
    n24
  );


  buf
  g59
  (
    n61,
    n19
  );


  buf
  g60
  (
    n117,
    n3
  );


  not
  g61
  (
    n153,
    n12
  );


  not
  g62
  (
    n92,
    n31
  );


  not
  g63
  (
    n122,
    n4
  );


  buf
  g64
  (
    n115,
    n10
  );


  buf
  g65
  (
    KeyWire_0_2,
    n2
  );


  buf
  g66
  (
    n35,
    n11
  );


  not
  g67
  (
    n95,
    n16
  );


  not
  g68
  (
    n67,
    n7
  );


  not
  g69
  (
    n86,
    n5
  );


  not
  g70
  (
    n123,
    n22
  );


  buf
  g71
  (
    n72,
    n24
  );


  not
  g72
  (
    n77,
    n31
  );


  not
  g73
  (
    n60,
    n28
  );


  not
  g74
  (
    n33,
    n20
  );


  not
  g75
  (
    n64,
    n21
  );


  buf
  g76
  (
    n130,
    n10
  );


  buf
  g77
  (
    n91,
    n22
  );


  buf
  g78
  (
    n148,
    n11
  );


  not
  g79
  (
    n145,
    n7
  );


  not
  g80
  (
    n121,
    n23
  );


  buf
  g81
  (
    n37,
    n17
  );


  buf
  g82
  (
    n109,
    n9
  );


  not
  g83
  (
    n84,
    n31
  );


  not
  g84
  (
    n108,
    n15
  );


  not
  g85
  (
    n51,
    n8
  );


  not
  g86
  (
    n80,
    n9
  );


  buf
  g87
  (
    n107,
    n30
  );


  not
  g88
  (
    n75,
    n8
  );


  buf
  g89
  (
    n131,
    n24
  );


  buf
  g90
  (
    n42,
    n2
  );


  not
  g91
  (
    n116,
    n2
  );


  not
  g92
  (
    n93,
    n1
  );


  buf
  g93
  (
    n73,
    n20
  );


  not
  g94
  (
    n94,
    n17
  );


  buf
  g95
  (
    n45,
    n13
  );


  buf
  g96
  (
    n39,
    n18
  );


  not
  g97
  (
    n139,
    n30
  );


  buf
  g98
  (
    n147,
    n19
  );


  not
  g99
  (
    n97,
    n9
  );


  not
  g100
  (
    n40,
    n27
  );


  buf
  g101
  (
    n136,
    n21
  );


  buf
  g102
  (
    n144,
    n15
  );


  buf
  g103
  (
    n58,
    n26
  );


  buf
  g104
  (
    n36,
    n20
  );


  not
  g105
  (
    n142,
    n27
  );


  not
  g106
  (
    n48,
    n4
  );


  not
  g107
  (
    n81,
    n14
  );


  buf
  g108
  (
    n140,
    n13
  );


  buf
  g109
  (
    n104,
    n23
  );


  buf
  g110
  (
    n146,
    n15
  );


  not
  g111
  (
    KeyWire_0_1,
    n19
  );


  buf
  g112
  (
    n158,
    n3
  );


  buf
  g113
  (
    n83,
    n27
  );


  not
  g114
  (
    n101,
    n16
  );


  buf
  g115
  (
    n56,
    n23
  );


  buf
  g116
  (
    n143,
    n1
  );


  not
  g117
  (
    n105,
    n22
  );


  buf
  g118
  (
    n52,
    n16
  );


  buf
  g119
  (
    n128,
    n5
  );


  not
  g120
  (
    n106,
    n8
  );


  buf
  g121
  (
    n47,
    n7
  );


  not
  g122
  (
    n79,
    n13
  );


  not
  g123
  (
    n159,
    n28
  );


  buf
  g124
  (
    n120,
    n10
  );


  buf
  g125
  (
    n43,
    n12
  );


  buf
  g126
  (
    n134,
    n12
  );


  not
  g127
  (
    n96,
    n30
  );


  not
  g128
  (
    n331,
    n33
  );


  buf
  g129
  (
    n204,
    n48
  );


  not
  g130
  (
    n203,
    n71
  );


  buf
  g131
  (
    n293,
    n78
  );


  not
  g132
  (
    n248,
    n59
  );


  not
  g133
  (
    n229,
    n65
  );


  buf
  g134
  (
    n241,
    n62
  );


  not
  g135
  (
    n339,
    n56
  );


  buf
  g136
  (
    n260,
    n51
  );


  not
  g137
  (
    n325,
    n62
  );


  not
  g138
  (
    n302,
    n76
  );


  not
  g139
  (
    n333,
    n44
  );


  not
  g140
  (
    n242,
    n58
  );


  buf
  g141
  (
    n181,
    n68
  );


  buf
  g142
  (
    n163,
    n65
  );


  not
  g143
  (
    n244,
    n51
  );


  not
  g144
  (
    n271,
    n55
  );


  buf
  g145
  (
    n323,
    n64
  );


  buf
  g146
  (
    n250,
    n72
  );


  buf
  g147
  (
    n224,
    n67
  );


  not
  g148
  (
    n329,
    n42
  );


  not
  g149
  (
    n295,
    n42
  );


  not
  g150
  (
    n274,
    n37
  );


  not
  g151
  (
    n263,
    n45
  );


  buf
  g152
  (
    n230,
    n64
  );


  buf
  g153
  (
    n200,
    n48
  );


  buf
  g154
  (
    n187,
    n77
  );


  not
  g155
  (
    n313,
    n53
  );


  buf
  g156
  (
    n310,
    n33
  );


  buf
  g157
  (
    n175,
    n34
  );


  not
  g158
  (
    n220,
    n78
  );


  buf
  g159
  (
    n183,
    n76
  );


  buf
  g160
  (
    n177,
    n58
  );


  not
  g161
  (
    n174,
    n47
  );


  buf
  g162
  (
    n179,
    n54
  );


  not
  g163
  (
    n235,
    n44
  );


  not
  g164
  (
    n164,
    n56
  );


  not
  g165
  (
    n268,
    n35
  );


  not
  g166
  (
    n321,
    n54
  );


  not
  g167
  (
    n236,
    n70
  );


  not
  g168
  (
    n275,
    n57
  );


  buf
  g169
  (
    n217,
    n52
  );


  not
  g170
  (
    n211,
    n35
  );


  buf
  g171
  (
    n249,
    n46
  );


  not
  g172
  (
    n286,
    n70
  );


  buf
  g173
  (
    n305,
    n71
  );


  buf
  g174
  (
    n343,
    n72
  );


  not
  g175
  (
    n195,
    n57
  );


  buf
  g176
  (
    n266,
    n40
  );


  buf
  g177
  (
    n269,
    n43
  );


  not
  g178
  (
    n334,
    n71
  );


  not
  g179
  (
    n223,
    n79
  );


  buf
  g180
  (
    n345,
    n45
  );


  not
  g181
  (
    n228,
    n52
  );


  not
  g182
  (
    n327,
    n33
  );


  buf
  g183
  (
    n283,
    n40
  );


  buf
  g184
  (
    n280,
    n57
  );


  buf
  g185
  (
    n189,
    n61
  );


  not
  g186
  (
    n287,
    n63
  );


  not
  g187
  (
    n185,
    n46
  );


  not
  g188
  (
    n259,
    n74
  );


  buf
  g189
  (
    n320,
    n61
  );


  not
  g190
  (
    n208,
    n38
  );


  not
  g191
  (
    n328,
    n47
  );


  not
  g192
  (
    n316,
    n48
  );


  buf
  g193
  (
    n319,
    n60
  );


  buf
  g194
  (
    n344,
    n61
  );


  not
  g195
  (
    n304,
    n45
  );


  not
  g196
  (
    n289,
    n71
  );


  buf
  g197
  (
    n272,
    n33
  );


  buf
  g198
  (
    n258,
    n49
  );


  buf
  g199
  (
    n337,
    n73
  );


  buf
  g200
  (
    n335,
    n59
  );


  not
  g201
  (
    n265,
    n67
  );


  not
  g202
  (
    n308,
    n68
  );


  buf
  g203
  (
    n225,
    n58
  );


  buf
  g204
  (
    n199,
    n69
  );


  buf
  g205
  (
    n178,
    n66
  );


  not
  g206
  (
    n276,
    n38
  );


  not
  g207
  (
    n300,
    n76
  );


  not
  g208
  (
    n197,
    n78
  );


  buf
  g209
  (
    n284,
    n56
  );


  buf
  g210
  (
    n218,
    n41
  );


  not
  g211
  (
    n166,
    n41
  );


  not
  g212
  (
    n253,
    n50
  );


  buf
  g213
  (
    n309,
    n69
  );


  buf
  g214
  (
    n307,
    n35
  );


  not
  g215
  (
    n221,
    n78
  );


  buf
  g216
  (
    n246,
    n39
  );


  buf
  g217
  (
    n296,
    n61
  );


  not
  g218
  (
    n173,
    n79
  );


  buf
  g219
  (
    n194,
    n52
  );


  not
  g220
  (
    n182,
    n60
  );


  not
  g221
  (
    n215,
    n59
  );


  not
  g222
  (
    n167,
    n50
  );


  not
  g223
  (
    n170,
    n34
  );


  buf
  g224
  (
    n162,
    n49
  );


  not
  g225
  (
    n226,
    n62
  );


  not
  g226
  (
    n292,
    n55
  );


  not
  g227
  (
    n330,
    n65
  );


  not
  g228
  (
    n238,
    n55
  );


  buf
  g229
  (
    n227,
    n40
  );


  not
  g230
  (
    n172,
    n63
  );


  not
  g231
  (
    n188,
    n75
  );


  not
  g232
  (
    n257,
    n56
  );


  not
  g233
  (
    n267,
    n39
  );


  not
  g234
  (
    n186,
    n34
  );


  buf
  g235
  (
    n326,
    n77
  );


  buf
  g236
  (
    n212,
    n44
  );


  not
  g237
  (
    n322,
    n36
  );


  not
  g238
  (
    n243,
    n70
  );


  not
  g239
  (
    n306,
    n69
  );


  not
  g240
  (
    n240,
    n73
  );


  not
  g241
  (
    n340,
    n55
  );


  not
  g242
  (
    n288,
    n53
  );


  buf
  g243
  (
    n234,
    n34
  );


  buf
  g244
  (
    n324,
    n51
  );


  not
  g245
  (
    n303,
    n67
  );


  not
  g246
  (
    n279,
    n36
  );


  not
  g247
  (
    n256,
    n70
  );


  buf
  g248
  (
    n202,
    n59
  );


  buf
  g249
  (
    n201,
    n65
  );


  buf
  g250
  (
    n315,
    n63
  );


  buf
  g251
  (
    n252,
    n60
  );


  buf
  g252
  (
    n233,
    n52
  );


  buf
  g253
  (
    n314,
    n60
  );


  not
  g254
  (
    n318,
    n74
  );


  buf
  g255
  (
    n277,
    n41
  );


  buf
  g256
  (
    n176,
    n64
  );


  not
  g257
  (
    n262,
    n66
  );


  not
  g258
  (
    n180,
    n42
  );


  buf
  g259
  (
    n206,
    n43
  );


  buf
  g260
  (
    n161,
    n73
  );


  not
  g261
  (
    n285,
    n77
  );


  buf
  g262
  (
    n346,
    n38
  );


  not
  g263
  (
    n297,
    n73
  );


  buf
  g264
  (
    n261,
    n66
  );


  buf
  g265
  (
    n245,
    n46
  );


  buf
  g266
  (
    n222,
    n68
  );


  buf
  g267
  (
    n198,
    n44
  );


  not
  g268
  (
    n281,
    n62
  );


  buf
  g269
  (
    n301,
    n75
  );


  not
  g270
  (
    n171,
    n42
  );


  not
  g271
  (
    n291,
    n38
  );


  not
  g272
  (
    n273,
    n37
  );


  not
  g273
  (
    n254,
    n36
  );


  buf
  g274
  (
    n332,
    n47
  );


  not
  g275
  (
    n169,
    n35
  );


  not
  g276
  (
    n278,
    n43
  );


  not
  g277
  (
    n270,
    n39
  );


  buf
  g278
  (
    n191,
    n47
  );


  buf
  g279
  (
    n264,
    n72
  );


  not
  g280
  (
    n210,
    n39
  );


  buf
  g281
  (
    n338,
    n37
  );


  not
  g282
  (
    n192,
    n66
  );


  not
  g283
  (
    n255,
    n58
  );


  not
  g284
  (
    n282,
    n57
  );


  not
  g285
  (
    n232,
    n77
  );


  buf
  g286
  (
    n290,
    n63
  );


  buf
  g287
  (
    n251,
    n67
  );


  buf
  g288
  (
    n209,
    n41
  );


  buf
  g289
  (
    n207,
    n53
  );


  not
  g290
  (
    n237,
    n50
  );


  not
  g291
  (
    n205,
    n51
  );


  not
  g292
  (
    n165,
    n54
  );


  not
  g293
  (
    n216,
    n74
  );


  buf
  g294
  (
    n219,
    n43
  );


  buf
  g295
  (
    n342,
    n69
  );


  not
  g296
  (
    n168,
    n45
  );


  not
  g297
  (
    n213,
    n75
  );


  not
  g298
  (
    n193,
    n76
  );


  buf
  g299
  (
    n214,
    n64
  );


  buf
  g300
  (
    n184,
    n53
  );


  buf
  g301
  (
    n190,
    n50
  );


  not
  g302
  (
    n311,
    n40
  );


  buf
  g303
  (
    n299,
    n54
  );


  buf
  g304
  (
    n298,
    n72
  );


  not
  g305
  (
    n196,
    n49
  );


  not
  g306
  (
    n341,
    n37
  );


  buf
  g307
  (
    n336,
    n46
  );


  not
  g308
  (
    n294,
    n75
  );


  not
  g309
  (
    n231,
    n74
  );


  buf
  g310
  (
    n317,
    n49
  );


  not
  g311
  (
    n239,
    n48
  );


  not
  g312
  (
    n312,
    n68
  );


  buf
  g313
  (
    n247,
    n36
  );


  not
  g314
  (
    n608,
    n211
  );


  buf
  g315
  (
    n442,
    n287
  );


  not
  g316
  (
    n582,
    n124
  );


  buf
  g317
  (
    n418,
    n103
  );


  not
  g318
  (
    n507,
    n154
  );


  buf
  g319
  (
    n531,
    n270
  );


  buf
  g320
  (
    n443,
    n129
  );


  buf
  g321
  (
    n530,
    n142
  );


  buf
  g322
  (
    n532,
    n130
  );


  not
  g323
  (
    n552,
    n279
  );


  buf
  g324
  (
    n491,
    n290
  );


  buf
  g325
  (
    n524,
    n136
  );


  not
  g326
  (
    n371,
    n257
  );


  not
  g327
  (
    n470,
    n88
  );


  buf
  g328
  (
    n449,
    n208
  );


  buf
  g329
  (
    n489,
    n90
  );


  buf
  g330
  (
    n368,
    n125
  );


  not
  g331
  (
    n607,
    n189
  );


  buf
  g332
  (
    n559,
    n256
  );


  not
  g333
  (
    n444,
    n288
  );


  buf
  g334
  (
    n410,
    n115
  );


  buf
  g335
  (
    n372,
    n258
  );


  buf
  g336
  (
    n569,
    n180
  );


  not
  g337
  (
    n541,
    n254
  );


  buf
  g338
  (
    n590,
    n114
  );


  buf
  g339
  (
    n595,
    n247
  );


  not
  g340
  (
    n415,
    n240
  );


  buf
  g341
  (
    n610,
    n295
  );


  not
  g342
  (
    n562,
    n236
  );


  buf
  g343
  (
    n563,
    n95
  );


  buf
  g344
  (
    n367,
    n195
  );


  not
  g345
  (
    n550,
    n274
  );


  not
  g346
  (
    n479,
    n203
  );


  buf
  g347
  (
    n589,
    n126
  );


  buf
  g348
  (
    n515,
    n282
  );


  not
  g349
  (
    n476,
    n159
  );


  not
  g350
  (
    n574,
    n143
  );


  buf
  g351
  (
    n370,
    n241
  );


  not
  g352
  (
    n396,
    n98
  );


  buf
  g353
  (
    n452,
    n289
  );


  not
  g354
  (
    n510,
    n288
  );


  not
  g355
  (
    n435,
    n110
  );


  buf
  g356
  (
    n437,
    n211
  );


  not
  g357
  (
    n616,
    n93
  );


  buf
  g358
  (
    n394,
    n80
  );


  buf
  g359
  (
    n596,
    n131
  );


  buf
  g360
  (
    n555,
    n210
  );


  buf
  g361
  (
    n518,
    n183
  );


  not
  g362
  (
    n487,
    n243
  );


  not
  g363
  (
    n619,
    n141
  );


  not
  g364
  (
    n440,
    n265
  );


  not
  g365
  (
    n480,
    n141
  );


  not
  g366
  (
    n409,
    n93
  );


  buf
  g367
  (
    n420,
    n254
  );


  buf
  g368
  (
    n473,
    n253
  );


  not
  g369
  (
    n511,
    n127
  );


  not
  g370
  (
    n427,
    n230
  );


  not
  g371
  (
    n355,
    n136
  );


  buf
  g372
  (
    n502,
    n258
  );


  not
  g373
  (
    n430,
    n202
  );


  buf
  g374
  (
    n587,
    n92
  );


  buf
  g375
  (
    n349,
    n89
  );


  buf
  g376
  (
    n542,
    n213
  );


  buf
  g377
  (
    n615,
    n284
  );


  not
  g378
  (
    n408,
    n221
  );


  buf
  g379
  (
    n392,
    n91
  );


  buf
  g380
  (
    n465,
    n121
  );


  not
  g381
  (
    n428,
    n218
  );


  buf
  g382
  (
    n389,
    n251
  );


  buf
  g383
  (
    n477,
    n289
  );


  not
  g384
  (
    n348,
    n96
  );


  buf
  g385
  (
    n434,
    n155
  );


  buf
  g386
  (
    n528,
    n101
  );


  not
  g387
  (
    n436,
    n138
  );


  buf
  g388
  (
    n441,
    n99
  );


  buf
  g389
  (
    n475,
    n218
  );


  not
  g390
  (
    n454,
    n286
  );


  not
  g391
  (
    n356,
    n280
  );


  buf
  g392
  (
    n488,
    n184
  );


  buf
  g393
  (
    n404,
    n149
  );


  buf
  g394
  (
    n463,
    n186
  );


  not
  g395
  (
    n591,
    n89
  );


  buf
  g396
  (
    n469,
    n272
  );


  buf
  g397
  (
    n593,
    n281
  );


  buf
  g398
  (
    n503,
    n132
  );


  not
  g399
  (
    n419,
    n139
  );


  not
  g400
  (
    n519,
    n81
  );


  buf
  g401
  (
    n433,
    n235
  );


  buf
  g402
  (
    n594,
    n231
  );


  buf
  g403
  (
    n579,
    n156
  );


  buf
  g404
  (
    n352,
    n256
  );


  buf
  g405
  (
    n377,
    n263
  );


  not
  g406
  (
    n557,
    n275
  );


  buf
  g407
  (
    n583,
    n115
  );


  not
  g408
  (
    n597,
    n235
  );


  buf
  g409
  (
    n405,
    n120
  );


  buf
  g410
  (
    n584,
    n188
  );


  not
  g411
  (
    n588,
    n81
  );


  not
  g412
  (
    n570,
    n117
  );


  not
  g413
  (
    n585,
    n205
  );


  not
  g414
  (
    n421,
    n110
  );


  not
  g415
  (
    n361,
    n118
  );


  buf
  g416
  (
    n453,
    n265
  );


  not
  g417
  (
    n397,
    n200
  );


  not
  g418
  (
    n412,
    n80
  );


  buf
  g419
  (
    n496,
    n106
  );


  not
  g420
  (
    n575,
    n145
  );


  buf
  g421
  (
    n380,
    n279
  );


  buf
  g422
  (
    n606,
    n118
  );


  not
  g423
  (
    n544,
    n130
  );


  buf
  g424
  (
    n572,
    n281
  );


  not
  g425
  (
    n536,
    n223
  );


  not
  g426
  (
    n383,
    n276
  );


  buf
  g427
  (
    n365,
    n251
  );


  buf
  g428
  (
    n450,
    n139
  );


  not
  g429
  (
    n603,
    n105
  );


  buf
  g430
  (
    n534,
    n107
  );


  not
  g431
  (
    n364,
    n205
  );


  not
  g432
  (
    n484,
    n114
  );


  not
  g433
  (
    n467,
    n113
  );


  buf
  g434
  (
    n546,
    n113
  );


  not
  g435
  (
    n540,
    n148
  );


  not
  g436
  (
    n390,
    n90
  );


  buf
  g437
  (
    n611,
    n246
  );


  not
  g438
  (
    n612,
    n273
  );


  buf
  g439
  (
    n353,
    n143
  );


  buf
  g440
  (
    n400,
    n107
  );


  buf
  g441
  (
    n369,
    n252
  );


  not
  g442
  (
    n567,
    n156
  );


  buf
  g443
  (
    n483,
    n144
  );


  not
  g444
  (
    n513,
    n285
  );


  buf
  g445
  (
    n547,
    n158
  );


  not
  g446
  (
    n388,
    n101
  );


  not
  g447
  (
    n517,
    n130
  );


  not
  g448
  (
    n432,
    n137
  );


  not
  g449
  (
    n514,
    n236
  );


  buf
  g450
  (
    n375,
    n247
  );


  not
  g451
  (
    n374,
    n92
  );


  buf
  g452
  (
    n499,
    n244
  );


  buf
  g453
  (
    n581,
    n84
  );


  buf
  g454
  (
    n521,
    n144
  );


  buf
  g455
  (
    n558,
    n245
  );


  not
  g456
  (
    n359,
    n98
  );


  buf
  g457
  (
    n573,
    n108
  );


  not
  g458
  (
    n598,
    n146
  );


  buf
  g459
  (
    n568,
    n85
  );


  buf
  g460
  (
    n527,
    n154
  );


  not
  g461
  (
    n577,
    n269
  );


  not
  g462
  (
    n347,
    n229
  );


  buf
  g463
  (
    n382,
    n145
  );


  not
  g464
  (
    n482,
    n257
  );


  buf
  g465
  (
    n578,
    n290
  );


  buf
  g466
  (
    n429,
    n134
  );


  not
  g467
  (
    n402,
    n263
  );


  buf
  g468
  (
    n509,
    n246
  );


  buf
  g469
  (
    n414,
    n130
  );


  not
  g470
  (
    n481,
    n87
  );


  not
  g471
  (
    n423,
    n133
  );


  not
  g472
  (
    n447,
    n234
  );


  buf
  g473
  (
    n529,
    n91
  );


  nor
  g474
  (
    n554,
    n292,
    n101,
    n90,
    n100
  );


  nor
  g475
  (
    n592,
    n296,
    n114,
    n177,
    n145
  );


  or
  g476
  (
    n399,
    n97,
    n277,
    n106,
    n185
  );


  nor
  g477
  (
    n537,
    n141,
    n198,
    n95,
    n127
  );


  xnor
  g478
  (
    n535,
    n261,
    n110,
    n138,
    n226
  );


  nand
  g479
  (
    n501,
    n224,
    n151,
    n79,
    n96
  );


  xnor
  g480
  (
    n354,
    n135,
    n132,
    n262,
    n198
  );


  and
  g481
  (
    n495,
    n121,
    n247,
    n81,
    n240
  );


  or
  g482
  (
    n520,
    n87,
    n181,
    n185,
    n115
  );


  xnor
  g483
  (
    n360,
    n282,
    n229,
    n102,
    n139
  );


  xor
  g484
  (
    n468,
    n90,
    n155,
    n183,
    n113
  );


  or
  g485
  (
    n600,
    n102,
    n293,
    n233,
    n210
  );


  nor
  g486
  (
    n466,
    n135,
    n125,
    n249,
    n284
  );


  nand
  g487
  (
    n508,
    n122,
    n137,
    n230,
    n81
  );


  and
  g488
  (
    n526,
    n270,
    n106,
    n107,
    n248
  );


  nor
  g489
  (
    n464,
    n228,
    n83,
    n151,
    n179
  );


  nor
  g490
  (
    n556,
    n212,
    n114,
    n136,
    n242
  );


  xor
  g491
  (
    n472,
    n148,
    n227,
    n184,
    n214
  );


  nor
  g492
  (
    n564,
    n112,
    n140,
    n157,
    n142
  );


  xor
  g493
  (
    n366,
    n116,
    n287,
    n283
  );


  nand
  g494
  (
    n500,
    n267,
    n111,
    n287,
    n192
  );


  xor
  g495
  (
    n586,
    n154,
    n194,
    n193,
    n273
  );


  nor
  g496
  (
    n460,
    n104,
    n201,
    n278,
    n217
  );


  xnor
  g497
  (
    n560,
    n233,
    n275,
    n142,
    n190
  );


  xor
  g498
  (
    n358,
    n268,
    n272,
    n278,
    n106
  );


  and
  g499
  (
    n457,
    n224,
    n103,
    n291,
    n134
  );


  xnor
  g500
  (
    n553,
    n294,
    n79,
    n128,
    n134
  );


  xor
  g501
  (
    n576,
    n182,
    n158,
    n115
  );


  nor
  g502
  (
    n492,
    n140,
    n132,
    n295,
    n197
  );


  nand
  g503
  (
    n494,
    n137,
    n225,
    n126,
    n279
  );


  xor
  g504
  (
    n566,
    n97,
    n89,
    n104,
    n290
  );


  nand
  g505
  (
    n406,
    n104,
    n112,
    n249,
    n262
  );


  nand
  g506
  (
    n545,
    n82,
    n244,
    n151,
    n105
  );


  nand
  g507
  (
    n571,
    n84,
    n269,
    n128,
    n131
  );


  xor
  g508
  (
    n373,
    n255,
    n199,
    n98,
    n249
  );


  xor
  g509
  (
    n613,
    n241,
    n264,
    n232,
    n121
  );


  nor
  g510
  (
    n471,
    n294,
    n296,
    n276,
    n128
  );


  or
  g511
  (
    n490,
    n269,
    n293,
    n239,
    n83
  );


  nand
  g512
  (
    n522,
    n237,
    n251,
    n207,
    n186
  );


  xor
  g513
  (
    n416,
    n255,
    n213,
    n120,
    n248
  );


  xnor
  g514
  (
    n381,
    n153,
    n191,
    n223,
    n96
  );


  xor
  g515
  (
    n474,
    n239,
    n286,
    n266,
    n117
  );


  xor
  g516
  (
    n618,
    n148,
    n103,
    n88,
    n86
  );


  nand
  g517
  (
    n533,
    n109,
    n84,
    n267,
    n129
  );


  and
  g518
  (
    n512,
    n149,
    n126,
    n87,
    n138
  );


  nand
  g519
  (
    n425,
    n209,
    n85,
    n242,
    n132
  );


  nor
  g520
  (
    n411,
    n111,
    n271,
    n144,
    n252
  );


  nand
  g521
  (
    n395,
    n291,
    n285,
    n284,
    n146
  );


  xnor
  g522
  (
    n431,
    n120,
    n189,
    n277,
    n85
  );


  nand
  g523
  (
    n580,
    n121,
    n82,
    n216,
    n125
  );


  nand
  g524
  (
    n561,
    n260,
    n119,
    n195,
    n110
  );


  xor
  g525
  (
    n357,
    n83,
    n138,
    n266,
    n259
  );


  nand
  g526
  (
    n378,
    n82,
    n94,
    n101,
    n149
  );


  xor
  g527
  (
    n549,
    n98,
    n212,
    n99,
    n147
  );


  xor
  g528
  (
    n505,
    n86,
    n262,
    n133,
    n144
  );


  xnor
  g529
  (
    n525,
    n158,
    n246,
    n257,
    n86
  );


  nor
  g530
  (
    n363,
    n153,
    n146,
    n143,
    n271
  );


  xor
  g531
  (
    n422,
    n91,
    n105,
    n120,
    n243
  );


  xnor
  g532
  (
    n461,
    n152,
    n260,
    n116,
    n202
  );


  or
  g533
  (
    n504,
    n252,
    n122,
    n295,
    n245
  );


  or
  g534
  (
    n403,
    n253,
    n95,
    n187,
    n125
  );


  and
  g535
  (
    n451,
    n150,
    n143,
    n153,
    n95
  );


  xnor
  g536
  (
    n448,
    n155,
    n237,
    n219,
    n197
  );


  and
  g537
  (
    n386,
    n228,
    n196,
    n234,
    n84
  );


  or
  g538
  (
    n497,
    n127,
    n219,
    n190,
    n118
  );


  xnor
  g539
  (
    n376,
    n275,
    n258,
    n221,
    n268
  );


  xnor
  g540
  (
    n506,
    n192,
    n127,
    n118,
    n199
  );


  nand
  g541
  (
    n362,
    n274,
    n281,
    n261,
    n100
  );


  nand
  g542
  (
    n614,
    n194,
    n292,
    n265,
    n150
  );


  or
  g543
  (
    n523,
    n232,
    n153,
    n93,
    n274
  );


  or
  g544
  (
    n458,
    n113,
    n244,
    n157,
    n250
  );


  nor
  g545
  (
    n393,
    n214,
    n286,
    n222,
    n282
  );


  and
  g546
  (
    n485,
    n159,
    n137,
    n294,
    n278
  );


  or
  g547
  (
    n401,
    n80,
    n141,
    n108,
    n260
  );


  and
  g548
  (
    n350,
    n225,
    n270,
    n83,
    n112
  );


  and
  g549
  (
    n417,
    n204,
    n291,
    n253,
    n261
  );


  nand
  g550
  (
    n424,
    n220,
    n243,
    n119,
    n104
  );


  xnor
  g551
  (
    n538,
    n111,
    n117,
    n92,
    n241
  );


  nand
  g552
  (
    n379,
    n135,
    n196,
    n248,
    n102
  );


  xnor
  g553
  (
    n462,
    n146,
    n94,
    n119
  );


  nor
  g554
  (
    n455,
    n123,
    n182,
    n107,
    n108
  );


  xnor
  g555
  (
    n609,
    n93,
    n250,
    n157,
    n124
  );


  xor
  g556
  (
    n565,
    n123,
    n191,
    n254,
    n82
  );


  xnor
  g557
  (
    n548,
    n216,
    n272,
    n129,
    n147
  );


  nand
  g558
  (
    n602,
    n208,
    n289,
    n207,
    n89
  );


  and
  g559
  (
    n617,
    n85,
    n135,
    n99,
    n86
  );


  nand
  g560
  (
    n498,
    n222,
    n88,
    n215,
    n80
  );


  and
  g561
  (
    n516,
    n259,
    n264,
    n126,
    n200
  );


  nor
  g562
  (
    n426,
    n152,
    n97,
    n123,
    n117
  );


  nand
  g563
  (
    n439,
    n148,
    n103,
    n187,
    n131
  );


  and
  g564
  (
    n445,
    n156,
    n288,
    n109,
    n87
  );


  or
  g565
  (
    n385,
    n250,
    n122,
    n152,
    n131
  );


  xor
  g566
  (
    n486,
    n255,
    n268,
    n112,
    n285
  );


  xor
  g567
  (
    n478,
    n109,
    n193,
    n116,
    n215
  );


  or
  g568
  (
    n446,
    n124,
    n178,
    n140,
    n271
  );


  xnor
  g569
  (
    n459,
    n155,
    n150,
    n283
  );


  nand
  g570
  (
    n413,
    n119,
    n129,
    n242,
    n256
  );


  xnor
  g571
  (
    n438,
    n152,
    n123,
    n111,
    n133
  );


  xnor
  g572
  (
    n391,
    n267,
    n217,
    n201,
    n276
  );


  nand
  g573
  (
    n351,
    n293,
    n128,
    n91,
    n97
  );


  nand
  g574
  (
    n456,
    n188,
    n100,
    n149,
    n151
  );


  xor
  g575
  (
    n604,
    n292,
    n245,
    n147,
    n263
  );


  xnor
  g576
  (
    n543,
    n159,
    n238,
    n259,
    n204
  );


  nand
  g577
  (
    n387,
    n116,
    n99,
    n96,
    n266
  );


  nor
  g578
  (
    n384,
    n100,
    n134,
    n209,
    n122
  );


  nand
  g579
  (
    n407,
    n139,
    n136,
    n92,
    n105
  );


  and
  g580
  (
    n601,
    n140,
    n206,
    n157,
    n264
  );


  and
  g581
  (
    n605,
    n226,
    n206,
    n156,
    n142
  );


  and
  g582
  (
    n493,
    n227,
    n109,
    n159,
    n154
  );


  and
  g583
  (
    n398,
    n238,
    n94,
    n133,
    n88
  );


  xor
  g584
  (
    n599,
    n203,
    n277,
    n124,
    n273
  );


  nor
  g585
  (
    n551,
    n231,
    n102,
    n220,
    n145
  );


  nand
  g586
  (
    n539,
    n147,
    n280,
    n108
  );


  not
  g587
  (
    n655,
    n361
  );


  buf
  g588
  (
    n654,
    n355
  );


  buf
  g589
  (
    n624,
    n383
  );


  buf
  g590
  (
    n659,
    n362
  );


  buf
  g591
  (
    n652,
    n360
  );


  buf
  g592
  (
    n642,
    n376
  );


  not
  g593
  (
    n648,
    n379
  );


  not
  g594
  (
    n622,
    n375
  );


  buf
  g595
  (
    KeyWire_0_13,
    n365
  );


  buf
  g596
  (
    n638,
    n351
  );


  buf
  g597
  (
    n626,
    n353
  );


  not
  g598
  (
    n651,
    n349
  );


  buf
  g599
  (
    n627,
    n386
  );


  not
  g600
  (
    n643,
    n369
  );


  not
  g601
  (
    n660,
    n374
  );


  not
  g602
  (
    n625,
    n370
  );


  buf
  g603
  (
    n641,
    n371
  );


  buf
  g604
  (
    n623,
    n388
  );


  not
  g605
  (
    n632,
    n350
  );


  not
  g606
  (
    n650,
    n373
  );


  buf
  g607
  (
    n637,
    n359
  );


  buf
  g608
  (
    n636,
    n378
  );


  not
  g609
  (
    n628,
    n368
  );


  buf
  g610
  (
    n646,
    n348
  );


  buf
  g611
  (
    n649,
    n372
  );


  buf
  g612
  (
    n657,
    n347
  );


  not
  g613
  (
    n656,
    n367
  );


  buf
  g614
  (
    n620,
    n354
  );


  not
  g615
  (
    n633,
    n352
  );


  not
  g616
  (
    n639,
    n387
  );


  not
  g617
  (
    n647,
    n358
  );


  not
  g618
  (
    n644,
    n363
  );


  buf
  g619
  (
    n640,
    n377
  );


  buf
  g620
  (
    n629,
    n382
  );


  not
  g621
  (
    n631,
    n357
  );


  not
  g622
  (
    n661,
    n385
  );


  buf
  g623
  (
    n634,
    n366
  );


  buf
  g624
  (
    n645,
    n364
  );


  not
  g625
  (
    n653,
    n356
  );


  buf
  g626
  (
    n621,
    n384
  );


  not
  g627
  (
    n630,
    n380
  );


  not
  g628
  (
    n635,
    n381
  );


  buf
  g629
  (
    n727,
    n620
  );


  not
  g630
  (
    n761,
    n649
  );


  buf
  g631
  (
    n704,
    n487
  );


  not
  g632
  (
    n746,
    n412
  );


  not
  g633
  (
    n747,
    n482
  );


  buf
  g634
  (
    n705,
    n460
  );


  not
  g635
  (
    n680,
    n479
  );


  not
  g636
  (
    n763,
    n654
  );


  not
  g637
  (
    n670,
    n623
  );


  buf
  g638
  (
    n716,
    n631
  );


  not
  g639
  (
    n718,
    n406
  );


  buf
  g640
  (
    n675,
    n629
  );


  not
  g641
  (
    n767,
    n428
  );


  buf
  g642
  (
    n698,
    n659
  );


  not
  g643
  (
    n699,
    n494
  );


  buf
  g644
  (
    n734,
    n391
  );


  buf
  g645
  (
    n684,
    n394
  );


  not
  g646
  (
    n742,
    n500
  );


  buf
  g647
  (
    n754,
    n627
  );


  buf
  g648
  (
    n773,
    n503
  );


  buf
  g649
  (
    n781,
    n431
  );


  buf
  g650
  (
    n772,
    n493
  );


  not
  g651
  (
    n725,
    n621
  );


  not
  g652
  (
    n715,
    n648
  );


  not
  g653
  (
    n723,
    n644
  );


  buf
  g654
  (
    n768,
    n450
  );


  not
  g655
  (
    n749,
    n441
  );


  buf
  g656
  (
    n710,
    n625
  );


  not
  g657
  (
    n757,
    n397
  );


  not
  g658
  (
    n735,
    n474
  );


  buf
  g659
  (
    n674,
    n415
  );


  not
  g660
  (
    n721,
    n644
  );


  not
  g661
  (
    n711,
    n443
  );


  not
  g662
  (
    n738,
    n659
  );


  buf
  g663
  (
    n726,
    n484
  );


  not
  g664
  (
    n744,
    n650
  );


  not
  g665
  (
    n697,
    n422
  );


  buf
  g666
  (
    n766,
    n449
  );


  buf
  g667
  (
    n717,
    n437
  );


  not
  g668
  (
    n682,
    n480
  );


  buf
  g669
  (
    n770,
    n398
  );


  not
  g670
  (
    n759,
    n399
  );


  not
  g671
  (
    n708,
    n409
  );


  buf
  g672
  (
    n732,
    n429
  );


  buf
  g673
  (
    n664,
    n447
  );


  buf
  g674
  (
    n758,
    n489
  );


  buf
  g675
  (
    n774,
    n632
  );


  not
  g676
  (
    n776,
    n462
  );


  buf
  g677
  (
    n692,
    n456
  );


  buf
  g678
  (
    KeyWire_0_4,
    n496
  );


  not
  g679
  (
    n683,
    n639
  );


  buf
  g680
  (
    n756,
    n435
  );


  not
  g681
  (
    n709,
    n625
  );


  not
  g682
  (
    n729,
    n626
  );


  buf
  g683
  (
    n700,
    n490
  );


  buf
  g684
  (
    n688,
    n628
  );


  buf
  g685
  (
    n740,
    n469
  );


  buf
  g686
  (
    n753,
    n621
  );


  not
  g687
  (
    n663,
    n622
  );


  not
  g688
  (
    n779,
    n402
  );


  or
  g689
  (
    n672,
    n476,
    n470,
    n643
  );


  xor
  g690
  (
    n771,
    n632,
    n466,
    n644
  );


  nor
  g691
  (
    n764,
    n463,
    n433,
    n650
  );


  xor
  g692
  (
    n669,
    n446,
    n423,
    n646
  );


  or
  g693
  (
    n695,
    n646,
    n629,
    n438
  );


  or
  g694
  (
    n681,
    n504,
    n392,
    n657
  );


  xor
  g695
  (
    n712,
    n645,
    n624,
    n486
  );


  xnor
  g696
  (
    n687,
    n408,
    n637,
    n471
  );


  and
  g697
  (
    n706,
    n419,
    n414,
    n626
  );


  nor
  g698
  (
    n666,
    n396,
    n622,
    n635
  );


  or
  g699
  (
    n728,
    n620,
    n652,
    n418
  );


  or
  g700
  (
    n714,
    n654,
    n401,
    n393
  );


  nand
  g701
  (
    n755,
    n641,
    n630,
    n404
  );


  nand
  g702
  (
    n769,
    n426,
    n461,
    n637
  );


  nor
  g703
  (
    n679,
    n472,
    n389,
    n459
  );


  xnor
  g704
  (
    n775,
    n651,
    n631,
    n465
  );


  or
  g705
  (
    n686,
    n656,
    n458,
    n395
  );


  or
  g706
  (
    n696,
    n636,
    n626,
    n468
  );


  xor
  g707
  (
    n777,
    n647,
    n634,
    n633
  );


  xnor
  g708
  (
    n713,
    n658,
    n507,
    n457
  );


  and
  g709
  (
    n737,
    n648,
    n656,
    n453
  );


  xor
  g710
  (
    n724,
    n467,
    n652,
    n628
  );


  nor
  g711
  (
    n668,
    n646,
    n623,
    n491
  );


  xor
  g712
  (
    n707,
    n464,
    n439,
    n645
  );


  nand
  g713
  (
    n741,
    n630,
    n651,
    n637
  );


  and
  g714
  (
    n739,
    n432,
    n657,
    n643
  );


  nand
  g715
  (
    n662,
    n647,
    n400,
    n653
  );


  nor
  g716
  (
    n752,
    n481,
    n417,
    n508
  );


  nor
  g717
  (
    n743,
    n655,
    n636,
    n640
  );


  or
  g718
  (
    n733,
    n483,
    n451,
    n440
  );


  and
  g719
  (
    n691,
    n407,
    n639,
    n649
  );


  xnor
  g720
  (
    n690,
    n623,
    n624,
    n657
  );


  xor
  g721
  (
    n720,
    n658,
    n448,
    n444
  );


  and
  g722
  (
    n677,
    n621,
    n454,
    n434
  );


  nand
  g723
  (
    n676,
    n655,
    n497,
    n654
  );


  nor
  g724
  (
    n736,
    n648,
    n642,
    n629
  );


  or
  g725
  (
    n778,
    n625,
    n405,
    n638
  );


  nor
  g726
  (
    n762,
    n410,
    n477,
    n424
  );


  and
  g727
  (
    n731,
    n633,
    n420,
    n442
  );


  and
  g728
  (
    n667,
    n638,
    n620,
    n632
  );


  xor
  g729
  (
    n748,
    n653,
    n641,
    n634
  );


  xnor
  g730
  (
    n678,
    n622,
    n488,
    n635
  );


  nand
  g731
  (
    n685,
    n498,
    n416,
    n390
  );


  xnor
  g732
  (
    n780,
    n492,
    n642,
    n403
  );


  nand
  g733
  (
    n722,
    n653,
    n647,
    n505
  );


  nor
  g734
  (
    n689,
    n645,
    n495,
    n485
  );


  nand
  g735
  (
    n765,
    n652,
    n436,
    n627
  );


  or
  g736
  (
    n760,
    n455,
    n445,
    n649
  );


  nor
  g737
  (
    n719,
    n640,
    n633,
    n473
  );


  nor
  g738
  (
    n701,
    n427,
    n475,
    n478
  );


  nand
  g739
  (
    n702,
    n628,
    n636,
    n655
  );


  xnor
  g740
  (
    n673,
    n630,
    n640,
    n425
  );


  or
  g741
  (
    n751,
    n650,
    n421,
    n639
  );


  and
  g742
  (
    n750,
    n635,
    n501,
    n430
  );


  xor
  g743
  (
    n745,
    n411,
    n499,
    n656
  );


  nor
  g744
  (
    n693,
    n643,
    n634,
    n642
  );


  nor
  g745
  (
    n730,
    n506,
    n624,
    n641
  );


  xor
  g746
  (
    n665,
    n452,
    n627,
    n651
  );


  and
  g747
  (
    n694,
    n631,
    n502,
    n413
  );


  xor
  g748
  (
    n703,
    n658,
    n659,
    n638
  );


  xor
  g749
  (
    n790,
    n330,
    n304,
    n311,
    n329
  );


  xnor
  g750
  (
    n810,
    n312,
    n300,
    n338,
    n662
  );


  or
  g751
  (
    n800,
    n336,
    n297,
    n680,
    n314
  );


  nor
  g752
  (
    n793,
    n303,
    n346,
    n695,
    n333
  );


  xor
  g753
  (
    n795,
    n298,
    n330,
    n343,
    n306
  );


  xnor
  g754
  (
    n802,
    n337,
    n686,
    n314,
    n318
  );


  and
  g755
  (
    n785,
    n696,
    n336,
    n666,
    n327
  );


  xnor
  g756
  (
    n799,
    n302,
    n309,
    n300,
    n310
  );


  xor
  g757
  (
    n809,
    n298,
    n328,
    n675,
    n324
  );


  nand
  g758
  (
    n801,
    n704,
    n320,
    n344,
    n331
  );


  nor
  g759
  (
    n798,
    n682,
    n338,
    n331,
    n707
  );


  nor
  g760
  (
    n797,
    n308,
    n683,
    n681,
    n708
  );


  xor
  g761
  (
    n794,
    n312,
    n303,
    n302,
    n335
  );


  nand
  g762
  (
    n829,
    n697,
    n318,
    n671,
    n304
  );


  xor
  g763
  (
    n821,
    n312,
    n345,
    n700,
    n324
  );


  nor
  g764
  (
    KeyWire_0_9,
    n332,
    n307,
    n667,
    n509
  );


  or
  g765
  (
    n811,
    n325,
    n332,
    n692,
    n330
  );


  xnor
  g766
  (
    n828,
    n301,
    n344,
    n314,
    n322
  );


  xor
  g767
  (
    n816,
    n313,
    n301,
    n337,
    n706
  );


  nand
  g768
  (
    n815,
    n321,
    n690,
    n342,
    n323
  );


  xnor
  g769
  (
    n813,
    n339,
    n332,
    n321,
    n305
  );


  nor
  g770
  (
    n817,
    n670,
    n337,
    n676,
    n694
  );


  xor
  g771
  (
    n792,
    n328,
    n334,
    n319,
    n299
  );


  xor
  g772
  (
    n806,
    n340,
    n344,
    n674,
    n326
  );


  xnor
  g773
  (
    n827,
    n313,
    n687,
    n688,
    n705
  );


  or
  g774
  (
    n805,
    n308,
    n709,
    n341,
    n342
  );


  xor
  g775
  (
    n822,
    n307,
    n320,
    n685,
    n298
  );


  nand
  g776
  (
    n788,
    n322,
    n340,
    n343,
    n335
  );


  or
  g777
  (
    n826,
    n663,
    n678,
    n300,
    n323
  );


  xnor
  g778
  (
    n789,
    n335,
    n345,
    n317,
    n339
  );


  xnor
  g779
  (
    n808,
    n664,
    n311,
    n702,
    n333
  );


  xor
  g780
  (
    n786,
    n334,
    n315,
    n309
  );


  or
  g781
  (
    n823,
    n693,
    n306,
    n329
  );


  xnor
  g782
  (
    n819,
    n310,
    n684,
    n304,
    n673
  );


  nand
  g783
  (
    n820,
    n308,
    n669,
    n323,
    n336
  );


  xnor
  g784
  (
    n830,
    n331,
    n299,
    n339,
    n703
  );


  and
  g785
  (
    n783,
    n672,
    n319,
    n305,
    n689
  );


  or
  g786
  (
    n796,
    n297,
    n317,
    n303,
    n333
  );


  xor
  g787
  (
    n824,
    n668,
    n321,
    n309,
    n318
  );


  xnor
  g788
  (
    n807,
    n325,
    n305,
    n334,
    n701
  );


  or
  g789
  (
    n818,
    n345,
    n691,
    n324,
    n341
  );


  xor
  g790
  (
    n803,
    n327,
    n297,
    n307,
    n302
  );


  or
  g791
  (
    n825,
    n329,
    n342,
    n665,
    n677
  );


  and
  g792
  (
    n784,
    n698,
    n296,
    n340,
    n320
  );


  xnor
  g793
  (
    n831,
    n316,
    n328,
    n299,
    n338
  );


  and
  g794
  (
    n782,
    n311,
    n327,
    n326,
    n317
  );


  xnor
  g795
  (
    n814,
    n301,
    n315,
    n319,
    n343
  );


  or
  g796
  (
    n791,
    n710,
    n326,
    n322,
    n341
  );


  xor
  g797
  (
    n804,
    n313,
    n310,
    n316
  );


  nand
  g798
  (
    n812,
    n711,
    n699,
    n679,
    n325
  );


  buf
  g799
  (
    n842,
    n565
  );


  buf
  g800
  (
    n888,
    n796
  );


  buf
  g801
  (
    n878,
    n795
  );


  buf
  g802
  (
    n889,
    n602
  );


  not
  g803
  (
    n844,
    n782
  );


  buf
  g804
  (
    n859,
    n566
  );


  buf
  g805
  (
    n854,
    n786
  );


  not
  g806
  (
    n874,
    n790
  );


  buf
  g807
  (
    n846,
    n608
  );


  buf
  g808
  (
    n840,
    n797
  );


  buf
  g809
  (
    n834,
    n559
  );


  not
  g810
  (
    n865,
    n586
  );


  buf
  g811
  (
    n864,
    n580
  );


  not
  g812
  (
    n881,
    n596
  );


  buf
  g813
  (
    n845,
    n795
  );


  not
  g814
  (
    n867,
    n712
  );


  buf
  g815
  (
    n858,
    n526
  );


  not
  g816
  (
    n838,
    n792
  );


  buf
  g817
  (
    n860,
    n796
  );


  not
  g818
  (
    n849,
    n521
  );


  not
  g819
  (
    n879,
    n594
  );


  buf
  g820
  (
    n850,
    n532
  );


  not
  g821
  (
    n877,
    n784
  );


  not
  g822
  (
    n856,
    n572
  );


  not
  g823
  (
    n873,
    n550
  );


  and
  g824
  (
    n866,
    n564,
    n569,
    n796
  );


  xnor
  g825
  (
    n851,
    n796,
    n605,
    n552,
    n535
  );


  and
  g826
  (
    n841,
    n563,
    n786,
    n588,
    n790
  );


  xnor
  g827
  (
    n876,
    n787,
    n795,
    n528,
    n589
  );


  xor
  g828
  (
    n884,
    n593,
    n579,
    n542,
    n567
  );


  and
  g829
  (
    n862,
    n603,
    n585,
    n788,
    n793
  );


  and
  g830
  (
    n872,
    n571,
    n544,
    n789,
    n520
  );


  xnor
  g831
  (
    n855,
    n561,
    n714,
    n797,
    n514
  );


  xor
  g832
  (
    n843,
    n530,
    n546,
    n788,
    n573
  );


  or
  g833
  (
    n871,
    n533,
    n537,
    n536,
    n551
  );


  and
  g834
  (
    n869,
    n787,
    n793,
    n590,
    n513
  );


  xnor
  g835
  (
    n880,
    n539,
    n578,
    n785,
    n555
  );


  and
  g836
  (
    n832,
    n789,
    n568,
    n548,
    n538
  );


  and
  g837
  (
    n870,
    n785,
    n782,
    n597,
    n613
  );


  and
  g838
  (
    n863,
    n790,
    n784,
    n609,
    n793
  );


  or
  g839
  (
    n891,
    n788,
    n547,
    n560,
    n529
  );


  xnor
  g840
  (
    n882,
    n599,
    n791,
    n519,
    n581
  );


  xnor
  g841
  (
    n883,
    n793,
    n527,
    n786,
    n787
  );


  nor
  g842
  (
    n885,
    n554,
    n788,
    n545,
    n595
  );


  xnor
  g843
  (
    n837,
    n574,
    n516,
    n524,
    n610
  );


  xor
  g844
  (
    n835,
    n517,
    n510,
    n525,
    n607
  );


  or
  g845
  (
    n875,
    n562,
    n791,
    n518,
    n556
  );


  nand
  g846
  (
    n861,
    n511,
    n540,
    n785,
    n794
  );


  and
  g847
  (
    n853,
    n794,
    n790,
    n543,
    n591
  );


  and
  g848
  (
    n857,
    n587,
    n592,
    n515,
    n582
  );


  nor
  g849
  (
    n890,
    n792,
    n612,
    n782,
    n797
  );


  and
  g850
  (
    n852,
    n601,
    n606,
    n557,
    n783
  );


  xnor
  g851
  (
    n886,
    n534,
    n604,
    n783,
    n576
  );


  or
  g852
  (
    n892,
    n789,
    n792,
    n512,
    n577
  );


  or
  g853
  (
    n868,
    n784,
    n523,
    n522,
    n787
  );


  xor
  g854
  (
    n847,
    n575,
    n795,
    n786,
    n553
  );


  nand
  g855
  (
    n839,
    n794,
    n598,
    n570,
    n558
  );


  xor
  g856
  (
    n848,
    n600,
    n791,
    n531,
    n789
  );


  xor
  g857
  (
    n836,
    n783,
    n611,
    n797,
    n583
  );


  nand
  g858
  (
    n833,
    n584,
    n792,
    n549,
    n791
  );


  nor
  g859
  (
    n887,
    n713,
    n541,
    n794,
    n785
  );


  xor
  g860
  (
    n910,
    n834,
    n835,
    n732,
    n740
  );


  xnor
  g861
  (
    n899,
    n738,
    n717,
    n834,
    n833
  );


  or
  g862
  (
    n902,
    n724,
    n798,
    n718
  );


  or
  g863
  (
    n903,
    n832,
    n738,
    n727,
    n835
  );


  or
  g864
  (
    n894,
    n723,
    n737,
    n739,
    n832
  );


  or
  g865
  (
    n895,
    n736,
    n660,
    n728,
    n835
  );


  and
  g866
  (
    n896,
    n725,
    n735,
    n833,
    n726
  );


  or
  g867
  (
    n893,
    n834,
    n743,
    n798
  );


  or
  g868
  (
    n909,
    n736,
    n660,
    n728
  );


  and
  g869
  (
    n900,
    n740,
    n661,
    n833
  );


  and
  g870
  (
    n908,
    n722,
    n734,
    n661,
    n833
  );


  and
  g871
  (
    n904,
    n743,
    n836,
    n733,
    n742
  );


  nand
  g872
  (
    n898,
    n715,
    n744,
    n732,
    n836
  );


  or
  g873
  (
    n897,
    n737,
    n741,
    n729,
    n739
  );


  nand
  g874
  (
    n901,
    n729,
    n836,
    n730,
    n742
  );


  xnor
  g875
  (
    n912,
    n741,
    n744,
    n731,
    n727
  );


  or
  g876
  (
    n906,
    n836,
    n837,
    n735,
    n730
  );


  nor
  g877
  (
    KeyWire_0_3,
    n835,
    n733,
    n834,
    n720
  );


  nand
  g878
  (
    n907,
    n721,
    n731,
    n660,
    n832
  );


  nand
  g879
  (
    n911,
    n716,
    n734,
    n719,
    n661
  );


  buf
  g880
  (
    n916,
    n747
  );


  not
  g881
  (
    n915,
    n905
  );


  not
  g882
  (
    n919,
    n900
  );


  buf
  g883
  (
    n913,
    n897
  );


  and
  g884
  (
    n914,
    n901,
    n899,
    n748,
    n749
  );


  and
  g885
  (
    n921,
    n751,
    n745,
    n746,
    n747
  );


  and
  g886
  (
    n917,
    n751,
    n745,
    n898,
    n750
  );


  xor
  g887
  (
    n918,
    n749,
    n752,
    n903,
    n750
  );


  or
  g888
  (
    n920,
    n746,
    n904,
    n748,
    n902
  );


  xor
  g889
  (
    n957,
    n814,
    n815,
    n813,
    n810
  );


  nor
  g890
  (
    n955,
    n918,
    n818,
    n914,
    n804
  );


  nand
  g891
  (
    n922,
    n804,
    n913,
    n917,
    n817
  );


  or
  g892
  (
    n951,
    n810,
    n817,
    n913,
    n921
  );


  nor
  g893
  (
    n949,
    n811,
    n815,
    n810,
    n916
  );


  nor
  g894
  (
    n952,
    n814,
    n916,
    n808,
    n801
  );


  nor
  g895
  (
    n931,
    n914,
    n811,
    n802,
    n803
  );


  nand
  g896
  (
    n932,
    n801,
    n824,
    n805,
    n806
  );


  nor
  g897
  (
    n943,
    n824,
    n819,
    n812,
    n822
  );


  or
  g898
  (
    n937,
    n802,
    n807,
    n819,
    n808
  );


  nor
  g899
  (
    n946,
    n800,
    n816,
    n913,
    n814
  );


  nand
  g900
  (
    n942,
    n801,
    n811,
    n816,
    n920
  );


  or
  g901
  (
    n936,
    n814,
    n805,
    n813,
    n810
  );


  nand
  g902
  (
    n940,
    n920,
    n803,
    n915,
    n806
  );


  and
  g903
  (
    n956,
    n818,
    n807,
    n808,
    n800
  );


  and
  g904
  (
    n941,
    n799,
    n812,
    n820,
    n813
  );


  nor
  g905
  (
    n935,
    n809,
    n917,
    n916,
    n821
  );


  and
  g906
  (
    n938,
    n920,
    n915,
    n799,
    n919
  );


  and
  g907
  (
    n925,
    n809,
    n918,
    n823,
    n807
  );


  xor
  g908
  (
    n948,
    n823,
    n802,
    n822
  );


  or
  g909
  (
    n939,
    n805,
    n812,
    n915,
    n809
  );


  nand
  g910
  (
    n929,
    n815,
    n919,
    n820
  );


  nand
  g911
  (
    n944,
    n813,
    n917,
    n799,
    n811
  );


  xor
  g912
  (
    n954,
    n825,
    n818,
    n918,
    n914
  );


  nor
  g913
  (
    n923,
    n917,
    n801,
    n804,
    n803
  );


  and
  g914
  (
    n924,
    n800,
    n918,
    n819,
    n820
  );


  or
  g915
  (
    n930,
    n800,
    n752,
    n817,
    n921
  );


  nor
  g916
  (
    n945,
    n753,
    n821,
    n914
  );


  and
  g917
  (
    n950,
    n805,
    n817,
    n815,
    n823
  );


  or
  g918
  (
    n953,
    n915,
    n816,
    n920,
    n913
  );


  nand
  g919
  (
    n926,
    n816,
    n821,
    n753,
    n812
  );


  nand
  g920
  (
    n927,
    n806,
    n808,
    n818,
    n804
  );


  and
  g921
  (
    n947,
    n803,
    n921,
    n807,
    n809
  );


  xor
  g922
  (
    n928,
    n820,
    n921,
    n806,
    n802
  );


  nand
  g923
  (
    n933,
    n919,
    n823,
    n824,
    n822
  );


  and
  g924
  (
    n934,
    n824,
    n819,
    n916,
    n799
  );


  and
  g925
  (
    n1014,
    n876,
    n843,
    n869,
    n928
  );


  xnor
  g926
  (
    n1003,
    n839,
    n856,
    n875,
    n867
  );


  xnor
  g927
  (
    n981,
    n850,
    n841,
    n937,
    n938
  );


  and
  g928
  (
    n983,
    n848,
    n875,
    n863,
    n844
  );


  xor
  g929
  (
    n1011,
    n853,
    n949,
    n889,
    n944
  );


  xnor
  g930
  (
    n1001,
    n838,
    n888,
    n883,
    n940
  );


  or
  g931
  (
    n1017,
    n863,
    n948,
    n945,
    n886
  );


  or
  g932
  (
    n1026,
    n842,
    n941,
    n888,
    n868
  );


  or
  g933
  (
    n993,
    n936,
    n855,
    n878
  );


  xnor
  g934
  (
    n986,
    n861,
    n932,
    n930,
    n945
  );


  xnor
  g935
  (
    n1009,
    n866,
    n841,
    n862,
    n846
  );


  and
  g936
  (
    n994,
    n859,
    n885,
    n875,
    n851
  );


  xnor
  g937
  (
    n1004,
    n870,
    n869,
    n857,
    n860
  );


  nand
  g938
  (
    n1024,
    n878,
    n841,
    n890,
    n845
  );


  xnor
  g939
  (
    n965,
    n862,
    n931,
    n847,
    n876
  );


  and
  g940
  (
    n1025,
    n879,
    n855,
    n876,
    n926
  );


  or
  g941
  (
    n1028,
    n843,
    n943,
    n935,
    n874
  );


  xor
  g942
  (
    n977,
    n852,
    n838,
    n879,
    n864
  );


  xor
  g943
  (
    n1005,
    n853,
    n856,
    n930,
    n852
  );


  nor
  g944
  (
    n968,
    n924,
    n838,
    n883,
    n881
  );


  nand
  g945
  (
    n1000,
    n859,
    n861,
    n937,
    n865
  );


  nand
  g946
  (
    n1021,
    n874,
    n840,
    n842,
    n947
  );


  nor
  g947
  (
    n961,
    n849,
    n928,
    n861,
    n883
  );


  nor
  g948
  (
    n974,
    n890,
    n875,
    n862,
    n837
  );


  xor
  g949
  (
    n1030,
    n924,
    n889,
    n943,
    n860
  );


  nor
  g950
  (
    n1012,
    n856,
    n881,
    n939,
    n864
  );


  nand
  g951
  (
    n997,
    n932,
    n938,
    n891,
    n863
  );


  xor
  g952
  (
    n978,
    n855,
    n845,
    n851,
    n868
  );


  and
  g953
  (
    n976,
    n935,
    n840,
    n939,
    n877
  );


  nor
  g954
  (
    n991,
    n871,
    n888,
    n950,
    n857
  );


  xnor
  g955
  (
    n1020,
    n882,
    n847,
    n858,
    n870
  );


  xnor
  g956
  (
    n1018,
    n884,
    n859,
    n891,
    n882
  );


  xnor
  g957
  (
    n989,
    n949,
    n844,
    n866,
    n838
  );


  nand
  g958
  (
    n980,
    n890,
    n945,
    n948,
    n942
  );


  and
  g959
  (
    n988,
    n869,
    n922,
    n848,
    n843
  );


  and
  g960
  (
    n975,
    n873,
    n840,
    n870,
    n889
  );


  nor
  g961
  (
    n1002,
    n880,
    n881,
    n940,
    n841
  );


  nand
  g962
  (
    n1019,
    n871,
    n858,
    n865,
    n849
  );


  xnor
  g963
  (
    n996,
    n844,
    n852,
    n944,
    n949
  );


  and
  g964
  (
    n1007,
    n942,
    n874,
    n950,
    n868
  );


  xor
  g965
  (
    n966,
    n837,
    n864,
    n839,
    n871
  );


  or
  g966
  (
    n979,
    n943,
    n863,
    n941,
    n946
  );


  or
  g967
  (
    n1015,
    n873,
    n845,
    n851,
    n860
  );


  nor
  g968
  (
    n1022,
    n947,
    n868,
    n933,
    n941
  );


  xnor
  g969
  (
    n969,
    n869,
    n940,
    n938,
    n854
  );


  or
  g970
  (
    n973,
    n936,
    n880,
    n864,
    n850
  );


  xor
  g971
  (
    n1029,
    n887,
    n926,
    n853,
    n867
  );


  nor
  g972
  (
    n971,
    n891,
    n888,
    n925,
    n877
  );


  xor
  g973
  (
    n1023,
    n882,
    n848,
    n887,
    n854
  );


  and
  g974
  (
    n1006,
    n839,
    n946,
    n850,
    n934
  );


  and
  g975
  (
    n1008,
    n847,
    n872,
    n923,
    n874
  );


  and
  g976
  (
    n982,
    n950,
    n933,
    n891,
    n844
  );


  xnor
  g977
  (
    n963,
    n854,
    n878,
    n853,
    n846
  );


  nor
  g978
  (
    n972,
    n872,
    n854,
    n849,
    n846
  );


  xor
  g979
  (
    n958,
    n877,
    n879,
    n866,
    n843
  );


  nor
  g980
  (
    n1027,
    n884,
    n885,
    n927,
    n939
  );


  nor
  g981
  (
    n959,
    n871,
    n858,
    n840,
    n872
  );


  xnor
  g982
  (
    n970,
    n946,
    n847,
    n887,
    n883
  );


  or
  g983
  (
    n990,
    n886,
    n884,
    n934,
    n859
  );


  xnor
  g984
  (
    n998,
    n865,
    n885,
    n837,
    n882
  );


  nand
  g985
  (
    n1013,
    n923,
    n873,
    n852,
    n944
  );


  xnor
  g986
  (
    n1016,
    n866,
    n925,
    n842,
    n942
  );


  or
  g987
  (
    n992,
    n880,
    n947,
    n929,
    n879
  );


  xnor
  g988
  (
    n987,
    n862,
    n922,
    n881,
    n858
  );


  and
  g989
  (
    n999,
    n860,
    n884,
    n846,
    n867
  );


  xor
  g990
  (
    n984,
    n929,
    n927,
    n880,
    n887
  );


  xor
  g991
  (
    n967,
    n845,
    n885,
    n861,
    n850
  );


  xor
  g992
  (
    n964,
    n876,
    n878,
    n877,
    n870
  );


  nor
  g993
  (
    n960,
    n857,
    n839,
    n886
  );


  xor
  g994
  (
    n985,
    n856,
    n848,
    n889,
    n842
  );


  and
  g995
  (
    n1010,
    n948,
    n873,
    n872,
    n931
  );


  or
  g996
  (
    n995,
    n849,
    n851,
    n936,
    n867
  );


  xnor
  g997
  (
    n962,
    n890,
    n857,
    n937,
    n865
  );


  not
  g998
  (
    n1077,
    n974
  );


  buf
  g999
  (
    n1065,
    n759
  );


  not
  g1000
  (
    n1034,
    n984
  );


  buf
  g1001
  (
    n1060,
    n911
  );


  buf
  g1002
  (
    n1080,
    n757
  );


  buf
  g1003
  (
    n1085,
    n827
  );


  not
  g1004
  (
    n1037,
    n828
  );


  buf
  g1005
  (
    n1051,
    n1011
  );


  not
  g1006
  (
    n1071,
    n754
  );


  not
  g1007
  (
    n1032,
    n908
  );


  buf
  g1008
  (
    n1056,
    n1016
  );


  not
  g1009
  (
    n1086,
    n975
  );


  buf
  g1010
  (
    n1061,
    n971
  );


  not
  g1011
  (
    n1041,
    n754
  );


  not
  g1012
  (
    n1053,
    n1020
  );


  not
  g1013
  (
    n1031,
    n967
  );


  not
  g1014
  (
    n1042,
    n826
  );


  not
  g1015
  (
    n1048,
    n825
  );


  buf
  g1016
  (
    n1045,
    n829
  );


  not
  g1017
  (
    n1093,
    n907
  );


  buf
  g1018
  (
    n1057,
    n1010
  );


  buf
  g1019
  (
    n1070,
    n758
  );


  not
  g1020
  (
    n1054,
    n1001
  );


  not
  g1021
  (
    n1064,
    n755
  );


  buf
  g1022
  (
    n1069,
    n1026
  );


  buf
  g1023
  (
    n1036,
    n761
  );


  not
  g1024
  (
    n1047,
    n828
  );


  not
  g1025
  (
    n1076,
    n764
  );


  not
  g1026
  (
    n1067,
    n764
  );


  buf
  g1027
  (
    n1079,
    n827
  );


  not
  g1028
  (
    n1058,
    n997
  );


  buf
  g1029
  (
    n1068,
    n1014
  );


  buf
  g1030
  (
    n1039,
    n983
  );


  not
  g1031
  (
    n1043,
    n757
  );


  buf
  g1032
  (
    n1081,
    n988
  );


  buf
  g1033
  (
    n1038,
    n826
  );


  buf
  g1034
  (
    n1084,
    n1012
  );


  buf
  g1035
  (
    n1050,
    n1007
  );


  buf
  g1036
  (
    n1062,
    n980
  );


  buf
  g1037
  (
    n1040,
    n1019
  );


  not
  g1038
  (
    n1083,
    n995
  );


  not
  g1039
  (
    n1066,
    n979
  );


  buf
  g1040
  (
    n1052,
    n770
  );


  buf
  g1041
  (
    n1033,
    n825
  );


  xor
  g1042
  (
    n1078,
    n999,
    n973,
    n1009,
    n978
  );


  and
  g1043
  (
    n1082,
    n756,
    n986,
    n758,
    n1022
  );


  nor
  g1044
  (
    n1046,
    n1015,
    n976,
    n910,
    n1027
  );


  xor
  g1045
  (
    n1049,
    n765,
    n756,
    n1017,
    n991
  );


  or
  g1046
  (
    n1075,
    n968,
    n1003,
    n759,
    n760
  );


  nand
  g1047
  (
    n1094,
    n990,
    n989,
    n1000,
    n987
  );


  xor
  g1048
  (
    n1055,
    n765,
    n763,
    n1004
  );


  nand
  g1049
  (
    n1072,
    n972,
    n827,
    n767,
    n906
  );


  or
  g1050
  (
    n1035,
    n1029,
    n985,
    n969,
    n826
  );


  or
  g1051
  (
    n1091,
    n767,
    n1030,
    n829,
    n768
  );


  and
  g1052
  (
    n1044,
    n1021,
    n826,
    n829,
    n977
  );


  nand
  g1053
  (
    n1074,
    n1024,
    n1028,
    n1002,
    n909
  );


  xnor
  g1054
  (
    n1063,
    n1006,
    n770,
    n828,
    n825
  );


  nand
  g1055
  (
    n1059,
    n998,
    n762,
    n1023,
    n994
  );


  xor
  g1056
  (
    n1092,
    n1018,
    n830,
    n1005,
    n827
  );


  nand
  g1057
  (
    n1089,
    n993,
    n996,
    n755,
    n981
  );


  and
  g1058
  (
    n1087,
    n766,
    n769,
    n762
  );


  and
  g1059
  (
    n1090,
    n761,
    n1025,
    n766,
    n828
  );


  or
  g1060
  (
    n1073,
    n1008,
    n768,
    n760,
    n982
  );


  nor
  g1061
  (
    n1088,
    n829,
    n992,
    n1013,
    n970
  );


  not
  g1062
  (
    n1159,
    n1052
  );


  not
  g1063
  (
    n1133,
    n1082
  );


  buf
  g1064
  (
    n1191,
    n1090
  );


  not
  g1065
  (
    n1342,
    n1046
  );


  not
  g1066
  (
    n1151,
    n1039
  );


  buf
  g1067
  (
    n1155,
    n1040
  );


  not
  g1068
  (
    n1265,
    n1056
  );


  buf
  g1069
  (
    n1317,
    n1075
  );


  buf
  g1070
  (
    n1282,
    n1032
  );


  buf
  g1071
  (
    n1242,
    n1093
  );


  buf
  g1072
  (
    n1225,
    n1042
  );


  not
  g1073
  (
    n1222,
    n1054
  );


  buf
  g1074
  (
    n1332,
    n1035
  );


  buf
  g1075
  (
    n1219,
    n1061
  );


  buf
  g1076
  (
    n1289,
    n1044
  );


  buf
  g1077
  (
    n1240,
    n1070
  );


  not
  g1078
  (
    n1212,
    n1055
  );


  buf
  g1079
  (
    n1156,
    n1034
  );


  buf
  g1080
  (
    n1308,
    n1043
  );


  not
  g1081
  (
    n1194,
    n1078
  );


  not
  g1082
  (
    n1261,
    n1092
  );


  buf
  g1083
  (
    n1182,
    n1065
  );


  buf
  g1084
  (
    n1276,
    n1038
  );


  not
  g1085
  (
    n1290,
    n1032
  );


  buf
  g1086
  (
    n1127,
    n1038
  );


  not
  g1087
  (
    n1295,
    n1089
  );


  not
  g1088
  (
    n1142,
    n1061
  );


  not
  g1089
  (
    n1246,
    n1091
  );


  not
  g1090
  (
    n1239,
    n1087
  );


  not
  g1091
  (
    n1196,
    n1043
  );


  buf
  g1092
  (
    n1237,
    n1037
  );


  not
  g1093
  (
    n1220,
    n1079
  );


  not
  g1094
  (
    n1108,
    n1058
  );


  not
  g1095
  (
    n1329,
    n1063
  );


  buf
  g1096
  (
    n1326,
    n1031
  );


  buf
  g1097
  (
    n1097,
    n1033
  );


  buf
  g1098
  (
    n1341,
    n1043
  );


  not
  g1099
  (
    n1331,
    n1069
  );


  not
  g1100
  (
    n1128,
    n1076
  );


  buf
  g1101
  (
    n1300,
    n1073
  );


  not
  g1102
  (
    n1333,
    n1059
  );


  not
  g1103
  (
    n1328,
    n1058
  );


  buf
  g1104
  (
    n1105,
    n1094
  );


  not
  g1105
  (
    n1173,
    n1064
  );


  not
  g1106
  (
    n1218,
    n1040
  );


  not
  g1107
  (
    n1186,
    n1081
  );


  not
  g1108
  (
    n1302,
    n1077
  );


  buf
  g1109
  (
    n1248,
    n1055
  );


  not
  g1110
  (
    n1176,
    n1071
  );


  not
  g1111
  (
    n1233,
    n1071
  );


  not
  g1112
  (
    n1313,
    n1084
  );


  buf
  g1113
  (
    n1161,
    n1093
  );


  buf
  g1114
  (
    n1198,
    n1059
  );


  not
  g1115
  (
    n1221,
    n1072
  );


  buf
  g1116
  (
    n1320,
    n1056
  );


  not
  g1117
  (
    n1287,
    n1068
  );


  not
  g1118
  (
    n1310,
    n1050
  );


  not
  g1119
  (
    n1203,
    n1045
  );


  not
  g1120
  (
    n1213,
    n1082
  );


  buf
  g1121
  (
    n1335,
    n1078
  );


  buf
  g1122
  (
    n1103,
    n1052
  );


  not
  g1123
  (
    n1149,
    n1042
  );


  buf
  g1124
  (
    n1279,
    n1083
  );


  buf
  g1125
  (
    n1228,
    n1059
  );


  not
  g1126
  (
    n1192,
    n1082
  );


  buf
  g1127
  (
    n1293,
    n1052
  );


  not
  g1128
  (
    n1263,
    n1085
  );


  not
  g1129
  (
    n1267,
    n1033
  );


  buf
  g1130
  (
    n1119,
    n1085
  );


  buf
  g1131
  (
    n1280,
    n1055
  );


  not
  g1132
  (
    n1325,
    n1031
  );


  buf
  g1133
  (
    n1136,
    n1035
  );


  not
  g1134
  (
    n1181,
    n1049
  );


  buf
  g1135
  (
    n1347,
    n1080
  );


  buf
  g1136
  (
    n1299,
    n1085
  );


  buf
  g1137
  (
    n1231,
    n1063
  );


  not
  g1138
  (
    n1109,
    n1033
  );


  not
  g1139
  (
    n1318,
    n1083
  );


  buf
  g1140
  (
    n1346,
    n1092
  );


  buf
  g1141
  (
    n1315,
    n1037
  );


  buf
  g1142
  (
    n1134,
    n1046
  );


  not
  g1143
  (
    n1122,
    n1060
  );


  buf
  g1144
  (
    n1324,
    n1066
  );


  buf
  g1145
  (
    n1146,
    n1053
  );


  not
  g1146
  (
    n1141,
    n1041
  );


  not
  g1147
  (
    n1338,
    n1048
  );


  not
  g1148
  (
    n1202,
    n1057
  );


  buf
  g1149
  (
    n1226,
    n1048
  );


  not
  g1150
  (
    n1157,
    n1047
  );


  buf
  g1151
  (
    n1185,
    n1068
  );


  buf
  g1152
  (
    n1135,
    n1075
  );


  not
  g1153
  (
    n1168,
    n1094
  );


  not
  g1154
  (
    n1232,
    n1077
  );


  not
  g1155
  (
    n1345,
    n1033
  );


  not
  g1156
  (
    n1166,
    n1054
  );


  not
  g1157
  (
    n1316,
    n1069
  );


  not
  g1158
  (
    n1207,
    n1072
  );


  not
  g1159
  (
    n1111,
    n1051
  );


  buf
  g1160
  (
    n1211,
    n1092
  );


  not
  g1161
  (
    n1188,
    n1064
  );


  buf
  g1162
  (
    n1130,
    n1066
  );


  not
  g1163
  (
    n1340,
    n1057
  );


  not
  g1164
  (
    n1336,
    n1062
  );


  not
  g1165
  (
    n1292,
    n1083
  );


  buf
  g1166
  (
    n1165,
    n1080
  );


  not
  g1167
  (
    n1264,
    n1088
  );


  buf
  g1168
  (
    n1337,
    n1046
  );


  buf
  g1169
  (
    n1210,
    n1046
  );


  not
  g1170
  (
    n1247,
    n1091
  );


  buf
  g1171
  (
    n1120,
    n1053
  );


  not
  g1172
  (
    n1230,
    n1060
  );


  buf
  g1173
  (
    n1095,
    n1076
  );


  buf
  g1174
  (
    n1216,
    n1045
  );


  not
  g1175
  (
    n1286,
    n1038
  );


  not
  g1176
  (
    n1164,
    n1066
  );


  not
  g1177
  (
    n1116,
    n1047
  );


  not
  g1178
  (
    n1102,
    n1073
  );


  not
  g1179
  (
    n1277,
    n1043
  );


  not
  g1180
  (
    n1307,
    n1076
  );


  buf
  g1181
  (
    n1137,
    n772
  );


  not
  g1182
  (
    n1256,
    n1060
  );


  not
  g1183
  (
    n1229,
    n1066
  );


  not
  g1184
  (
    n1174,
    n1089
  );


  not
  g1185
  (
    n1281,
    n1077
  );


  not
  g1186
  (
    n1139,
    n1051
  );


  buf
  g1187
  (
    n1348,
    n1078
  );


  not
  g1188
  (
    n1140,
    n1058
  );


  not
  g1189
  (
    n1170,
    n771
  );


  not
  g1190
  (
    n1169,
    n1044
  );


  buf
  g1191
  (
    n1209,
    n773
  );


  buf
  g1192
  (
    n1180,
    n1090
  );


  not
  g1193
  (
    n1143,
    n1062
  );


  buf
  g1194
  (
    n1273,
    n1087
  );


  not
  g1195
  (
    n1104,
    n1034
  );


  not
  g1196
  (
    n1150,
    n1090
  );


  not
  g1197
  (
    n1124,
    n1047
  );


  buf
  g1198
  (
    n1309,
    n1091
  );


  buf
  g1199
  (
    n1254,
    n1031
  );


  not
  g1200
  (
    n1262,
    n1038
  );


  not
  g1201
  (
    n1189,
    n773
  );


  not
  g1202
  (
    n1350,
    n1070
  );


  not
  g1203
  (
    n1339,
    n1067
  );


  not
  g1204
  (
    n1271,
    n1058
  );


  not
  g1205
  (
    n1251,
    n1049
  );


  not
  g1206
  (
    n1301,
    n1075
  );


  buf
  g1207
  (
    n1270,
    n1037
  );


  buf
  g1208
  (
    n1100,
    n1051
  );


  not
  g1209
  (
    n1125,
    n1067
  );


  buf
  g1210
  (
    n1201,
    n1032
  );


  not
  g1211
  (
    n1115,
    n1071
  );


  not
  g1212
  (
    n1129,
    n1065
  );


  buf
  g1213
  (
    n1330,
    n1072
  );


  not
  g1214
  (
    n1311,
    n1088
  );


  not
  g1215
  (
    n1208,
    n1067
  );


  not
  g1216
  (
    n1183,
    n1086
  );


  buf
  g1217
  (
    n1154,
    n1085
  );


  buf
  g1218
  (
    n1096,
    n1065
  );


  not
  g1219
  (
    n1344,
    n1049
  );


  not
  g1220
  (
    n1145,
    n1048
  );


  not
  g1221
  (
    n1117,
    n1082
  );


  buf
  g1222
  (
    n1190,
    n1078
  );


  not
  g1223
  (
    n1195,
    n1089
  );


  not
  g1224
  (
    n1243,
    n1031
  );


  not
  g1225
  (
    n1227,
    n1088
  );


  not
  g1226
  (
    n1314,
    n1064
  );


  buf
  g1227
  (
    n1234,
    n1086
  );


  buf
  g1228
  (
    n1241,
    n1090
  );


  buf
  g1229
  (
    n1312,
    n1041
  );


  buf
  g1230
  (
    n1187,
    n1039
  );


  buf
  g1231
  (
    n1238,
    n1091
  );


  not
  g1232
  (
    n1178,
    n1079
  );


  not
  g1233
  (
    n1193,
    n1055
  );


  not
  g1234
  (
    n1250,
    n1084
  );


  not
  g1235
  (
    n1235,
    n1056
  );


  buf
  g1236
  (
    n1138,
    n1086
  );


  buf
  g1237
  (
    n1275,
    n1070
  );


  buf
  g1238
  (
    n1285,
    n1048
  );


  not
  g1239
  (
    n1304,
    n1047
  );


  buf
  g1240
  (
    n1306,
    n1087
  );


  buf
  g1241
  (
    n1321,
    n1049
  );


  not
  g1242
  (
    n1132,
    n1077
  );


  not
  g1243
  (
    n1205,
    n1062
  );


  buf
  g1244
  (
    n1147,
    n1079
  );


  buf
  g1245
  (
    n1148,
    n1041
  );


  not
  g1246
  (
    n1126,
    n1036
  );


  not
  g1247
  (
    n1249,
    n1069
  );


  buf
  g1248
  (
    n1131,
    n1044
  );


  not
  g1249
  (
    n1305,
    n1041
  );


  not
  g1250
  (
    n1172,
    n1074
  );


  not
  g1251
  (
    n1274,
    n1054
  );


  buf
  g1252
  (
    n1123,
    n1042
  );


  not
  g1253
  (
    n1294,
    n1074
  );


  not
  g1254
  (
    n1245,
    n1074
  );


  buf
  g1255
  (
    n1199,
    n772
  );


  not
  g1256
  (
    n1278,
    n1045
  );


  buf
  g1257
  (
    n1303,
    n1040
  );


  buf
  g1258
  (
    n1197,
    n1072
  );


  not
  g1259
  (
    n1260,
    n1081
  );


  buf
  g1260
  (
    n1291,
    n1042
  );


  buf
  g1261
  (
    n1283,
    n1084
  );


  not
  g1262
  (
    n1171,
    n1057
  );


  buf
  g1263
  (
    n1252,
    n1032
  );


  buf
  g1264
  (
    n1175,
    n1035
  );


  not
  g1265
  (
    n1215,
    n1065
  );


  buf
  g1266
  (
    n1284,
    n1064
  );


  buf
  g1267
  (
    n1322,
    n1073
  );


  buf
  g1268
  (
    n1223,
    n1057
  );


  not
  g1269
  (
    n1114,
    n1040
  );


  buf
  g1270
  (
    n1259,
    n1081
  );


  buf
  g1271
  (
    n1244,
    n1053
  );


  buf
  g1272
  (
    n1163,
    n1089
  );


  buf
  g1273
  (
    n1152,
    n1039
  );


  buf
  g1274
  (
    n1269,
    n1054
  );


  not
  g1275
  (
    n1113,
    n1059
  );


  not
  g1276
  (
    n1121,
    n1079
  );


  not
  g1277
  (
    n1144,
    n1074
  );


  buf
  g1278
  (
    n1217,
    n1087
  );


  not
  g1279
  (
    KeyWire_0_14,
    n1050
  );


  not
  g1280
  (
    n1343,
    n1063
  );


  not
  g1281
  (
    n1204,
    n1053
  );


  not
  g1282
  (
    n1258,
    n1037
  );


  buf
  g1283
  (
    n1349,
    n1067
  );


  not
  g1284
  (
    n1298,
    n1070
  );


  not
  g1285
  (
    n1160,
    n1051
  );


  not
  g1286
  (
    n1272,
    n1062
  );


  not
  g1287
  (
    n1098,
    n1092
  );


  not
  g1288
  (
    n1253,
    n1084
  );


  buf
  g1289
  (
    n1323,
    n1036
  );


  buf
  g1290
  (
    n1200,
    n1044
  );


  buf
  g1291
  (
    n1099,
    n1039
  );


  buf
  g1292
  (
    n1106,
    n1083
  );


  buf
  g1293
  (
    n1334,
    n1061
  );


  not
  g1294
  (
    n1112,
    n1050
  );


  not
  g1295
  (
    n1297,
    n1036
  );


  not
  g1296
  (
    n1319,
    n1045
  );


  buf
  g1297
  (
    n1206,
    n1088
  );


  not
  g1298
  (
    n1266,
    n1094
  );


  not
  g1299
  (
    n1101,
    n1034
  );


  not
  g1300
  (
    n1296,
    n1036
  );


  buf
  g1301
  (
    n1327,
    n1069
  );


  buf
  g1302
  (
    n1167,
    n1063
  );


  not
  g1303
  (
    n1257,
    n1093
  );


  buf
  g1304
  (
    n1236,
    n1073
  );


  buf
  g1305
  (
    n1177,
    n1035
  );


  not
  g1306
  (
    n1214,
    n1052
  );


  buf
  g1307
  (
    n1118,
    n1061
  );


  buf
  g1308
  (
    n1179,
    n1093
  );


  not
  g1309
  (
    n1162,
    n1086
  );


  not
  g1310
  (
    n1107,
    n1068
  );


  not
  g1311
  (
    n1268,
    n1080
  );


  buf
  g1312
  (
    n1255,
    n771
  );


  buf
  g1313
  (
    n1288,
    n1050
  );


  not
  g1314
  (
    n1110,
    n1080
  );


  not
  g1315
  (
    n1158,
    n1075
  );


  or
  g1316
  (
    n1224,
    n1068,
    n1094,
    n1060,
    n1034
  );


  and
  g1317
  (
    n1184,
    n1076,
    n1056,
    n1071,
    n1081
  );


  not
  g1318
  (
    n1364,
    n1141
  );


  not
  g1319
  (
    n1396,
    n1161
  );


  buf
  g1320
  (
    n1354,
    n1136
  );


  not
  g1321
  (
    n1612,
    n1124
  );


  buf
  g1322
  (
    n1504,
    n1130
  );


  buf
  g1323
  (
    n1374,
    n1120
  );


  buf
  g1324
  (
    n1419,
    n1113
  );


  not
  g1325
  (
    n1573,
    n1150
  );


  not
  g1326
  (
    n1484,
    n1115
  );


  buf
  g1327
  (
    n1506,
    n1170
  );


  buf
  g1328
  (
    n1556,
    n1102
  );


  buf
  g1329
  (
    n1530,
    n1147
  );


  buf
  g1330
  (
    n1498,
    n1146
  );


  not
  g1331
  (
    n1388,
    n1098
  );


  not
  g1332
  (
    KeyWire_0_11,
    n780
  );


  buf
  g1333
  (
    n1464,
    n1118
  );


  not
  g1334
  (
    n1439,
    n1102
  );


  not
  g1335
  (
    n1480,
    n346
  );


  not
  g1336
  (
    n1550,
    n1102
  );


  buf
  g1337
  (
    n1647,
    n1114
  );


  buf
  g1338
  (
    n1355,
    n1160
  );


  buf
  g1339
  (
    n1602,
    n1131
  );


  not
  g1340
  (
    n1361,
    n1108
  );


  not
  g1341
  (
    n1427,
    n1161
  );


  buf
  g1342
  (
    n1594,
    n1170
  );


  buf
  g1343
  (
    n1524,
    n1144
  );


  buf
  g1344
  (
    n1485,
    n1112
  );


  not
  g1345
  (
    n1539,
    n1158
  );


  buf
  g1346
  (
    n1406,
    n1111
  );


  not
  g1347
  (
    n1589,
    n1095
  );


  buf
  g1348
  (
    n1366,
    n617
  );


  buf
  g1349
  (
    KeyWire_0_15,
    n1166
  );


  not
  g1350
  (
    n1353,
    n1165
  );


  buf
  g1351
  (
    n1554,
    n778
  );


  buf
  g1352
  (
    n1389,
    n1139
  );


  not
  g1353
  (
    n1508,
    n1109
  );


  buf
  g1354
  (
    n1569,
    n1095
  );


  not
  g1355
  (
    n1648,
    n1148
  );


  buf
  g1356
  (
    n1462,
    n1125
  );


  not
  g1357
  (
    n1395,
    n1114
  );


  not
  g1358
  (
    n1566,
    n1145
  );


  not
  g1359
  (
    n1571,
    n778
  );


  not
  g1360
  (
    KeyWire_0_8,
    n1111
  );


  buf
  g1361
  (
    n1629,
    n1169
  );


  buf
  g1362
  (
    n1563,
    n953
  );


  not
  g1363
  (
    n1449,
    n1162
  );


  buf
  g1364
  (
    n1471,
    n781
  );


  buf
  g1365
  (
    n1616,
    n1141
  );


  not
  g1366
  (
    n1555,
    n1128
  );


  buf
  g1367
  (
    n1436,
    n1107
  );


  buf
  g1368
  (
    n1620,
    n1166
  );


  not
  g1369
  (
    n1630,
    n775
  );


  buf
  g1370
  (
    n1520,
    n1132
  );


  not
  g1371
  (
    n1523,
    n1099
  );


  not
  g1372
  (
    n1625,
    n956
  );


  not
  g1373
  (
    n1450,
    n1162
  );


  buf
  g1374
  (
    n1398,
    n1135
  );


  not
  g1375
  (
    KeyWire_0_7,
    n160
  );


  not
  g1376
  (
    n1577,
    n1103
  );


  not
  g1377
  (
    n1372,
    n1152
  );


  not
  g1378
  (
    n1392,
    n1139
  );


  buf
  g1379
  (
    n1433,
    n1149
  );


  not
  g1380
  (
    n1386,
    n1128
  );


  not
  g1381
  (
    n1548,
    n892
  );


  not
  g1382
  (
    n1601,
    n1147
  );


  not
  g1383
  (
    KeyWire_0_12,
    n1098
  );


  buf
  g1384
  (
    n1631,
    n1115
  );


  not
  g1385
  (
    n1410,
    n1121
  );


  buf
  g1386
  (
    n1380,
    n952
  );


  not
  g1387
  (
    n1624,
    n1103
  );


  not
  g1388
  (
    n1603,
    n1156
  );


  not
  g1389
  (
    n1460,
    n1097
  );


  not
  g1390
  (
    n1444,
    n1157
  );


  not
  g1391
  (
    n1515,
    n1142
  );


  not
  g1392
  (
    n1635,
    n1127
  );


  buf
  g1393
  (
    n1422,
    n1142
  );


  buf
  g1394
  (
    n1512,
    n1153
  );


  buf
  g1395
  (
    n1509,
    n346
  );


  buf
  g1396
  (
    n1617,
    n1111
  );


  not
  g1397
  (
    n1399,
    n1167
  );


  not
  g1398
  (
    n1584,
    n1105
  );


  buf
  g1399
  (
    n1579,
    n830
  );


  not
  g1400
  (
    n1356,
    n1134
  );


  not
  g1401
  (
    n1409,
    n1144
  );


  buf
  g1402
  (
    n1588,
    n1101
  );


  not
  g1403
  (
    n1543,
    n1116
  );


  not
  g1404
  (
    n1496,
    n1129
  );


  buf
  g1405
  (
    n1455,
    n1119
  );


  buf
  g1406
  (
    n1442,
    n1106
  );


  not
  g1407
  (
    n1487,
    n779
  );


  not
  g1408
  (
    n1475,
    n1146
  );


  buf
  g1409
  (
    n1611,
    n1126
  );


  not
  g1410
  (
    n1465,
    n1100
  );


  buf
  g1411
  (
    n1572,
    n1096
  );


  not
  g1412
  (
    n1453,
    n1130
  );


  buf
  g1413
  (
    n1382,
    n1152
  );


  buf
  g1414
  (
    n1413,
    n1134
  );


  not
  g1415
  (
    n1549,
    n957
  );


  buf
  g1416
  (
    n1521,
    n1145
  );


  buf
  g1417
  (
    n1459,
    n1124
  );


  buf
  g1418
  (
    n1478,
    n1114
  );


  buf
  g1419
  (
    n1593,
    n1133
  );


  buf
  g1420
  (
    n1514,
    n1110
  );


  not
  g1421
  (
    n1637,
    n774
  );


  not
  g1422
  (
    n1638,
    n1155
  );


  buf
  g1423
  (
    n1477,
    n1122
  );


  buf
  g1424
  (
    n1619,
    n1171
  );


  not
  g1425
  (
    n1608,
    n1099
  );


  buf
  g1426
  (
    n1476,
    n1138
  );


  not
  g1427
  (
    n1610,
    n1169
  );


  not
  g1428
  (
    n1446,
    n1153
  );


  not
  g1429
  (
    n1456,
    n1096
  );


  buf
  g1430
  (
    n1488,
    n780
  );


  buf
  g1431
  (
    n1605,
    n1118
  );


  buf
  g1432
  (
    n1431,
    n1122
  );


  buf
  g1433
  (
    n1373,
    n954
  );


  not
  g1434
  (
    n1614,
    n1159
  );


  not
  g1435
  (
    n1551,
    n1112
  );


  buf
  g1436
  (
    n1536,
    n1109
  );


  buf
  g1437
  (
    n1621,
    n953
  );


  not
  g1438
  (
    n1385,
    n1109
  );


  not
  g1439
  (
    n1502,
    n1158
  );


  not
  g1440
  (
    n1447,
    n1136
  );


  not
  g1441
  (
    n1408,
    n1119
  );


  not
  g1442
  (
    n1639,
    n1154
  );


  not
  g1443
  (
    n1371,
    n1095
  );


  buf
  g1444
  (
    n1495,
    n1152
  );


  not
  g1445
  (
    n1578,
    n1134
  );


  buf
  g1446
  (
    n1636,
    n1166
  );


  buf
  g1447
  (
    n1559,
    n1123
  );


  not
  g1448
  (
    n1404,
    n1137
  );


  not
  g1449
  (
    n1434,
    n831
  );


  buf
  g1450
  (
    n1576,
    n1143
  );


  not
  g1451
  (
    n1424,
    n1134
  );


  not
  g1452
  (
    n1586,
    n1109
  );


  not
  g1453
  (
    n1393,
    n1141
  );


  buf
  g1454
  (
    n1599,
    n1135
  );


  buf
  g1455
  (
    n1640,
    n1124
  );


  buf
  g1456
  (
    n1469,
    n1149
  );


  not
  g1457
  (
    n1390,
    n956
  );


  buf
  g1458
  (
    n1547,
    n1129
  );


  not
  g1459
  (
    n1405,
    n1116
  );


  not
  g1460
  (
    n1360,
    n1151
  );


  buf
  g1461
  (
    n1545,
    n615
  );


  not
  g1462
  (
    n1500,
    n1120
  );


  not
  g1463
  (
    n1486,
    n1126
  );


  buf
  g1464
  (
    n1416,
    n1128
  );


  not
  g1465
  (
    n1527,
    n1147
  );


  not
  g1466
  (
    n1560,
    n1133
  );


  buf
  g1467
  (
    n1468,
    n1107
  );


  buf
  g1468
  (
    n1583,
    n1107
  );


  buf
  g1469
  (
    n1622,
    n1138
  );


  buf
  g1470
  (
    n1582,
    n1150
  );


  buf
  g1471
  (
    n1600,
    n1143
  );


  not
  g1472
  (
    n1466,
    n1097
  );


  not
  g1473
  (
    n1497,
    n1161
  );


  not
  g1474
  (
    n1597,
    n1123
  );


  buf
  g1475
  (
    n1632,
    n1115
  );


  not
  g1476
  (
    n1362,
    n1112
  );


  not
  g1477
  (
    n1457,
    n830
  );


  not
  g1478
  (
    n1649,
    n1152
  );


  not
  g1479
  (
    n1526,
    n955
  );


  buf
  g1480
  (
    n1452,
    n1106
  );


  not
  g1481
  (
    n1542,
    n831
  );


  not
  g1482
  (
    n1378,
    n1099
  );


  not
  g1483
  (
    n1580,
    n951
  );


  buf
  g1484
  (
    n1558,
    n1097
  );


  buf
  g1485
  (
    n1428,
    n775
  );


  not
  g1486
  (
    n1618,
    n892
  );


  buf
  g1487
  (
    n1592,
    n1117
  );


  buf
  g1488
  (
    n1623,
    n831
  );


  buf
  g1489
  (
    n1463,
    n1167
  );


  buf
  g1490
  (
    n1546,
    n1115
  );


  buf
  g1491
  (
    n1585,
    n1104
  );


  not
  g1492
  (
    n1552,
    n1124
  );


  buf
  g1493
  (
    n1414,
    n1164
  );


  not
  g1494
  (
    n1626,
    n952
  );


  buf
  g1495
  (
    n1567,
    n1140
  );


  not
  g1496
  (
    n1606,
    n1116
  );


  buf
  g1497
  (
    n1633,
    n1139
  );


  not
  g1498
  (
    n1493,
    n1153
  );


  not
  g1499
  (
    n1651,
    n1117
  );


  not
  g1500
  (
    n1489,
    n1125
  );


  not
  g1501
  (
    n1383,
    n1129
  );


  not
  g1502
  (
    n1642,
    n1159
  );


  buf
  g1503
  (
    n1634,
    n779
  );


  not
  g1504
  (
    n1517,
    n1169
  );


  buf
  g1505
  (
    n1426,
    n1100
  );


  buf
  g1506
  (
    n1369,
    n1105
  );


  not
  g1507
  (
    n1575,
    n1122
  );


  buf
  g1508
  (
    n1375,
    n1143
  );


  not
  g1509
  (
    n1490,
    n1149
  );


  not
  g1510
  (
    n1458,
    n1113
  );


  buf
  g1511
  (
    n1531,
    n1126
  );


  buf
  g1512
  (
    n1607,
    n1120
  );


  not
  g1513
  (
    n1430,
    n831
  );


  buf
  g1514
  (
    n1363,
    n1138
  );


  not
  g1515
  (
    n1604,
    n1137
  );


  buf
  g1516
  (
    n1441,
    n912
  );


  not
  g1517
  (
    n1370,
    n1106
  );


  not
  g1518
  (
    n1401,
    n1098
  );


  buf
  g1519
  (
    n1454,
    n1104
  );


  buf
  g1520
  (
    n1381,
    n1169
  );


  buf
  g1521
  (
    n1533,
    n1118
  );


  buf
  g1522
  (
    n1544,
    n1153
  );


  not
  g1523
  (
    n1568,
    n1127
  );


  not
  g1524
  (
    n1535,
    n1095
  );


  not
  g1525
  (
    n1359,
    n1157
  );


  buf
  g1526
  (
    n1519,
    n1143
  );


  not
  g1527
  (
    n1423,
    n1114
  );


  not
  g1528
  (
    n1513,
    n776
  );


  not
  g1529
  (
    n1445,
    n776
  );


  buf
  g1530
  (
    n1596,
    n1163
  );


  not
  g1531
  (
    n1472,
    n1110
  );


  buf
  g1532
  (
    n1397,
    n1103
  );


  not
  g1533
  (
    n1411,
    n1146
  );


  not
  g1534
  (
    n1451,
    n1096
  );


  buf
  g1535
  (
    n1562,
    n1140
  );


  not
  g1536
  (
    n1412,
    n1160
  );


  buf
  g1537
  (
    n1609,
    n1107
  );


  buf
  g1538
  (
    n1570,
    n1163
  );


  not
  g1539
  (
    n1420,
    n1130
  );


  not
  g1540
  (
    n1473,
    n1167
  );


  buf
  g1541
  (
    n1587,
    n1139
  );


  not
  g1542
  (
    n1627,
    n1121
  );


  not
  g1543
  (
    n1357,
    n1113
  );


  buf
  g1544
  (
    n1507,
    n1145
  );


  not
  g1545
  (
    n1650,
    n1106
  );


  buf
  g1546
  (
    n1491,
    n1168
  );


  buf
  g1547
  (
    n1481,
    n1142
  );


  buf
  g1548
  (
    n1499,
    n1155
  );


  not
  g1549
  (
    n1503,
    n1161
  );


  buf
  g1550
  (
    n1553,
    n1164
  );


  not
  g1551
  (
    n1516,
    n1148
  );


  not
  g1552
  (
    n1641,
    n1150
  );


  not
  g1553
  (
    n1501,
    n1160
  );


  buf
  g1554
  (
    n1407,
    n1170
  );


  buf
  g1555
  (
    n1628,
    n1159
  );


  buf
  g1556
  (
    n1438,
    n1151
  );


  not
  g1557
  (
    n1479,
    n957
  );


  buf
  g1558
  (
    n1421,
    n1151
  );


  buf
  g1559
  (
    n1432,
    n955
  );


  buf
  g1560
  (
    n1541,
    n1168
  );


  not
  g1561
  (
    n1402,
    n1164
  );


  buf
  g1562
  (
    n1394,
    n953
  );


  not
  g1563
  (
    n1425,
    n1096
  );


  buf
  g1564
  (
    n1352,
    n1150
  );


  buf
  g1565
  (
    n1525,
    n1110
  );


  not
  g1566
  (
    n1522,
    n1119
  );


  not
  g1567
  (
    n1391,
    n1140
  );


  not
  g1568
  (
    n1595,
    n1102
  );


  buf
  g1569
  (
    n1467,
    n1156
  );


  not
  g1570
  (
    n1415,
    n1108
  );


  not
  g1571
  (
    n1376,
    n1101
  );


  not
  g1572
  (
    n1492,
    n951
  );


  buf
  g1573
  (
    n1400,
    n614
  );


  buf
  g1574
  (
    KeyWire_0_6,
    n1101
  );


  buf
  g1575
  (
    n1435,
    n1126
  );


  not
  g1576
  (
    n1537,
    n1117
  );


  not
  g1577
  (
    n1557,
    n1125
  );


  not
  g1578
  (
    n1574,
    n957
  );


  buf
  g1579
  (
    n1528,
    n777
  );


  buf
  g1580
  (
    n1448,
    n1171
  );


  buf
  g1581
  (
    n1494,
    n1112
  );


  buf
  g1582
  (
    n1565,
    n1113
  );


  buf
  g1583
  (
    n1532,
    n1132
  );


  not
  g1584
  (
    n1598,
    n1154
  );


  not
  g1585
  (
    n1368,
    n1123
  );


  not
  g1586
  (
    n1482,
    n1119
  );


  not
  g1587
  (
    n1538,
    n777
  );


  buf
  g1588
  (
    KeyWire_0_5,
    n954
  );


  buf
  g1589
  (
    n1615,
    n1117
  );


  not
  g1590
  (
    n1518,
    n1155
  );


  not
  g1591
  (
    n1417,
    n1111
  );


  not
  g1592
  (
    n1358,
    n1157
  );


  buf
  g1593
  (
    n1483,
    n951
  );


  not
  g1594
  (
    n1429,
    n1118
  );


  not
  g1595
  (
    n1377,
    n1105
  );


  not
  g1596
  (
    n1403,
    n1158
  );


  buf
  g1597
  (
    n1474,
    n781
  );


  and
  g1598
  (
    n1387,
    n1159,
    n1146,
    n1141,
    n1156
  );


  xor
  g1599
  (
    n1564,
    n1167,
    n1137,
    n774,
    n1136
  );


  nand
  g1600
  (
    n1365,
    n1144,
    n1142,
    n1132,
    n1136
  );


  or
  g1601
  (
    n1461,
    n1147,
    n1156,
    n1154,
    n1101
  );


  xnor
  g1602
  (
    KeyWire_0_10,
    n1149,
    n1105,
    n1168,
    n1125
  );


  nand
  g1603
  (
    n1384,
    n830,
    n1138,
    n1104
  );


  nor
  g1604
  (
    n1440,
    n1165,
    n1144,
    n1155,
    n1170
  );


  nor
  g1605
  (
    n1529,
    n160,
    n1110,
    n1120,
    n616
  );


  and
  g1606
  (
    n1418,
    n1158,
    n1133,
    n952,
    n160
  );


  and
  g1607
  (
    n1643,
    n1166,
    n1151,
    n1145,
    n892
  );


  nand
  g1608
  (
    n1443,
    n1129,
    n1133,
    n1116,
    n1098
  );


  xor
  g1609
  (
    n1470,
    n1121,
    n1165,
    n1099,
    n1127
  );


  or
  g1610
  (
    n1379,
    n1122,
    n1100,
    n1128,
    n1160
  );


  nand
  g1611
  (
    n1590,
    n1154,
    n1137,
    n1127,
    n1097
  );


  nand
  g1612
  (
    n1367,
    n1108,
    n1135,
    n1164,
    n1148
  );


  or
  g1613
  (
    n1540,
    n1163,
    n954,
    n1131,
    n1108
  );


  and
  g1614
  (
    n1613,
    n1123,
    n1162,
    n1100
  );


  xnor
  g1615
  (
    n1511,
    n1130,
    n1168,
    n955,
    n1131
  );


  or
  g1616
  (
    n1534,
    n892,
    n1135,
    n1132,
    n1148
  );


  or
  g1617
  (
    n1437,
    n1103,
    n1131,
    n1163,
    n1140
  );


  or
  g1618
  (
    n1505,
    n1121,
    n956,
    n1157,
    n1165
  );


  or
  g1619
  (
    n1713,
    n1627,
    n1176
  );


  xor
  g1620
  (
    n1834,
    n1253,
    n1295
  );


  xnor
  g1621
  (
    n1889,
    n1367,
    n1288
  );


  xor
  g1622
  (
    n1811,
    n1625,
    n1631
  );


  nand
  g1623
  (
    n1692,
    n1271,
    n1293
  );


  xnor
  g1624
  (
    n1867,
    n1191,
    n1382,
    n1206,
    n1230
  );


  or
  g1625
  (
    n1727,
    n1181,
    n1270,
    n1391,
    n1298
  );


  xnor
  g1626
  (
    n1810,
    n1257,
    n1502,
    n1493,
    n1411
  );


  nand
  g1627
  (
    n1804,
    n1468,
    n1338,
    n1210,
    n1319
  );


  nand
  g1628
  (
    n1896,
    n1218,
    n1465,
    n1268,
    n1301
  );


  xor
  g1629
  (
    n1933,
    n1360,
    n1430,
    n1262,
    n1288
  );


  or
  g1630
  (
    n1908,
    n1602,
    n1451,
    n1224,
    n1646
  );


  nand
  g1631
  (
    n1919,
    n1222,
    n1533,
    n1318,
    n1254
  );


  xnor
  g1632
  (
    n1738,
    n1315,
    n1459,
    n1252,
    n1225
  );


  and
  g1633
  (
    n1931,
    n1347,
    n1349,
    n1199,
    n1598
  );


  or
  g1634
  (
    n1895,
    n1205,
    n1179,
    n1245,
    n1256
  );


  nor
  g1635
  (
    n1735,
    n1259,
    n1422,
    n1549,
    n1236
  );


  and
  g1636
  (
    n1687,
    n1223,
    n1348,
    n1618,
    n1631
  );


  nor
  g1637
  (
    n1877,
    n1575,
    n1364,
    n1570,
    n1198
  );


  nand
  g1638
  (
    n1654,
    n1535,
    n1487,
    n1264,
    n1247
  );


  xnor
  g1639
  (
    n1802,
    n1175,
    n1629,
    n1610,
    n1222
  );


  nand
  g1640
  (
    n1677,
    n1241,
    n1246,
    n1392,
    n1435
  );


  xnor
  g1641
  (
    n1803,
    n1607,
    n1331,
    n1208,
    n1268
  );


  or
  g1642
  (
    n1756,
    n1340,
    n1621,
    n1179,
    n1221
  );


  or
  g1643
  (
    n1824,
    n1322,
    n1196,
    n1265,
    n1243
  );


  or
  g1644
  (
    n1830,
    n1240,
    n1599,
    n1538,
    n1302
  );


  xor
  g1645
  (
    n1904,
    n1269,
    n1286,
    n1339,
    n1501
  );


  and
  g1646
  (
    n1717,
    n1174,
    n1643,
    n1226,
    n1349
  );


  and
  g1647
  (
    n1697,
    n1284,
    n1321,
    n1238,
    n1455
  );


  or
  g1648
  (
    n1890,
    n1280,
    n1304,
    n1426,
    n1516
  );


  or
  g1649
  (
    n1920,
    n1563,
    n1243,
    n1526,
    n1447
  );


  or
  g1650
  (
    n1917,
    n1190,
    n1283,
    n1212,
    n1220
  );


  nand
  g1651
  (
    n1840,
    n1186,
    n1216,
    n1200,
    n1287
  );


  xor
  g1652
  (
    n1750,
    n1587,
    n1618,
    n1349,
    n1201
  );


  xnor
  g1653
  (
    n1854,
    n1223,
    n1216,
    n1233,
    n1291
  );


  or
  g1654
  (
    n1884,
    n1542,
    n1202,
    n1309,
    n1299
  );


  nand
  g1655
  (
    n1859,
    n1325,
    n1542,
    n1581,
    n1571
  );


  and
  g1656
  (
    n1792,
    n1284,
    n1587,
    n1252,
    n1576
  );


  or
  g1657
  (
    n1669,
    n1197,
    n1579,
    n1286,
    n1211
  );


  xor
  g1658
  (
    n1716,
    n1292,
    n1244,
    n1424,
    n1180
  );


  and
  g1659
  (
    n1746,
    n1554,
    n1449,
    n1358,
    n1472
  );


  and
  g1660
  (
    n1674,
    n1547,
    n1417,
    n1176,
    n1216
  );


  nand
  g1661
  (
    n1764,
    n1420,
    n1198,
    n1208,
    n1621
  );


  or
  g1662
  (
    n1790,
    n1644,
    n1228,
    n1195,
    n1186
  );


  nor
  g1663
  (
    n1652,
    n1205,
    n1540,
    n1597,
    n1337
  );


  or
  g1664
  (
    n1894,
    n1323,
    n1215,
    n1399,
    n1303
  );


  or
  g1665
  (
    n1762,
    n1185,
    n1578,
    n1627,
    n1194
  );


  nor
  g1666
  (
    n1852,
    n1346,
    n1637,
    n1340,
    n1603
  );


  or
  g1667
  (
    n1843,
    n1187,
    n1567,
    n1223,
    n1552
  );


  xor
  g1668
  (
    n1748,
    n1329,
    n1240,
    n1540,
    n1312
  );


  xor
  g1669
  (
    n1733,
    n1456,
    n1172,
    n1419,
    n1193
  );


  nor
  g1670
  (
    n1671,
    n1546,
    n1461,
    n1616,
    n1593
  );


  xnor
  g1671
  (
    n1696,
    n1274,
    n1580,
    n1638,
    n1334
  );


  xor
  g1672
  (
    n1845,
    n1291,
    n1494,
    n1277,
    n1350
  );


  and
  g1673
  (
    n1729,
    n1479,
    n1406,
    n1269,
    n1612
  );


  and
  g1674
  (
    n1875,
    n1189,
    n1341,
    n1371,
    n1323
  );


  xor
  g1675
  (
    n1722,
    n1234,
    n1286,
    n1275,
    n1529
  );


  nand
  g1676
  (
    n1685,
    n1250,
    n1278,
    n1336,
    n1171
  );


  nand
  g1677
  (
    n1797,
    n1513,
    n1553,
    n1259,
    n1243
  );


  nor
  g1678
  (
    n1848,
    n1197,
    n1244,
    n1189,
    n1332
  );


  xor
  g1679
  (
    n1666,
    n1236,
    n1244,
    n1217,
    n1546
  );


  xor
  g1680
  (
    n1712,
    n1298,
    n1605,
    n1445,
    n1242
  );


  nand
  g1681
  (
    n1778,
    n1248,
    n1569,
    n1317,
    n1288
  );


  and
  g1682
  (
    n1771,
    n1277,
    n1550,
    n1649,
    n1283
  );


  nand
  g1683
  (
    n1751,
    n1650,
    n1336,
    n1267,
    n1186
  );


  nand
  g1684
  (
    n1715,
    n1192,
    n1335,
    n1207,
    n1251
  );


  xor
  g1685
  (
    n1846,
    n1279,
    n1324,
    n1243,
    n1647
  );


  xor
  g1686
  (
    n1780,
    n1213,
    n1639,
    n1568,
    n1188
  );


  nor
  g1687
  (
    n1873,
    n1385,
    n1577,
    n1551,
    n1314
  );


  or
  g1688
  (
    n1839,
    n1281,
    n1262,
    n1195,
    n1218
  );


  xnor
  g1689
  (
    n1885,
    n1555,
    n1208,
    n1440,
    n1596
  );


  nand
  g1690
  (
    n1740,
    n1266,
    n1238,
    n1172,
    n1633
  );


  and
  g1691
  (
    n1849,
    n1598,
    n1390,
    n1608,
    n1318
  );


  xnor
  g1692
  (
    n1863,
    n1315,
    n1327,
    n1640,
    n1184
  );


  or
  g1693
  (
    n1928,
    n1294,
    n1590,
    n1272,
    n1350
  );


  xor
  g1694
  (
    n1711,
    n1594,
    n1299,
    n1312,
    n1211
  );


  nor
  g1695
  (
    n1822,
    n1297,
    n1444,
    n1527,
    n1254
  );


  nand
  g1696
  (
    n1864,
    n1251,
    n1230,
    n1550,
    n1192
  );


  nand
  g1697
  (
    n1660,
    n1345,
    n1326,
    n1321,
    n1193
  );


  xor
  g1698
  (
    n1903,
    n1596,
    n1376,
    n1290,
    n1626
  );


  or
  g1699
  (
    n1847,
    n1384,
    n1204,
    n1221,
    n1295
  );


  or
  g1700
  (
    n1878,
    n1226,
    n1477,
    n1267,
    n1316
  );


  and
  g1701
  (
    n1888,
    n1344,
    n1614,
    n1443,
    n1327
  );


  xor
  g1702
  (
    n1892,
    n1231,
    n1327,
    n1250,
    n1308
  );


  or
  g1703
  (
    n1857,
    n1279,
    n1271,
    n1562,
    n1346
  );


  xnor
  g1704
  (
    n1865,
    n1612,
    n1434,
    n1256,
    n1309
  );


  nand
  g1705
  (
    n1719,
    n1316,
    n1475,
    n1600,
    n1223
  );


  nand
  g1706
  (
    n1680,
    n1191,
    n1531,
    n1270,
    n1374
  );


  nor
  g1707
  (
    n1815,
    n1273,
    n1244,
    n1327,
    n1340
  );


  and
  g1708
  (
    n1708,
    n1232,
    n1474,
    n1320,
    n1263
  );


  nor
  g1709
  (
    n1765,
    n1261,
    n1204,
    n1218,
    n1642
  );


  xor
  g1710
  (
    n1667,
    n1259,
    n1563,
    n1219,
    n1568
  );


  nor
  g1711
  (
    n1682,
    n1348,
    n1330,
    n1416,
    n1202
  );


  xnor
  g1712
  (
    n1714,
    n1350,
    n1308,
    n1270,
    n1423
  );


  nand
  g1713
  (
    n1786,
    n1274,
    n1305,
    n1566,
    n1574
  );


  nor
  g1714
  (
    n1883,
    n1203,
    n1383,
    n1496,
    n1249
  );


  xor
  g1715
  (
    n1731,
    n1481,
    n1213,
    n1573,
    n1337
  );


  or
  g1716
  (
    n1862,
    n1307,
    n1395,
    n1324,
    n1293
  );


  nand
  g1717
  (
    n1791,
    n1614,
    n1208,
    n1242,
    n1448
  );


  xnor
  g1718
  (
    n1684,
    n1258,
    n1336,
    n1279
  );


  nand
  g1719
  (
    n1755,
    n1381,
    n1316,
    n1620,
    n1184
  );


  and
  g1720
  (
    n1800,
    n1324,
    n1201,
    n1256,
    n1304
  );


  and
  g1721
  (
    n1930,
    n1281,
    n1649,
    n1225,
    n1490
  );


  xor
  g1722
  (
    n1835,
    n1190,
    n1300,
    n1272,
    n1641
  );


  nor
  g1723
  (
    n1679,
    n1585,
    n1397,
    n1173,
    n1204
  );


  or
  g1724
  (
    n1906,
    n1495,
    n1403,
    n1373,
    n1177
  );


  nand
  g1725
  (
    n1709,
    n1595,
    n1549,
    n1305,
    n1319
  );


  nor
  g1726
  (
    n1912,
    n1182,
    n1646,
    n1305,
    n1272
  );


  xnor
  g1727
  (
    n1837,
    n1273,
    n1184,
    n1354,
    n1398
  );


  and
  g1728
  (
    n1747,
    n1560,
    n1233,
    n1275,
    n1438
  );


  and
  g1729
  (
    n1730,
    n1175,
    n1615,
    n1588,
    n1604
  );


  nor
  g1730
  (
    n1785,
    n1431,
    n1293,
    n1264,
    n1269
  );


  xor
  g1731
  (
    n1703,
    n1258,
    n1331,
    n1302,
    n1328
  );


  nand
  g1732
  (
    n1720,
    n1582,
    n1262,
    n1242,
    n1349
  );


  nand
  g1733
  (
    n1818,
    n1339,
    n1561,
    n1484,
    n1464
  );


  nor
  g1734
  (
    n1869,
    n1321,
    n1263,
    n1343,
    n1375
  );


  nand
  g1735
  (
    n1916,
    n1193,
    n1648,
    n1285,
    n1278
  );


  nand
  g1736
  (
    n1825,
    n1589,
    n1310,
    n1368,
    n1630
  );


  xor
  g1737
  (
    n1882,
    n1571,
    n1184,
    n1418,
    n1644
  );


  xor
  g1738
  (
    n1900,
    n1210,
    n1269,
    n1557,
    n1548
  );


  xor
  g1739
  (
    n1808,
    n1648,
    n1203,
    n1266,
    n1335
  );


  nor
  g1740
  (
    n1773,
    n1207,
    n1307,
    n1603,
    n1215
  );


  or
  g1741
  (
    n1768,
    n1638,
    n1251,
    n1510,
    n1558
  );


  and
  g1742
  (
    n1793,
    n1466,
    n1282,
    n1637,
    n1225
  );


  and
  g1743
  (
    n1898,
    n1341,
    n1362,
    n1264,
    n1179
  );


  and
  g1744
  (
    n1718,
    n1345,
    n1452,
    n1237,
    n1255
  );


  and
  g1745
  (
    n1861,
    n1228,
    n1304,
    n1326,
    n1314
  );


  nand
  g1746
  (
    n1876,
    n1592,
    n1252,
    n1273,
    n1209
  );


  and
  g1747
  (
    n1723,
    n1213,
    n1635,
    n1338,
    n1551
  );


  nor
  g1748
  (
    n1787,
    n1567,
    n1640,
    n1219,
    n1522
  );


  or
  g1749
  (
    n1705,
    n1559,
    n1387,
    n1181,
    n1604
  );


  xnor
  g1750
  (
    n1925,
    n1343,
    n1232,
    n1306,
    n1497
  );


  xnor
  g1751
  (
    n1910,
    n1583,
    n1185,
    n1203,
    n1409
  );


  xor
  g1752
  (
    n1659,
    n1572,
    n1485,
    n1258,
    n1247
  );


  xnor
  g1753
  (
    n1907,
    n1289,
    n1199,
    n1508,
    n1365
  );


  nand
  g1754
  (
    n1820,
    n1293,
    n1601,
    n1191,
    n1338
  );


  or
  g1755
  (
    n1686,
    n1177,
    n1189,
    n1498,
    n1295
  );


  xor
  g1756
  (
    n1655,
    n1183,
    n1471,
    n1347,
    n1322
  );


  and
  g1757
  (
    n1743,
    n1565,
    n1235,
    n1492,
    n1347
  );


  or
  g1758
  (
    n1668,
    n1334,
    n1476,
    n1308,
    n1339
  );


  nand
  g1759
  (
    n1741,
    n1237,
    n1330,
    n1311,
    n1187
  );


  or
  g1760
  (
    n1770,
    n1228,
    n1297,
    n1341,
    n1266
  );


  xnor
  g1761
  (
    n1656,
    n1400,
    n1217,
    n1333,
    n1436
  );


  nor
  g1762
  (
    n1812,
    n1279,
    n1276,
    n1318,
    n1410
  );


  or
  g1763
  (
    n1763,
    n1249,
    n1317,
    n1286,
    n1222
  );


  and
  g1764
  (
    n1827,
    n1333,
    n1335,
    n1172,
    n1599
  );


  nor
  g1765
  (
    n1689,
    n1199,
    n1623,
    n1363,
    n1389
  );


  or
  g1766
  (
    n1658,
    n1331,
    n1408,
    n1200,
    n1544
  );


  nor
  g1767
  (
    n1798,
    n1194,
    n1241,
    n1582,
    n1313
  );


  xnor
  g1768
  (
    n1683,
    n1482,
    n1624,
    n1275,
    n1346
  );


  or
  g1769
  (
    n1886,
    n1241,
    n1266,
    n1180,
    n1556
  );


  nor
  g1770
  (
    n1922,
    n1632,
    n1307,
    n1246,
    n1296
  );


  nor
  g1771
  (
    n1758,
    n1523,
    n1317,
    n1331,
    n1290
  );


  xnor
  g1772
  (
    n1657,
    n1359,
    n1181,
    n1229,
    n1205
  );


  nor
  g1773
  (
    n1879,
    n1611,
    n1287,
    n1235,
    n1366
  );


  xor
  g1774
  (
    n1901,
    n1232,
    n1314,
    n1521,
    n1317
  );


  nor
  g1775
  (
    n1871,
    n1532,
    n1350,
    n1272,
    n1217
  );


  and
  g1776
  (
    n1672,
    n1344,
    n1217,
    n1234,
    n1320
  );


  nor
  g1777
  (
    n1844,
    n1348,
    n1173,
    n1589,
    n1342
  );


  and
  g1778
  (
    n1831,
    n1287,
    n1200,
    n1203,
    n1558
  );


  nor
  g1779
  (
    n1914,
    n1229,
    n1388,
    n1597,
    n1301
  );


  xor
  g1780
  (
    n1734,
    n1310,
    n1326,
    n1281,
    n1210
  );


  nand
  g1781
  (
    n1935,
    n1469,
    n1480,
    n1488,
    n1261
  );


  nor
  g1782
  (
    n1742,
    n1348,
    n1285,
    n1559,
    n1183
  );


  nor
  g1783
  (
    n1860,
    n1230,
    n1178,
    n1507,
    n1292
  );


  or
  g1784
  (
    n1784,
    n1536,
    n1248,
    n1219,
    n1294
  );


  xor
  g1785
  (
    n1782,
    n1214,
    n1277,
    n1564,
    n1478
  );


  nor
  g1786
  (
    n1868,
    n1220,
    n1378,
    n1177,
    n1641
  );


  nor
  g1787
  (
    n1813,
    n1594,
    n1188,
    n1216,
    n1517
  );


  nor
  g1788
  (
    n1921,
    n1226,
    n1427,
    n1187,
    n1602
  );


  and
  g1789
  (
    n1927,
    n1341,
    n1302,
    n1609,
    n1323
  );


  or
  g1790
  (
    n1829,
    n1311,
    n1425,
    n1306,
    n1209
  );


  or
  g1791
  (
    n1700,
    n1324,
    n1463,
    n1591,
    n1296
  );


  xor
  g1792
  (
    n1691,
    n1231,
    n1547,
    n1428,
    n1180
  );


  and
  g1793
  (
    n1681,
    n1450,
    n1271,
    n1414,
    n1247
  );


  or
  g1794
  (
    n1752,
    n1514,
    n1569,
    n1626,
    n1625
  );


  nor
  g1795
  (
    n1833,
    n1633,
    n1229,
    n1233,
    n1239
  );


  xnor
  g1796
  (
    n1779,
    n1642,
    n1322,
    n1467,
    n1185
  );


  or
  g1797
  (
    n1745,
    n1259,
    n1290,
    n1257,
    n1305
  );


  nor
  g1798
  (
    n1766,
    n1647,
    n1178,
    n1212,
    n1191
  );


  xnor
  g1799
  (
    n1856,
    n1607,
    n1619,
    n1329,
    n1309
  );


  and
  g1800
  (
    n1832,
    n1292,
    n1613,
    n1310,
    n1294
  );


  xor
  g1801
  (
    n1805,
    n1611,
    n1296,
    n1544,
    n1421
  );


  nand
  g1802
  (
    n1781,
    n1282,
    n1628,
    n1296,
    n1268
  );


  or
  g1803
  (
    n1725,
    n1289,
    n1302,
    n1572,
    n1337
  );


  xor
  g1804
  (
    n1902,
    n1263,
    n1325,
    n1393,
    n1312
  );


  and
  g1805
  (
    n1721,
    n1189,
    n1174,
    n1240,
    n1630
  );


  and
  g1806
  (
    n1788,
    n1528,
    n1209,
    n1271,
    n1330
  );


  or
  g1807
  (
    n1934,
    n1173,
    n1511,
    n1340,
    n1457
  );


  xor
  g1808
  (
    n1851,
    n1345,
    n1210,
    n1462,
    n1316
  );


  nand
  g1809
  (
    n1688,
    n1181,
    n1273,
    n1323,
    n1311
  );


  and
  g1810
  (
    n1929,
    n1636,
    n1377,
    n1584,
    n1174
  );


  xor
  g1811
  (
    n1694,
    n1545,
    n1192,
    n1294,
    n1329
  );


  and
  g1812
  (
    n1704,
    n1446,
    n1261,
    n1247,
    n1215
  );


  and
  g1813
  (
    n1838,
    n1303,
    n1556,
    n1206,
    n1442
  );


  xnor
  g1814
  (
    n1905,
    n1239,
    n1407,
    n1255,
    n1454
  );


  xnor
  g1815
  (
    n1662,
    n1283,
    n1277,
    n1352,
    n1193
  );


  or
  g1816
  (
    n1663,
    n1206,
    n1634,
    n1519,
    n1175
  );


  and
  g1817
  (
    n1855,
    n1298,
    n1342,
    n1228,
    n1226
  );


  and
  g1818
  (
    n1707,
    n1332,
    n1282,
    n1328,
    n1234
  );


  nand
  g1819
  (
    n1913,
    n1285,
    n1543,
    n1227,
    n1574
  );


  or
  g1820
  (
    n1665,
    n1288,
    n1345,
    n1315,
    n1576
  );


  or
  g1821
  (
    n1932,
    n1192,
    n1586,
    n1332,
    n1608
  );


  nand
  g1822
  (
    n1728,
    n1473,
    n1562,
    n1251,
    n1301
  );


  xnor
  g1823
  (
    n1874,
    n1224,
    n1617,
    n1307,
    n1212
  );


  xnor
  g1824
  (
    n1673,
    n1372,
    n1312,
    n1541,
    n1622
  );


  nand
  g1825
  (
    n1821,
    n1301,
    n1380,
    n1588,
    n1254
  );


  nor
  g1826
  (
    n1783,
    n1263,
    n1636,
    n1617,
    n1579
  );


  and
  g1827
  (
    n1816,
    n1541,
    n1214,
    n1554,
    n1275
  );


  xor
  g1828
  (
    n1866,
    n1174,
    n1276,
    n1248,
    n1214
  );


  nor
  g1829
  (
    n1695,
    n1319,
    n1289,
    n1237,
    n1429
  );


  and
  g1830
  (
    n1795,
    n1278,
    n1353,
    n1202,
    n1267
  );


  nand
  g1831
  (
    n1767,
    n1321,
    n1236,
    n1235,
    n1592
  );


  xor
  g1832
  (
    n1858,
    n1234,
    n1342,
    n1356,
    n1183
  );


  and
  g1833
  (
    n1776,
    n1308,
    n1245,
    n1261,
    n1609
  );


  or
  g1834
  (
    n1826,
    n1314,
    n1176,
    n1242,
    n1441
  );


  nor
  g1835
  (
    n1853,
    n1322,
    n1270,
    n1333,
    n1291
  );


  nor
  g1836
  (
    n1698,
    n1326,
    n1555,
    n1188,
    n1186
  );


  xnor
  g1837
  (
    n1870,
    n1415,
    n1282,
    n1343,
    n1591
  );


  and
  g1838
  (
    n1749,
    n1311,
    n1204,
    n1328,
    n1402
  );


  xnor
  g1839
  (
    n1807,
    n1530,
    n1586,
    n1584,
    n1320
  );


  xor
  g1840
  (
    n1926,
    n1183,
    n1396,
    n1284,
    n1583
  );


  nor
  g1841
  (
    n1724,
    n1566,
    n1218,
    n1267,
    n1553
  );


  and
  g1842
  (
    n1678,
    n1632,
    n1460,
    n1255,
    n1347
  );


  and
  g1843
  (
    n1923,
    n1231,
    n1194,
    n1458,
    n1483
  );


  or
  g1844
  (
    n1732,
    n1197,
    n1287,
    n1285,
    n1280
  );


  nor
  g1845
  (
    n1911,
    n1334,
    n1361,
    n1173,
    n1209
  );


  and
  g1846
  (
    n1760,
    n1178,
    n1564,
    n1334,
    n1593
  );


  xnor
  g1847
  (
    n1675,
    n1211,
    n1239,
    n1254,
    n1175
  );


  xor
  g1848
  (
    n1676,
    n1578,
    n1299,
    n1229,
    n1620
  );


  xor
  g1849
  (
    n1769,
    n1306,
    n1539,
    n1297,
    n1240
  );


  and
  g1850
  (
    n1872,
    n1249,
    n1236,
    n1338,
    n1300
  );


  nand
  g1851
  (
    n1841,
    n1265,
    n1643,
    n1355,
    n1320
  );


  or
  g1852
  (
    n1737,
    n1503,
    n1188,
    n1238,
    n1537
  );


  nor
  g1853
  (
    n1836,
    n1245,
    n1344,
    n1227,
    n1525
  );


  and
  g1854
  (
    n1772,
    n1211,
    n1573,
    n1585,
    n1187
  );


  nand
  g1855
  (
    n1744,
    n1257,
    n1199,
    n1258,
    n1313
  );


  nor
  g1856
  (
    n1909,
    n1190,
    n1299,
    n1575,
    n1265
  );


  xor
  g1857
  (
    n1789,
    n1303,
    n1198,
    n1520,
    n1628
  );


  or
  g1858
  (
    n1736,
    n1278,
    n1605,
    n1329,
    n1212
  );


  xnor
  g1859
  (
    n1842,
    n1198,
    n1412,
    n1600,
    n1645
  );


  and
  g1860
  (
    n1661,
    n1227,
    n1518,
    n1225,
    n1500
  );


  and
  g1861
  (
    n1881,
    n1274,
    n1313,
    n1509,
    n1610
  );


  nor
  g1862
  (
    n1775,
    n1201,
    n1230,
    n1196,
    n1231
  );


  or
  g1863
  (
    n1828,
    n1232,
    n1241,
    n1202,
    n1570
  );


  and
  g1864
  (
    n1774,
    n1245,
    n1595,
    n1257,
    n1601
  );


  or
  g1865
  (
    n1806,
    n1280,
    n1437,
    n1577,
    n1224
  );


  or
  g1866
  (
    n1936,
    n1539,
    n1176,
    n1504,
    n1246
  );


  and
  g1867
  (
    n1761,
    n1512,
    n1250,
    n1506,
    n1260
  );


  xor
  g1868
  (
    n1701,
    n1171,
    n1295,
    n1239,
    n1623
  );


  nor
  g1869
  (
    n1915,
    n1561,
    n1253,
    n1335,
    n1246
  );


  nor
  g1870
  (
    n1702,
    n1224,
    n1557,
    n1179,
    n1325
  );


  or
  g1871
  (
    n1880,
    n1180,
    n1276,
    n1260,
    n1250
  );


  nor
  g1872
  (
    n1817,
    n1178,
    n1325,
    n1433,
    n1639
  );


  nor
  g1873
  (
    n1693,
    n1580,
    n1337,
    n1306,
    n1260
  );


  nor
  g1874
  (
    n1670,
    n1268,
    n1543,
    n1291,
    n1284
  );


  and
  g1875
  (
    n1850,
    n1214,
    n1297,
    n1303,
    n1545
  );


  xor
  g1876
  (
    n1819,
    n1613,
    n1206,
    n1255,
    n1221
  );


  and
  g1877
  (
    n1706,
    n1194,
    n1343,
    n1252,
    n1264
  );


  xnor
  g1878
  (
    n1897,
    n1524,
    n1262,
    n1439,
    n1565
  );


  or
  g1879
  (
    n1653,
    n1195,
    n1237,
    n1344,
    n1339
  );


  xor
  g1880
  (
    n1664,
    n1207,
    n1342,
    n1309,
    n1394
  );


  or
  g1881
  (
    n1814,
    n1629,
    n1196,
    n1197,
    n1499
  );


  nand
  g1882
  (
    n1893,
    n1298,
    n1182,
    n1470,
    n1190
  );


  nand
  g1883
  (
    n1726,
    n1238,
    n1634,
    n1207,
    n1172
  );


  and
  g1884
  (
    n1809,
    n1379,
    n1606,
    n1233,
    n1276
  );


  xnor
  g1885
  (
    n1891,
    n1635,
    n1369,
    n1205,
    n1215
  );


  xor
  g1886
  (
    n1823,
    n1235,
    n1219,
    n1315,
    n1292
  );


  or
  g1887
  (
    n1924,
    n1248,
    n1453,
    n1328,
    n1182
  );


  or
  g1888
  (
    n1699,
    n1290,
    n1220,
    n1357,
    n1274
  );


  and
  g1889
  (
    n1799,
    n1489,
    n1622,
    n1249,
    n1201
  );


  and
  g1890
  (
    n1794,
    n1505,
    n1318,
    n1491,
    n1624
  );


  xnor
  g1891
  (
    n1899,
    n1280,
    n1289,
    n1581,
    n1300
  );


  nand
  g1892
  (
    n1757,
    n1548,
    n1222,
    n1386,
    n1606
  );


  nor
  g1893
  (
    n1759,
    n1413,
    n1552,
    n1330,
    n1283
  );


  and
  g1894
  (
    n1777,
    n1220,
    n1310,
    n1370,
    n1650
  );


  xnor
  g1895
  (
    n1754,
    n1332,
    n1560,
    n1195,
    n1304
  );


  or
  g1896
  (
    n1753,
    n1182,
    n1486,
    n1227,
    n1196
  );


  xor
  g1897
  (
    n1796,
    n1313,
    n1534,
    n1432,
    n1200
  );


  or
  g1898
  (
    n1710,
    n1319,
    n1256,
    n1615,
    n1619
  );


  nor
  g1899
  (
    n1739,
    n1300,
    n1281,
    n1405,
    n1590
  );


  nand
  g1900
  (
    n1887,
    n1213,
    n1221,
    n1253
  );


  and
  g1901
  (
    n1801,
    n1333,
    n1265,
    n1346,
    n1401
  );


  xnor
  g1902
  (
    n1918,
    n1351,
    n1185,
    n1616,
    n1515
  );


  xnor
  g1903
  (
    n1690,
    n1177,
    n1404,
    n1260,
    n1645
  );


  xor
  g1904
  (
    n1964,
    n1733,
    n1767,
    n1745,
    n1699
  );


  xnor
  g1905
  (
    n1968,
    n1654,
    n1709,
    n1764,
    n1723
  );


  and
  g1906
  (
    n1966,
    n1737,
    n1781,
    n1683,
    n1710
  );


  and
  g1907
  (
    n1942,
    n1729,
    n1681,
    n1760,
    n1782
  );


  nor
  g1908
  (
    n1953,
    n1720,
    n1742,
    n1675,
    n1778
  );


  xnor
  g1909
  (
    n1944,
    n1722,
    n1713,
    n1670,
    n1653
  );


  nand
  g1910
  (
    n1957,
    n1665,
    n1652,
    n1669,
    n1712
  );


  or
  g1911
  (
    n1946,
    n1695,
    n1735,
    n1739,
    n1765
  );


  xor
  g1912
  (
    n1940,
    n1685,
    n1711,
    n1730,
    n1783
  );


  xnor
  g1913
  (
    n1938,
    n1751,
    n1750,
    n1721,
    n1775
  );


  nand
  g1914
  (
    n1962,
    n1757,
    n1756,
    n1655,
    n1771
  );


  or
  g1915
  (
    n1937,
    n1668,
    n1719,
    n1731,
    n1659
  );


  or
  g1916
  (
    n1941,
    n1700,
    n1740,
    n1662,
    n1776
  );


  xor
  g1917
  (
    n1963,
    n1738,
    n1785,
    n1706,
    n1688
  );


  xnor
  g1918
  (
    n1952,
    n1703,
    n1770,
    n1747,
    n1746
  );


  or
  g1919
  (
    n1956,
    n1741,
    n1761,
    n1656,
    n1680
  );


  or
  g1920
  (
    n1961,
    n1671,
    n1718,
    n1690,
    n1724
  );


  nor
  g1921
  (
    n1950,
    n1697,
    n1743,
    n1715,
    n1777
  );


  and
  g1922
  (
    n1943,
    n1678,
    n1784,
    n1780,
    n1657
  );


  or
  g1923
  (
    n1949,
    n1734,
    n1772,
    n1755,
    n1663
  );


  nor
  g1924
  (
    n1959,
    n1661,
    n1726,
    n1707,
    n1768
  );


  nand
  g1925
  (
    n1970,
    n1701,
    n1677,
    n1727,
    n1651
  );


  xor
  g1926
  (
    n1955,
    n1679,
    n1673,
    n1774,
    n1704
  );


  xor
  g1927
  (
    n1969,
    n1779,
    n1666,
    n1694,
    n1664
  );


  and
  g1928
  (
    n1958,
    n1773,
    n1651,
    n1660,
    n1732
  );


  nand
  g1929
  (
    n1951,
    n1762,
    n1754,
    n1748,
    n1687
  );


  xnor
  g1930
  (
    n1954,
    n1708,
    n1672,
    n1716,
    n1702
  );


  or
  g1931
  (
    n1948,
    n1692,
    n1684,
    n1758,
    n1693
  );


  nand
  g1932
  (
    KeyWire_0_0,
    n1698,
    n1689,
    n1725,
    n1686
  );


  or
  g1933
  (
    n1965,
    n1763,
    n1691,
    n1696,
    n1759
  );


  or
  g1934
  (
    n1939,
    n1717,
    n1752,
    n1769,
    n1766
  );


  xor
  g1935
  (
    n1945,
    n1753,
    n1658,
    n1705,
    n1676
  );


  nand
  g1936
  (
    n1947,
    n1714,
    n1744,
    n1667,
    n1682
  );


  nor
  g1937
  (
    n1967,
    n1728,
    n1736,
    n1749,
    n1674
  );


  xnor
  g1938
  (
    n1996,
    n1852,
    n1835,
    n1955,
    n1957
  );


  or
  g1939
  (
    n1985,
    n1942,
    n1854,
    n1954,
    n1822
  );


  or
  g1940
  (
    n2003,
    n1941,
    n1867,
    n1958,
    n1952
  );


  nand
  g1941
  (
    n1991,
    n1799,
    n1792,
    n1877,
    n1851
  );


  xor
  g1942
  (
    n1993,
    n1949,
    n1808,
    n1811,
    n1848
  );


  or
  g1943
  (
    n1982,
    n1853,
    n1857,
    n1875,
    n1850
  );


  xor
  g1944
  (
    n1987,
    n1815,
    n1810,
    n1796,
    n1879
  );


  xnor
  g1945
  (
    n2002,
    n1951,
    n1790,
    n1863,
    n1964
  );


  nor
  g1946
  (
    n1981,
    n1832,
    n1880,
    n1940,
    n1946
  );


  nand
  g1947
  (
    n1983,
    n1819,
    n1787,
    n1884,
    n1836
  );


  and
  g1948
  (
    n1995,
    n1807,
    n1806,
    n1801,
    n1814
  );


  and
  g1949
  (
    n1992,
    n1948,
    n1834,
    n1859,
    n1849
  );


  xnor
  g1950
  (
    n1976,
    n1829,
    n1959,
    n1786,
    n1858
  );


  nand
  g1951
  (
    n1998,
    n1825,
    n1864,
    n1874,
    n1789
  );


  nand
  g1952
  (
    n1988,
    n1800,
    n1883,
    n1813,
    n1860
  );


  and
  g1953
  (
    n1979,
    n1969,
    n1960,
    n1947,
    n1847
  );


  nor
  g1954
  (
    n1971,
    n1966,
    n1837,
    n1950,
    n1818
  );


  xor
  g1955
  (
    n1984,
    n1841,
    n1826,
    n1868,
    n1838
  );


  nor
  g1956
  (
    n2000,
    n1961,
    n1816,
    n1823,
    n1827
  );


  xor
  g1957
  (
    n1990,
    n1794,
    n1791,
    n1965,
    n1809
  );


  nand
  g1958
  (
    n1980,
    n1881,
    n1956,
    n1812,
    n1803
  );


  or
  g1959
  (
    n1975,
    n1871,
    n1817,
    n1830,
    n1970
  );


  nor
  g1960
  (
    n1973,
    n1831,
    n1967,
    n1802,
    n1963
  );


  xnor
  g1961
  (
    n1974,
    n1804,
    n1872,
    n1788,
    n1828
  );


  xor
  g1962
  (
    n1994,
    n1855,
    n1845,
    n1962,
    n1844
  );


  xor
  g1963
  (
    n2001,
    n1882,
    n1842,
    n1856,
    n1938
  );


  nand
  g1964
  (
    n1972,
    n1870,
    n1878,
    n1833,
    n1839
  );


  xnor
  g1965
  (
    n1989,
    n1861,
    n1869,
    n1876,
    n1873
  );


  xnor
  g1966
  (
    n1986,
    n1866,
    n1805,
    n1824,
    n1843
  );


  and
  g1967
  (
    n1997,
    n1795,
    n1953,
    n1865,
    n1846
  );


  nand
  g1968
  (
    n1978,
    n1793,
    n1820,
    n1840,
    n1821
  );


  nand
  g1969
  (
    n1977,
    n1943,
    n1798,
    n1944,
    n1862
  );


  or
  g1970
  (
    n1999,
    n1968,
    n1945,
    n1797,
    n1939
  );


  nand
  g1971
  (
    n2008,
    n1975,
    n1901,
    n1924,
    n1909
  );


  xnor
  g1972
  (
    n2010,
    n1918,
    n1903,
    n1934,
    n1893
  );


  or
  g1973
  (
    n2014,
    n1887,
    n1917,
    n1907,
    n1888
  );


  nand
  g1974
  (
    n2004,
    n1892,
    n1915,
    n1910,
    n1889
  );


  or
  g1975
  (
    n2021,
    n1902,
    n1891,
    n1971,
    n1912
  );


  and
  g1976
  (
    n2020,
    n1894,
    n618,
    n1983,
    n1990
  );


  xor
  g1977
  (
    n2018,
    n1988,
    n1906,
    n1992,
    n1899
  );


  and
  g1978
  (
    n2016,
    n1980,
    n1987,
    n1885,
    n1935
  );


  xnor
  g1979
  (
    n2006,
    n1977,
    n1925,
    n1900,
    n1922
  );


  xnor
  g1980
  (
    n2005,
    n1886,
    n1931,
    n1897,
    n1981
  );


  xor
  g1981
  (
    n2013,
    n1929,
    n1890,
    n1979,
    n1923
  );


  nor
  g1982
  (
    n2022,
    n1927,
    n1898,
    n1986,
    n1933
  );


  or
  g1983
  (
    n2009,
    n1913,
    n1908,
    n1905,
    n1982
  );


  nor
  g1984
  (
    n2019,
    n1991,
    n1973,
    n1930,
    n1920
  );


  nor
  g1985
  (
    n2015,
    n1921,
    n1984,
    n1926,
    n1896
  );


  and
  g1986
  (
    n2011,
    n1972,
    n1928,
    n1914,
    n1989
  );


  nand
  g1987
  (
    n2017,
    n1936,
    n1895,
    n1976,
    n1916
  );


  nor
  g1988
  (
    n2012,
    n1985,
    n619,
    n1978,
    n1919
  );


  xor
  g1989
  (
    n2007,
    n1911,
    n1932,
    n1904,
    n1974
  );


  nand
  g1990
  (
    n2028,
    n2002,
    n2015,
    n2003,
    n1997
  );


  nor
  g1991
  (
    n2027,
    n1994,
    n1998,
    n2001,
    n2014
  );


  nor
  g1992
  (
    n2030,
    n2022,
    n1995,
    n2004,
    n1993
  );


  nand
  g1993
  (
    n2023,
    n2013,
    n2012,
    n2008,
    n2020
  );


  nor
  g1994
  (
    n2029,
    n2000,
    n2006,
    n2017,
    n2011
  );


  and
  g1995
  (
    n2025,
    n2021,
    n2019,
    n2003,
    n2010
  );


  nor
  g1996
  (
    n2024,
    n160,
    n2007,
    n1996,
    n2016
  );


  xnor
  g1997
  (
    n2026,
    n2009,
    n2005,
    n1999,
    n2018
  );


  or
  g1998
  (
    n2032,
    n2025,
    n2026,
    n2023,
    n2029
  );


  nor
  g1999
  (
    n2031,
    n2027,
    n2030,
    n2024,
    n2028
  );


  xor
  KeyGate_0_0
  (
    n1960,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n135,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n138,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n905,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n671,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1646,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1351,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1510,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1581,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n787,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n1645,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1561,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n1591,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n658,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1153,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1644,
    KeyNOTWire_0_15
  );


endmodule

