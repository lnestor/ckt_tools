module MyXor(A, B, C);

input A, B;
output C;

xor XOR1(C, A, B);

endmodule

