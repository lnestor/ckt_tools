// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_834_381 written by SynthGen on 2021/05/24 19:48:31
module Stat_834_381( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31,
 n177, n183, n175, n176, n192, n194, n181, n186,
 n196, n189, n590, n597, n587, n840, n852, n854,
 n860, n861, n865);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31;

output n177, n183, n175, n176, n192, n194, n181, n186,
 n196, n189, n590, n597, n587, n840, n852, n854,
 n860, n861, n865;

wire n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n178,
 n179, n180, n182, n184, n185, n187, n188, n190,
 n191, n193, n195, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n588, n589, n591, n592, n593, n594, n595,
 n596, n598, n599, n600, n601, n602, n603, n604,
 n605, n606, n607, n608, n609, n610, n611, n612,
 n613, n614, n615, n616, n617, n618, n619, n620,
 n621, n622, n623, n624, n625, n626, n627, n628,
 n629, n630, n631, n632, n633, n634, n635, n636,
 n637, n638, n639, n640, n641, n642, n643, n644,
 n645, n646, n647, n648, n649, n650, n651, n652,
 n653, n654, n655, n656, n657, n658, n659, n660,
 n661, n662, n663, n664, n665, n666, n667, n668,
 n669, n670, n671, n672, n673, n674, n675, n676,
 n677, n678, n679, n680, n681, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n758, n759, n760, n761, n762, n763, n764,
 n765, n766, n767, n768, n769, n770, n771, n772,
 n773, n774, n775, n776, n777, n778, n779, n780,
 n781, n782, n783, n784, n785, n786, n787, n788,
 n789, n790, n791, n792, n793, n794, n795, n796,
 n797, n798, n799, n800, n801, n802, n803, n804,
 n805, n806, n807, n808, n809, n810, n811, n812,
 n813, n814, n815, n816, n817, n818, n819, n820,
 n821, n822, n823, n824, n825, n826, n827, n828,
 n829, n830, n831, n832, n833, n834, n835, n836,
 n837, n838, n839, n841, n842, n843, n844, n845,
 n846, n847, n848, n849, n850, n851, n853, n855,
 n856, n857, n858, n859, n862, n863, n864;

not  g0 (n64, n9);
not  g1 (n33, n25);
not  g2 (n47, n23);
not  g3 (n83, n3);
not  g4 (n61, n8);
buf  g5 (n74, n12);
not  g6 (n77, n27);
buf  g7 (n49, n30);
not  g8 (n93, n25);
not  g9 (n34, n10);
buf  g10 (n106, n14);
buf  g11 (n105, n5);
buf  g12 (n92, n10);
not  g13 (n78, n15);
not  g14 (n109, n13);
not  g15 (n69, n6);
not  g16 (n118, n10);
buf  g17 (n44, n20);
not  g18 (n97, n31);
not  g19 (n68, n30);
not  g20 (n96, n14);
buf  g21 (n115, n5);
buf  g22 (n98, n27);
buf  g23 (n42, n18);
buf  g24 (n95, n19);
buf  g25 (n41, n12);
buf  g26 (n123, n5);
not  g27 (n122, n6);
buf  g28 (n54, n21);
buf  g29 (n50, n26);
buf  g30 (n103, n15);
buf  g31 (n101, n16);
not  g32 (n121, n20);
buf  g33 (n84, n4);
buf  g34 (n38, n11);
buf  g35 (n37, n29);
not  g36 (n85, n24);
buf  g37 (n51, n16);
not  g38 (n46, n31);
buf  g39 (n32, n3);
not  g40 (n53, n1);
not  g41 (n90, n18);
not  g42 (n110, n17);
not  g43 (n35, n27);
buf  g44 (n89, n7);
not  g45 (n56, n28);
buf  g46 (n111, n2);
buf  g47 (n102, n30);
not  g48 (n100, n31);
not  g49 (n72, n6);
not  g50 (n71, n2);
not  g51 (n60, n4);
not  g52 (n79, n13);
not  g53 (n108, n7);
not  g54 (n65, n9);
buf  g55 (n91, n1);
buf  g56 (n63, n17);
buf  g57 (n99, n26);
buf  g58 (n66, n8);
buf  g59 (n45, n13);
not  g60 (n57, n28);
buf  g61 (n82, n25);
buf  g62 (n70, n4);
buf  g63 (n39, n1);
buf  g64 (n117, n21);
buf  g65 (n58, n17);
not  g66 (n59, n7);
buf  g67 (n114, n24);
not  g68 (n107, n19);
not  g69 (n86, n22);
buf  g70 (n67, n22);
buf  g71 (n76, n23);
buf  g72 (n52, n16);
buf  g73 (n62, n21);
not  g74 (n113, n11);
not  g75 (n55, n3);
not  g76 (n104, n20);
buf  g77 (n81, n19);
buf  g78 (n119, n22);
buf  g79 (n40, n12);
buf  g80 (n87, n2);
not  g81 (n112, n18);
not  g82 (n94, n8);
not  g83 (n36, n28);
buf  g84 (n120, n26);
buf  g85 (n73, n15);
not  g86 (n124, n29);
not  g87 (n75, n29);
buf  g88 (n48, n24);
not  g89 (n116, n11);
not  g90 (n80, n14);
buf  g91 (n88, n9);
not  g92 (n43, n23);
buf  g93 (n170, n41);
not  g94 (n145, n59);
not  g95 (n160, n79);
buf  g96 (n159, n55);
not  g97 (n136, n49);
buf  g98 (n167, n59);
not  g99 (n157, n44);
buf  g100 (n152, n73);
buf  g101 (n132, n76);
nand g102 (n137, n60, n62);
or   g103 (n171, n58, n62, n84, n80);
nand g104 (n133, n77, n51, n74);
xnor g105 (n149, n44, n52, n58, n87);
nor  g106 (n166, n76, n32, n68, n81);
xnor g107 (n150, n61, n32, n46, n54);
xnor g108 (n165, n37, n86, n36, n87);
and  g109 (n155, n43, n69, n64, n40);
xor  g110 (n172, n51, n64, n63, n86);
xor  g111 (n144, n49, n70, n45, n60);
xor  g112 (n128, n80, n75, n50);
nand g113 (n158, n57, n43, n42, n66);
xnor g114 (n127, n41, n72, n83, n74);
xor  g115 (n139, n35, n72, n85, n67);
nor  g116 (n151, n67, n85, n77, n65);
xor  g117 (n129, n73, n78, n50, n39);
and  g118 (n135, n71, n66, n36, n62);
xor  g119 (n156, n44, n40, n79, n33);
or   g120 (n126, n63, n85, n71, n84);
nor  g121 (n163, n82, n48, n46, n84);
and  g122 (n148, n48, n35, n82, n56);
xnor g123 (n162, n69, n64, n53, n49);
and  g124 (n154, n61, n55, n72, n78);
or   g125 (n169, n71, n39, n37, n35);
xnor g126 (n168, n83, n55, n33, n76);
nand g127 (n141, n47, n81, n51, n50);
or   g128 (n164, n48, n38);
and  g129 (n138, n37, n56, n34, n79);
or   g130 (n134, n39, n61, n34, n57);
nand g131 (n173, n33, n69, n36, n60);
xor  g132 (n146, n47, n65, n45, n56);
xnor g133 (n143, n57, n83, n54, n80);
or   g134 (n142, n43, n75, n86, n59);
xor  g135 (n130, n82, n52, n70);
or   g136 (n161, n70, n77, n67, n66);
or   g137 (n125, n41, n46, n42);
xor  g138 (n153, n40, n78, n65, n32);
and  g139 (n147, n47, n58, n53, n68);
nand g140 (n140, n53, n45, n81, n54);
or   g141 (n131, n73, n68, n34, n63);
not  g142 (n197, n126);
not  g143 (n194, n140);
buf  g144 (n195, n133);
buf  g145 (n174, n152);
not  g146 (n181, n128);
buf  g147 (n200, n146);
buf  g148 (n180, n138);
buf  g149 (n182, n127);
not  g150 (n198, n145);
not  g151 (n183, n141);
not  g152 (n178, n139);
buf  g153 (n189, n137);
not  g154 (n185, n142);
buf  g155 (n201, n136);
buf  g156 (n190, n149);
buf  g157 (n184, n129);
buf  g158 (n193, n125);
buf  g159 (n177, n144);
not  g160 (n179, n130);
buf  g161 (n187, n143);
buf  g162 (n186, n134);
buf  g163 (n196, n132);
not  g164 (n199, n151);
buf  g165 (n176, n148);
buf  g166 (n192, n147);
not  g167 (n188, n131);
not  g168 (n191, n135);
buf  g169 (n175, n150);
not  g170 (n205, n89);
not  g171 (n210, n89);
buf  g172 (n213, n197);
buf  g173 (n206, n198);
not  g174 (n216, n190);
buf  g175 (n207, n192);
not  g176 (n215, n191);
not  g177 (n204, n193);
not  g178 (n212, n186);
buf  g179 (n203, n187);
buf  g180 (n219, n201);
not  g181 (n209, n194);
buf  g182 (n208, n195);
not  g183 (n214, n199);
nor  g184 (n218, n89, n88);
nor  g185 (n211, n196, n88, n188, n90);
nand g186 (n217, n184, n200, n90, n88);
and  g187 (n202, n189, n87, n185, n90);
buf  g188 (n223, n208);
not  g189 (n222, n202);
and  g190 (n220, n206, n209);
xnor g191 (n227, n203, n210);
and  g192 (n228, n209, n206, n204, n205);
and  g193 (n226, n203, n205, n209, n210);
nor  g194 (n225, n208, n211, n210, n202);
xor  g195 (n229, n207, n206, n211, n208);
xnor g196 (n221, n204, n202, n207, n211);
nor  g197 (n224, n203, n205, n204, n207);
buf  g198 (n236, n226);
buf  g199 (n231, n227);
not  g200 (n234, n225);
not  g201 (n230, n222);
buf  g202 (n232, n221);
buf  g203 (n238, n224);
buf  g204 (n237, n223);
not  g205 (n235, n228);
not  g206 (n233, n220);
not  g207 (n240, n235);
not  g208 (n241, n236);
not  g209 (n247, n232);
not  g210 (n239, n231);
not  g211 (n254, n232);
not  g212 (n257, n235);
buf  g213 (n255, n236);
buf  g214 (n243, n234);
not  g215 (n251, n233);
buf  g216 (n242, n233);
buf  g217 (n244, n232);
buf  g218 (n245, n230);
not  g219 (n246, n234);
not  g220 (n250, n230);
not  g221 (n248, n231);
buf  g222 (n256, n231);
buf  g223 (n249, n234);
not  g224 (n252, n233);
buf  g225 (n253, n235);
buf  g226 (n258, n230);
buf  g227 (n272, n244);
not  g228 (n264, n212);
not  g229 (n285, n216);
not  g230 (n283, n251);
not  g231 (n280, n246);
buf  g232 (n259, n242);
buf  g233 (n282, n258);
not  g234 (n278, n249);
not  g235 (n267, n213);
not  g236 (n274, n243);
buf  g237 (n269, n249);
not  g238 (n270, n153);
xor  g239 (n276, n216, n255, n239, n248);
xor  g240 (n260, n244, n256, n240, n248);
xor  g241 (n281, n215, n241, n250, n252);
xnor g242 (n265, n154, n241, n250, n156);
or   g243 (n262, n215, n253, n244, n251);
nor  g244 (n273, n243, n248, n241, n254);
or   g245 (n271, n254, n245, n216, n257);
and  g246 (n266, n247, n252, n251, n249);
nand g247 (n287, n213, n213, n246, n240);
xnor g248 (n275, n157, n215, n256, n254);
xnor g249 (n279, n214, n155, n239, n258);
nor  g250 (n263, n252, n258, n214, n250);
or   g251 (n277, n257, n257, n242, n253);
nand g252 (n284, n253, n245, n242, n214);
and  g253 (n261, n246, n256, n255, n245);
and  g254 (n286, n239, n247, n243, n212);
xor  g255 (n268, n212, n247, n240, n255);
buf  g256 (n302, n264);
buf  g257 (n308, n263);
buf  g258 (n301, n271);
not  g259 (n298, n277);
not  g260 (n289, n275);
buf  g261 (n290, n276);
not  g262 (n294, n273);
buf  g263 (n300, n274);
not  g264 (n297, n265);
not  g265 (n309, n266);
not  g266 (n292, n261);
not  g267 (n304, n260);
not  g268 (n296, n270);
buf  g269 (n293, n278);
not  g270 (n305, n276);
buf  g271 (n306, n277);
buf  g272 (n307, n267);
not  g273 (n295, n272);
buf  g274 (n303, n268);
buf  g275 (n299, n275);
not  g276 (n310, n262);
buf  g277 (n291, n259);
buf  g278 (n288, n278);
buf  g279 (n311, n269);
not  g280 (n319, n288);
not  g281 (n325, n290);
buf  g282 (n320, n289);
not  g283 (n326, n292);
buf  g284 (n313, n290);
not  g285 (n321, n295);
buf  g286 (n312, n289);
buf  g287 (n317, n288);
not  g288 (n323, n290);
not  g289 (n316, n296);
nor  g290 (n318, n294, n293, n295);
xnor g291 (n322, n294, n296, n292, n295);
xnor g292 (n324, n291, n293, n288, n297);
xnor g293 (n315, n291, n289, n296, n292);
nor  g294 (n314, n291, n294, n297);
not  g295 (n331, n322);
buf  g296 (n345, n312);
buf  g297 (n342, n316);
buf  g298 (n338, n321);
buf  g299 (n335, n313);
not  g300 (n343, n324);
buf  g301 (n328, n321);
buf  g302 (n339, n318);
buf  g303 (n337, n323);
buf  g304 (n340, n323);
not  g305 (n344, n325);
not  g306 (n332, n325);
not  g307 (n327, n317);
not  g308 (n336, n326);
not  g309 (n330, n314);
buf  g310 (n329, n315);
buf  g311 (n333, n324);
buf  g312 (n341, n320);
buf  g313 (n334, n322);
buf  g314 (n346, n319);
buf  g315 (n359, n346);
buf  g316 (n362, n343);
not  g317 (n361, n93);
buf  g318 (n348, n95);
not  g319 (n368, n238);
buf  g320 (n352, n100);
buf  g321 (n353, n94);
not  g322 (n369, n96);
buf  g323 (n351, n101);
buf  g324 (n364, n328);
nor  g325 (n355, n342, n237);
and  g326 (n354, n336, n329, n99, n327);
nor  g327 (n366, n94, n99, n339, n344);
and  g328 (n370, n331, n330, n101, n237);
xnor g329 (n365, n96, n333, n100, n101);
xnor g330 (n349, n345, n103, n97, n343);
nor  g331 (n367, n338, n99, n92, n102);
or   g332 (n357, n332, n96, n92, n97);
and  g333 (n347, n340, n91, n102, n97);
nor  g334 (n372, n236, n103, n93, n238);
or   g335 (n363, n94, n335, n346, n342);
nand g336 (n371, n344, n334, n98, n95);
nor  g337 (n360, n93, n237, n103, n238);
or   g338 (n356, n98, n95, n341, n102);
nand g339 (n350, n345, n91, n337);
and  g340 (n358, n98, n92, n100, n341);
buf  g341 (n373, n301);
not  g342 (n375, n303);
buf  g343 (n393, n299);
buf  g344 (n418, n368);
not  g345 (n415, n302);
not  g346 (n403, n302);
not  g347 (n389, n104);
buf  g348 (n376, n350);
buf  g349 (n387, n302);
not  g350 (n402, n355);
buf  g351 (n416, n349);
buf  g352 (n411, n218);
buf  g353 (n392, n362);
not  g354 (n413, n367);
buf  g355 (n412, n303);
buf  g356 (n381, n300);
not  g357 (n408, n219);
buf  g358 (n386, n363);
not  g359 (n390, n219);
buf  g360 (n400, n359);
not  g361 (n420, n303);
not  g362 (n417, n358);
buf  g363 (n394, n105);
not  g364 (n414, n354);
not  g365 (n382, n368);
buf  g366 (n378, n298);
not  g367 (n391, n218);
buf  g368 (n406, n356);
not  g369 (n384, n369);
not  g370 (n401, n370);
nand g371 (n424, n217, n351, n106);
nor  g372 (n383, n371, n347, n108);
and  g373 (n385, n217, n105, n360);
nor  g374 (n374, n219, n108, n369);
xnor g375 (n422, n357, n352, n300);
xnor g376 (n419, n356, n106, n347);
nor  g377 (n379, n107, n364);
and  g378 (n410, n298, n355, n371);
nand g379 (n397, n353, n107, n108);
or   g380 (n396, n360, n300, n217);
nor  g381 (n398, n104, n354, n366);
xor  g382 (n388, n106, n365, n362);
nand g383 (n395, n351, n104, n348);
xnor g384 (n409, n105, n361, n218);
nor  g385 (n423, n357, n298, n109);
nor  g386 (n399, n301, n358, n367);
and  g387 (n407, n301, n361, n372);
nand g388 (n421, n299, n107, n359);
and  g389 (n380, n370, n352, n372);
and  g390 (n377, n365, n363, n366);
nor  g391 (n404, n349, n350, n299);
xor  g392 (n405, n353, n348, n109);
buf  g393 (n468, n390);
not  g394 (n427, n413);
buf  g395 (n443, n404);
buf  g396 (n511, n380);
not  g397 (n448, n380);
buf  g398 (n469, n410);
not  g399 (n487, n390);
buf  g400 (n545, n385);
buf  g401 (n445, n401);
buf  g402 (n562, n379);
buf  g403 (n461, n389);
buf  g404 (n464, n391);
not  g405 (n442, n399);
not  g406 (n564, n399);
not  g407 (n539, n393);
not  g408 (n538, n409);
not  g409 (n555, n417);
buf  g410 (n561, n379);
not  g411 (n536, n403);
not  g412 (n513, n408);
not  g413 (n466, n381);
buf  g414 (n432, n415);
not  g415 (n475, n382);
not  g416 (n566, n400);
buf  g417 (n472, n415);
not  g418 (n494, n402);
buf  g419 (n485, n417);
not  g420 (n527, n398);
not  g421 (n535, n407);
not  g422 (n517, n400);
buf  g423 (n462, n397);
buf  g424 (n565, n392);
not  g425 (n433, n413);
not  g426 (n543, n397);
not  g427 (n530, n406);
not  g428 (n456, n406);
not  g429 (n471, n376);
buf  g430 (n467, n416);
buf  g431 (n457, n404);
buf  g432 (n495, n394);
not  g433 (n544, n378);
buf  g434 (n516, n414);
not  g435 (n463, n409);
not  g436 (n453, n384);
not  g437 (n506, n389);
not  g438 (n431, n393);
buf  g439 (n449, n396);
not  g440 (n434, n376);
not  g441 (n512, n383);
not  g442 (n437, n402);
not  g443 (n482, n375);
not  g444 (n502, n410);
buf  g445 (n438, n396);
not  g446 (n473, n381);
buf  g447 (n440, n412);
buf  g448 (n515, n373);
buf  g449 (n501, n404);
buf  g450 (n531, n411);
not  g451 (n558, n417);
buf  g452 (n490, n398);
not  g453 (n533, n419);
not  g454 (n550, n377);
buf  g455 (n508, n373);
not  g456 (n521, n405);
not  g457 (n559, n401);
not  g458 (n505, n382);
buf  g459 (n476, n403);
buf  g460 (n478, n403);
not  g461 (n548, n387);
not  g462 (n451, n384);
buf  g463 (n509, n418);
not  g464 (n481, n391);
buf  g465 (n557, n397);
not  g466 (n452, n411);
not  g467 (n454, n374);
buf  g468 (n522, n378);
buf  g469 (n524, n405);
not  g470 (n503, n416);
buf  g471 (n491, n392);
buf  g472 (n430, n398);
not  g473 (n534, n395);
buf  g474 (n514, n418);
not  g475 (n529, n386);
buf  g476 (n426, n412);
buf  g477 (n542, n419);
buf  g478 (n553, n380);
not  g479 (n504, n413);
buf  g480 (n450, n393);
not  g481 (n435, n420);
not  g482 (n460, n374);
buf  g483 (n519, n375);
not  g484 (n439, n399);
not  g485 (n477, n394);
buf  g486 (n540, n388);
buf  g487 (n479, n412);
not  g488 (n441, n386);
buf  g489 (n554, n389);
not  g490 (n486, n382);
buf  g491 (n549, n383);
buf  g492 (n458, n406);
buf  g493 (n520, n414);
not  g494 (n560, n401);
not  g495 (n470, n390);
not  g496 (n444, n375);
buf  g497 (n436, n408);
not  g498 (n541, n388);
buf  g499 (n447, n387);
not  g500 (n551, n416);
buf  g501 (n455, n411);
not  g502 (n489, n376);
not  g503 (n499, n407);
buf  g504 (n429, n415);
not  g505 (n507, n419);
buf  g506 (n525, n379);
not  g507 (n497, n384);
buf  g508 (n484, n395);
not  g509 (n492, n378);
buf  g510 (n459, n374);
buf  g511 (n563, n396);
not  g512 (n537, n385);
buf  g513 (n474, n402);
not  g514 (n552, n418);
buf  g515 (n523, n383);
not  g516 (n500, n409);
not  g517 (n547, n377);
not  g518 (n480, n386);
not  g519 (n532, n385);
not  g520 (n546, n407);
buf  g521 (n526, n395);
buf  g522 (n496, n373);
buf  g523 (n465, n408);
not  g524 (n518, n387);
not  g525 (n528, n410);
buf  g526 (n493, n381);
buf  g527 (n498, n391);
buf  g528 (n488, n394);
not  g529 (n425, n377);
not  g530 (n556, n400);
not  g531 (n446, n388);
buf  g532 (n428, n414);
buf  g533 (n483, n392);
buf  g534 (n510, n405);
buf  g535 (n578, n436);
not  g536 (n568, n427);
buf  g537 (n574, n435);
not  g538 (n576, n428);
not  g539 (n572, n438);
not  g540 (n577, n434);
buf  g541 (n570, n432);
not  g542 (n575, n430);
buf  g543 (n571, n437);
nor  g544 (n580, n426, n437, n429);
nand g545 (n573, n434, n429, n433, n431);
xnor g546 (n579, n428, n438, n430, n432);
nor  g547 (n567, n426, n427, n436, n431);
or   g548 (n569, n425, n425, n433, n435);
xor  g549 (n597, n446, n443, n579);
or   g550 (n591, n578, n571, n439, n569);
nand g551 (n594, n447, n574, n567, n445);
and  g552 (n593, n568, n571, n572, n569);
xnor g553 (n595, n578, n568, n577);
and  g554 (n598, n569, n576, n570, n446);
or   g555 (n586, n567, n574, n439);
or   g556 (n584, n110, n579, n567, n444);
nor  g557 (n583, n580, n578, n577, n576);
nand g558 (n581, n579, n573, n110, n440);
or   g559 (n582, n447, n575, n576);
nor  g560 (n590, n448, n572, n570, n580);
xnor g561 (n585, n109, n579, n578, n575);
xnor g562 (n592, n576, n442, n440, n570);
xnor g563 (n587, n441, n442, n444, n580);
xor  g564 (n596, n575, n111, n573);
xnor g565 (n589, n445, n580, n577);
and  g566 (n588, n572, n571, n110, n441);
buf  g567 (n602, n592);
not  g568 (n613, n587);
not  g569 (n601, n590);
buf  g570 (n611, n596);
not  g571 (n609, n597);
buf  g572 (n612, n585);
not  g573 (n608, n593);
buf  g574 (n610, n584);
not  g575 (n599, n589);
not  g576 (n600, n588);
not  g577 (n604, n586);
buf  g578 (n607, n591);
not  g579 (n605, n595);
not  g580 (n603, n111);
or   g581 (n606, n594, n598);
xor  g582 (n652, n466, n498, n487);
nand g583 (n662, n599, n483, n456, n601);
and  g584 (n638, n612, n472, n606, n502);
nand g585 (n620, n478, n492, n509, n493);
and  g586 (n621, n485, n448, n606, n601);
nor  g587 (n635, n609, n495, n490, n610);
nand g588 (n632, n458, n602, n506, n607);
nand g589 (n616, n471, n602, n603, n501);
xor  g590 (n648, n613, n497, n304, n599);
or   g591 (n642, n457, n473, n496, n604);
xor  g592 (n647, n482, n456, n612, n304);
xnor g593 (n637, n453, n499, n493, n506);
nand g594 (n660, n304, n500, n484, n476);
nand g595 (n619, n492, n496, n477, n475);
and  g596 (n655, n611, n491, n490, n487);
or   g597 (n640, n478, n472, n508, n449);
nand g598 (n653, n305, n504, n454, n505);
nand g599 (n624, n607, n449, n450, n600);
nor  g600 (n631, n455, n603, n479, n488);
xor  g601 (n644, n494, n475, n465, n605);
or   g602 (n622, n604, n502, n613, n496);
and  g603 (n649, n610, n458, n509, n499);
nor  g604 (n651, n450, n468, n501, n504);
xnor g605 (n643, n474, n451, n459, n489);
or   g606 (n656, n493, n457, n507, n506);
nand g607 (n614, n491, n503, n602, n467);
xor  g608 (n615, n611, n486, n489, n607);
nand g609 (n636, n495, n500, n507, n461);
xnor g610 (n623, n476, n494, n468, n500);
nor  g611 (n626, n611, n505, n600, n601);
xor  g612 (n654, n471, n499, n610, n606);
and  g613 (n630, n599, n613, n484, n464);
xor  g614 (n625, n609, n466, n463, n477);
and  g615 (n659, n507, n480, n470, n464);
or   g616 (n645, n503, n454, n467, n460);
and  g617 (n646, n608, n462, n501, n612);
nor  g618 (n641, n603, n460, n605, n498);
or   g619 (n633, n459, n504, n488, n495);
xnor g620 (n618, n481, n485, n469, n608);
and  g621 (n657, n452, n481, n473, n502);
xnor g622 (n639, n470, n489, n455, n505);
or   g623 (n658, n451, n482, n483, n611);
nand g624 (n634, n604, n508, n474, n453);
xor  g625 (n650, n605, n508, n490, n612);
nor  g626 (n617, n465, n461, n463, n479);
xnor g627 (n627, n480, n494, n497, n452);
nand g628 (n628, n469, n609, n491, n462);
xnor g629 (n629, n608, n497, n492, n610);
nand g630 (n661, n486, n503, n613, n600);
or   g631 (n700, n645, n531, n117, n617);
xor  g632 (n717, n539, n555, n650, n111);
or   g633 (n698, n518, n662, n658, n529);
nand g634 (n670, n625, n639, n647, n517);
or   g635 (n694, n538, n546, n639, n541);
and  g636 (n709, n537, n654, n633, n645);
xor  g637 (n676, n622, n531, n114, n519);
xnor g638 (n715, n626, n513, n115, n116);
nand g639 (n672, n620, n648, n531, n638);
nand g640 (n739, n545, n646, n533, n523);
nor  g641 (n663, n521, n620, n510, n549);
xnor g642 (n678, n513, n619, n541, n642);
xnor g643 (n691, n637, n638, n520, n646);
or   g644 (n701, n556, n656, n555);
and  g645 (n683, n642, n420, n651, n614);
xnor g646 (n696, n634, n524, n512, n616);
xor  g647 (n667, n641, n525, n650, n516);
or   g648 (n737, n615, n618, n113, n625);
nor  g649 (n723, n546, n621, n533, n515);
nor  g650 (n679, n661, n545, n112, n641);
or   g651 (n689, n659, n550, n622, n657);
and  g652 (n680, n654, n615, n634, n625);
xnor g653 (n684, n516, n550, n545, n636);
nor  g654 (n703, n534, n420, n547, n523);
nand g655 (n695, n629, n525, n535);
and  g656 (n736, n618, n624, n650, n631);
xor  g657 (n688, n540, n643, n554, n543);
xor  g658 (n735, n624, n635, n645, n513);
xor  g659 (n732, n113, n647, n619, n511);
nor  g660 (n674, n656, n644, n623, n528);
nor  g661 (n729, n522, n547, n516, n633);
nor  g662 (n675, n116, n552, n640, n626);
or   g663 (n666, n640, n114, n536, n526);
nor  g664 (n693, n653, n511, n518, n548);
nor  g665 (n710, n529, n655, n617, n648);
nor  g666 (n681, n551, n651, n547, n660);
xor  g667 (n721, n649, n542, n662);
nor  g668 (n692, n636, n662, n525, n551);
nand g669 (n685, n649, n517, n514, n526);
xnor g670 (n707, n652, n115, n616, n628);
nand g671 (n724, n661, n628, n634, n631);
and  g672 (n690, n522, n655, n627, n537);
xnor g673 (n708, n540, n532, n112, n549);
xor  g674 (n699, n517, n658, n524, n530);
and  g675 (n719, n648, n640, n512, n553);
and  g676 (n671, n550, n637, n642, n655);
xor  g677 (n726, n643, n512, n631, n515);
and  g678 (n668, n532, n552, n548, n649);
xnor g679 (n714, n526, n115, n623, n549);
or   g680 (n665, n538, n534, n639, n515);
nor  g681 (n702, n537, n519, n615, n632);
nand g682 (n704, n657, n544, n541, n546);
nor  g683 (n677, n646, n659, n621, n653);
nor  g684 (n731, n527, n536, n618, n651);
nand g685 (n728, n520, n556, n533, n626);
xor  g686 (n682, n629, n654, n658, n511);
or   g687 (n738, n628, n622, n112, n530);
and  g688 (n725, n551, n629, n630, n616);
xnor g689 (n673, n114, n528, n553, n635);
nor  g690 (n686, n633, n535, n552, n527);
xor  g691 (n734, n621, n544, n528, n521);
nor  g692 (n669, n614, n620, n518, n660);
nor  g693 (n687, n532, n540, n659, n638);
nor  g694 (n697, n660, n644, n627, n519);
xor  g695 (n727, n636, n637, n530, n553);
nor  g696 (n711, n539, n521, n623, n617);
xor  g697 (n733, n632, n635, n661, n652);
and  g698 (n722, n643, n630, n527);
nor  g699 (n706, n544, n652, n641, n644);
and  g700 (n705, n627, n534, n556, n523);
xnor g701 (n720, n619, n624, n522, n554);
nor  g702 (n730, n520, n539, n647, n632);
xor  g703 (n664, n554, n509, n548, n538);
and  g704 (n718, n510, n542, n555, n113);
xor  g705 (n713, n657, n543, n614, n653);
or   g706 (n716, n529, n543, n116, n536);
nand g707 (n712, n524, n514, n510);
or   g708 (n744, n683, n676, n665, n685);
nand g709 (n743, n672, n673, n670, n666);
or   g710 (n741, n667, n674, n664, n677);
and  g711 (n742, n668, n691, n679, n684);
nor  g712 (n745, n678, n688, n681, n689);
nand g713 (n747, n663, n686, n671, n692);
xor  g714 (n746, n669, n680, n682, n690);
xnor g715 (n740, n694, n675, n687, n693);
buf  g716 (n758, n743);
buf  g717 (n750, n743);
not  g718 (n748, n741);
not  g719 (n751, n746);
not  g720 (n757, n746);
not  g721 (n753, n742);
not  g722 (n766, n741);
buf  g723 (n759, n740);
buf  g724 (n755, n742);
not  g725 (n760, n743);
not  g726 (n765, n741);
not  g727 (n764, n744);
not  g728 (n752, n159);
buf  g729 (n754, n745);
and  g730 (n768, n745, n118);
xnor g731 (n767, n119, n743, n118, n747);
xnor g732 (n756, n695, n696, n747, n746);
xnor g733 (n761, n117, n744, n747, n742);
xor  g734 (n763, n744, n747, n746, n119);
nor  g735 (n749, n745, n158, n740, n117);
or   g736 (n769, n744, n742, n741, n119);
nand g737 (n762, n745, n740, n697, n118);
buf  g738 (n790, n768);
not  g739 (n785, n769);
buf  g740 (n774, n285);
buf  g741 (n788, n560);
buf  g742 (n784, n761);
buf  g743 (n771, n759);
and  g744 (n792, n284, n120, n559, n749);
xnor g745 (n782, n758, n120, n422, n757);
and  g746 (n779, n765, n283, n120, n423);
and  g747 (n791, n759, n422, n760);
xnor g748 (n776, n754, n557, n763, n285);
nand g749 (n786, n558, n766, n762);
or   g750 (n777, n750, n559, n560, n765);
xnor g751 (n787, n557, n422, n558, n282);
nand g752 (n775, n762, n286, n748, n421);
xor  g753 (n770, n283, n764, n121, n768);
xor  g754 (n783, n764, n761, n763, n561);
xnor g755 (n780, n769, n280, n281, n279);
and  g756 (n773, n755, n557, n558, n286);
nor  g757 (n772, n752, n281, n756, n767);
nand g758 (n789, n280, n282, n305, n421);
nor  g759 (n781, n767, n279, n284, n560);
nor  g760 (n778, n753, n751, n421, n559);
buf  g761 (n799, n770);
buf  g762 (n802, n779);
buf  g763 (n797, n776);
buf  g764 (n798, n777);
not  g765 (n800, n774);
buf  g766 (n795, n775);
buf  g767 (n794, n773);
buf  g768 (n793, n772);
not  g769 (n796, n778);
buf  g770 (n801, n771);
nor  g771 (n806, n793, n712, n160, n306);
xnor g772 (n818, n729, n800, n715, n727);
or   g773 (n821, n307, n792, n121, n802);
xor  g774 (n809, n795, n170, n736, n229);
and  g775 (n824, n561, n121, n308, n725);
or   g776 (n822, n166, n788, n800, n306);
or   g777 (n810, n739, n796, n167, n562);
nor  g778 (n815, n798, n782, n307, n733);
and  g779 (n805, n307, n801, n797);
and  g780 (n811, n171, n711, n699, n722);
nor  g781 (n812, n306, n787, n789, n802);
xnor g782 (n820, n793, n717, n703, n563);
or   g783 (n827, n709, n802, n737, n162);
nor  g784 (n819, n735, n308, n704, n706);
xor  g785 (n828, n718, n783, n786, n796);
nor  g786 (n817, n172, n720, n702, n705);
or   g787 (n804, n563, n710, n780, n790);
or   g788 (n832, n561, n799, n796, n173);
xnor g789 (n813, n714, n700, n164, n728);
nand g790 (n829, n784, n721, n708, n799);
nand g791 (n830, n781, n795, n169, n732);
or   g792 (n807, n161, n793, n798, n785);
and  g793 (n816, n730, n724, n738, n726);
and  g794 (n808, n562, n168, n163, n698);
xor  g795 (n825, n308, n701, n562, n723);
nand g796 (n823, n794, n563, n801, n305);
nor  g797 (n814, n800, n165, n731, n713);
nand g798 (n831, n719, n716, n795, n794);
or   g799 (n803, n707, n797, n794, n734);
and  g800 (n826, n791, n799, n798, n797);
not  g801 (n834, n804);
not  g802 (n833, n803);
and  g803 (n837, n807, n812, n806, n805);
or   g804 (n836, n808, n809, n810, n813);
xnor g805 (n835, n811, n833, n834);
not  g806 (n840, n836);
nand g807 (n842, n122, n836, n837);
or   g808 (n841, n424, n564, n836, n837);
xor  g809 (n839, n835, n564, n814);
or   g810 (n838, n815, n835, n565, n423);
xnor g811 (n843, n835, n423, n837, n816);
nand g812 (n844, n122, n839, n819, n817);
and  g813 (n846, n818, n841, n824, n565);
and  g814 (n845, n843, n820, n821, n122);
and  g815 (n847, n822, n823, n840, n842);
or   g816 (n849, n825, n847);
xor  g817 (n848, n845, n826, n123, n828);
and  g818 (n850, n846, n123, n827, n844);
buf  g819 (n851, n829);
or   g820 (n852, n848, n849, n124, n123);
or   g821 (n853, n852, n309);
and  g822 (n855, n853, n124, n424);
or   g823 (n854, n853, n287, n124);
nand g824 (n856, n855, n310);
xnor g825 (n858, n856, n326, n311);
xor  g826 (n857, n856, n311);
buf  g827 (n859, n850);
buf  g828 (n860, n858);
or   g829 (n861, n858, n857);
and  g830 (n862, n566, n566, n861, n565);
buf  g831 (n863, n862);
and  g832 (n864, n830, n862, n831);
xor  g833 (n865, n832, n566, n864, n863);
endmodule
