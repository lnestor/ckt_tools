

module Stat_2476_35_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n945,
  n954,
  n942,
  n951,
  n946,
  n965,
  n959,
  n950,
  n962,
  n964,
  n967,
  n966,
  n949,
  n960,
  n963,
  n943,
  n958,
  n957,
  n955,
  n956,
  n947,
  n961,
  n968,
  n971,
  n1022,
  n1086,
  n1085,
  n2508,
  n2512,
  n2513,
  n2510,
  n2514,
  n2516,
  n2515,
  n2509,
  n2518,
  n2511,
  n2519,
  n2517,
  n2507,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input n33;input n34;input n35;input n36;input n37;input n38;input n39;input n40;input n41;input n42;input n43;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n945;output n954;output n942;output n951;output n946;output n965;output n959;output n950;output n962;output n964;output n967;output n966;output n949;output n960;output n963;output n943;output n958;output n957;output n955;output n956;output n947;output n961;output n968;output n971;output n1022;output n1086;output n1085;output n2508;output n2512;output n2513;output n2510;output n2514;output n2516;output n2515;output n2509;output n2518;output n2511;output n2519;output n2517;output n2507;
  wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n944;wire n948;wire n952;wire n953;wire n969;wire n970;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  buf
  g0
  (
    n61,
    n16
  );


  buf
  g1
  (
    n176,
    n14
  );


  not
  g2
  (
    n200,
    n9
  );


  buf
  g3
  (
    n207,
    n27
  );


  not
  g4
  (
    n148,
    n12
  );


  buf
  g5
  (
    n156,
    n1
  );


  buf
  g6
  (
    n85,
    n43
  );


  not
  g7
  (
    n55,
    n21
  );


  not
  g8
  (
    n92,
    n20
  );


  buf
  g9
  (
    n69,
    n27
  );


  not
  g10
  (
    n122,
    n12
  );


  buf
  g11
  (
    n150,
    n14
  );


  buf
  g12
  (
    n173,
    n8
  );


  buf
  g13
  (
    n158,
    n21
  );


  not
  g14
  (
    n91,
    n43
  );


  buf
  g15
  (
    n131,
    n23
  );


  not
  g16
  (
    n179,
    n10
  );


  not
  g17
  (
    n209,
    n38
  );


  not
  g18
  (
    n64,
    n17
  );


  buf
  g19
  (
    n174,
    n38
  );


  not
  g20
  (
    n165,
    n37
  );


  buf
  g21
  (
    n115,
    n37
  );


  buf
  g22
  (
    n172,
    n3
  );


  not
  g23
  (
    n101,
    n18
  );


  not
  g24
  (
    n177,
    n35
  );


  not
  g25
  (
    n65,
    n36
  );


  not
  g26
  (
    n86,
    n32
  );


  buf
  g27
  (
    n75,
    n4
  );


  not
  g28
  (
    n153,
    n12
  );


  not
  g29
  (
    n159,
    n31
  );


  not
  g30
  (
    n168,
    n29
  );


  not
  g31
  (
    n183,
    n28
  );


  buf
  g32
  (
    n121,
    n3
  );


  not
  g33
  (
    n45,
    n42
  );


  not
  g34
  (
    n98,
    n34
  );


  buf
  g35
  (
    n74,
    n36
  );


  not
  g36
  (
    n175,
    n29
  );


  not
  g37
  (
    n178,
    n26
  );


  not
  g38
  (
    n215,
    n11
  );


  not
  g39
  (
    n184,
    n38
  );


  not
  g40
  (
    n196,
    n5
  );


  buf
  g41
  (
    n81,
    n21
  );


  not
  g42
  (
    n77,
    n25
  );


  buf
  g43
  (
    n66,
    n24
  );


  buf
  g44
  (
    n180,
    n3
  );


  buf
  g45
  (
    n154,
    n31
  );


  buf
  g46
  (
    n181,
    n22
  );


  not
  g47
  (
    n202,
    n15
  );


  buf
  g48
  (
    n161,
    n19
  );


  not
  g49
  (
    n141,
    n17
  );


  not
  g50
  (
    n132,
    n31
  );


  not
  g51
  (
    n104,
    n34
  );


  not
  g52
  (
    n166,
    n22
  );


  buf
  g53
  (
    n164,
    n32
  );


  not
  g54
  (
    n108,
    n12
  );


  buf
  g55
  (
    n56,
    n6
  );


  not
  g56
  (
    n146,
    n16
  );


  buf
  g57
  (
    n193,
    n42
  );


  buf
  g58
  (
    n95,
    n4
  );


  not
  g59
  (
    n201,
    n35
  );


  not
  g60
  (
    n208,
    n7
  );


  buf
  g61
  (
    n99,
    n18
  );


  not
  g62
  (
    n53,
    n23
  );


  not
  g63
  (
    n136,
    n26
  );


  not
  g64
  (
    n130,
    n23
  );


  not
  g65
  (
    n44,
    n17
  );


  buf
  g66
  (
    n70,
    n16
  );


  buf
  g67
  (
    n67,
    n36
  );


  not
  g68
  (
    n52,
    n25
  );


  buf
  g69
  (
    n90,
    n10
  );


  buf
  g70
  (
    n214,
    n15
  );


  not
  g71
  (
    n171,
    n43
  );


  buf
  g72
  (
    n155,
    n36
  );


  not
  g73
  (
    n138,
    n26
  );


  buf
  g74
  (
    n71,
    n5
  );


  buf
  g75
  (
    n169,
    n17
  );


  not
  g76
  (
    n89,
    n34
  );


  not
  g77
  (
    n113,
    n13
  );


  not
  g78
  (
    n129,
    n39
  );


  buf
  g79
  (
    n112,
    n25
  );


  not
  g80
  (
    n87,
    n32
  );


  not
  g81
  (
    n100,
    n40
  );


  not
  g82
  (
    n162,
    n30
  );


  buf
  g83
  (
    n189,
    n19
  );


  not
  g84
  (
    n49,
    n26
  );


  buf
  g85
  (
    n47,
    n6
  );


  buf
  g86
  (
    n139,
    n5
  );


  not
  g87
  (
    n106,
    n27
  );


  buf
  g88
  (
    n57,
    n38
  );


  not
  g89
  (
    n120,
    n3
  );


  not
  g90
  (
    n72,
    n27
  );


  buf
  g91
  (
    n96,
    n35
  );


  buf
  g92
  (
    n78,
    n13
  );


  buf
  g93
  (
    n134,
    n30
  );


  not
  g94
  (
    n182,
    n19
  );


  buf
  g95
  (
    n211,
    n29
  );


  buf
  g96
  (
    n195,
    n2
  );


  buf
  g97
  (
    n212,
    n29
  );


  buf
  g98
  (
    n163,
    n13
  );


  not
  g99
  (
    n167,
    n30
  );


  not
  g100
  (
    n188,
    n40
  );


  buf
  g101
  (
    n137,
    n13
  );


  not
  g102
  (
    n88,
    n1
  );


  buf
  g103
  (
    n107,
    n4
  );


  not
  g104
  (
    n83,
    n41
  );


  buf
  g105
  (
    n140,
    n10
  );


  buf
  g106
  (
    n60,
    n5
  );


  not
  g107
  (
    n144,
    n15
  );


  buf
  g108
  (
    n187,
    n21
  );


  buf
  g109
  (
    n82,
    n20
  );


  buf
  g110
  (
    n210,
    n8
  );


  not
  g111
  (
    n58,
    n37
  );


  buf
  g112
  (
    n205,
    n18
  );


  buf
  g113
  (
    n203,
    n30
  );


  not
  g114
  (
    n133,
    n37
  );


  buf
  g115
  (
    n143,
    n42
  );


  not
  g116
  (
    n152,
    n1
  );


  buf
  g117
  (
    n194,
    n18
  );


  not
  g118
  (
    n213,
    n42
  );


  buf
  g119
  (
    n63,
    n19
  );


  not
  g120
  (
    n157,
    n32
  );


  buf
  g121
  (
    n197,
    n43
  );


  not
  g122
  (
    n151,
    n22
  );


  buf
  g123
  (
    n128,
    n6
  );


  not
  g124
  (
    n46,
    n4
  );


  buf
  g125
  (
    n198,
    n2
  );


  not
  g126
  (
    KeyWire_0_12,
    n9
  );


  buf
  g127
  (
    n147,
    n33
  );


  buf
  g128
  (
    n84,
    n7
  );


  not
  g129
  (
    n116,
    n10
  );


  buf
  g130
  (
    n80,
    n9
  );


  not
  g131
  (
    n79,
    n28
  );


  not
  g132
  (
    n76,
    n14
  );


  not
  g133
  (
    n142,
    n11
  );


  not
  g134
  (
    n48,
    n31
  );


  buf
  g135
  (
    n103,
    n2
  );


  buf
  g136
  (
    n190,
    n24
  );


  buf
  g137
  (
    n145,
    n34
  );


  not
  g138
  (
    n117,
    n39
  );


  buf
  g139
  (
    n110,
    n9
  );


  buf
  g140
  (
    n186,
    n2
  );


  buf
  g141
  (
    n149,
    n6
  );


  not
  g142
  (
    n109,
    n41
  );


  not
  g143
  (
    n73,
    n8
  );


  not
  g144
  (
    n119,
    n8
  );


  buf
  g145
  (
    n206,
    n35
  );


  buf
  g146
  (
    KeyWire_0_29,
    n20
  );


  buf
  g147
  (
    n51,
    n14
  );


  not
  g148
  (
    n170,
    n39
  );


  not
  g149
  (
    n97,
    n16
  );


  not
  g150
  (
    n111,
    n15
  );


  buf
  g151
  (
    n127,
    n40
  );


  not
  g152
  (
    n114,
    n1
  );


  buf
  g153
  (
    n62,
    n11
  );


  not
  g154
  (
    n125,
    n28
  );


  not
  g155
  (
    n126,
    n33
  );


  buf
  g156
  (
    n102,
    n24
  );


  buf
  g157
  (
    n123,
    n33
  );


  not
  g158
  (
    n160,
    n20
  );


  not
  g159
  (
    n191,
    n41
  );


  buf
  g160
  (
    n185,
    n7
  );


  not
  g161
  (
    n204,
    n24
  );


  not
  g162
  (
    n105,
    n41
  );


  not
  g163
  (
    n118,
    n11
  );


  buf
  g164
  (
    n93,
    n40
  );


  buf
  g165
  (
    n135,
    n23
  );


  not
  g166
  (
    n124,
    n7
  );


  not
  g167
  (
    n94,
    n22
  );


  buf
  g168
  (
    n54,
    n28
  );


  buf
  g169
  (
    n59,
    n25
  );


  buf
  g170
  (
    n199,
    n39
  );


  buf
  g171
  (
    n192,
    n33
  );


  not
  g172
  (
    n564,
    n93
  );


  not
  g173
  (
    n645,
    n44
  );


  buf
  g174
  (
    n628,
    n183
  );


  buf
  g175
  (
    n722,
    n121
  );


  buf
  g176
  (
    n562,
    n98
  );


  not
  g177
  (
    KeyWire_0_9,
    n140
  );


  not
  g178
  (
    n570,
    n178
  );


  buf
  g179
  (
    n732,
    n58
  );


  buf
  g180
  (
    n430,
    n94
  );


  buf
  g181
  (
    n475,
    n183
  );


  not
  g182
  (
    n383,
    n52
  );


  not
  g183
  (
    n657,
    n92
  );


  buf
  g184
  (
    n452,
    n60
  );


  not
  g185
  (
    n282,
    n88
  );


  not
  g186
  (
    n523,
    n111
  );


  not
  g187
  (
    n574,
    n52
  );


  buf
  g188
  (
    n377,
    n124
  );


  buf
  g189
  (
    n420,
    n45
  );


  not
  g190
  (
    n539,
    n171
  );


  buf
  g191
  (
    n422,
    n191
  );


  buf
  g192
  (
    n476,
    n128
  );


  not
  g193
  (
    n274,
    n104
  );


  buf
  g194
  (
    n290,
    n141
  );


  not
  g195
  (
    n315,
    n165
  );


  not
  g196
  (
    n498,
    n143
  );


  not
  g197
  (
    n800,
    n120
  );


  buf
  g198
  (
    n543,
    n112
  );


  buf
  g199
  (
    n723,
    n180
  );


  buf
  g200
  (
    n260,
    n80
  );


  not
  g201
  (
    n292,
    n117
  );


  buf
  g202
  (
    n264,
    n71
  );


  not
  g203
  (
    n697,
    n98
  );


  buf
  g204
  (
    n537,
    n136
  );


  not
  g205
  (
    n644,
    n139
  );


  buf
  g206
  (
    n629,
    n57
  );


  buf
  g207
  (
    n656,
    n138
  );


  buf
  g208
  (
    n768,
    n131
  );


  not
  g209
  (
    n527,
    n89
  );


  not
  g210
  (
    n649,
    n81
  );


  not
  g211
  (
    n509,
    n67
  );


  buf
  g212
  (
    n558,
    n46
  );


  buf
  g213
  (
    n680,
    n176
  );


  buf
  g214
  (
    n789,
    n68
  );


  buf
  g215
  (
    n677,
    n180
  );


  buf
  g216
  (
    n682,
    n140
  );


  buf
  g217
  (
    n469,
    n185
  );


  buf
  g218
  (
    n388,
    n183
  );


  not
  g219
  (
    n251,
    n151
  );


  buf
  g220
  (
    n286,
    n76
  );


  buf
  g221
  (
    n707,
    n58
  );


  buf
  g222
  (
    n672,
    n99
  );


  buf
  g223
  (
    n709,
    n159
  );


  not
  g224
  (
    n615,
    n94
  );


  buf
  g225
  (
    n600,
    n68
  );


  buf
  g226
  (
    n437,
    n86
  );


  buf
  g227
  (
    n595,
    n65
  );


  buf
  g228
  (
    n363,
    n128
  );


  buf
  g229
  (
    n733,
    n170
  );


  not
  g230
  (
    n798,
    n163
  );


  not
  g231
  (
    n386,
    n140
  );


  buf
  g232
  (
    n725,
    n79
  );


  buf
  g233
  (
    n505,
    n59
  );


  not
  g234
  (
    n436,
    n102
  );


  buf
  g235
  (
    n354,
    n189
  );


  not
  g236
  (
    n227,
    n79
  );


  not
  g237
  (
    n427,
    n115
  );


  buf
  g238
  (
    n333,
    n125
  );


  not
  g239
  (
    n791,
    n150
  );


  buf
  g240
  (
    n216,
    n52
  );


  buf
  g241
  (
    n581,
    n87
  );


  not
  g242
  (
    n783,
    n77
  );


  not
  g243
  (
    n696,
    n172
  );


  not
  g244
  (
    n235,
    n59
  );


  buf
  g245
  (
    n765,
    n172
  );


  not
  g246
  (
    n337,
    n165
  );


  not
  g247
  (
    n488,
    n88
  );


  not
  g248
  (
    n610,
    n127
  );


  not
  g249
  (
    n357,
    n79
  );


  not
  g250
  (
    n511,
    n134
  );


  buf
  g251
  (
    n770,
    n147
  );


  not
  g252
  (
    n473,
    n61
  );


  not
  g253
  (
    n460,
    n62
  );


  not
  g254
  (
    n234,
    n175
  );


  not
  g255
  (
    n651,
    n51
  );


  not
  g256
  (
    n233,
    n56
  );


  buf
  g257
  (
    n730,
    n151
  );


  buf
  g258
  (
    n321,
    n106
  );


  buf
  g259
  (
    n409,
    n133
  );


  buf
  g260
  (
    n394,
    n60
  );


  buf
  g261
  (
    n326,
    n97
  );


  not
  g262
  (
    n503,
    n54
  );


  buf
  g263
  (
    n506,
    n176
  );


  not
  g264
  (
    n501,
    n103
  );


  buf
  g265
  (
    n494,
    n168
  );


  not
  g266
  (
    n784,
    n85
  );


  not
  g267
  (
    n777,
    n89
  );


  not
  g268
  (
    n246,
    n86
  );


  buf
  g269
  (
    n398,
    n100
  );


  not
  g270
  (
    n761,
    n144
  );


  buf
  g271
  (
    n555,
    n125
  );


  not
  g272
  (
    n492,
    n68
  );


  buf
  g273
  (
    n793,
    n65
  );


  not
  g274
  (
    n332,
    n148
  );


  buf
  g275
  (
    n642,
    n186
  );


  not
  g276
  (
    n706,
    n133
  );


  buf
  g277
  (
    n454,
    n99
  );


  not
  g278
  (
    n284,
    n48
  );


  buf
  g279
  (
    n466,
    n95
  );


  buf
  g280
  (
    n384,
    n106
  );


  not
  g281
  (
    n755,
    n77
  );


  buf
  g282
  (
    n392,
    n138
  );


  not
  g283
  (
    n297,
    n175
  );


  buf
  g284
  (
    n464,
    n152
  );


  buf
  g285
  (
    n450,
    n161
  );


  buf
  g286
  (
    n218,
    n167
  );


  buf
  g287
  (
    n459,
    n140
  );


  not
  g288
  (
    n263,
    n49
  );


  not
  g289
  (
    n510,
    n95
  );


  not
  g290
  (
    n481,
    n137
  );


  buf
  g291
  (
    n228,
    n130
  );


  buf
  g292
  (
    n620,
    n170
  );


  buf
  g293
  (
    n325,
    n74
  );


  buf
  g294
  (
    n425,
    n85
  );


  not
  g295
  (
    n419,
    n72
  );


  buf
  g296
  (
    n355,
    n111
  );


  buf
  g297
  (
    n257,
    n78
  );


  not
  g298
  (
    n391,
    n81
  );


  buf
  g299
  (
    n385,
    n110
  );


  not
  g300
  (
    n666,
    n164
  );


  not
  g301
  (
    n772,
    n119
  );


  not
  g302
  (
    n801,
    n108
  );


  buf
  g303
  (
    n623,
    n136
  );


  buf
  g304
  (
    n300,
    n172
  );


  buf
  g305
  (
    n229,
    n155
  );


  buf
  g306
  (
    n463,
    n124
  );


  not
  g307
  (
    n631,
    n159
  );


  not
  g308
  (
    n368,
    n71
  );


  buf
  g309
  (
    n625,
    n186
  );


  not
  g310
  (
    n547,
    n56
  );


  not
  g311
  (
    n411,
    n188
  );


  buf
  g312
  (
    n708,
    n80
  );


  not
  g313
  (
    n445,
    n107
  );


  not
  g314
  (
    n240,
    n120
  );


  buf
  g315
  (
    n710,
    n181
  );


  buf
  g316
  (
    n626,
    n103
  );


  not
  g317
  (
    n739,
    n178
  );


  not
  g318
  (
    n804,
    n75
  );


  not
  g319
  (
    n529,
    n181
  );


  not
  g320
  (
    n599,
    n167
  );


  not
  g321
  (
    n609,
    n69
  );


  buf
  g322
  (
    n467,
    n164
  );


  buf
  g323
  (
    n557,
    n174
  );


  buf
  g324
  (
    n270,
    n84
  );


  not
  g325
  (
    n489,
    n46
  );


  not
  g326
  (
    n277,
    n122
  );


  not
  g327
  (
    n359,
    n139
  );


  buf
  g328
  (
    n681,
    n82
  );


  not
  g329
  (
    n622,
    n46
  );


  not
  g330
  (
    n731,
    n84
  );


  not
  g331
  (
    n340,
    n184
  );


  buf
  g332
  (
    n688,
    n103
  );


  not
  g333
  (
    n532,
    n185
  );


  not
  g334
  (
    n780,
    n89
  );


  buf
  g335
  (
    n456,
    n135
  );


  buf
  g336
  (
    n571,
    n84
  );


  not
  g337
  (
    n592,
    n166
  );


  buf
  g338
  (
    n561,
    n150
  );


  buf
  g339
  (
    n639,
    n57
  );


  buf
  g340
  (
    n429,
    n166
  );


  not
  g341
  (
    n724,
    n49
  );


  buf
  g342
  (
    n735,
    n139
  );


  buf
  g343
  (
    n718,
    n143
  );


  not
  g344
  (
    n573,
    n118
  );


  not
  g345
  (
    n245,
    n147
  );


  buf
  g346
  (
    n338,
    n71
  );


  not
  g347
  (
    n309,
    n53
  );


  buf
  g348
  (
    n775,
    n122
  );


  buf
  g349
  (
    n444,
    n109
  );


  buf
  g350
  (
    n787,
    n108
  );


  not
  g351
  (
    n641,
    n72
  );


  not
  g352
  (
    n367,
    n181
  );


  buf
  g353
  (
    n758,
    n51
  );


  buf
  g354
  (
    n546,
    n118
  );


  buf
  g355
  (
    n273,
    n102
  );


  not
  g356
  (
    n378,
    n121
  );


  not
  g357
  (
    n410,
    n152
  );


  not
  g358
  (
    n514,
    n83
  );


  buf
  g359
  (
    n586,
    n159
  );


  not
  g360
  (
    n749,
    n178
  );


  not
  g361
  (
    n345,
    n154
  );


  buf
  g362
  (
    n285,
    n66
  );


  buf
  g363
  (
    n685,
    n92
  );


  not
  g364
  (
    n675,
    n114
  );


  buf
  g365
  (
    n742,
    n113
  );


  buf
  g366
  (
    n379,
    n188
  );


  buf
  g367
  (
    n462,
    n144
  );


  buf
  g368
  (
    n364,
    n129
  );


  not
  g369
  (
    n289,
    n150
  );


  buf
  g370
  (
    n699,
    n174
  );


  not
  g371
  (
    KeyWire_0_0,
    n70
  );


  buf
  g372
  (
    n671,
    n185
  );


  not
  g373
  (
    n711,
    n66
  );


  buf
  g374
  (
    n375,
    n183
  );


  buf
  g375
  (
    n556,
    n57
  );


  not
  g376
  (
    n582,
    n64
  );


  not
  g377
  (
    n438,
    n48
  );


  buf
  g378
  (
    n305,
    n127
  );


  buf
  g379
  (
    n576,
    n190
  );


  not
  g380
  (
    n605,
    n117
  );


  buf
  g381
  (
    n371,
    n149
  );


  buf
  g382
  (
    n404,
    n133
  );


  buf
  g383
  (
    n797,
    n155
  );


  buf
  g384
  (
    n588,
    n130
  );


  buf
  g385
  (
    n295,
    n44
  );


  buf
  g386
  (
    n266,
    n119
  );


  not
  g387
  (
    n608,
    n131
  );


  buf
  g388
  (
    n312,
    n105
  );


  not
  g389
  (
    n241,
    n182
  );


  not
  g390
  (
    n343,
    n61
  );


  not
  g391
  (
    n676,
    n67
  );


  not
  g392
  (
    n540,
    n109
  );


  not
  g393
  (
    n773,
    n106
  );


  buf
  g394
  (
    n579,
    n142
  );


  buf
  g395
  (
    n254,
    n46
  );


  buf
  g396
  (
    n705,
    n117
  );


  not
  g397
  (
    n655,
    n62
  );


  not
  g398
  (
    n316,
    n179
  );


  buf
  g399
  (
    n238,
    n135
  );


  buf
  g400
  (
    n413,
    n120
  );


  buf
  g401
  (
    n549,
    n113
  );


  not
  g402
  (
    n474,
    n184
  );


  not
  g403
  (
    n796,
    n123
  );


  buf
  g404
  (
    n778,
    n190
  );


  not
  g405
  (
    n399,
    n142
  );


  not
  g406
  (
    n261,
    n105
  );


  buf
  g407
  (
    n390,
    n133
  );


  not
  g408
  (
    n740,
    n76
  );


  buf
  g409
  (
    n689,
    n49
  );


  buf
  g410
  (
    n446,
    n65
  );


  not
  g411
  (
    n434,
    n188
  );


  buf
  g412
  (
    n304,
    n147
  );


  buf
  g413
  (
    n575,
    n177
  );


  buf
  g414
  (
    n374,
    n88
  );


  buf
  g415
  (
    n403,
    n155
  );


  not
  g416
  (
    n243,
    n171
  );


  not
  g417
  (
    n360,
    n127
  );


  not
  g418
  (
    n560,
    n89
  );


  not
  g419
  (
    n314,
    n169
  );


  buf
  g420
  (
    n439,
    n153
  );


  not
  g421
  (
    n667,
    n113
  );


  not
  g422
  (
    n351,
    n63
  );


  not
  g423
  (
    n678,
    n61
  );


  buf
  g424
  (
    n334,
    n67
  );


  buf
  g425
  (
    n415,
    n173
  );


  buf
  g426
  (
    n294,
    n101
  );


  buf
  g427
  (
    n530,
    n97
  );


  not
  g428
  (
    n265,
    n78
  );


  not
  g429
  (
    n665,
    n132
  );


  buf
  g430
  (
    n774,
    n130
  );


  not
  g431
  (
    n376,
    n173
  );


  not
  g432
  (
    n550,
    n143
  );


  buf
  g433
  (
    n652,
    n53
  );


  buf
  g434
  (
    n366,
    n107
  );


  not
  g435
  (
    n504,
    n78
  );


  buf
  g436
  (
    n479,
    n91
  );


  not
  g437
  (
    n759,
    n99
  );


  not
  g438
  (
    n442,
    n169
  );


  not
  g439
  (
    n482,
    n102
  );


  not
  g440
  (
    n353,
    n153
  );


  buf
  g441
  (
    n616,
    n98
  );


  buf
  g442
  (
    n643,
    n132
  );


  not
  g443
  (
    n692,
    n50
  );


  not
  g444
  (
    n647,
    n85
  );


  buf
  g445
  (
    n451,
    n168
  );


  not
  g446
  (
    n660,
    n47
  );


  buf
  g447
  (
    n283,
    n64
  );


  not
  g448
  (
    n223,
    n131
  );


  not
  g449
  (
    n598,
    n170
  );


  not
  g450
  (
    n350,
    n104
  );


  buf
  g451
  (
    n544,
    n55
  );


  buf
  g452
  (
    n328,
    n151
  );


  buf
  g453
  (
    n373,
    n145
  );


  not
  g454
  (
    n719,
    n107
  );


  not
  g455
  (
    n342,
    n128
  );


  not
  g456
  (
    n458,
    n136
  );


  not
  g457
  (
    n322,
    n154
  );


  buf
  g458
  (
    n568,
    n175
  );


  not
  g459
  (
    n636,
    n157
  );


  not
  g460
  (
    n317,
    n85
  );


  buf
  g461
  (
    n247,
    n71
  );


  buf
  g462
  (
    n585,
    n144
  );


  not
  g463
  (
    n589,
    n189
  );


  not
  g464
  (
    n301,
    n184
  );


  not
  g465
  (
    n307,
    n97
  );


  not
  g466
  (
    n745,
    n167
  );


  buf
  g467
  (
    n221,
    n148
  );


  buf
  g468
  (
    n237,
    n110
  );


  not
  g469
  (
    n776,
    n163
  );


  not
  g470
  (
    n365,
    n75
  );


  buf
  g471
  (
    n669,
    n49
  );


  buf
  g472
  (
    n471,
    n142
  );


  not
  g473
  (
    n470,
    n81
  );


  not
  g474
  (
    n278,
    n166
  );


  buf
  g475
  (
    n408,
    n158
  );


  not
  g476
  (
    n418,
    n119
  );


  not
  g477
  (
    n248,
    n99
  );


  buf
  g478
  (
    n306,
    n79
  );


  not
  g479
  (
    n617,
    n65
  );


  not
  g480
  (
    n635,
    n156
  );


  buf
  g481
  (
    n563,
    n76
  );


  buf
  g482
  (
    n449,
    n90
  );


  buf
  g483
  (
    n344,
    n100
  );


  not
  g484
  (
    n741,
    n63
  );


  not
  g485
  (
    n769,
    n182
  );


  not
  g486
  (
    n412,
    n104
  );


  buf
  g487
  (
    n472,
    n147
  );


  not
  g488
  (
    n684,
    n44
  );


  buf
  g489
  (
    n662,
    n149
  );


  buf
  g490
  (
    n794,
    n162
  );


  not
  g491
  (
    n299,
    n167
  );


  not
  g492
  (
    n703,
    n59
  );


  not
  g493
  (
    n728,
    n64
  );


  buf
  g494
  (
    n502,
    n186
  );


  not
  g495
  (
    n424,
    n62
  );


  buf
  g496
  (
    n737,
    n48
  );


  not
  g497
  (
    n490,
    n141
  );


  not
  g498
  (
    n551,
    n108
  );


  not
  g499
  (
    n650,
    n60
  );


  not
  g500
  (
    n358,
    n105
  );


  buf
  g501
  (
    n634,
    n117
  );


  not
  g502
  (
    n593,
    n158
  );


  buf
  g503
  (
    n583,
    n177
  );


  not
  g504
  (
    n538,
    n76
  );


  not
  g505
  (
    n487,
    n135
  );


  buf
  g506
  (
    n714,
    n95
  );


  buf
  g507
  (
    n242,
    n154
  );


  buf
  g508
  (
    n762,
    n96
  );


  not
  g509
  (
    n552,
    n63
  );


  not
  g510
  (
    n381,
    n52
  );


  buf
  g511
  (
    n621,
    n134
  );


  buf
  g512
  (
    n781,
    n158
  );


  not
  g513
  (
    n754,
    n51
  );


  buf
  g514
  (
    n432,
    n68
  );


  buf
  g515
  (
    n441,
    n122
  );


  buf
  g516
  (
    n632,
    n105
  );


  buf
  g517
  (
    n674,
    n157
  );


  not
  g518
  (
    n319,
    n174
  );


  buf
  g519
  (
    n361,
    n112
  );


  not
  g520
  (
    n303,
    n69
  );


  buf
  g521
  (
    n799,
    n115
  );


  not
  g522
  (
    n395,
    n84
  );


  not
  g523
  (
    n496,
    n149
  );


  not
  g524
  (
    KeyWire_0_10,
    n131
  );


  not
  g525
  (
    n533,
    n78
  );


  buf
  g526
  (
    n746,
    n50
  );


  not
  g527
  (
    n790,
    n107
  );


  not
  g528
  (
    n569,
    n169
  );


  not
  g529
  (
    n726,
    n80
  );


  buf
  g530
  (
    n406,
    n135
  );


  not
  g531
  (
    n694,
    n179
  );


  buf
  g532
  (
    n785,
    n181
  );


  not
  g533
  (
    n486,
    n86
  );


  buf
  g534
  (
    n517,
    n134
  );


  buf
  g535
  (
    n603,
    n111
  );


  not
  g536
  (
    n795,
    n64
  );


  not
  g537
  (
    KeyWire_0_13,
    n161
  );


  buf
  g538
  (
    n638,
    n73
  );


  not
  g539
  (
    n528,
    n100
  );


  not
  g540
  (
    n602,
    n115
  );


  not
  g541
  (
    n701,
    n90
  );


  not
  g542
  (
    n302,
    n96
  );


  buf
  g543
  (
    n276,
    n165
  );


  not
  g544
  (
    n461,
    n116
  );


  not
  g545
  (
    n686,
    n90
  );


  not
  g546
  (
    n330,
    n55
  );


  buf
  g547
  (
    n531,
    n168
  );


  not
  g548
  (
    n271,
    n56
  );


  buf
  g549
  (
    n516,
    n58
  );


  not
  g550
  (
    n594,
    n153
  );


  buf
  g551
  (
    n545,
    n57
  );


  not
  g552
  (
    n515,
    n136
  );


  not
  g553
  (
    n423,
    n123
  );


  buf
  g554
  (
    n715,
    n69
  );


  buf
  g555
  (
    n447,
    n162
  );


  not
  g556
  (
    n559,
    n53
  );


  not
  g557
  (
    n567,
    n158
  );


  buf
  g558
  (
    n499,
    n125
  );


  not
  g559
  (
    n262,
    n72
  );


  not
  g560
  (
    n465,
    n118
  );


  buf
  g561
  (
    n673,
    n110
  );


  not
  g562
  (
    n750,
    n153
  );


  buf
  g563
  (
    n249,
    n114
  );


  not
  g564
  (
    n721,
    n60
  );


  buf
  g565
  (
    n329,
    n104
  );


  not
  g566
  (
    n226,
    n91
  );


  not
  g567
  (
    n663,
    n70
  );


  buf
  g568
  (
    n766,
    n54
  );


  not
  g569
  (
    n803,
    n182
  );


  not
  g570
  (
    n572,
    n83
  );


  buf
  g571
  (
    n782,
    n83
  );


  buf
  g572
  (
    n607,
    n191
  );


  not
  g573
  (
    n630,
    n82
  );


  not
  g574
  (
    n346,
    n74
  );


  buf
  g575
  (
    n281,
    n176
  );


  buf
  g576
  (
    n727,
    n91
  );


  not
  g577
  (
    n440,
    n165
  );


  not
  g578
  (
    n653,
    n175
  );


  not
  g579
  (
    KeyWire_0_5,
    n114
  );


  buf
  g580
  (
    n397,
    n123
  );


  buf
  g581
  (
    n318,
    n127
  );


  buf
  g582
  (
    n339,
    n54
  );


  buf
  g583
  (
    n507,
    n145
  );


  buf
  g584
  (
    n779,
    n161
  );


  buf
  g585
  (
    n231,
    n148
  );


  not
  g586
  (
    n275,
    n144
  );


  not
  g587
  (
    n613,
    n55
  );


  not
  g588
  (
    n253,
    n96
  );


  not
  g589
  (
    n584,
    n186
  );


  buf
  g590
  (
    n313,
    n61
  );


  not
  g591
  (
    n405,
    n159
  );


  not
  g592
  (
    n443,
    n122
  );


  not
  g593
  (
    n747,
    n116
  );


  not
  g594
  (
    n614,
    n151
  );


  not
  g595
  (
    n646,
    n53
  );


  not
  g596
  (
    n704,
    n95
  );


  buf
  g597
  (
    n580,
    n96
  );


  not
  g598
  (
    n788,
    n173
  );


  buf
  g599
  (
    n396,
    n113
  );


  not
  g600
  (
    n590,
    n58
  );


  buf
  g601
  (
    n512,
    n87
  );


  buf
  g602
  (
    n348,
    n155
  );


  not
  g603
  (
    n744,
    n62
  );


  not
  g604
  (
    n256,
    n73
  );


  buf
  g605
  (
    n659,
    n121
  );


  buf
  g606
  (
    n389,
    n87
  );


  not
  g607
  (
    n335,
    n81
  );


  buf
  g608
  (
    n734,
    n141
  );


  not
  g609
  (
    n690,
    n44
  );


  not
  g610
  (
    n280,
    n82
  );


  not
  g611
  (
    n751,
    n174
  );


  buf
  g612
  (
    n414,
    n123
  );


  buf
  g613
  (
    n393,
    n119
  );


  buf
  g614
  (
    n597,
    n189
  );


  not
  g615
  (
    n491,
    n160
  );


  not
  g616
  (
    n520,
    n112
  );


  buf
  g617
  (
    n288,
    n187
  );


  buf
  g618
  (
    n500,
    n103
  );


  buf
  g619
  (
    n258,
    n74
  );


  buf
  g620
  (
    n485,
    n48
  );


  not
  g621
  (
    n700,
    n66
  );


  buf
  g622
  (
    n272,
    n156
  );


  buf
  g623
  (
    n455,
    n161
  );


  not
  g624
  (
    n480,
    n149
  );


  buf
  g625
  (
    n596,
    n55
  );


  buf
  g626
  (
    n372,
    n125
  );


  not
  g627
  (
    n627,
    n187
  );


  not
  g628
  (
    n287,
    n185
  );


  not
  g629
  (
    n542,
    n137
  );


  buf
  g630
  (
    n591,
    n73
  );


  not
  g631
  (
    n417,
    n137
  );


  buf
  g632
  (
    n767,
    n114
  );


  buf
  g633
  (
    n323,
    n146
  );


  not
  g634
  (
    n347,
    n142
  );


  not
  g635
  (
    n637,
    n180
  );


  not
  g636
  (
    n757,
    n180
  );


  buf
  g637
  (
    n535,
    n145
  );


  not
  g638
  (
    n521,
    n93
  );


  not
  g639
  (
    n513,
    n98
  );


  not
  g640
  (
    n401,
    n101
  );


  buf
  g641
  (
    n421,
    n152
  );


  not
  g642
  (
    n756,
    n132
  );


  buf
  g643
  (
    n668,
    n56
  );


  not
  g644
  (
    n407,
    n130
  );


  not
  g645
  (
    n341,
    n102
  );


  buf
  g646
  (
    n268,
    n77
  );


  buf
  g647
  (
    n250,
    n152
  );


  buf
  g648
  (
    n457,
    n187
  );


  not
  g649
  (
    n518,
    n129
  );


  buf
  g650
  (
    n664,
    n116
  );


  buf
  g651
  (
    n717,
    n50
  );


  buf
  g652
  (
    n748,
    n154
  );


  buf
  g653
  (
    n493,
    n164
  );


  buf
  g654
  (
    KeyWire_0_24,
    n83
  );


  not
  g655
  (
    n416,
    n92
  );


  buf
  g656
  (
    n519,
    n184
  );


  not
  g657
  (
    n640,
    n118
  );


  buf
  g658
  (
    n661,
    n124
  );


  not
  g659
  (
    n606,
    n94
  );


  not
  g660
  (
    n698,
    n166
  );


  buf
  g661
  (
    n648,
    n72
  );


  buf
  g662
  (
    n217,
    n190
  );


  buf
  g663
  (
    n525,
    n91
  );


  not
  g664
  (
    n320,
    n182
  );


  not
  g665
  (
    n548,
    n63
  );


  not
  g666
  (
    n554,
    n176
  );


  not
  g667
  (
    n716,
    n138
  );


  not
  g668
  (
    n729,
    n126
  );


  buf
  g669
  (
    n497,
    n47
  );


  not
  g670
  (
    n693,
    n129
  );


  not
  g671
  (
    n453,
    n162
  );


  buf
  g672
  (
    n658,
    n111
  );


  not
  g673
  (
    n370,
    n164
  );


  not
  g674
  (
    n578,
    n146
  );


  not
  g675
  (
    n468,
    n101
  );


  buf
  g676
  (
    n771,
    n110
  );


  buf
  g677
  (
    n536,
    n146
  );


  buf
  g678
  (
    n524,
    n82
  );


  buf
  g679
  (
    n601,
    n112
  );


  buf
  g680
  (
    n232,
    n177
  );


  buf
  g681
  (
    n448,
    n157
  );


  not
  g682
  (
    n380,
    n157
  );


  not
  g683
  (
    n477,
    n45
  );


  not
  g684
  (
    n611,
    n187
  );


  buf
  g685
  (
    n433,
    n88
  );


  not
  g686
  (
    n764,
    n179
  );


  buf
  g687
  (
    n269,
    n75
  );


  not
  g688
  (
    n670,
    n59
  );


  buf
  g689
  (
    n352,
    n134
  );


  buf
  g690
  (
    n220,
    n139
  );


  buf
  g691
  (
    n713,
    n108
  );


  not
  g692
  (
    n565,
    n45
  );


  buf
  g693
  (
    n291,
    n50
  );


  buf
  g694
  (
    n349,
    n124
  );


  buf
  g695
  (
    n296,
    n87
  );


  not
  g696
  (
    n239,
    n177
  );


  not
  g697
  (
    n387,
    n148
  );


  not
  g698
  (
    n541,
    n126
  );


  not
  g699
  (
    n743,
    n70
  );


  buf
  g700
  (
    n752,
    n132
  );


  buf
  g701
  (
    n526,
    n109
  );


  not
  g702
  (
    n508,
    n170
  );


  not
  g703
  (
    KeyWire_0_11,
    n80
  );


  buf
  g704
  (
    n219,
    n120
  );


  not
  g705
  (
    n426,
    n160
  );


  not
  g706
  (
    n428,
    n66
  );


  not
  g707
  (
    n702,
    n138
  );


  not
  g708
  (
    n252,
    n109
  );


  not
  g709
  (
    n738,
    n163
  );


  not
  g710
  (
    n435,
    n137
  );


  not
  g711
  (
    n566,
    n106
  );


  not
  g712
  (
    n222,
    n75
  );


  buf
  g713
  (
    n587,
    n129
  );


  not
  g714
  (
    n331,
    n145
  );


  buf
  g715
  (
    n604,
    n169
  );


  buf
  g716
  (
    n478,
    n77
  );


  not
  g717
  (
    n267,
    n121
  );


  not
  g718
  (
    n753,
    n73
  );


  not
  g719
  (
    n230,
    n90
  );


  buf
  g720
  (
    n687,
    n92
  );


  not
  g721
  (
    n244,
    n93
  );


  not
  g722
  (
    KeyWire_0_1,
    n128
  );


  not
  g723
  (
    n298,
    n191
  );


  buf
  g724
  (
    n760,
    n156
  );


  not
  g725
  (
    n633,
    n162
  );


  not
  g726
  (
    n695,
    n100
  );


  buf
  g727
  (
    n720,
    n94
  );


  not
  g728
  (
    n400,
    n67
  );


  buf
  g729
  (
    n308,
    n160
  );


  buf
  g730
  (
    n618,
    n178
  );


  not
  g731
  (
    n327,
    n97
  );


  not
  g732
  (
    n522,
    n69
  );


  not
  g733
  (
    n553,
    n54
  );


  buf
  g734
  (
    n362,
    n45
  );


  not
  g735
  (
    n369,
    n179
  );


  not
  g736
  (
    n483,
    n143
  );


  not
  g737
  (
    n683,
    n70
  );


  not
  g738
  (
    n679,
    n189
  );


  not
  g739
  (
    n259,
    n86
  );


  buf
  g740
  (
    n293,
    n116
  );


  not
  g741
  (
    n792,
    n141
  );


  not
  g742
  (
    n495,
    n160
  );


  not
  g743
  (
    n763,
    n101
  );


  not
  g744
  (
    n236,
    n93
  );


  buf
  g745
  (
    n311,
    n168
  );


  buf
  g746
  (
    n431,
    n115
  );


  not
  g747
  (
    n534,
    n163
  );


  buf
  g748
  (
    n736,
    n126
  );


  not
  g749
  (
    n255,
    n126
  );


  buf
  g750
  (
    n279,
    n47
  );


  not
  g751
  (
    n612,
    n171
  );


  buf
  g752
  (
    n402,
    n51
  );


  buf
  g753
  (
    n484,
    n173
  );


  buf
  g754
  (
    n712,
    n47
  );


  buf
  g755
  (
    n577,
    n172
  );


  not
  g756
  (
    n324,
    n190
  );


  not
  g757
  (
    n619,
    n74
  );


  not
  g758
  (
    n336,
    n171
  );


  nor
  g759
  (
    n224,
    n150,
    n188
  );


  and
  g760
  (
    n624,
    n146,
    n156
  );


  buf
  g761
  (
    n806,
    n216
  );


  not
  g762
  (
    n805,
    n216
  );


  xor
  g763
  (
    n807,
    n805,
    n216,
    n217
  );


  not
  g764
  (
    n809,
    n807
  );


  buf
  g765
  (
    n808,
    n807
  );


  buf
  g766
  (
    n811,
    n191
  );


  nor
  g767
  (
    n810,
    n192,
    n808
  );


  and
  g768
  (
    n813,
    n811,
    n222,
    n217,
    n218
  );


  and
  g769
  (
    n814,
    n222,
    n218,
    n219,
    n220
  );


  nand
  g770
  (
    n818,
    n221,
    n810,
    n811
  );


  xnor
  g771
  (
    n812,
    n221,
    n811,
    n217,
    n220
  );


  and
  g772
  (
    n816,
    n219,
    n218,
    n221
  );


  xor
  g773
  (
    n815,
    n220,
    n221,
    n217,
    n810
  );


  and
  g774
  (
    n817,
    n810,
    n219,
    n220
  );


  buf
  g775
  (
    KeyWire_0_16,
    n224
  );


  not
  g776
  (
    n838,
    n223
  );


  not
  g777
  (
    n830,
    n813
  );


  buf
  g778
  (
    n824,
    n806
  );


  not
  g779
  (
    n823,
    n222
  );


  not
  g780
  (
    n831,
    n816
  );


  not
  g781
  (
    n835,
    n224
  );


  not
  g782
  (
    n827,
    n223
  );


  not
  g783
  (
    n825,
    n813
  );


  not
  g784
  (
    n821,
    n816
  );


  buf
  g785
  (
    n828,
    n812
  );


  buf
  g786
  (
    n820,
    n223
  );


  not
  g787
  (
    n833,
    n814
  );


  buf
  g788
  (
    n832,
    n815
  );


  buf
  g789
  (
    n822,
    n814
  );


  buf
  g790
  (
    n837,
    n224
  );


  nor
  g791
  (
    n836,
    n222,
    n813,
    n814,
    n815
  );


  xnor
  g792
  (
    n834,
    n813,
    n812,
    n815,
    n223
  );


  and
  g793
  (
    n819,
    n815,
    n811,
    n817,
    n814
  );


  or
  g794
  (
    n826,
    n224,
    n817,
    n816
  );


  buf
  g795
  (
    n857,
    n828
  );


  buf
  g796
  (
    n848,
    n819
  );


  buf
  g797
  (
    n872,
    n822
  );


  buf
  g798
  (
    n851,
    n194
  );


  not
  g799
  (
    n871,
    n807
  );


  buf
  g800
  (
    n870,
    n836
  );


  not
  g801
  (
    n840,
    n831
  );


  not
  g802
  (
    n867,
    n820
  );


  buf
  g803
  (
    n849,
    n193
  );


  buf
  g804
  (
    n842,
    n835
  );


  nand
  g805
  (
    n861,
    n830,
    n819,
    n808,
    n837
  );


  xnor
  g806
  (
    n852,
    n820,
    n837,
    n824,
    n807
  );


  xnor
  g807
  (
    n850,
    n837,
    n826,
    n194,
    n817
  );


  nand
  g808
  (
    n859,
    n818,
    n809,
    n832,
    n836
  );


  nand
  g809
  (
    n847,
    n832,
    n827,
    n833,
    n820
  );


  xor
  g810
  (
    n864,
    n809,
    n821,
    n808,
    n834
  );


  xor
  g811
  (
    n853,
    n834,
    n194,
    n826,
    n827
  );


  xnor
  g812
  (
    n865,
    n192,
    n820,
    n831,
    n830
  );


  xnor
  g813
  (
    n839,
    n821,
    n838,
    n825,
    n193
  );


  nand
  g814
  (
    n854,
    n833,
    n828,
    n809,
    n838
  );


  nand
  g815
  (
    n868,
    n836,
    n837,
    n195,
    n832
  );


  xnor
  g816
  (
    n869,
    n826,
    n830,
    n822,
    n828
  );


  and
  g817
  (
    n846,
    n833,
    n836,
    n824,
    n195
  );


  nor
  g818
  (
    n866,
    n194,
    n834,
    n823,
    n829
  );


  nor
  g819
  (
    n860,
    n821,
    n826,
    n827,
    n838
  );


  nand
  g820
  (
    n862,
    n817,
    n831,
    n823,
    n825
  );


  xnor
  g821
  (
    n856,
    n822,
    n818,
    n819,
    n831
  );


  or
  g822
  (
    n855,
    n809,
    n829,
    n823
  );


  nand
  g823
  (
    n863,
    n193,
    n825,
    n824,
    n821
  );


  xnor
  g824
  (
    n844,
    n823,
    n830,
    n828,
    n833
  );


  xnor
  g825
  (
    n841,
    n829,
    n827,
    n192,
    n835
  );


  or
  g826
  (
    n843,
    n825,
    n822,
    n193,
    n834
  );


  and
  g827
  (
    n858,
    n838,
    n819,
    n832,
    n818
  );


  nor
  g828
  (
    n845,
    n818,
    n835,
    n824
  );


  not
  g829
  (
    n874,
    n840
  );


  buf
  g830
  (
    n876,
    n842
  );


  not
  g831
  (
    n873,
    n841
  );


  buf
  g832
  (
    n875,
    n839
  );


  not
  g833
  (
    n883,
    n873
  );


  not
  g834
  (
    n878,
    n861
  );


  buf
  g835
  (
    n892,
    n875
  );


  not
  g836
  (
    n882,
    n843
  );


  not
  g837
  (
    n885,
    n844
  );


  buf
  g838
  (
    n887,
    n874
  );


  buf
  g839
  (
    n890,
    n875
  );


  buf
  g840
  (
    n877,
    n851
  );


  xnor
  g841
  (
    n880,
    n874,
    n853,
    n875,
    n847
  );


  xnor
  g842
  (
    n889,
    n874,
    n876,
    n845
  );


  or
  g843
  (
    n888,
    n859,
    n860,
    n858,
    n856
  );


  or
  g844
  (
    n884,
    n860,
    n848,
    n857,
    n861
  );


  or
  g845
  (
    n891,
    n873,
    n873,
    n874,
    n854
  );


  or
  g846
  (
    n879,
    n860,
    n875,
    n876,
    n861
  );


  xnor
  g847
  (
    n886,
    n876,
    n850,
    n846,
    n873
  );


  or
  g848
  (
    n881,
    n849,
    n860,
    n855,
    n852
  );


  not
  g849
  (
    n923,
    n877
  );


  not
  g850
  (
    n908,
    n883
  );


  not
  g851
  (
    n917,
    n881
  );


  not
  g852
  (
    n901,
    n877
  );


  not
  g853
  (
    n912,
    n878
  );


  not
  g854
  (
    n899,
    n880
  );


  buf
  g855
  (
    n911,
    n878
  );


  not
  g856
  (
    n906,
    n879
  );


  not
  g857
  (
    n902,
    n878
  );


  not
  g858
  (
    n913,
    n879
  );


  not
  g859
  (
    n894,
    n879
  );


  not
  g860
  (
    n905,
    n882
  );


  buf
  g861
  (
    n903,
    n883
  );


  buf
  g862
  (
    n904,
    n878
  );


  not
  g863
  (
    n919,
    n884
  );


  buf
  g864
  (
    n907,
    n883
  );


  buf
  g865
  (
    n922,
    n882
  );


  not
  g866
  (
    n916,
    n884
  );


  buf
  g867
  (
    n915,
    n881
  );


  buf
  g868
  (
    n895,
    n882
  );


  not
  g869
  (
    n920,
    n884
  );


  buf
  g870
  (
    n909,
    n877
  );


  not
  g871
  (
    n898,
    n881
  );


  buf
  g872
  (
    n896,
    n880
  );


  buf
  g873
  (
    n893,
    n880
  );


  buf
  g874
  (
    n918,
    n883
  );


  buf
  g875
  (
    n924,
    n882
  );


  not
  g876
  (
    n914,
    n877
  );


  buf
  g877
  (
    n900,
    n879
  );


  buf
  g878
  (
    n910,
    n884
  );


  not
  g879
  (
    n921,
    n880
  );


  buf
  g880
  (
    n897,
    n881
  );


  not
  g881
  (
    n928,
    n893
  );


  not
  g882
  (
    n929,
    n894
  );


  buf
  g883
  (
    n925,
    n893
  );


  buf
  g884
  (
    n927,
    n885
  );


  xnor
  g885
  (
    n926,
    n885,
    n893
  );


  buf
  g886
  (
    n931,
    n925
  );


  not
  g887
  (
    n930,
    n925
  );


  not
  g888
  (
    n932,
    n925
  );


  not
  g889
  (
    n941,
    n926
  );


  buf
  g890
  (
    n940,
    n931
  );


  not
  g891
  (
    n939,
    n932
  );


  not
  g892
  (
    n938,
    n925
  );


  not
  g893
  (
    n933,
    n931
  );


  not
  g894
  (
    n936,
    n926
  );


  nand
  g895
  (
    n935,
    n932,
    n926,
    n927
  );


  nor
  g896
  (
    n934,
    n927,
    n931,
    n930,
    n932
  );


  xor
  g897
  (
    n937,
    n932,
    n931,
    n225
  );


  xnor
  g898
  (
    n945,
    n892,
    n935
  );


  nor
  g899
  (
    n955,
    n902,
    n890
  );


  nand
  g900
  (
    n948,
    n888,
    n897
  );


  xor
  g901
  (
    n942,
    n889,
    n939
  );


  not
  g902
  (
    n946,
    n901
  );


  xnor
  g903
  (
    n963,
    n899,
    n933,
    n900
  );


  xor
  g904
  (
    n957,
    n898,
    n895,
    n885,
    n937
  );


  xor
  g905
  (
    n947,
    n897,
    n903,
    n894
  );


  nand
  g906
  (
    n944,
    n886,
    n890,
    n892,
    n936
  );


  nor
  g907
  (
    n959,
    n885,
    n933,
    n899,
    n900
  );


  or
  g908
  (
    n965,
    n935,
    n888,
    n936,
    n933
  );


  or
  g909
  (
    n960,
    n902,
    n933,
    n896,
    n937
  );


  or
  g910
  (
    n956,
    n937,
    n895,
    n896,
    n890
  );


  nor
  g911
  (
    n967,
    n887,
    n886,
    n890,
    n891
  );


  nand
  g912
  (
    n958,
    n934,
    n935,
    n902,
    n195
  );


  xor
  g913
  (
    n949,
    n934,
    n902,
    n889,
    n938
  );


  nand
  g914
  (
    n954,
    n887,
    n937,
    n889,
    n897
  );


  xnor
  g915
  (
    n962,
    n896,
    n936,
    n888,
    n891
  );


  or
  g916
  (
    n964,
    n939,
    n887,
    n886,
    n901
  );


  xor
  g917
  (
    n968,
    n891,
    n898,
    n894,
    n888
  );


  xor
  g918
  (
    n961,
    n898,
    n892,
    n895,
    n938
  );


  nor
  g919
  (
    n951,
    n901,
    n934,
    n935,
    n938
  );


  nor
  g920
  (
    n953,
    n886,
    n889,
    n892,
    n898
  );


  nor
  g921
  (
    n943,
    n896,
    n894,
    n900,
    n903
  );


  and
  g922
  (
    n952,
    n899,
    n899,
    n897,
    n900
  );


  xnor
  g923
  (
    n950,
    n936,
    n887,
    n938,
    n939
  );


  xnor
  g924
  (
    n966,
    n934,
    n903,
    n891,
    n895
  );


  not
  g925
  (
    n969,
    n965
  );


  not
  g926
  (
    n971,
    n969
  );


  buf
  g927
  (
    n970,
    n969
  );


  not
  g928
  (
    n972,
    n971
  );


  or
  g929
  (
    n976,
    n972,
    n940,
    n941
  );


  and
  g930
  (
    n974,
    n196,
    n940,
    n972
  );


  xnor
  g931
  (
    n973,
    n195,
    n939,
    n972,
    n941
  );


  and
  g932
  (
    n975,
    n941,
    n941,
    n196,
    n972
  );


  buf
  g933
  (
    n990,
    n974
  );


  buf
  g934
  (
    n987,
    n226
  );


  buf
  g935
  (
    n982,
    n226
  );


  not
  g936
  (
    n978,
    n975
  );


  buf
  g937
  (
    n992,
    n974
  );


  or
  g938
  (
    n984,
    n863,
    n227,
    n968,
    n229
  );


  nand
  g939
  (
    n985,
    n976,
    n976,
    n228,
    n966
  );


  nor
  g940
  (
    n983,
    n228,
    n863,
    n967,
    n230
  );


  xnor
  g941
  (
    n979,
    n973,
    n229,
    n861
  );


  xnor
  g942
  (
    n988,
    n974,
    n225,
    n863,
    n862
  );


  or
  g943
  (
    n980,
    n862,
    n227,
    n863,
    n976
  );


  or
  g944
  (
    n981,
    n973,
    n230,
    n975,
    n226
  );


  xor
  g945
  (
    n986,
    n973,
    n228,
    n976,
    n862
  );


  and
  g946
  (
    n989,
    n229,
    n228,
    n226,
    n862
  );


  xnor
  g947
  (
    n977,
    n973,
    n974,
    n227,
    n975
  );


  or
  g948
  (
    n991,
    n975,
    n230,
    n227,
    n225
  );


  not
  g949
  (
    n1009,
    n992
  );


  not
  g950
  (
    n1008,
    n981
  );


  xor
  g951
  (
    n1006,
    n991,
    n986,
    n987,
    n983
  );


  xor
  g952
  (
    n996,
    n981,
    n982,
    n985,
    n977
  );


  and
  g953
  (
    n999,
    n990,
    n983,
    n988
  );


  xor
  g954
  (
    n997,
    n987,
    n985,
    n980
  );


  xor
  g955
  (
    n993,
    n982,
    n992,
    n197,
    n989
  );


  xnor
  g956
  (
    n1000,
    n980,
    n979,
    n989,
    n982
  );


  xnor
  g957
  (
    n1001,
    n986,
    n197,
    n978,
    n981
  );


  xor
  g958
  (
    n994,
    n978,
    n196,
    n986,
    n197
  );


  nor
  g959
  (
    n995,
    n989,
    n991,
    n864,
    n992
  );


  xor
  g960
  (
    n1011,
    n981,
    n988,
    n197,
    n984
  );


  nor
  g961
  (
    n1004,
    n980,
    n984,
    n979,
    n864
  );


  nand
  g962
  (
    n1010,
    n987,
    n977,
    n864
  );


  xnor
  g963
  (
    n1005,
    n978,
    n985,
    n984,
    n990
  );


  nor
  g964
  (
    n1002,
    n978,
    n977,
    n980,
    n983
  );


  nand
  g965
  (
    n1012,
    n979,
    n984,
    n198,
    n987
  );


  nand
  g966
  (
    n1007,
    n991,
    n990,
    n986
  );


  nor
  g967
  (
    n998,
    n991,
    n988,
    n982,
    n196
  );


  nand
  g968
  (
    n1003,
    n989,
    n979,
    n988,
    n992
  );


  xor
  g969
  (
    n1016,
    n996,
    n1000,
    n997,
    n998
  );


  or
  g970
  (
    n1014,
    n996,
    n1001,
    n1002,
    n998
  );


  and
  g971
  (
    n1019,
    n999,
    n1000,
    n997,
    n1002
  );


  nor
  g972
  (
    n1013,
    n995,
    n996
  );


  xnor
  g973
  (
    n1017,
    n1000,
    n998,
    n997,
    n1001
  );


  and
  g974
  (
    n1020,
    n997,
    n995,
    n999,
    n1001
  );


  and
  g975
  (
    n1018,
    n999,
    n999,
    n1002,
    n995
  );


  xnor
  g976
  (
    n1015,
    n1002,
    n1001,
    n1000,
    n998
  );


  or
  g977
  (
    n1023,
    n1006,
    n1003,
    n1005,
    n1015
  );


  xnor
  g978
  (
    n1022,
    n1006,
    n1003,
    n1004,
    n1007
  );


  nand
  g979
  (
    n1024,
    n1014,
    n1003,
    n1005
  );


  xor
  g980
  (
    n1021,
    n1013,
    n1004,
    n1005,
    n1006
  );


  and
  g981
  (
    n1025,
    n1007,
    n1004,
    n1018,
    n1006
  );


  or
  g982
  (
    n1026,
    n1004,
    n1016,
    n1003,
    n1017
  );


  or
  g983
  (
    n1030,
    n1019,
    n1007,
    n904,
    n1025
  );


  nand
  g984
  (
    n1028,
    n904,
    n1020,
    n1007,
    n1024
  );


  xnor
  g985
  (
    KeyWire_0_23,
    n904,
    n230,
    n1022,
    n864
  );


  nor
  g986
  (
    n1027,
    n1023,
    n231,
    n865
  );


  buf
  g987
  (
    n1034,
    n1030
  );


  not
  g988
  (
    n1033,
    n1028
  );


  buf
  g989
  (
    n1031,
    n1027
  );


  not
  g990
  (
    n1035,
    n1030
  );


  buf
  g991
  (
    n1037,
    n1030
  );


  buf
  g992
  (
    n1036,
    n1030
  );


  nor
  g993
  (
    n1032,
    n1008,
    n1029
  );


  or
  g994
  (
    n1038,
    n1009,
    n1031,
    n1011
  );


  nand
  g995
  (
    n1042,
    n1031,
    n1011,
    n1010,
    n1009
  );


  nand
  g996
  (
    n1039,
    n1031,
    n1009,
    n1010
  );


  xor
  g997
  (
    n1041,
    n1010,
    n1008,
    n1011
  );


  and
  g998
  (
    n1040,
    n1008,
    n1031,
    n1010,
    n1032
  );


  and
  g999
  (
    n1043,
    n869,
    n928,
    n1038,
    n866
  );


  xor
  g1000
  (
    n1045,
    n867,
    n1034,
    n868,
    n869
  );


  nor
  g1001
  (
    n1049,
    n1033,
    n1042,
    n1035,
    n866
  );


  nor
  g1002
  (
    n1055,
    n1042,
    n866,
    n1037
  );


  nor
  g1003
  (
    n1059,
    n865,
    n869,
    n928,
    n1038
  );


  xor
  g1004
  (
    n1056,
    n1042,
    n870,
    n1039,
    n1041
  );


  nor
  g1005
  (
    n1060,
    n867,
    n1032,
    n1035,
    n868
  );


  xnor
  g1006
  (
    n1058,
    n1036,
    n867,
    n929,
    n1039
  );


  xnor
  g1007
  (
    n1052,
    n870,
    n1040,
    n928,
    n927
  );


  xnor
  g1008
  (
    n1050,
    n871,
    n1039,
    n1034,
    n1037
  );


  xnor
  g1009
  (
    n1054,
    n1032,
    n1037,
    n1040,
    n1034
  );


  nor
  g1010
  (
    n1048,
    n927,
    n1034,
    n1035,
    n1041
  );


  xor
  g1011
  (
    n1053,
    n1041,
    n1032,
    n1039,
    n868
  );


  nand
  g1012
  (
    n1047,
    n928,
    n868,
    n870,
    n1036
  );


  or
  g1013
  (
    n1044,
    n1037,
    n1033,
    n865,
    n1040
  );


  nand
  g1014
  (
    n1051,
    n1033,
    n1041,
    n1040,
    n1042
  );


  or
  g1015
  (
    n1046,
    n1035,
    n869,
    n865,
    n867
  );


  xor
  g1016
  (
    n1057,
    n1033,
    n1036,
    n870
  );


  buf
  g1017
  (
    n1071,
    n1059
  );


  buf
  g1018
  (
    n1078,
    n871
  );


  buf
  g1019
  (
    n1076,
    n1012
  );


  buf
  g1020
  (
    n1063,
    n871
  );


  not
  g1021
  (
    n1074,
    n1043
  );


  not
  g1022
  (
    n1075,
    n1056
  );


  not
  g1023
  (
    n1065,
    n1048
  );


  buf
  g1024
  (
    n1094,
    n1059
  );


  buf
  g1025
  (
    n1086,
    n872
  );


  buf
  g1026
  (
    n1067,
    n872
  );


  not
  g1027
  (
    n1087,
    n198
  );


  buf
  g1028
  (
    n1089,
    n1051
  );


  buf
  g1029
  (
    n1072,
    n1044
  );


  buf
  g1030
  (
    n1085,
    n1056
  );


  buf
  g1031
  (
    n1082,
    n929
  );


  buf
  g1032
  (
    n1092,
    n1054
  );


  buf
  g1033
  (
    n1088,
    n1012
  );


  not
  g1034
  (
    n1061,
    n871
  );


  buf
  g1035
  (
    n1064,
    n1060
  );


  not
  g1036
  (
    n1096,
    n1057
  );


  buf
  g1037
  (
    n1077,
    n1055
  );


  buf
  g1038
  (
    n1068,
    n1049
  );


  not
  g1039
  (
    n1093,
    n1055
  );


  not
  g1040
  (
    n1079,
    n1053
  );


  not
  g1041
  (
    n1080,
    n1057
  );


  not
  g1042
  (
    KeyWire_0_21,
    n231
  );


  not
  g1043
  (
    n1070,
    n1046
  );


  buf
  g1044
  (
    n1062,
    n1012
  );


  not
  g1045
  (
    n1091,
    n1052
  );


  buf
  g1046
  (
    n1084,
    n1056
  );


  xor
  g1047
  (
    n1073,
    n1055,
    n1058
  );


  nand
  g1048
  (
    n1081,
    n198,
    n1060,
    n1057,
    n1026
  );


  and
  g1049
  (
    n1069,
    n1055,
    n1059,
    n1047,
    n1060
  );


  or
  g1050
  (
    n1095,
    n1058,
    n1050,
    n1056,
    n1059
  );


  xnor
  g1051
  (
    n1066,
    n1057,
    n929,
    n1045,
    n1058
  );


  nand
  g1052
  (
    n1083,
    n1058,
    n929,
    n1012,
    n1060
  );


  buf
  g1053
  (
    n1121,
    n1071
  );


  buf
  g1054
  (
    n1120,
    n1067
  );


  not
  g1055
  (
    n1131,
    n1063
  );


  not
  g1056
  (
    n1103,
    n1073
  );


  buf
  g1057
  (
    n1144,
    n1068
  );


  buf
  g1058
  (
    n1124,
    n1070
  );


  buf
  g1059
  (
    n1122,
    n1076
  );


  not
  g1060
  (
    n1114,
    n1065
  );


  buf
  g1061
  (
    n1112,
    n1068
  );


  buf
  g1062
  (
    n1159,
    n1066
  );


  buf
  g1063
  (
    n1158,
    n1072
  );


  buf
  g1064
  (
    n1100,
    n1065
  );


  buf
  g1065
  (
    n1130,
    n1067
  );


  buf
  g1066
  (
    n1138,
    n1063
  );


  buf
  g1067
  (
    n1104,
    n1069
  );


  not
  g1068
  (
    n1156,
    n1075
  );


  not
  g1069
  (
    n1145,
    n1072
  );


  buf
  g1070
  (
    n1101,
    n1073
  );


  buf
  g1071
  (
    n1119,
    n1075
  );


  buf
  g1072
  (
    n1149,
    n1070
  );


  buf
  g1073
  (
    n1126,
    n1077
  );


  buf
  g1074
  (
    n1154,
    n1066
  );


  buf
  g1075
  (
    n1137,
    n1076
  );


  not
  g1076
  (
    n1133,
    n1061
  );


  buf
  g1077
  (
    n1098,
    n1072
  );


  buf
  g1078
  (
    n1109,
    n1063
  );


  buf
  g1079
  (
    n1160,
    n1068
  );


  buf
  g1080
  (
    n1129,
    n1067
  );


  buf
  g1081
  (
    n1115,
    n1073
  );


  not
  g1082
  (
    n1102,
    n1065
  );


  buf
  g1083
  (
    n1152,
    n1075
  );


  buf
  g1084
  (
    n1153,
    n1064
  );


  buf
  g1085
  (
    n1147,
    n1061
  );


  buf
  g1086
  (
    n1140,
    n1062
  );


  buf
  g1087
  (
    n1107,
    n1065
  );


  not
  g1088
  (
    n1127,
    n1073
  );


  not
  g1089
  (
    n1118,
    n1069
  );


  buf
  g1090
  (
    n1146,
    n1074
  );


  not
  g1091
  (
    n1110,
    n1066
  );


  buf
  g1092
  (
    n1117,
    n1064
  );


  not
  g1093
  (
    n1157,
    n1068
  );


  not
  g1094
  (
    n1150,
    n1070
  );


  not
  g1095
  (
    n1106,
    n1076
  );


  not
  g1096
  (
    n1128,
    n1064
  );


  not
  g1097
  (
    n1105,
    n1069
  );


  buf
  g1098
  (
    n1143,
    n1071
  );


  not
  g1099
  (
    n1141,
    n1071
  );


  buf
  g1100
  (
    n1132,
    n1066
  );


  not
  g1101
  (
    n1155,
    n1070
  );


  not
  g1102
  (
    n1142,
    n1072
  );


  not
  g1103
  (
    n1099,
    n1062
  );


  not
  g1104
  (
    n1123,
    n1064
  );


  not
  g1105
  (
    n1113,
    n1062
  );


  not
  g1106
  (
    n1116,
    n1071
  );


  not
  g1107
  (
    n1139,
    n1074
  );


  buf
  g1108
  (
    n1148,
    n1062
  );


  not
  g1109
  (
    n1108,
    n1075
  );


  buf
  g1110
  (
    n1125,
    n1077
  );


  buf
  g1111
  (
    n1135,
    n1074
  );


  buf
  g1112
  (
    n1136,
    n1069
  );


  not
  g1113
  (
    n1151,
    n1074
  );


  not
  g1114
  (
    n1111,
    n1067
  );


  buf
  g1115
  (
    n1097,
    n1076
  );


  not
  g1116
  (
    n1134,
    n1063
  );


  not
  g1117
  (
    n1225,
    n1088
  );


  buf
  g1118
  (
    n1316,
    n1115
  );


  buf
  g1119
  (
    n1229,
    n1157
  );


  buf
  g1120
  (
    n1162,
    n1108
  );


  buf
  g1121
  (
    n1191,
    n910
  );


  buf
  g1122
  (
    n1174,
    n1120
  );


  buf
  g1123
  (
    n1184,
    n1160
  );


  buf
  g1124
  (
    n1180,
    n1079
  );


  buf
  g1125
  (
    n1201,
    n1132
  );


  not
  g1126
  (
    n1352,
    n922
  );


  not
  g1127
  (
    n1236,
    n1082
  );


  buf
  g1128
  (
    n1347,
    n908
  );


  not
  g1129
  (
    n1173,
    n200
  );


  buf
  g1130
  (
    n1290,
    n1089
  );


  buf
  g1131
  (
    n1405,
    n919
  );


  not
  g1132
  (
    n1376,
    n1086
  );


  buf
  g1133
  (
    n1371,
    n1105
  );


  buf
  g1134
  (
    n1228,
    n917
  );


  not
  g1135
  (
    n1338,
    n1153
  );


  buf
  g1136
  (
    n1194,
    n1157
  );


  buf
  g1137
  (
    n1343,
    n920
  );


  buf
  g1138
  (
    n1409,
    n1148
  );


  not
  g1139
  (
    n1329,
    n1105
  );


  buf
  g1140
  (
    n1232,
    n208
  );


  not
  g1141
  (
    n1262,
    n1151
  );


  buf
  g1142
  (
    n1275,
    n1125
  );


  not
  g1143
  (
    n1164,
    n206
  );


  not
  g1144
  (
    n1357,
    n1080
  );


  not
  g1145
  (
    n1339,
    n1126
  );


  not
  g1146
  (
    n1259,
    n205
  );


  buf
  g1147
  (
    n1287,
    n212
  );


  buf
  g1148
  (
    n1374,
    n913
  );


  buf
  g1149
  (
    n1332,
    n911
  );


  buf
  g1150
  (
    n1285,
    n920
  );


  not
  g1151
  (
    n1326,
    n1111
  );


  not
  g1152
  (
    n1383,
    n921
  );


  buf
  g1153
  (
    n1234,
    n1149
  );


  not
  g1154
  (
    n1395,
    n918
  );


  not
  g1155
  (
    n1257,
    n918
  );


  buf
  g1156
  (
    n1381,
    n1111
  );


  buf
  g1157
  (
    n1226,
    n1111
  );


  buf
  g1158
  (
    n1212,
    n1136
  );


  buf
  g1159
  (
    n1227,
    n202
  );


  buf
  g1160
  (
    n1208,
    n1137
  );


  buf
  g1161
  (
    n1166,
    n1131
  );


  buf
  g1162
  (
    n1192,
    n200
  );


  buf
  g1163
  (
    n1384,
    n1083
  );


  buf
  g1164
  (
    n1344,
    n1106
  );


  buf
  g1165
  (
    n1355,
    n1127
  );


  not
  g1166
  (
    n1261,
    n1159
  );


  buf
  g1167
  (
    n1392,
    n1099
  );


  buf
  g1168
  (
    n1190,
    n1143
  );


  buf
  g1169
  (
    n1248,
    n1106
  );


  not
  g1170
  (
    n1266,
    n1148
  );


  buf
  g1171
  (
    n1312,
    n1145
  );


  not
  g1172
  (
    n1235,
    n1141
  );


  not
  g1173
  (
    n1411,
    n1118
  );


  buf
  g1174
  (
    n1350,
    n1081
  );


  not
  g1175
  (
    n1375,
    n1097
  );


  not
  g1176
  (
    n1233,
    n204
  );


  buf
  g1177
  (
    n1325,
    n1139
  );


  buf
  g1178
  (
    n1380,
    n1114
  );


  not
  g1179
  (
    n1303,
    n915
  );


  not
  g1180
  (
    n1373,
    n209
  );


  not
  g1181
  (
    n1291,
    n1137
  );


  not
  g1182
  (
    n1243,
    n923
  );


  buf
  g1183
  (
    n1361,
    n1134
  );


  buf
  g1184
  (
    n1378,
    n913
  );


  buf
  g1185
  (
    n1366,
    n1093
  );


  buf
  g1186
  (
    n1283,
    n1104
  );


  not
  g1187
  (
    n1245,
    n1120
  );


  not
  g1188
  (
    n1394,
    n207
  );


  not
  g1189
  (
    n1181,
    n1108
  );


  not
  g1190
  (
    n1237,
    n1122
  );


  not
  g1191
  (
    n1367,
    n1083
  );


  buf
  g1192
  (
    n1274,
    n1160
  );


  buf
  g1193
  (
    n1295,
    n207
  );


  buf
  g1194
  (
    n1305,
    n215
  );


  not
  g1195
  (
    n1284,
    n912
  );


  not
  g1196
  (
    n1300,
    n1096
  );


  buf
  g1197
  (
    n1319,
    n1143
  );


  buf
  g1198
  (
    n1175,
    n212
  );


  buf
  g1199
  (
    n1337,
    n1104
  );


  not
  g1200
  (
    n1340,
    n1150
  );


  not
  g1201
  (
    n1199,
    n1137
  );


  buf
  g1202
  (
    n1256,
    n908
  );


  buf
  g1203
  (
    n1252,
    n1091
  );


  buf
  g1204
  (
    n1265,
    n1149
  );


  not
  g1205
  (
    n1216,
    n1105
  );


  buf
  g1206
  (
    n1218,
    n208
  );


  buf
  g1207
  (
    n1186,
    n1121
  );


  not
  g1208
  (
    n1410,
    n1081
  );


  buf
  g1209
  (
    n1389,
    n1128
  );


  not
  g1210
  (
    n1296,
    n1131
  );


  buf
  g1211
  (
    n1416,
    n1140
  );


  not
  g1212
  (
    n1203,
    n1118
  );


  buf
  g1213
  (
    n1297,
    n202
  );


  buf
  g1214
  (
    n1177,
    n1131
  );


  buf
  g1215
  (
    n1210,
    n1130
  );


  buf
  g1216
  (
    n1314,
    n1122
  );


  not
  g1217
  (
    n1187,
    n211
  );


  not
  g1218
  (
    n1349,
    n1080
  );


  not
  g1219
  (
    n1358,
    n1120
  );


  buf
  g1220
  (
    n1204,
    n1098
  );


  not
  g1221
  (
    n1293,
    n908
  );


  buf
  g1222
  (
    n1353,
    n1124
  );


  buf
  g1223
  (
    n1396,
    n1129
  );


  not
  g1224
  (
    n1306,
    n1084
  );


  buf
  g1225
  (
    n1271,
    n200
  );


  buf
  g1226
  (
    n1264,
    n1095
  );


  not
  g1227
  (
    n1289,
    n1096
  );


  not
  g1228
  (
    n1231,
    n1144
  );


  buf
  g1229
  (
    n1205,
    n1086
  );


  not
  g1230
  (
    n1255,
    n920
  );


  not
  g1231
  (
    n1168,
    n907
  );


  not
  g1232
  (
    n1249,
    n210
  );


  buf
  g1233
  (
    n1189,
    n205
  );


  not
  g1234
  (
    n1336,
    n909
  );


  not
  g1235
  (
    n1185,
    n209
  );


  not
  g1236
  (
    n1412,
    n904
  );


  buf
  g1237
  (
    n1360,
    n914
  );


  not
  g1238
  (
    n1279,
    n912
  );


  not
  g1239
  (
    n1213,
    n1117
  );


  not
  g1240
  (
    n1278,
    n917
  );


  buf
  g1241
  (
    n1372,
    n1080
  );


  not
  g1242
  (
    n1224,
    n213
  );


  buf
  g1243
  (
    n1391,
    n1158
  );


  buf
  g1244
  (
    n1292,
    n906
  );


  buf
  g1245
  (
    n1345,
    n1143
  );


  not
  g1246
  (
    n1330,
    n906
  );


  buf
  g1247
  (
    n1400,
    n1094
  );


  not
  g1248
  (
    n1320,
    n1095
  );


  not
  g1249
  (
    n1379,
    n208
  );


  buf
  g1250
  (
    n1258,
    n1101
  );


  not
  g1251
  (
    n1183,
    n1133
  );


  buf
  g1252
  (
    n1348,
    n909
  );


  buf
  g1253
  (
    n1388,
    n906
  );


  buf
  g1254
  (
    n1220,
    n1138
  );


  buf
  g1255
  (
    n1341,
    n1135
  );


  not
  g1256
  (
    n1301,
    n1117
  );


  buf
  g1257
  (
    n1382,
    n1157
  );


  buf
  g1258
  (
    n1167,
    n1121
  );


  buf
  g1259
  (
    n1215,
    n1090
  );


  not
  g1260
  (
    n1351,
    n1119
  );


  not
  g1261
  (
    n1246,
    n911
  );


  not
  g1262
  (
    n1403,
    n1085
  );


  not
  g1263
  (
    n1322,
    n1139
  );


  buf
  g1264
  (
    n1402,
    n1128
  );


  buf
  g1265
  (
    n1222,
    n1129
  );


  buf
  g1266
  (
    n1407,
    n202
  );


  not
  g1267
  (
    n1318,
    n1144
  );


  not
  g1268
  (
    n1196,
    n1126
  );


  buf
  g1269
  (
    n1404,
    n1126
  );


  buf
  g1270
  (
    n1364,
    n1156
  );


  buf
  g1271
  (
    n1298,
    n1092
  );


  buf
  g1272
  (
    n1398,
    n1140
  );


  buf
  g1273
  (
    n1178,
    n1137
  );


  buf
  g1274
  (
    n1268,
    n1149
  );


  buf
  g1275
  (
    n1365,
    n1086
  );


  buf
  g1276
  (
    n1219,
    n1081
  );


  buf
  g1277
  (
    n1327,
    n911
  );


  buf
  g1278
  (
    n1324,
    n1153
  );


  not
  g1279
  (
    n1172,
    n1152
  );


  not
  g1280
  (
    n1281,
    n1079
  );


  buf
  g1281
  (
    n1335,
    n1147
  );


  buf
  g1282
  (
    n1334,
    n1120
  );


  buf
  g1283
  (
    n1299,
    n1115
  );


  buf
  g1284
  (
    n1304,
    n910
  );


  buf
  g1285
  (
    n1317,
    n1151
  );


  not
  g1286
  (
    n1214,
    n1086
  );


  buf
  g1287
  (
    n1333,
    n1102
  );


  not
  g1288
  (
    n1406,
    n923
  );


  not
  g1289
  (
    n1221,
    n204
  );


  not
  g1290
  (
    n1368,
    n1156
  );


  not
  g1291
  (
    n1182,
    n215
  );


  not
  g1292
  (
    KeyWire_0_15,
    n207
  );


  buf
  g1293
  (
    n1359,
    n1145
  );


  not
  g1294
  (
    n1390,
    n1106
  );


  not
  g1295
  (
    n1195,
    n1142
  );


  not
  g1296
  (
    n1313,
    n1159
  );


  buf
  g1297
  (
    n1244,
    n1107
  );


  nor
  g1298
  (
    n1288,
    n921,
    n1097,
    n1084,
    n1110
  );


  nor
  g1299
  (
    n1165,
    n215,
    n1155,
    n1101,
    n1093
  );


  and
  g1300
  (
    n1323,
    n1148,
    n214,
    n1154,
    n1090
  );


  nor
  g1301
  (
    n1193,
    n1138,
    n1134,
    n1103,
    n1116
  );


  xor
  g1302
  (
    n1200,
    n211,
    n1144,
    n1152,
    n1123
  );


  or
  g1303
  (
    n1415,
    n1145,
    n1125,
    n905,
    n1087
  );


  xnor
  g1304
  (
    n1310,
    n1142,
    n1116,
    n1152,
    n918
  );


  and
  g1305
  (
    n1211,
    n1106,
    n916,
    n199
  );


  nand
  g1306
  (
    n1399,
    n1077,
    n1154,
    n1092,
    n1127
  );


  nor
  g1307
  (
    n1346,
    n1153,
    n1122,
    n919,
    n201
  );


  xor
  g1308
  (
    n1207,
    n1134,
    n1122,
    n1121,
    n1083
  );


  nor
  g1309
  (
    n1209,
    n912,
    n210,
    n914,
    n1084
  );


  nor
  g1310
  (
    n1277,
    n1128,
    n1160,
    n213,
    n924
  );


  nor
  g1311
  (
    n1269,
    n1092,
    n1078,
    n1100
  );


  nor
  g1312
  (
    n1230,
    n1085,
    n919,
    n1158,
    n205
  );


  xnor
  g1313
  (
    n1408,
    n905,
    n1098,
    n915,
    n203
  );


  xor
  g1314
  (
    n1223,
    n1141,
    n201,
    n907,
    n1129
  );


  and
  g1315
  (
    n1387,
    n1087,
    n204,
    n1117,
    n1159
  );


  or
  g1316
  (
    n1282,
    n908,
    n1113,
    n1082,
    n1125
  );


  and
  g1317
  (
    n1188,
    n200,
    n211,
    n1085,
    n1087
  );


  or
  g1318
  (
    n1239,
    n1112,
    n921,
    n1111,
    n1152
  );


  nor
  g1319
  (
    n1385,
    n1103,
    n916,
    n1142,
    n1090
  );


  and
  g1320
  (
    n1331,
    n205,
    n203,
    n201,
    n1091
  );


  xnor
  g1321
  (
    n1397,
    n204,
    n214,
    n1089,
    n1108
  );


  xnor
  g1322
  (
    n1217,
    n214,
    n1155,
    n917,
    n909
  );


  or
  g1323
  (
    n1363,
    n922,
    n1095,
    n1102,
    n1078
  );


  nor
  g1324
  (
    n1242,
    n199,
    n1146,
    n1154,
    n1147
  );


  nand
  g1325
  (
    n1251,
    n1115,
    n920,
    n1160,
    n1097
  );


  xor
  g1326
  (
    n1267,
    n211,
    n914,
    n1108,
    n1099
  );


  nand
  g1327
  (
    n1393,
    n213,
    n918,
    n1124,
    n1107
  );


  xor
  g1328
  (
    n1276,
    n1133,
    n1081,
    n1089,
    n1113
  );


  nand
  g1329
  (
    n1250,
    n1103,
    n915,
    n1136,
    n1147
  );


  xor
  g1330
  (
    n1170,
    n202,
    n1097,
    n1093,
    n1132
  );


  xnor
  g1331
  (
    n1202,
    n201,
    n1134,
    n1103,
    n212
  );


  or
  g1332
  (
    n1362,
    n1126,
    n207,
    n905,
    n1118
  );


  xor
  g1333
  (
    n1263,
    n1119,
    n1131,
    n199,
    n1096
  );


  or
  g1334
  (
    n1179,
    n1149,
    n206,
    n912,
    n1129
  );


  or
  g1335
  (
    n1302,
    n1150,
    n1098,
    n1080,
    n1113
  );


  xor
  g1336
  (
    n1308,
    n1155,
    n1100,
    n1089,
    n1143
  );


  or
  g1337
  (
    n1328,
    n210,
    n909,
    n1146,
    n1084
  );


  and
  g1338
  (
    n1273,
    n1141,
    n1110,
    n1104,
    n208
  );


  and
  g1339
  (
    n1307,
    n1141,
    n1132,
    n1109,
    n1130
  );


  or
  g1340
  (
    n1247,
    n1095,
    n1148,
    n1158,
    n1101
  );


  nand
  g1341
  (
    n1401,
    n1140,
    n1135,
    n1159,
    n1124
  );


  xnor
  g1342
  (
    n1240,
    n1079,
    n1140,
    n1107,
    n1151
  );


  nand
  g1343
  (
    n1163,
    n199,
    n1116,
    n911,
    n1128
  );


  xnor
  g1344
  (
    n1294,
    n1147,
    n203,
    n1136,
    n1104
  );


  nor
  g1345
  (
    n1386,
    n1130,
    n922,
    n1127,
    n1094
  );


  nand
  g1346
  (
    n1369,
    n198,
    n1125,
    n1135,
    n1100
  );


  nand
  g1347
  (
    n1197,
    n1135,
    n1092,
    n907,
    n1101
  );


  nand
  g1348
  (
    n1311,
    n916,
    n1113,
    n1124,
    n1100
  );


  nor
  g1349
  (
    n1414,
    n1109,
    n1110,
    n1145,
    n906
  );


  and
  g1350
  (
    n1176,
    n1114,
    n1154,
    n910,
    n917
  );


  nor
  g1351
  (
    n1286,
    n1136,
    n212,
    n1155,
    n1157
  );


  xor
  g1352
  (
    n1171,
    n913,
    n1112,
    n1098,
    n1146
  );


  or
  g1353
  (
    n1315,
    n1099,
    n914,
    n1123,
    n1158
  );


  xnor
  g1354
  (
    n1169,
    n209,
    n923,
    n1096,
    n905
  );


  and
  g1355
  (
    n1241,
    n1077,
    n1094,
    n1110,
    n1093
  );


  nand
  g1356
  (
    n1161,
    n1094,
    n206,
    n1112,
    n1088
  );


  nand
  g1357
  (
    n1377,
    n1121,
    n1139,
    n1082,
    n1150
  );


  and
  g1358
  (
    n1321,
    n1102,
    n1091,
    n203,
    n1142
  );


  xnor
  g1359
  (
    n1280,
    n1079,
    n1156,
    n206,
    n1132
  );


  nor
  g1360
  (
    n1253,
    n1119,
    n1123,
    n1088,
    n1127
  );


  nor
  g1361
  (
    n1198,
    n1078,
    n913,
    n1109,
    n1102
  );


  xnor
  g1362
  (
    n1370,
    n1133,
    n919,
    n1117,
    n922
  );


  xnor
  g1363
  (
    n1309,
    n1118,
    n1144,
    n1088,
    n1138
  );


  nand
  g1364
  (
    n1413,
    n210,
    n907,
    n1083,
    n1105
  );


  nand
  g1365
  (
    n1206,
    n1090,
    n1114,
    n1091,
    n921
  );


  nand
  g1366
  (
    KeyWire_0_22,
    n1146,
    n1087,
    n915,
    n1114
  );


  nand
  g1367
  (
    n1354,
    n1119,
    n215,
    n1112,
    n1156
  );


  xnor
  g1368
  (
    n1254,
    n1138,
    n1109,
    n1107,
    n910
  );


  and
  g1369
  (
    n1270,
    n209,
    n1151,
    n1082,
    n1150
  );


  nand
  g1370
  (
    n1356,
    n213,
    n1139,
    n1130,
    n1153
  );


  nor
  g1371
  (
    n1238,
    n1123,
    n1115,
    n1099,
    n1133
  );


  or
  g1372
  (
    n1260,
    n923,
    n1085,
    n214,
    n1116
  );


  xor
  g1373
  (
    n1782,
    n1416,
    n770,
    n1351,
    n744
  );


  xnor
  g1374
  (
    n2235,
    n382,
    n1386,
    n1379,
    n1168
  );


  xor
  g1375
  (
    n1738,
    n1340,
    n241,
    n475,
    n471
  );


  xnor
  g1376
  (
    n1741,
    n262,
    n498,
    n233,
    n1227
  );


  or
  g1377
  (
    n1643,
    n1187,
    n394,
    n1268,
    n1221
  );


  and
  g1378
  (
    n1899,
    n1190,
    n287,
    n643,
    n734
  );


  or
  g1379
  (
    KeyWire_0_26,
    n1400,
    n406,
    n1350,
    n1170
  );


  and
  g1380
  (
    n1824,
    n541,
    n658,
    n1225,
    n346
  );


  nand
  g1381
  (
    n1596,
    n690,
    n470,
    n720,
    n239
  );


  xor
  g1382
  (
    n1719,
    n283,
    n441,
    n788,
    n536
  );


  nand
  g1383
  (
    n1884,
    n524,
    n777,
    n1285,
    n593
  );


  or
  g1384
  (
    n1549,
    n682,
    n575,
    n1228,
    n665
  );


  and
  g1385
  (
    KeyWire_0_4,
    n780,
    n1264,
    n413,
    n1357
  );


  and
  g1386
  (
    n2191,
    n389,
    n687,
    n611,
    n361
  );


  xnor
  g1387
  (
    n1595,
    n566,
    n656,
    n1173,
    n1409
  );


  nor
  g1388
  (
    n1720,
    n1260,
    n1340,
    n688,
    n363
  );


  xor
  g1389
  (
    n2122,
    n482,
    n1186,
    n1406,
    n362
  );


  nor
  g1390
  (
    n1902,
    n287,
    n695,
    n263,
    n363
  );


  xnor
  g1391
  (
    n1835,
    n434,
    n1365,
    n322,
    n637
  );


  xor
  g1392
  (
    n1739,
    n607,
    n1232,
    n375,
    n403
  );


  xor
  g1393
  (
    n1635,
    n744,
    n1239,
    n475,
    n1376
  );


  nor
  g1394
  (
    n2054,
    n352,
    n1415,
    n749,
    n733
  );


  nand
  g1395
  (
    n1992,
    n280,
    n249,
    n371,
    n1215
  );


  nor
  g1396
  (
    n1918,
    n391,
    n1257,
    n434,
    n660
  );


  nand
  g1397
  (
    n1925,
    n1384,
    n1348,
    n311,
    n1388
  );


  and
  g1398
  (
    n2143,
    n1377,
    n1282,
    n246,
    n804
  );


  nand
  g1399
  (
    n2146,
    n439,
    n293,
    n794,
    n1193
  );


  xnor
  g1400
  (
    n1496,
    n1214,
    n235,
    n1354,
    n1413
  );


  and
  g1401
  (
    n1502,
    n337,
    n776,
    n637,
    n475
  );


  xnor
  g1402
  (
    KeyWire_0_14,
    n365,
    n251,
    n549,
    n629
  );


  nor
  g1403
  (
    n1795,
    n696,
    n690,
    n489,
    n570
  );


  and
  g1404
  (
    n1750,
    n1217,
    n1169,
    n768,
    n391
  );


  xor
  g1405
  (
    n1690,
    n788,
    n502,
    n462,
    n500
  );


  or
  g1406
  (
    n2032,
    n345,
    n268,
    n415,
    n428
  );


  and
  g1407
  (
    n2167,
    n1347,
    n593,
    n1313,
    n1258
  );


  or
  g1408
  (
    n2211,
    n515,
    n787,
    n530,
    n801
  );


  xnor
  g1409
  (
    n1685,
    n1278,
    n1292,
    n661,
    n1171
  );


  nor
  g1410
  (
    n1933,
    n793,
    n1228,
    n1186,
    n1355
  );


  xnor
  g1411
  (
    n1715,
    n408,
    n583,
    n1233,
    n622
  );


  xor
  g1412
  (
    n2150,
    n1398,
    n749,
    n710,
    n238
  );


  or
  g1413
  (
    n1453,
    n341,
    n646,
    n1393,
    n1370
  );


  xor
  g1414
  (
    n1430,
    n642,
    n1315,
    n481,
    n601
  );


  or
  g1415
  (
    n1575,
    n278,
    n679,
    n456,
    n1322
  );


  xnor
  g1416
  (
    n1514,
    n1161,
    n1205,
    n653,
    n719
  );


  xnor
  g1417
  (
    n1988,
    n603,
    n604,
    n501,
    n240
  );


  or
  g1418
  (
    n2185,
    n302,
    n522,
    n1390,
    n1392
  );


  or
  g1419
  (
    n1996,
    n1396,
    n398,
    n592,
    n1386
  );


  or
  g1420
  (
    n2117,
    n272,
    n592,
    n273,
    n1218
  );


  xnor
  g1421
  (
    n1626,
    n1318,
    n1349,
    n1255,
    n258
  );


  xnor
  g1422
  (
    n1631,
    n495,
    n492,
    n701,
    n1286
  );


  or
  g1423
  (
    KeyWire_0_6,
    n397,
    n1329,
    n438,
    n645
  );


  xor
  g1424
  (
    n2036,
    n342,
    n510,
    n427,
    n1394
  );


  nand
  g1425
  (
    n1511,
    n328,
    n345,
    n473,
    n528
  );


  nor
  g1426
  (
    n1718,
    n487,
    n1400,
    n402,
    n600
  );


  xnor
  g1427
  (
    n1493,
    n327,
    n1226,
    n513,
    n1202
  );


  xor
  g1428
  (
    n1510,
    n796,
    n1334,
    n1374,
    n1294
  );


  xnor
  g1429
  (
    n1602,
    n638,
    n550,
    n1280,
    n585
  );


  xnor
  g1430
  (
    n2075,
    n1335,
    n420,
    n1234,
    n290
  );


  and
  g1431
  (
    n2096,
    n924,
    n531,
    n584,
    n1217
  );


  xor
  g1432
  (
    n1584,
    n709,
    n647,
    n872,
    n1288
  );


  xor
  g1433
  (
    n1498,
    n411,
    n543,
    n522,
    n553
  );


  nand
  g1434
  (
    n1500,
    n751,
    n802,
    n1269,
    n1163
  );


  nor
  g1435
  (
    n1763,
    n439,
    n294,
    n1314,
    n1383
  );


  nor
  g1436
  (
    n2018,
    n1206,
    n524,
    n1210,
    n451
  );


  and
  g1437
  (
    n1732,
    n1359,
    n466,
    n300,
    n718
  );


  or
  g1438
  (
    n2179,
    n626,
    n1185,
    n658,
    n1323
  );


  nand
  g1439
  (
    n2225,
    n750,
    n545,
    n526,
    n541
  );


  xnor
  g1440
  (
    n1445,
    n1172,
    n1358,
    n622,
    n479
  );


  and
  g1441
  (
    KeyWire_0_3,
    n289,
    n491,
    n489,
    n680
  );


  or
  g1442
  (
    n1564,
    n1185,
    n1293,
    n295,
    n1307
  );


  or
  g1443
  (
    n1943,
    n787,
    n734,
    n687,
    n253
  );


  nor
  g1444
  (
    n1759,
    n1231,
    n421,
    n1352,
    n1411
  );


  nor
  g1445
  (
    n1658,
    n670,
    n493,
    n501,
    n454
  );


  nor
  g1446
  (
    n2215,
    n698,
    n581,
    n320,
    n613
  );


  or
  g1447
  (
    n1600,
    n1257,
    n330,
    n484,
    n299
  );


  nor
  g1448
  (
    n1634,
    n771,
    n1334,
    n493,
    n1301
  );


  and
  g1449
  (
    n2240,
    n440,
    n800,
    n1251,
    n470
  );


  nor
  g1450
  (
    n1885,
    n362,
    n1354,
    n1362,
    n674
  );


  xnor
  g1451
  (
    n2184,
    n1300,
    n692,
    n260,
    n1364
  );


  nand
  g1452
  (
    n2133,
    n797,
    n699,
    n746,
    n377
  );


  or
  g1453
  (
    n1560,
    n519,
    n274,
    n676,
    n474
  );


  nor
  g1454
  (
    n2025,
    n1300,
    n557,
    n1397,
    n314
  );


  and
  g1455
  (
    n1994,
    n779,
    n689,
    n610,
    n357
  );


  nor
  g1456
  (
    n1494,
    n1198,
    n1211,
    n425,
    n730
  );


  or
  g1457
  (
    n2031,
    n1187,
    n799,
    n736,
    n511
  );


  xnor
  g1458
  (
    n1893,
    n1376,
    n717,
    n365,
    n1366
  );


  and
  g1459
  (
    n2228,
    n405,
    n565,
    n763,
    n796
  );


  nor
  g1460
  (
    n1665,
    n697,
    n516,
    n715,
    n1268
  );


  and
  g1461
  (
    n1915,
    n400,
    n1335,
    n334,
    n1319
  );


  and
  g1462
  (
    n2090,
    n579,
    n540,
    n1299,
    n1294
  );


  nor
  g1463
  (
    n1804,
    n335,
    n361,
    n452,
    n616
  );


  or
  g1464
  (
    n1946,
    n1326,
    n496,
    n293,
    n1362
  );


  nand
  g1465
  (
    n2124,
    n384,
    n545,
    n1215,
    n333
  );


  or
  g1466
  (
    n1481,
    n377,
    n590,
    n1363,
    n329
  );


  nand
  g1467
  (
    KeyWire_0_30,
    n571,
    n452,
    n420,
    n372
  );


  or
  g1468
  (
    KeyWire_0_8,
    n491,
    n498,
    n1336,
    n487
  );


  and
  g1469
  (
    n2014,
    n274,
    n647,
    n581,
    n1375
  );


  xnor
  g1470
  (
    n1431,
    n1225,
    n305,
    n486,
    n1253
  );


  nor
  g1471
  (
    n1477,
    n769,
    n477,
    n505,
    n1163
  );


  xnor
  g1472
  (
    n1855,
    n1351,
    n1243,
    n528,
    n1364
  );


  nor
  g1473
  (
    n1766,
    n642,
    n393,
    n1188,
    n492
  );


  xor
  g1474
  (
    n1958,
    n342,
    n496,
    n297,
    n684
  );


  xor
  g1475
  (
    n1426,
    n590,
    n1213,
    n759,
    n548
  );


  nor
  g1476
  (
    n1859,
    n1181,
    n1202,
    n1293,
    n1275
  );


  nor
  g1477
  (
    n1819,
    n343,
    n758,
    n761,
    n281
  );


  or
  g1478
  (
    n1615,
    n1345,
    n1348,
    n335,
    n642
  );


  nand
  g1479
  (
    n2227,
    n1371,
    n1246,
    n470,
    n1191
  );


  nor
  g1480
  (
    n2151,
    n639,
    n664,
    n236,
    n1252
  );


  xor
  g1481
  (
    n1423,
    n688,
    n232,
    n724,
    n626
  );


  nor
  g1482
  (
    n1694,
    n1356,
    n291,
    n631,
    n551
  );


  and
  g1483
  (
    n1667,
    n1276,
    n338,
    n474,
    n719
  );


  xnor
  g1484
  (
    n2012,
    n267,
    n341,
    n270,
    n1219
  );


  nand
  g1485
  (
    n1748,
    n348,
    n1207,
    n763,
    n494
  );


  nand
  g1486
  (
    n2026,
    n571,
    n302,
    n1369,
    n455
  );


  nor
  g1487
  (
    n1794,
    n437,
    n1196,
    n1166,
    n419
  );


  nand
  g1488
  (
    n1757,
    n575,
    n675,
    n648,
    n383
  );


  and
  g1489
  (
    n1546,
    n655,
    n286,
    n783,
    n324
  );


  nand
  g1490
  (
    n1834,
    n1228,
    n498,
    n407,
    n567
  );


  and
  g1491
  (
    n2186,
    n662,
    n1298,
    n469,
    n1192
  );


  nand
  g1492
  (
    n2058,
    n1196,
    n493,
    n612,
    n350
  );


  nor
  g1493
  (
    n1836,
    n1275,
    n1401,
    n641,
    n1378
  );


  and
  g1494
  (
    n1673,
    n318,
    n630,
    n1267,
    n431
  );


  xor
  g1495
  (
    n2206,
    n532,
    n1245,
    n500,
    n234
  );


  or
  g1496
  (
    n1917,
    n1209,
    n632,
    n559,
    n478
  );


  nor
  g1497
  (
    n1463,
    n1242,
    n1325,
    n253,
    n343
  );


  xnor
  g1498
  (
    n1568,
    n241,
    n1328,
    n289,
    n612
  );


  and
  g1499
  (
    n1588,
    n1413,
    n354,
    n1375,
    n625
  );


  and
  g1500
  (
    n1533,
    n1359,
    n573,
    n331,
    n1285
  );


  or
  g1501
  (
    n2077,
    n1344,
    n465,
    n1220,
    n298
  );


  and
  g1502
  (
    n1805,
    n650,
    n1392,
    n487,
    n277
  );


  and
  g1503
  (
    n2155,
    n613,
    n321,
    n325,
    n1393
  );


  or
  g1504
  (
    n1870,
    n529,
    n1367,
    n252,
    n603
  );


  and
  g1505
  (
    n2130,
    n1324,
    n397,
    n481,
    n497
  );


  or
  g1506
  (
    n2224,
    n1305,
    n476,
    n376,
    n538
  );


  and
  g1507
  (
    n1961,
    n513,
    n386,
    n650,
    n326
  );


  xnor
  g1508
  (
    n1882,
    n566,
    n529,
    n1210,
    n1168
  );


  xnor
  g1509
  (
    n1434,
    n1229,
    n271,
    n254,
    n315
  );


  nor
  g1510
  (
    n2027,
    n451,
    n1233,
    n595,
    n691
  );


  xnor
  g1511
  (
    n2009,
    n379,
    n513,
    n449,
    n793
  );


  xnor
  g1512
  (
    n2246,
    n1271,
    n508,
    n762,
    n1399
  );


  xor
  g1513
  (
    n1581,
    n1287,
    n353,
    n624,
    n422
  );


  xnor
  g1514
  (
    n1781,
    n1350,
    n370,
    n517,
    n294
  );


  or
  g1515
  (
    n1991,
    n681,
    n555,
    n629,
    n582
  );


  or
  g1516
  (
    n1540,
    n240,
    n1327,
    n1310,
    n455
  );


  and
  g1517
  (
    n1528,
    n1222,
    n744,
    n1213,
    n615
  );


  nor
  g1518
  (
    n2222,
    n394,
    n760,
    n1382,
    n1221
  );


  xor
  g1519
  (
    n1427,
    n494,
    n1222,
    n800,
    n614
  );


  nand
  g1520
  (
    n1490,
    n317,
    n1249,
    n434,
    n508
  );


  nand
  g1521
  (
    n1627,
    n732,
    n753,
    n623,
    n1167
  );


  or
  g1522
  (
    n2231,
    n400,
    n736,
    n1255,
    n452
  );


  and
  g1523
  (
    n1971,
    n804,
    n514,
    n1324,
    n742
  );


  or
  g1524
  (
    n2135,
    n337,
    n503,
    n296,
    n280
  );


  xnor
  g1525
  (
    n2020,
    n656,
    n464,
    n350,
    n287
  );


  or
  g1526
  (
    n2223,
    n506,
    n1282,
    n363,
    n359
  );


  or
  g1527
  (
    n1823,
    n1248,
    n457,
    n313,
    n610
  );


  xor
  g1528
  (
    n1471,
    n785,
    n298,
    n1409,
    n276
  );


  xor
  g1529
  (
    n2016,
    n1394,
    n1274,
    n403,
    n651
  );


  nor
  g1530
  (
    n1812,
    n438,
    n568,
    n523,
    n1268
  );


  and
  g1531
  (
    n1957,
    n311,
    n248,
    n249,
    n1390
  );


  nor
  g1532
  (
    n1497,
    n471,
    n776,
    n1295,
    n1231
  );


  and
  g1533
  (
    n2178,
    n1316,
    n564,
    n1271,
    n618
  );


  xor
  g1534
  (
    n1826,
    n442,
    n546,
    n1171,
    n620
  );


  nor
  g1535
  (
    KeyWire_0_17,
    n681,
    n271,
    n430,
    n245
  );


  nor
  g1536
  (
    n2171,
    n417,
    n1308,
    n700,
    n439
  );


  nand
  g1537
  (
    n1976,
    n398,
    n476,
    n242,
    n525
  );


  and
  g1538
  (
    n2092,
    n616,
    n1204,
    n251,
    n574
  );


  xor
  g1539
  (
    n1796,
    n1248,
    n1273,
    n597,
    n732
  );


  and
  g1540
  (
    n1811,
    n754,
    n620,
    n275,
    n801
  );


  nand
  g1541
  (
    n2049,
    n1230,
    n764,
    n426,
    n1278
  );


  and
  g1542
  (
    n1742,
    n329,
    n618,
    n1356,
    n713
  );


  nor
  g1543
  (
    n1903,
    n784,
    n752,
    n571,
    n743
  );


  or
  g1544
  (
    n1587,
    n1201,
    n1264,
    n497,
    n409
  );


  and
  g1545
  (
    n1534,
    n1265,
    n1357,
    n1411,
    n1307
  );


  xor
  g1546
  (
    n1504,
    n418,
    n1269,
    n284,
    n324
  );


  nand
  g1547
  (
    n1519,
    n461,
    n1311,
    n504,
    n1333
  );


  nor
  g1548
  (
    n2079,
    n341,
    n803,
    n1206,
    n242
  );


  or
  g1549
  (
    n2069,
    n347,
    n354,
    n672,
    n696
  );


  xnor
  g1550
  (
    n1810,
    n711,
    n1272,
    n605,
    n1299
  );


  nand
  g1551
  (
    n1865,
    n461,
    n778,
    n691,
    n1207
  );


  nor
  g1552
  (
    n1561,
    n415,
    n467,
    n598,
    n792
  );


  nor
  g1553
  (
    n1707,
    n1290,
    n518,
    n785,
    n524
  );


  xnor
  g1554
  (
    n1825,
    n1336,
    n731,
    n1317,
    n1163
  );


  and
  g1555
  (
    n1669,
    n548,
    n651,
    n1277,
    n473
  );


  xnor
  g1556
  (
    n1466,
    n1273,
    n1203,
    n522,
    n339
  );


  or
  g1557
  (
    n1524,
    n453,
    n1174,
    n1296,
    n274
  );


  and
  g1558
  (
    n1613,
    n1320,
    n1391,
    n392,
    n1388
  );


  or
  g1559
  (
    n1422,
    n617,
    n509,
    n737,
    n284
  );


  xnor
  g1560
  (
    n2145,
    n337,
    n313,
    n557,
    n791
  );


  xor
  g1561
  (
    n2107,
    n498,
    n445,
    n441,
    n456
  );


  or
  g1562
  (
    n1458,
    n1333,
    n1173,
    n301,
    n1397
  );


  xnor
  g1563
  (
    n1601,
    n390,
    n549,
    n1401,
    n546
  );


  xnor
  g1564
  (
    n1590,
    n470,
    n738,
    n599,
    n1204
  );


  xor
  g1565
  (
    n1576,
    n1180,
    n380,
    n437,
    n658
  );


  nor
  g1566
  (
    n1492,
    n1193,
    n763,
    n428,
    n1297
  );


  or
  g1567
  (
    n1959,
    n619,
    n1277,
    n244,
    n630
  );


  nor
  g1568
  (
    n1711,
    n517,
    n447,
    n646,
    n639
  );


  xor
  g1569
  (
    n1926,
    n795,
    n1261,
    n589,
    n670
  );


  xor
  g1570
  (
    n1905,
    n349,
    n402,
    n1396,
    n360
  );


  xnor
  g1571
  (
    n2165,
    n1188,
    n1319,
    n239,
    n1387
  );


  nor
  g1572
  (
    n1704,
    n534,
    n516,
    n326,
    n753
  );


  and
  g1573
  (
    n2216,
    n440,
    n290,
    n773,
    n1286
  );


  nand
  g1574
  (
    n1934,
    n1343,
    n243,
    n1177,
    n502
  );


  xor
  g1575
  (
    n2236,
    n393,
    n1312,
    n652,
    n304
  );


  xnor
  g1576
  (
    n1815,
    n1200,
    n1335,
    n694,
    n398
  );


  nor
  g1577
  (
    n1728,
    n380,
    n246,
    n587,
    n476
  );


  or
  g1578
  (
    n2212,
    n463,
    n721,
    n696,
    n504
  );


  xor
  g1579
  (
    n2102,
    n538,
    n1342,
    n1179,
    n1313
  );


  xnor
  g1580
  (
    n1773,
    n599,
    n608,
    n730,
    n278
  );


  nand
  g1581
  (
    n2226,
    n1266,
    n1164,
    n1353,
    n378
  );


  and
  g1582
  (
    n1563,
    n762,
    n778,
    n1288,
    n1328
  );


  and
  g1583
  (
    n1850,
    n556,
    n514,
    n339,
    n770
  );


  xor
  g1584
  (
    n1963,
    n648,
    n1398,
    n1286,
    n750
  );


  nor
  g1585
  (
    n1623,
    n735,
    n1330,
    n755,
    n1358
  );


  or
  g1586
  (
    n1436,
    n1209,
    n480,
    n279,
    n686
  );


  nor
  g1587
  (
    n2000,
    n1364,
    n344,
    n246,
    n655
  );


  xor
  g1588
  (
    n1867,
    n300,
    n700,
    n679,
    n590
  );


  or
  g1589
  (
    n1842,
    n740,
    n668,
    n1171,
    n325
  );


  nand
  g1590
  (
    n1969,
    n1200,
    n522,
    n466,
    n1377
  );


  xnor
  g1591
  (
    n1603,
    n709,
    n1307,
    n715,
    n768
  );


  or
  g1592
  (
    n1898,
    n1281,
    n1370,
    n789,
    n1397
  );


  and
  g1593
  (
    n1580,
    n1283,
    n631,
    n332,
    n387
  );


  xor
  g1594
  (
    n1432,
    n774,
    n523,
    n437,
    n722
  );


  nor
  g1595
  (
    n1809,
    n492,
    n369,
    n543,
    n689
  );


  or
  g1596
  (
    n1696,
    n1297,
    n571,
    n1381,
    n372
  );


  xor
  g1597
  (
    n1760,
    n410,
    n708,
    n628,
    n450
  );


  and
  g1598
  (
    n1443,
    n649,
    n1414,
    n775,
    n1164
  );


  or
  g1599
  (
    n1425,
    n1207,
    n606,
    n561,
    n1403
  );


  xnor
  g1600
  (
    n2040,
    n567,
    n1399,
    n596,
    n776
  );


  or
  g1601
  (
    n1931,
    n752,
    n792,
    n260,
    n568
  );


  xnor
  g1602
  (
    n1952,
    n1387,
    n314,
    n355,
    n718
  );


  xor
  g1603
  (
    n2213,
    n1191,
    n253,
    n729,
    n441
  );


  nor
  g1604
  (
    n1614,
    n1202,
    n307,
    n245,
    n410
  );


  or
  g1605
  (
    n2210,
    n1293,
    n1338,
    n1246,
    n1164
  );


  nand
  g1606
  (
    n1983,
    n701,
    n551,
    n464,
    n1167
  );


  nor
  g1607
  (
    n2042,
    n569,
    n499,
    n434,
    n248
  );


  xor
  g1608
  (
    n1752,
    n292,
    n660,
    n1262,
    n1286
  );


  and
  g1609
  (
    n1472,
    n636,
    n507,
    n1214,
    n603
  );


  nand
  g1610
  (
    n1641,
    n621,
    n708,
    n1247,
    n442
  );


  xor
  g1611
  (
    n1740,
    n769,
    n1162,
    n1174,
    n475
  );


  nand
  g1612
  (
    n1455,
    n561,
    n728,
    n1389,
    n1398
  );


  nor
  g1613
  (
    n2111,
    n448,
    n566,
    n1197,
    n1233
  );


  xnor
  g1614
  (
    n1892,
    n383,
    n375,
    n269,
    n720
  );


  xor
  g1615
  (
    n1936,
    n1224,
    n509,
    n1249,
    n1385
  );


  and
  g1616
  (
    n1827,
    n704,
    n536,
    n297,
    n713
  );


  xor
  g1617
  (
    n1828,
    n451,
    n607,
    n747,
    n1211
  );


  xor
  g1618
  (
    n1890,
    n412,
    n1343,
    n745,
    n558
  );


  xor
  g1619
  (
    n1522,
    n446,
    n468,
    n487,
    n1235
  );


  or
  g1620
  (
    n1444,
    n372,
    n395,
    n669,
    n428
  );


  nand
  g1621
  (
    n1878,
    n650,
    n1291,
    n418,
    n1337
  );


  nor
  g1622
  (
    n1947,
    n373,
    n404,
    n1243,
    n336
  );


  nand
  g1623
  (
    n1505,
    n1368,
    n407,
    n600,
    n680
  );


  xnor
  g1624
  (
    n1817,
    n1315,
    n1288,
    n1303,
    n1374
  );


  and
  g1625
  (
    n1841,
    n670,
    n1175,
    n739
  );


  xnor
  g1626
  (
    n1770,
    n667,
    n1394,
    n784,
    n1341
  );


  nor
  g1627
  (
    n1468,
    n722,
    n1407,
    n1261,
    n1327
  );


  and
  g1628
  (
    n1799,
    n594,
    n580,
    n1385,
    n644
  );


  nand
  g1629
  (
    n1659,
    n252,
    n582,
    n1236,
    n798
  );


  xnor
  g1630
  (
    n1869,
    n563,
    n1331,
    n641,
    n546
  );


  xor
  g1631
  (
    n1677,
    n700,
    n1190,
    n531,
    n1381
  );


  nand
  g1632
  (
    n1814,
    n1365,
    n714,
    n488,
    n260
  );


  xor
  g1633
  (
    n1632,
    n1210,
    n336,
    n754,
    n355
  );


  nor
  g1634
  (
    n1922,
    n350,
    n1383,
    n288,
    n255
  );


  nor
  g1635
  (
    n2193,
    n680,
    n1269,
    n1237,
    n1323
  );


  nand
  g1636
  (
    n1526,
    n264,
    n1232,
    n271,
    n562
  );


  or
  g1637
  (
    n1706,
    n1294,
    n758,
    n657,
    n1187
  );


  nor
  g1638
  (
    n1713,
    n322,
    n1308,
    n738,
    n1325
  );


  nor
  g1639
  (
    n1661,
    n499,
    n1238,
    n467,
    n583
  );


  and
  g1640
  (
    n1749,
    n1353,
    n1260,
    n427,
    n262
  );


  xor
  g1641
  (
    n1640,
    n304,
    n573,
    n286,
    n485
  );


  or
  g1642
  (
    n1990,
    n1355,
    n592,
    n1198,
    n466
  );


  or
  g1643
  (
    n1897,
    n1194,
    n282,
    n446,
    n1312
  );


  nor
  g1644
  (
    n1439,
    n559,
    n366,
    n537,
    n1340
  );


  and
  g1645
  (
    n2134,
    n384,
    n374,
    n1404,
    n385
  );


  nor
  g1646
  (
    n1998,
    n433,
    n1363,
    n413,
    n1343
  );


  or
  g1647
  (
    n2080,
    n1367,
    n526,
    n512,
    n1363
  );


  xor
  g1648
  (
    n2086,
    n568,
    n349,
    n418,
    n1299
  );


  or
  g1649
  (
    n1531,
    n254,
    n544,
    n1219,
    n1303
  );


  xor
  g1650
  (
    n1465,
    n1384,
    n299,
    n597,
    n1354
  );


  and
  g1651
  (
    n1985,
    n436,
    n510,
    n1239,
    n291
  );


  nor
  g1652
  (
    n2061,
    n1207,
    n352,
    n322,
    n1400
  );


  nor
  g1653
  (
    n1896,
    n504,
    n654,
    n673,
    n774
  );


  and
  g1654
  (
    n1442,
    n235,
    n555,
    n1345,
    n423
  );


  xor
  g1655
  (
    n2052,
    n1306,
    n1360,
    n609,
    n1183
  );


  and
  g1656
  (
    n1583,
    n721,
    n1368,
    n1219,
    n1212
  );


  or
  g1657
  (
    n1567,
    n1168,
    n723,
    n537,
    n625
  );


  nor
  g1658
  (
    n2001,
    n709,
    n1299,
    n604,
    n305
  );


  nand
  g1659
  (
    n1978,
    n318,
    n433,
    n546,
    n431
  );


  xor
  g1660
  (
    n2157,
    n1319,
    n609,
    n1379,
    n286
  );


  nor
  g1661
  (
    n1876,
    n1405,
    n1161,
    n1332,
    n250
  );


  nand
  g1662
  (
    n2153,
    n595,
    n1175,
    n1169,
    n537
  );


  nor
  g1663
  (
    n2154,
    n390,
    n607,
    n698,
    n482
  );


  and
  g1664
  (
    n1683,
    n1337,
    n1305,
    n371,
    n450
  );


  nor
  g1665
  (
    n1457,
    n1211,
    n678,
    n1172,
    n602
  );


  nor
  g1666
  (
    n1675,
    n1225,
    n521,
    n1192,
    n488
  );


  xnor
  g1667
  (
    n1907,
    n1321,
    n460,
    n272,
    n1415
  );


  nor
  g1668
  (
    n2047,
    n1369,
    n485,
    n1241,
    n728
  );


  xnor
  g1669
  (
    n1599,
    n457,
    n265,
    n239,
    n1256
  );


  nand
  g1670
  (
    n1512,
    n373,
    n669,
    n668,
    n1361
  );


  nor
  g1671
  (
    n1593,
    n1287,
    n1321,
    n1165,
    n384
  );


  and
  g1672
  (
    n1813,
    n1317,
    n1340,
    n803,
    n525
  );


  nand
  g1673
  (
    n2200,
    n381,
    n1170,
    n405,
    n659
  );


  nand
  g1674
  (
    n2139,
    n780,
    n374,
    n460,
    n626
  );


  nor
  g1675
  (
    n2169,
    n1278,
    n1392,
    n1325,
    n711
  );


  xor
  g1676
  (
    n1911,
    n745,
    n725,
    n1289,
    n558
  );


  and
  g1677
  (
    n1598,
    n717,
    n655,
    n545,
    n422
  );


  nand
  g1678
  (
    n1647,
    n718,
    n587,
    n536,
    n684
  );


  nand
  g1679
  (
    n1591,
    n579,
    n1401,
    n1346,
    n1276
  );


  nor
  g1680
  (
    n2189,
    n473,
    n359,
    n390,
    n739
  );


  xnor
  g1681
  (
    n1532,
    n1277,
    n299,
    n792,
    n652
  );


  or
  g1682
  (
    n1474,
    n1257,
    n553,
    n369,
    n739
  );


  xor
  g1683
  (
    n1778,
    n255,
    n1310,
    n1402,
    n761
  );


  nand
  g1684
  (
    n1592,
    n276,
    n502,
    n333,
    n1242
  );


  xnor
  g1685
  (
    n1930,
    n595,
    n401,
    n634,
    n448
  );


  or
  g1686
  (
    n1914,
    n779,
    n625,
    n745,
    n370
  );


  and
  g1687
  (
    n1672,
    n752,
    n1332,
    n282,
    n411
  );


  xor
  g1688
  (
    n1995,
    n640,
    n1289,
    n588,
    n363
  );


  xor
  g1689
  (
    n1803,
    n313,
    n425,
    n791,
    n481
  );


  xnor
  g1690
  (
    n1780,
    n772,
    n447,
    n691,
    n1331
  );


  or
  g1691
  (
    n1662,
    n692,
    n1328,
    n290,
    n1272
  );


  xor
  g1692
  (
    n1572,
    n544,
    n663,
    n605,
    n1330
  );


  and
  g1693
  (
    n1609,
    n301,
    n1208,
    n1414,
    n1239
  );


  xor
  g1694
  (
    n2053,
    n308,
    n645,
    n333,
    n1330
  );


  xor
  g1695
  (
    n1527,
    n1182,
    n1215,
    n643,
    n781
  );


  and
  g1696
  (
    n1687,
    n348,
    n798,
    n243,
    n628
  );


  or
  g1697
  (
    n1538,
    n1313,
    n1237,
    n608,
    n1306
  );


  and
  g1698
  (
    n1518,
    n421,
    n706,
    n673,
    n356
  );


  nor
  g1699
  (
    n1944,
    n1252,
    n742,
    n1391,
    n1197
  );


  xnor
  g1700
  (
    n1523,
    n1280,
    n551,
    n785,
    n259
  );


  xor
  g1701
  (
    n2230,
    n443,
    n465,
    n360,
    n726
  );


  xor
  g1702
  (
    n1579,
    n1289,
    n405,
    n376,
    n1396
  );


  and
  g1703
  (
    n1840,
    n644,
    n777,
    n683,
    n258
  );


  xor
  g1704
  (
    n2024,
    n765,
    n654,
    n532,
    n686
  );


  nand
  g1705
  (
    n1503,
    n627,
    n638,
    n653,
    n1368
  );


  xnor
  g1706
  (
    n2028,
    n775,
    n722,
    n562,
    n737
  );


  or
  g1707
  (
    n1636,
    n1259,
    n347,
    n1167,
    n351
  );


  nor
  g1708
  (
    n1837,
    n378,
    n1380,
    n324,
    n743
  );


  or
  g1709
  (
    n1558,
    n746,
    n639,
    n755,
    n698
  );


  or
  g1710
  (
    n2008,
    n295,
    n278,
    n352,
    n1387
  );


  nor
  g1711
  (
    n1703,
    n697,
    n1401,
    n1267,
    n740
  );


  nor
  g1712
  (
    n1948,
    n584,
    n385,
    n298,
    n501
  );


  and
  g1713
  (
    n2103,
    n733,
    n717,
    n1267,
    n1407
  );


  and
  g1714
  (
    n1729,
    n385,
    n798,
    n516,
    n652
  );


  and
  g1715
  (
    n1637,
    n1187,
    n1249,
    n1258,
    n483
  );


  xnor
  g1716
  (
    n1552,
    n706,
    n316,
    n398,
    n246
  );


  and
  g1717
  (
    n2084,
    n424,
    n517,
    n1290
  );


  nand
  g1718
  (
    n1831,
    n1297,
    n712,
    n1197,
    n373
  );


  nor
  g1719
  (
    n1765,
    n303,
    n1310,
    n585,
    n447
  );


  xnor
  g1720
  (
    n1866,
    n1292,
    n1320,
    n418,
    n1382
  );


  xnor
  g1721
  (
    n2076,
    n430,
    n1393,
    n1295,
    n653
  );


  or
  g1722
  (
    n2164,
    n724,
    n767,
    n1244,
    n268
  );


  nand
  g1723
  (
    n1565,
    n338,
    n550,
    n685,
    n372
  );


  or
  g1724
  (
    n1589,
    n644,
    n530,
    n346,
    n495
  );


  nand
  g1725
  (
    n1721,
    n542,
    n1274,
    n248,
    n252
  );


  xor
  g1726
  (
    n2190,
    n462,
    n499,
    n611,
    n796
  );


  xor
  g1727
  (
    n1774,
    n612,
    n327,
    n637,
    n1189
  );


  or
  g1728
  (
    n1838,
    n1261,
    n660,
    n1397,
    n324
  );


  nor
  g1729
  (
    n1606,
    n578,
    n577,
    n629,
    n420
  );


  or
  g1730
  (
    n1862,
    n1347,
    n714,
    n586,
    n245
  );


  xor
  g1731
  (
    n2093,
    n685,
    n604,
    n472,
    n686
  );


  nand
  g1732
  (
    n2089,
    n550,
    n1352,
    n576,
    n1182
  );


  or
  g1733
  (
    n2044,
    n1220,
    n388,
    n567,
    n415
  );


  nor
  g1734
  (
    n1499,
    n621,
    n1330,
    n583,
    n412
  );


  nand
  g1735
  (
    n2199,
    n417,
    n362,
    n515,
    n556
  );


  or
  g1736
  (
    n1785,
    n1193,
    n270,
    n724,
    n451
  );


  nand
  g1737
  (
    n1999,
    n1196,
    n1229,
    n599,
    n1281
  );


  nand
  g1738
  (
    n1951,
    n465,
    n1183,
    n519,
    n1181
  );


  xor
  g1739
  (
    n1806,
    n688,
    n1395,
    n761,
    n539
  );


  or
  g1740
  (
    n1864,
    n448,
    n1339,
    n1359,
    n644
  );


  or
  g1741
  (
    n2129,
    n791,
    n392,
    n606,
    n1342
  );


  xnor
  g1742
  (
    n2207,
    n347,
    n1190,
    n323,
    n376
  );


  nor
  g1743
  (
    n2082,
    n1216,
    n773,
    n507,
    n266
  );


  nor
  g1744
  (
    n1744,
    n471,
    n627,
    n309,
    n317
  );


  nor
  g1745
  (
    n2205,
    n236,
    n1326,
    n584,
    n1239
  );


  nor
  g1746
  (
    n2170,
    n1407,
    n1412,
    n1339,
    n759
  );


  or
  g1747
  (
    n2046,
    n1321,
    n756,
    n1195,
    n619
  );


  xnor
  g1748
  (
    n2132,
    n256,
    n467,
    n245,
    n553
  );


  xnor
  g1749
  (
    n1639,
    n401,
    n1344,
    n748,
    n512
  );


  xnor
  g1750
  (
    n1830,
    n769,
    n344,
    n676,
    n378
  );


  nor
  g1751
  (
    n1970,
    n494,
    n532,
    n497,
    n1310
  );


  or
  g1752
  (
    n2003,
    n1253,
    n277,
    n345,
    n1166
  );


  xnor
  g1753
  (
    n2029,
    n567,
    n1233,
    n735,
    n614
  );


  nor
  g1754
  (
    n2037,
    n389,
    n634,
    n1409,
    n739
  );


  and
  g1755
  (
    n1642,
    n1316,
    n238,
    n308,
    n494
  );


  or
  g1756
  (
    n1428,
    n1250,
    n704,
    n247,
    n453
  );


  nand
  g1757
  (
    n1910,
    n1238,
    n764,
    n1309,
    n564
  );


  nand
  g1758
  (
    n2104,
    n266,
    n285,
    n1265,
    n609
  );


  xor
  g1759
  (
    n2094,
    n585,
    n573,
    n1362,
    n1244
  );


  xnor
  g1760
  (
    n1450,
    n407,
    n477,
    n382,
    n249
  );


  or
  g1761
  (
    n1495,
    n292,
    n1331,
    n640,
    n493
  );


  nor
  g1762
  (
    n1743,
    n1392,
    n386,
    n746,
    n485
  );


  xnor
  g1763
  (
    n1419,
    n531,
    n1322,
    n579,
    n443
  );


  or
  g1764
  (
    n1491,
    n518,
    n663,
    n263,
    n387
  );


  xnor
  g1765
  (
    n2004,
    n284,
    n668,
    n463,
    n1265
  );


  nand
  g1766
  (
    n1989,
    n754,
    n247,
    n1346,
    n1258
  );


  xor
  g1767
  (
    n1845,
    n342,
    n320,
    n1245,
    n790
  );


  xnor
  g1768
  (
    n1480,
    n266,
    n234,
    n1178,
    n1250
  );


  nand
  g1769
  (
    n1923,
    n1256,
    n275,
    n1223,
    n303
  );


  nand
  g1770
  (
    n1965,
    n726,
    n1204,
    n344,
    n1247
  );


  xor
  g1771
  (
    KeyWire_0_28,
    n356,
    n481,
    n482,
    n692
  );


  and
  g1772
  (
    n1577,
    n706,
    n328,
    n269,
    n505
  );


  and
  g1773
  (
    n1972,
    n625,
    n659,
    n327,
    n924
  );


  xnor
  g1774
  (
    n1790,
    n285,
    n444,
    n705,
    n364
  );


  and
  g1775
  (
    n1784,
    n653,
    n379,
    n730,
    n1213
  );


  nand
  g1776
  (
    n1544,
    n1324,
    n772,
    n309,
    n1408
  );


  or
  g1777
  (
    n1555,
    n1284,
    n741,
    n687,
    n361
  );


  xor
  g1778
  (
    n1982,
    n684,
    n638,
    n589,
    n733
  );


  nand
  g1779
  (
    n1501,
    n1245,
    n1219,
    n491,
    n1230
  );


  and
  g1780
  (
    n1429,
    n1243,
    n558,
    n1367,
    n237
  );


  xnor
  g1781
  (
    n1653,
    n465,
    n1338,
    n768,
    n506
  );


  nand
  g1782
  (
    n2119,
    n1225,
    n334,
    n252,
    n601
  );


  nand
  g1783
  (
    n2045,
    n1234,
    n613,
    n768,
    n435
  );


  or
  g1784
  (
    n2176,
    n514,
    n1335,
    n535,
    n1341
  );


  or
  g1785
  (
    n1521,
    n371,
    n542,
    n510,
    n673
  );


  nor
  g1786
  (
    n1802,
    n1338,
    n1178,
    n560,
    n1242
  );


  nand
  g1787
  (
    n1473,
    n686,
    n664,
    n495,
    n340
  );


  nor
  g1788
  (
    n1987,
    n728,
    n539,
    n761,
    n660
  );


  nand
  g1789
  (
    n2041,
    n614,
    n509,
    n1304,
    n416
  );


  xnor
  g1790
  (
    n1452,
    n277,
    n1261,
    n569,
    n468
  );


  and
  g1791
  (
    n1776,
    n445,
    n450,
    n421,
    n358
  );


  nor
  g1792
  (
    n1515,
    n1200,
    n780,
    n543,
    n396
  );


  xor
  g1793
  (
    n1921,
    n782,
    n552,
    n566,
    n1411
  );


  xor
  g1794
  (
    n1668,
    n557,
    n637,
    n609,
    n1208
  );


  and
  g1795
  (
    n1697,
    n435,
    n667,
    n570,
    n1229
  );


  xnor
  g1796
  (
    n2100,
    n1297,
    n1380,
    n663,
    n330
  );


  xnor
  g1797
  (
    n1682,
    n801,
    n618,
    n1333,
    n428
  );


  xor
  g1798
  (
    n2098,
    n1382,
    n1176,
    n701,
    n1216
  );


  and
  g1799
  (
    n2101,
    n321,
    n515,
    n1347,
    n765
  );


  nand
  g1800
  (
    n1912,
    n323,
    n626,
    n798,
    n725
  );


  xnor
  g1801
  (
    n1791,
    n1316,
    n591,
    n1339,
    n758
  );


  xnor
  g1802
  (
    n2159,
    n1241,
    n1379,
    n1388,
    n670
  );


  xnor
  g1803
  (
    n2158,
    n469,
    n1398,
    n377,
    n445
  );


  xor
  g1804
  (
    n2217,
    n731,
    n232,
    n349,
    n268
  );


  nand
  g1805
  (
    n1554,
    n432,
    n751,
    n640,
    n438
  );


  nor
  g1806
  (
    n1984,
    n1184,
    n1185,
    n1281,
    n1349
  );


  xor
  g1807
  (
    n1945,
    n1204,
    n1348,
    n654,
    n1289
  );


  xor
  g1808
  (
    n2085,
    n1243,
    n685,
    n1362,
    n479
  );


  or
  g1809
  (
    n2019,
    n315,
    n423,
    n1179,
    n459
  );


  nor
  g1810
  (
    n1821,
    n616,
    n310,
    n1358,
    n258
  );


  nand
  g1811
  (
    n1679,
    n1413,
    n1236,
    n331,
    n429
  );


  or
  g1812
  (
    n1758,
    n489,
    n1214,
    n623
  );


  nand
  g1813
  (
    n2065,
    n500,
    n729,
    n574,
    n436
  );


  xnor
  g1814
  (
    n1769,
    n1170,
    n235,
    n1318,
    n394
  );


  nand
  g1815
  (
    n2232,
    n272,
    n257,
    n793,
    n683
  );


  nor
  g1816
  (
    n1680,
    n1264,
    n381,
    n1169,
    n799
  );


  and
  g1817
  (
    n1462,
    n679,
    n715,
    n1210,
    n496
  );


  nand
  g1818
  (
    n1756,
    n1314,
    n1314,
    n771,
    n1252
  );


  nor
  g1819
  (
    n1787,
    n399,
    n766,
    n1226,
    n525
  );


  nand
  g1820
  (
    n1833,
    n771,
    n1346,
    n729,
    n378
  );


  nor
  g1821
  (
    n2174,
    n461,
    n598,
    n539,
    n1205
  );


  xor
  g1822
  (
    n2201,
    n1366,
    n250,
    n1370,
    n627
  );


  nor
  g1823
  (
    n1816,
    n1323,
    n1384,
    n621,
    n439
  );


  xor
  g1824
  (
    n2106,
    n1324,
    n1209,
    n397,
    n1178
  );


  xnor
  g1825
  (
    n2074,
    n473,
    n547,
    n632,
    n247
  );


  or
  g1826
  (
    n1767,
    n585,
    n331,
    n579,
    n366
  );


  xnor
  g1827
  (
    n1857,
    n1205,
    n330,
    n689,
    n593
  );


  xnor
  g1828
  (
    n1953,
    n294,
    n665,
    n339,
    n486
  );


  nor
  g1829
  (
    n2051,
    n1280,
    n707,
    n782,
    n261
  );


  xnor
  g1830
  (
    n1624,
    n1162,
    n779,
    n577,
    n716
  );


  nor
  g1831
  (
    KeyWire_0_25,
    n784,
    n368,
    n749,
    n513
  );


  and
  g1832
  (
    n2071,
    n1267,
    n520,
    n454,
    n321
  );


  or
  g1833
  (
    n2088,
    n1271,
    n316,
    n588,
    n365
  );


  xor
  g1834
  (
    n1908,
    n273,
    n1368,
    n1381,
    n1374
  );


  nor
  g1835
  (
    n1977,
    n1191,
    n273,
    n262,
    n787
  );


  xor
  g1836
  (
    n2121,
    n1273,
    n669,
    n297,
    n562
  );


  and
  g1837
  (
    n1920,
    n666,
    n1350,
    n256,
    n348
  );


  and
  g1838
  (
    n1786,
    n715,
    n610,
    n402,
    n676
  );


  xnor
  g1839
  (
    n2113,
    n1408,
    n360,
    n704,
    n293
  );


  and
  g1840
  (
    n2181,
    n295,
    n1345,
    n535,
    n1246
  );


  xnor
  g1841
  (
    n1726,
    n369,
    n1175,
    n799,
    n1388
  );


  and
  g1842
  (
    n2137,
    n457,
    n323,
    n328,
    n1199
  );


  or
  g1843
  (
    n2221,
    n1317,
    n296,
    n659,
    n757
  );


  nor
  g1844
  (
    n1722,
    n366,
    n695,
    n1179,
    n390
  );


  xor
  g1845
  (
    n1798,
    n463,
    n501,
    n358,
    n1223
  );


  and
  g1846
  (
    n2066,
    n1254,
    n1185,
    n790,
    n735
  );


  and
  g1847
  (
    n1935,
    n620,
    n725,
    n777,
    n602
  );


  and
  g1848
  (
    n1734,
    n340,
    n540,
    n559,
    n1375
  );


  xnor
  g1849
  (
    n1916,
    n742,
    n1415,
    n361,
    n464
  );


  and
  g1850
  (
    n1863,
    n785,
    n749,
    n1262,
    n703
  );


  and
  g1851
  (
    n1949,
    n1260,
    n561,
    n472,
    n722
  );


  or
  g1852
  (
    n1547,
    n568,
    n1336,
    n547,
    n393
  );


  xor
  g1853
  (
    n1913,
    n1309,
    n1217,
    n713,
    n442
  );


  nand
  g1854
  (
    n1582,
    n433,
    n669,
    n773,
    n1197
  );


  nand
  g1855
  (
    n1844,
    n436,
    n1162,
    n1228,
    n1184
  );


  nand
  g1856
  (
    n2149,
    n723,
    n413,
    n484,
    n564
  );


  or
  g1857
  (
    n1461,
    n270,
    n528,
    n1255,
    n429
  );


  or
  g1858
  (
    n1895,
    n1180,
    n1327,
    n733,
    n318
  );


  or
  g1859
  (
    n2073,
    n623,
    n693,
    n507,
    n612
  );


  or
  g1860
  (
    n1625,
    n610,
    n1224,
    n479,
    n720
  );


  or
  g1861
  (
    n1605,
    n1235,
    n275,
    n608,
    n714
  );


  and
  g1862
  (
    n1822,
    n243,
    n708,
    n1284,
    n1279
  );


  xnor
  g1863
  (
    n1861,
    n1247,
    n538,
    n1407,
    n781
  );


  nand
  g1864
  (
    n2110,
    n601,
    n1161,
    n440,
    n716
  );


  xnor
  g1865
  (
    n1848,
    n261,
    n1246,
    n595,
    n666
  );


  nand
  g1866
  (
    n2097,
    n628,
    n301,
    n794,
    n770
  );


  nand
  g1867
  (
    n1604,
    n1412,
    n427,
    n1380,
    n547
  );


  xnor
  g1868
  (
    n1446,
    n759,
    n281,
    n1301,
    n723
  );


  nand
  g1869
  (
    n1611,
    n529,
    n597,
    n319,
    n242
  );


  or
  g1870
  (
    n2064,
    n1240,
    n395,
    n536,
    n371
  );


  xnor
  g1871
  (
    n1877,
    n599,
    n241,
    n740,
    n1277
  );


  or
  g1872
  (
    n2067,
    n1399,
    n627,
    n266,
    n1181
  );


  nand
  g1873
  (
    n1557,
    n1188,
    n1339,
    n776,
    n296
  );


  nand
  g1874
  (
    n1708,
    n478,
    n274,
    n453,
    n1173
  );


  and
  g1875
  (
    n1441,
    n600,
    n272,
    n682,
    n410
  );


  nor
  g1876
  (
    n2013,
    n1367,
    n804,
    n1259,
    n766
  );


  nand
  g1877
  (
    n1705,
    n374,
    n352,
    n1274,
    n554
  );


  or
  g1878
  (
    n1654,
    n480,
    n1222,
    n383,
    n583
  );


  xnor
  g1879
  (
    n1612,
    n705,
    n611,
    n456,
    n533
  );


  nand
  g1880
  (
    n1793,
    n444,
    n737,
    n1291,
    n279
  );


  xor
  g1881
  (
    n1839,
    n289,
    n765,
    n1403,
    n693
  );


  nand
  g1882
  (
    n2244,
    n276,
    n642,
    n1377,
    n775
  );


  nor
  g1883
  (
    n1929,
    n326,
    n1338,
    n256,
    n1215
  );


  xnor
  g1884
  (
    n2072,
    n511,
    n773,
    n409,
    n332
  );


  or
  g1885
  (
    n2220,
    n1229,
    n354,
    n286,
    n435
  );


  xnor
  g1886
  (
    n1880,
    n1334,
    n1352,
    n780,
    n336
  );


  and
  g1887
  (
    n1709,
    n1177,
    n427,
    n355,
    n1161
  );


  nand
  g1888
  (
    n1578,
    n464,
    n782,
    n605,
    n1296
  );


  nor
  g1889
  (
    n2234,
    n667,
    n675,
    n1329,
    n367
  );


  xnor
  g1890
  (
    KeyWire_0_27,
    n678,
    n472,
    n762,
    n691
  );


  nand
  g1891
  (
    n2237,
    n1251,
    n1165,
    n634,
    n490
  );


  and
  g1892
  (
    n1543,
    n1411,
    n1329,
    n646,
    n285
  );


  and
  g1893
  (
    n2188,
    n524,
    n315,
    n1211,
    n617
  );


  and
  g1894
  (
    n2087,
    n512,
    n717,
    n306,
    n604
  );


  and
  g1895
  (
    n1792,
    n259,
    n534,
    n260,
    n802
  );


  or
  g1896
  (
    n1849,
    n1315,
    n711,
    n1223,
    n1182
  );


  or
  g1897
  (
    n2243,
    n647,
    n317,
    n336,
    n742
  );


  xnor
  g1898
  (
    n2140,
    n356,
    n403,
    n661,
    n619
  );


  xor
  g1899
  (
    n2034,
    n736,
    n1288,
    n381,
    n601
  );


  nand
  g1900
  (
    n1747,
    n682,
    n754,
    n663,
    n1236
  );


  or
  g1901
  (
    n1710,
    n678,
    n382,
    n1279,
    n1300
  );


  and
  g1902
  (
    n1650,
    n1232,
    n1332,
    n1272,
    n560
  );


  xnor
  g1903
  (
    n2038,
    n1263,
    n1205,
    n654,
    n549
  );


  nand
  g1904
  (
    n1617,
    n519,
    n638,
    n1343,
    n622
  );


  xnor
  g1905
  (
    n1768,
    n1305,
    n364,
    n319,
    n396
  );


  or
  g1906
  (
    n2166,
    n1366,
    n569,
    n483,
    n1222
  );


  xor
  g1907
  (
    n1968,
    n496,
    n391,
    n705,
    n783
  );


  xor
  g1908
  (
    n1666,
    n256,
    n364,
    n681,
    n772
  );


  xor
  g1909
  (
    n1941,
    n1373,
    n747,
    n593,
    n554
  );


  nor
  g1910
  (
    n1847,
    n1195,
    n310,
    n292
  );


  xnor
  g1911
  (
    n2081,
    n288,
    n795,
    n232,
    n1301
  );


  nand
  g1912
  (
    n1417,
    n1396,
    n393,
    n301,
    n586
  );


  xor
  g1913
  (
    n1464,
    n436,
    n549,
    n681,
    n656
  );


  xnor
  g1914
  (
    n2208,
    n778,
    n1404,
    n702,
    n640
  );


  xnor
  g1915
  (
    n1712,
    n453,
    n617,
    n683,
    n788
  );


  and
  g1916
  (
    n1421,
    n426,
    n1351,
    n702,
    n419
  );


  nor
  g1917
  (
    n2030,
    n435,
    n1287,
    n423,
    n1325
  );


  xor
  g1918
  (
    n2055,
    n1266,
    n237,
    n312,
    n1353
  );


  nand
  g1919
  (
    n1485,
    n1326,
    n572,
    n412,
    n588
  );


  nor
  g1920
  (
    n1789,
    n1183,
    n1230,
    n374,
    n531
  );


  or
  g1921
  (
    n1437,
    n790,
    n456,
    n542,
    n344
  );


  nand
  g1922
  (
    n2114,
    n396,
    n251,
    n261,
    n1282
  );


  nor
  g1923
  (
    n2125,
    n1258,
    n587,
    n258,
    n526
  );


  or
  g1924
  (
    n1886,
    n703,
    n234,
    n343,
    n800
  );


  and
  g1925
  (
    n1702,
    n235,
    n295,
    n596,
    n581
  );


  xor
  g1926
  (
    n1674,
    n283,
    n652,
    n478,
    n1318
  );


  xor
  g1927
  (
    n1894,
    n400,
    n454,
    n1244,
    n1403
  );


  and
  g1928
  (
    n1868,
    n1372,
    n310,
    n651,
    n560
  );


  nand
  g1929
  (
    n1820,
    n1256,
    n462,
    n774,
    n635
  );


  xor
  g1930
  (
    n1559,
    n535,
    n1177,
    n527,
    n268
  );


  xor
  g1931
  (
    n1858,
    n541,
    n290,
    n236,
    n559
  );


  nand
  g1932
  (
    n1919,
    n1399,
    n1220,
    n615,
    n1387
  );


  xnor
  g1933
  (
    n1751,
    n1235,
    n247,
    n747,
    n1199
  );


  nor
  g1934
  (
    n2039,
    n365,
    n402,
    n578,
    n448
  );


  xnor
  g1935
  (
    n1993,
    n1255,
    n657,
    n1250,
    n1321
  );


  nand
  g1936
  (
    n1986,
    n1303,
    n302,
    n576,
    n1360
  );


  and
  g1937
  (
    n1548,
    n1403,
    n511,
    n565,
    n697
  );


  nor
  g1938
  (
    n1681,
    n1295,
    n572,
    n1199,
    n389
  );


  or
  g1939
  (
    n1714,
    n1201,
    n1217,
    n639,
    n455
  );


  xor
  g1940
  (
    n2007,
    n629,
    n523,
    n320,
    n552
  );


  and
  g1941
  (
    n2116,
    n1166,
    n1331,
    n323,
    n597
  );


  xor
  g1942
  (
    n2015,
    n422,
    n616,
    n504,
    n499
  );


  or
  g1943
  (
    n2017,
    n1240,
    n1377,
    n675,
    n1206
  );


  xor
  g1944
  (
    n1883,
    n574,
    n242,
    n278,
    n261
  );


  nand
  g1945
  (
    n1622,
    n594,
    n429,
    n1268,
    n317
  );


  xnor
  g1946
  (
    n2128,
    n307,
    n385,
    n586,
    n309
  );


  xnor
  g1947
  (
    n1801,
    n565,
    n795,
    n528,
    n750
  );


  xnor
  g1948
  (
    n1762,
    n767,
    n416,
    n1200,
    n1378
  );


  nor
  g1949
  (
    n1891,
    n734,
    n474,
    n572,
    n578
  );


  xor
  g1950
  (
    n1853,
    n672,
    n1298,
    n279,
    n299
  );


  and
  g1951
  (
    n1638,
    n665,
    n404,
    n1284,
    n563
  );


  and
  g1952
  (
    n1775,
    n444,
    n443,
    n315,
    n1199
  );


  and
  g1953
  (
    n1772,
    n594,
    n580,
    n1391,
    n539
  );


  and
  g1954
  (
    n1646,
    n611,
    n753,
    n787,
    n521
  );


  nand
  g1955
  (
    n2209,
    n545,
    n338,
    n239,
    n1256
  );


  xor
  g1956
  (
    n1956,
    n556,
    n1341,
    n582,
    n1348
  );


  xnor
  g1957
  (
    n2168,
    n695,
    n479,
    n396,
    n1198
  );


  or
  g1958
  (
    n1691,
    n1290,
    n438,
    n305,
    n1189
  );


  xnor
  g1959
  (
    n1800,
    n276,
    n1311,
    n424,
    n333
  );


  nand
  g1960
  (
    n1657,
    n319,
    n1364,
    n1273,
    n1385
  );


  xnor
  g1961
  (
    n2033,
    n688,
    n633,
    n342,
    n237
  );


  nand
  g1962
  (
    n2138,
    n792,
    n1283,
    n373,
    n760
  );


  and
  g1963
  (
    n1888,
    n530,
    n331,
    n1375,
    n561
  );


  or
  g1964
  (
    n1807,
    n358,
    n716,
    n1336,
    n1303
  );


  xnor
  g1965
  (
    n2147,
    n1234,
    n370,
    n1365,
    n1171
  );


  or
  g1966
  (
    n1901,
    n678,
    n796,
    n355,
    n751
  );


  xnor
  g1967
  (
    n2183,
    n1191,
    n514,
    n502,
    n518
  );


  or
  g1968
  (
    n1788,
    n641,
    n458,
    n1389,
    n755
  );


  and
  g1969
  (
    n1566,
    n1221,
    n1337,
    n1259,
    n540
  );


  or
  g1970
  (
    n2057,
    n1226,
    n400,
    n762,
    n281
  );


  nand
  g1971
  (
    n1779,
    n631,
    n748,
    n544,
    n683
  );


  and
  g1972
  (
    n1954,
    n1307,
    n1309,
    n580,
    n680
  );


  xnor
  g1973
  (
    n1684,
    n1404,
    n1355,
    n527,
    n756
  );


  xnor
  g1974
  (
    n2006,
    n1309,
    n645,
    n1179,
    n1186
  );


  nand
  g1975
  (
    n1475,
    n391,
    n458,
    n1365,
    n666
  );


  xor
  g1976
  (
    n2002,
    n358,
    n303,
    n789,
    n705
  );


  or
  g1977
  (
    n1854,
    n1178,
    n1349,
    n414,
    n1165
  );


  or
  g1978
  (
    n1456,
    n288,
    n1173,
    n356,
    n736
  );


  nor
  g1979
  (
    n2229,
    n1166,
    n415,
    n233,
    n253
  );


  nor
  g1980
  (
    n1871,
    n1165,
    n243,
    n1293,
    n731
  );


  xnor
  g1981
  (
    n1846,
    n1351,
    n563,
    n311,
    n1194
  );


  nor
  g1982
  (
    n1438,
    n1322,
    n1201,
    n602,
    n1241
  );


  nor
  g1983
  (
    n2022,
    n727,
    n1323,
    n484,
    n497
  );


  xor
  g1984
  (
    n2108,
    n409,
    n558,
    n270,
    n574
  );


  xnor
  g1985
  (
    n1418,
    n533,
    n384,
    n1285,
    n622
  );


  xor
  g1986
  (
    KeyWire_0_20,
    n509,
    n774,
    n1226,
    n1404
  );


  xnor
  g1987
  (
    n2195,
    n406,
    n1302,
    n1189,
    n562
  );


  xnor
  g1988
  (
    n1660,
    n368,
    n395,
    n410,
    n587
  );


  and
  g1989
  (
    n1973,
    n530,
    n375,
    n576,
    n537
  );


  nor
  g1990
  (
    n1940,
    n763,
    n791,
    n1306,
    n420
  );


  nand
  g1991
  (
    n1539,
    n433,
    n1306,
    n1376,
    n655
  );


  or
  g1992
  (
    n2131,
    n329,
    n297,
    n786,
    n341
  );


  or
  g1993
  (
    n2241,
    n1253,
    n417,
    n250,
    n362
  );


  or
  g1994
  (
    n1764,
    n1232,
    n334,
    n437,
    n534
  );


  or
  g1995
  (
    n1570,
    n1412,
    n605,
    n699,
    n1270
  );


  and
  g1996
  (
    n1451,
    n267,
    n259,
    n460,
    n1405
  );


  xor
  g1997
  (
    n1484,
    n1254,
    n1378,
    n781,
    n417
  );


  nand
  g1998
  (
    n2214,
    n1317,
    n1263,
    n786,
    n1315
  );


  xor
  g1999
  (
    n1551,
    n1180,
    n306,
    n707,
    n1172
  );


  and
  g2000
  (
    n2182,
    n624,
    n592,
    n237,
    n424
  );


  nor
  g2001
  (
    n1928,
    n419,
    n1181,
    n443,
    n1264
  );


  nor
  g2002
  (
    n2163,
    n1245,
    n786,
    n1212,
    n1349
  );


  xor
  g2003
  (
    n1872,
    n468,
    n800,
    n380,
    n314
  );


  xnor
  g2004
  (
    n2198,
    n714,
    n255,
    n1201,
    n671
  );


  and
  g2005
  (
    n2172,
    n495,
    n1196,
    n580,
    n1280
  );


  nor
  g2006
  (
    n1629,
    n349,
    n444,
    n308,
    n710
  );


  nor
  g2007
  (
    n1873,
    n477,
    n516,
    n707,
    n1195
  );


  and
  g2008
  (
    n1664,
    n527,
    n630,
    n1180,
    n573
  );


  xnor
  g2009
  (
    n1630,
    n334,
    n1333,
    n319,
    n1235
  );


  and
  g2010
  (
    n2192,
    n469,
    n657,
    n1227,
    n1320
  );


  xor
  g2011
  (
    n1513,
    n386,
    n584,
    n588,
    n1344
  );


  and
  g2012
  (
    n1700,
    n728,
    n557,
    n745,
    n1278
  );


  xor
  g2013
  (
    n1541,
    n399,
    n1329,
    n704,
    n624
  );


  xor
  g2014
  (
    n1727,
    n515,
    n661,
    n367,
    n757
  );


  nand
  g2015
  (
    n1932,
    n1287,
    n335,
    n724,
    n1212
  );


  or
  g2016
  (
    n2059,
    n1285,
    n565,
    n570,
    n340
  );


  and
  g2017
  (
    n1571,
    n662,
    n1359,
    n1291,
    n1298
  );


  xnor
  g2018
  (
    n1967,
    n690,
    n624,
    n716,
    n666
  );


  or
  g2019
  (
    n1753,
    n1236,
    n249,
    n1322,
    n518
  );


  or
  g2020
  (
    n2118,
    n1248,
    n750,
    n411,
    n283
  );


  and
  g2021
  (
    n1509,
    n1279,
    n802,
    n357,
    n651
  );


  xnor
  g2022
  (
    n1649,
    n343,
    n589,
    n294,
    n1184
  );


  xnor
  g2023
  (
    n1448,
    n1270,
    n632,
    n392,
    n731
  );


  and
  g2024
  (
    n1676,
    n1341,
    n672,
    n281,
    n234
  );


  nor
  g2025
  (
    n2238,
    n1314,
    n313,
    n732,
    n674
  );


  nand
  g2026
  (
    n1843,
    n327,
    n735,
    n614,
    n738
  );


  and
  g2027
  (
    n2203,
    n1412,
    n388,
    n520,
    n664
  );


  nand
  g2028
  (
    n2099,
    n635,
    n1254,
    n721,
    n633
  );


  nor
  g2029
  (
    n1874,
    n1380,
    n693,
    n1209,
    n447
  );


  xor
  g2030
  (
    KeyWire_0_7,
    n527,
    n490,
    n383,
    n511
  );


  or
  g2031
  (
    n1585,
    n643,
    n778,
    n232,
    n512
  );


  nand
  g2032
  (
    n2068,
    n326,
    n1360,
    n1378,
    n404
  );


  nor
  g2033
  (
    n1950,
    n650,
    n575,
    n1327,
    n649
  );


  xnor
  g2034
  (
    n1435,
    n786,
    n1182,
    n332,
    n305
  );


  xor
  g2035
  (
    n1628,
    n408,
    n520,
    n547,
    n633
  );


  and
  g2036
  (
    n1460,
    n700,
    n544,
    n406,
    n1357
  );


  xor
  g2037
  (
    n1797,
    n713,
    n658,
    n318,
    n564
  );


  nand
  g2038
  (
    n1960,
    n449,
    n641,
    n329,
    n376
  );


  and
  g2039
  (
    n1688,
    n682,
    n603,
    n703,
    n1240
  );


  nand
  g2040
  (
    n1608,
    n784,
    n1176,
    n1337,
    n265
  );


  or
  g2041
  (
    n2043,
    n508,
    n325,
    n748
  );


  or
  g2042
  (
    n1449,
    n1383,
    n503,
    n615,
    n656
  );


  or
  g2043
  (
    n1927,
    n692,
    n679,
    n1169,
    n1416
  );


  nor
  g2044
  (
    n2242,
    n630,
    n664,
    n1372,
    n729
  );


  or
  g2045
  (
    n1829,
    n337,
    n1372,
    n485,
    n710
  );


  xor
  g2046
  (
    n2233,
    n254,
    n738,
    n409,
    n1395
  );


  and
  g2047
  (
    n1486,
    n631,
    n795,
    n1334,
    n505
  );


  xor
  g2048
  (
    n1645,
    n520,
    n421,
    n1373,
    n238
  );


  xor
  g2049
  (
    n1467,
    n446,
    n1172,
    n1203,
    n1363
  );


  or
  g2050
  (
    n2141,
    n648,
    n1406,
    n1275,
    n1304
  );


  nor
  g2051
  (
    n2112,
    n1361,
    n490,
    n591,
    n755
  );


  xor
  g2052
  (
    n1938,
    n1382,
    n1355,
    n1170,
    n264
  );


  or
  g2053
  (
    n2083,
    n662,
    n311,
    n775,
    n532
  );


  xor
  g2054
  (
    n2127,
    n322,
    n316,
    n1279,
    n1227
  );


  and
  g2055
  (
    n2011,
    n1276,
    n1269,
    n404,
    n1395
  );


  xor
  g2056
  (
    n1545,
    n241,
    n801,
    n804,
    n671
  );


  xor
  g2057
  (
    n1955,
    n463,
    n1312,
    n271,
    n387
  );


  xor
  g2058
  (
    n1909,
    n553,
    n694,
    n1216
  );


  xnor
  g2059
  (
    n1698,
    n702,
    n1320,
    n1227,
    n707
  );


  nand
  g2060
  (
    n1530,
    n280,
    n540,
    n454,
    n712
  );


  or
  g2061
  (
    n1745,
    n695,
    n1410,
    n1402,
    n613
  );


  nand
  g2062
  (
    n1730,
    n772,
    n267,
    n255,
    n727
  );


  xnor
  g2063
  (
    n2175,
    n1370,
    n1410,
    n760,
    n741
  );


  xnor
  g2064
  (
    n1535,
    n429,
    n1270,
    n521,
    n1371
  );


  nand
  g2065
  (
    n1470,
    n1254,
    n1408,
    n789,
    n606
  );


  and
  g2066
  (
    n2023,
    n766,
    n388,
    n335,
    n359
  );


  xnor
  g2067
  (
    n1777,
    n727,
    n388,
    n1311,
    n1163
  );


  nor
  g2068
  (
    n2136,
    n1183,
    n607,
    n460,
    n432
  );


  and
  g2069
  (
    n1900,
    n483,
    n1281,
    n1284,
    n1313
  );


  xnor
  g2070
  (
    n2010,
    n1408,
    n382,
    n788,
    n753
  );


  nand
  g2071
  (
    n1962,
    n381,
    n1202,
    n346,
    n548
  );


  nand
  g2072
  (
    n1506,
    n1386,
    n461,
    n368,
    n449
  );


  nand
  g2073
  (
    n1618,
    n277,
    n1332,
    n416,
    n430
  );


  or
  g2074
  (
    n1663,
    n924,
    n357,
    n1240,
    n468
  );


  nor
  g2075
  (
    n1433,
    n781,
    n1265,
    n414,
    n387
  );


  nor
  g2076
  (
    n1553,
    n1298,
    n1381,
    n1262,
    n635
  );


  xnor
  g2077
  (
    n2095,
    n533,
    n633,
    n1274,
    n489
  );


  xor
  g2078
  (
    n1479,
    n620,
    n332,
    n248,
    n756
  );


  nor
  g2079
  (
    n1483,
    n1176,
    n591,
    n1194,
    n732
  );


  nand
  g2080
  (
    n1860,
    n575,
    n685,
    n309,
    n306
  );


  nand
  g2081
  (
    n1939,
    n1212,
    n1174,
    n1162,
    n1400
  );


  or
  g2082
  (
    n1924,
    n600,
    n556,
    n1237,
    n264
  );


  xor
  g2083
  (
    n2109,
    n399,
    n1250,
    n1218
  );


  xor
  g2084
  (
    n2219,
    n1366,
    n397,
    n712,
    n1218
  );


  nand
  g2085
  (
    n1651,
    n263,
    n643,
    n508,
    n455
  );


  and
  g2086
  (
    n2239,
    n265,
    n699,
    n1190,
    n790
  );


  xor
  g2087
  (
    n2050,
    n740,
    n771,
    n264,
    n1393
  );


  nor
  g2088
  (
    n1670,
    n1224,
    n452,
    n635,
    n555
  );


  and
  g2089
  (
    n2120,
    n474,
    n690,
    n364,
    n257
  );


  nand
  g2090
  (
    n1536,
    n1216,
    n476,
    n467,
    n1386
  );


  nor
  g2091
  (
    n1542,
    n623,
    n543,
    n472,
    n667
  );


  or
  g2092
  (
    n1621,
    n672,
    n1308,
    n594,
    n414
  );


  xor
  g2093
  (
    n2156,
    n360,
    n648,
    n1383,
    n797
  );


  nand
  g2094
  (
    n2194,
    n636,
    n394,
    n727,
    n1379
  );


  nor
  g2095
  (
    n1671,
    n289,
    n254,
    n1311,
    n370
  );


  nand
  g2096
  (
    n1652,
    n440,
    n368,
    n426,
    n432
  );


  and
  g2097
  (
    n2048,
    n529,
    n367,
    n450,
    n596
  );


  xnor
  g2098
  (
    n2173,
    n1296,
    n480,
    n291,
    n770
  );


  xnor
  g2099
  (
    n1852,
    n647,
    n581,
    n1167,
    n1356
  );


  or
  g2100
  (
    n1695,
    n1195,
    n1221,
    n312,
    n1361
  );


  or
  g2101
  (
    n1420,
    n1174,
    n500,
    n307,
    n1344
  );


  nor
  g2102
  (
    n1469,
    n719,
    n291,
    n486,
    n725
  );


  xor
  g2103
  (
    n1644,
    n285,
    n422,
    n1316,
    n590
  );


  xnor
  g2104
  (
    n1716,
    n312,
    n288,
    n1238,
    n1237
  );


  xor
  g2105
  (
    n2123,
    n1208,
    n661,
    n445,
    n783
  );


  xor
  g2106
  (
    n1755,
    n1302,
    n459,
    n492,
    n1410
  );


  xnor
  g2107
  (
    n1746,
    n346,
    n602,
    n395,
    n353
  );


  or
  g2108
  (
    n2056,
    n783,
    n469,
    n671,
    n560
  );


  nor
  g2109
  (
    n1693,
    n673,
    n552,
    n240,
    n789
  );


  xnor
  g2110
  (
    n1689,
    n665,
    n426,
    n577,
    n359
  );


  xor
  g2111
  (
    n1686,
    n1415,
    n1262,
    n482,
    n1259
  );


  nand
  g2112
  (
    n2177,
    n507,
    n310,
    n351
  );


  nor
  g2113
  (
    n1537,
    n419,
    n1164,
    n872,
    n677
  );


  and
  g2114
  (
    n1489,
    n1176,
    n389,
    n541,
    n330
  );


  nor
  g2115
  (
    n1569,
    n257,
    n1270,
    n676,
    n338
  );


  and
  g2116
  (
    n1736,
    n645,
    n267,
    n1342,
    n367
  );


  xor
  g2117
  (
    n1980,
    n304,
    n1244,
    n300,
    n563
  );


  nand
  g2118
  (
    n2202,
    n280,
    n1305,
    n1188,
    n1272
  );


  or
  g2119
  (
    n1851,
    n251,
    n696,
    n1220,
    n510
  );


  and
  g2120
  (
    n1701,
    n671,
    n710,
    n486,
    n636
  );


  or
  g2121
  (
    n1508,
    n1371,
    n709,
    n425,
    n703
  );


  xnor
  g2122
  (
    n2005,
    n782,
    n759,
    n521,
    n1413
  );


  xnor
  g2123
  (
    n1597,
    n1318,
    n314,
    n490,
    n525
  );


  xnor
  g2124
  (
    n2162,
    n287,
    n366,
    n675,
    n1208
  );


  or
  g2125
  (
    n1574,
    n706,
    n353,
    n720,
    n634
  );


  and
  g2126
  (
    n1997,
    n304,
    n302,
    n233,
    n1353
  );


  nor
  g2127
  (
    n2060,
    n751,
    n1390,
    n1213,
    n721
  );


  xor
  g2128
  (
    n2197,
    n379,
    n1276,
    n307,
    n694
  );


  or
  g2129
  (
    n1737,
    n414,
    n1290,
    n503,
    n743
  );


  nand
  g2130
  (
    n1818,
    n718,
    n1252,
    n1260,
    n1410
  );


  or
  g2131
  (
    n2148,
    n238,
    n636,
    n1234,
    n1319
  );


  or
  g2132
  (
    n1517,
    n345,
    n1282,
    n282,
    n1357
  );


  xnor
  g2133
  (
    n1754,
    n441,
    n752,
    n505,
    n1390
  );


  xnor
  g2134
  (
    n1594,
    n621,
    n279,
    n687,
    n578
  );


  xor
  g2135
  (
    n1476,
    n269,
    n1328,
    n233,
    n797
  );


  nand
  g2136
  (
    n2196,
    n726,
    n684,
    n1242,
    n1350
  );


  nand
  g2137
  (
    n1981,
    n1184,
    n577,
    n618,
    n406
  );


  or
  g2138
  (
    n2204,
    n1238,
    n471,
    n503,
    n1230
  );


  or
  g2139
  (
    n1610,
    n353,
    n799,
    n542,
    n572
  );


  xor
  g2140
  (
    n1723,
    n734,
    n757,
    n554,
    n1296
  );


  or
  g2141
  (
    n1525,
    n730,
    n765,
    n596,
    n1360
  );


  or
  g2142
  (
    n2091,
    n1283,
    n1358,
    n1354,
    n1292
  );


  and
  g2143
  (
    n1656,
    n1385,
    n379,
    n298,
    n1405
  );


  xnor
  g2144
  (
    n2035,
    n1302,
    n764,
    n1304,
    n244
  );


  xor
  g2145
  (
    n1889,
    n570,
    n617,
    n1224,
    n1247
  );


  and
  g2146
  (
    n1964,
    n380,
    n1308,
    n1414,
    n793
  );


  nand
  g2147
  (
    n1562,
    n462,
    n1253,
    n1394,
    n408
  );


  nand
  g2148
  (
    n2160,
    n231,
    n719,
    n1189,
    n1302
  );


  xor
  g2149
  (
    n1771,
    n1263,
    n283,
    n377,
    n347
  );


  xnor
  g2150
  (
    n1678,
    n340,
    n1301,
    n240,
    n693
  );


  nor
  g2151
  (
    n1556,
    n1168,
    n458,
    n308,
    n263
  );


  xor
  g2152
  (
    n1586,
    n466,
    n555,
    n741,
    n446
  );


  nor
  g2153
  (
    n1731,
    n1372,
    n275,
    n767,
    n1203
  );


  nor
  g2154
  (
    n1725,
    n701,
    n523,
    n689,
    n488
  );


  or
  g2155
  (
    n2245,
    n551,
    n1186,
    n802,
    n488
  );


  and
  g2156
  (
    n1488,
    n306,
    n708,
    n1291,
    n569
  );


  xnor
  g2157
  (
    n2218,
    n1371,
    n1374,
    n459,
    n723
  );


  nand
  g2158
  (
    n1487,
    n766,
    n699,
    n491,
    n423
  );


  xor
  g2159
  (
    n1699,
    n1369,
    n608,
    n744,
    n1257
  );


  nand
  g2160
  (
    n1856,
    n1292,
    n747,
    n425,
    n757
  );


  xnor
  g2161
  (
    n1937,
    n1406,
    n449,
    n432,
    n548
  );


  and
  g2162
  (
    n1879,
    n657,
    n769,
    n526,
    n677
  );


  nand
  g2163
  (
    n1783,
    n459,
    n702,
    n478,
    n1198
  );


  nor
  g2164
  (
    n2144,
    n668,
    n1342,
    n632,
    n412
  );


  nor
  g2165
  (
    n1808,
    n535,
    n506,
    n748,
    n348
  );


  nor
  g2166
  (
    n1733,
    n1266,
    n259,
    n413,
    n1177
  );


  xnor
  g2167
  (
    n1573,
    n1223,
    n244,
    n662,
    n1283
  );


  nor
  g2168
  (
    n1692,
    n586,
    n1206,
    n1251,
    n257
  );


  or
  g2169
  (
    n1507,
    n1395,
    n1271,
    n1312,
    n591
  );


  or
  g2170
  (
    n1979,
    n407,
    n1373,
    n328,
    n552
  );


  and
  g2171
  (
    n1478,
    n619,
    n408,
    n646,
    n779
  );


  and
  g2172
  (
    n1942,
    n442,
    n1248,
    n697,
    n764
  );


  and
  g2173
  (
    n2021,
    n244,
    n582,
    n726,
    n1347
  );


  or
  g2174
  (
    n2063,
    n1389,
    n284,
    n351,
    n1194
  );


  xnor
  g2175
  (
    n1440,
    n401,
    n300,
    n533,
    n615
  );


  or
  g2176
  (
    n1516,
    n1192,
    n794,
    n431,
    n1361
  );


  nor
  g2177
  (
    n1904,
    n1369,
    n477,
    n320,
    n273
  );


  and
  g2178
  (
    n2152,
    n741,
    n354,
    n339,
    n1391
  );


  xor
  g2179
  (
    n1974,
    n1249,
    n712,
    n1300,
    n483
  );


  nand
  g2180
  (
    n1529,
    n1384,
    n777,
    n399,
    n534
  );


  xor
  g2181
  (
    n1619,
    n375,
    n350,
    n677,
    n649
  );


  xor
  g2182
  (
    n1717,
    n674,
    n803,
    n1409,
    n1326
  );


  xor
  g2183
  (
    n2115,
    n250,
    n1295,
    n386,
    n1373
  );


  xor
  g2184
  (
    n1482,
    n1345,
    n1263,
    n1192,
    n1231
  );


  nor
  g2185
  (
    n1875,
    n1414,
    n677,
    n1294,
    n794
  );


  xnor
  g2186
  (
    n1616,
    n1241,
    n767,
    n411,
    n265
  );


  and
  g2187
  (
    n1454,
    n296,
    n316,
    n1304,
    n797
  );


  or
  g2188
  (
    n2180,
    n519,
    n484,
    n1402,
    n1356
  );


  xor
  g2189
  (
    n1447,
    n606,
    n554,
    n424,
    n321
  );


  and
  g2190
  (
    n1459,
    n431,
    n416,
    n430,
    n674
  );


  nor
  g2191
  (
    n1832,
    n598,
    n628,
    n1405,
    n803
  );


  xnor
  g2192
  (
    n1633,
    n760,
    n1402,
    n1346,
    n1203
  );


  nand
  g2193
  (
    n2070,
    n369,
    n659,
    n1389,
    n506
  );


  xor
  g2194
  (
    n2187,
    n756,
    n1231,
    n1251,
    n589
  );


  xor
  g2195
  (
    n1761,
    n598,
    n282,
    n1352,
    n746
  );


  nor
  g2196
  (
    n1735,
    n312,
    n401,
    n405,
    n457
  );


  nand
  g2197
  (
    n1887,
    n711,
    n293,
    n403,
    n357
  );


  xor
  g2198
  (
    n2161,
    n698,
    n758,
    n1275,
    n1266
  );


  xnor
  g2199
  (
    n1724,
    n458,
    n1376,
    n480,
    n303
  );


  nor
  g2200
  (
    n1607,
    n737,
    n538,
    n743,
    n236
  );


  and
  g2201
  (
    n2105,
    n1193,
    n269,
    n262,
    n576
  );


  nand
  g2202
  (
    n1520,
    n1406,
    n649,
    n392,
    n550
  );


  or
  g2203
  (
    n2421,
    n2104,
    n1495,
    n1747,
    n2071
  );


  and
  g2204
  (
    n2451,
    n2081,
    n1501,
    n1704,
    n1433
  );


  or
  g2205
  (
    n2288,
    n1936,
    n1891,
    n2091,
    n2227
  );


  and
  g2206
  (
    n2298,
    n2012,
    n1718,
    n2222,
    n1825
  );


  xnor
  g2207
  (
    n2377,
    n1550,
    n2028,
    n1442,
    n1448
  );


  or
  g2208
  (
    n2440,
    n1693,
    n1795,
    n2230,
    n1672
  );


  and
  g2209
  (
    n2386,
    n1881,
    n1549,
    n2168,
    n2148
  );


  and
  g2210
  (
    n2268,
    n1450,
    n1451,
    n2120,
    n1979
  );


  nand
  g2211
  (
    n2318,
    n2080,
    n1768,
    n1711,
    n1972
  );


  nand
  g2212
  (
    n2394,
    n1681,
    n1909,
    n1680,
    n1830
  );


  xnor
  g2213
  (
    n2380,
    n2201,
    n1560,
    n1749,
    n1797
  );


  and
  g2214
  (
    n2427,
    n1705,
    n2037,
    n2161,
    n1806
  );


  nand
  g2215
  (
    n2343,
    n2233,
    n1659,
    n2180,
    n2149
  );


  xnor
  g2216
  (
    n2338,
    n1484,
    n1742,
    n2049,
    n1883
  );


  or
  g2217
  (
    n2374,
    n2139,
    n2239,
    n1842,
    n1476
  );


  xor
  g2218
  (
    n2247,
    n2066,
    n1460,
    n2034,
    n1733
  );


  nor
  g2219
  (
    n2415,
    n1843,
    n2153,
    n1618,
    n1464
  );


  and
  g2220
  (
    n2317,
    n2185,
    n1669,
    n1922,
    n2134
  );


  nor
  g2221
  (
    n2357,
    n1572,
    n2062,
    n1939,
    n1973
  );


  xor
  g2222
  (
    n2341,
    n1430,
    n1773,
    n1639,
    n1521
  );


  nor
  g2223
  (
    n2365,
    n1631,
    n1661,
    n2099,
    n1919
  );


  xnor
  g2224
  (
    n2311,
    n1528,
    n2061,
    n1697,
    n1997
  );


  nor
  g2225
  (
    n2324,
    n1757,
    n1911,
    n1569,
    n1895
  );


  or
  g2226
  (
    n2260,
    n2205,
    n1422,
    n1581,
    n1703
  );


  xnor
  g2227
  (
    n2414,
    n1860,
    n1723,
    n1850,
    n1709
  );


  xnor
  g2228
  (
    n2340,
    n1579,
    n1473,
    n1898,
    n1905
  );


  xor
  g2229
  (
    n2301,
    n1966,
    n1882,
    n1421,
    n2110
  );


  or
  g2230
  (
    n2356,
    n1533,
    n2242,
    n1598,
    n1727
  );


  xor
  g2231
  (
    n2399,
    n2084,
    n2143,
    n1957,
    n1548
  );


  xnor
  g2232
  (
    n2306,
    n1621,
    n1991,
    n1947,
    n1531
  );


  nand
  g2233
  (
    n2335,
    n1760,
    n1525,
    n1457,
    n1461
  );


  xnor
  g2234
  (
    n2334,
    n1417,
    n1506,
    n1468,
    n1852
  );


  xor
  g2235
  (
    n2291,
    n1959,
    n1726,
    n1804,
    n1950
  );


  or
  g2236
  (
    n2253,
    n1761,
    n1846,
    n1787,
    n1910
  );


  or
  g2237
  (
    n2350,
    n1876,
    n1532,
    n2109,
    n1519
  );


  xnor
  g2238
  (
    n2434,
    n1914,
    n2232,
    n1724,
    n2141
  );


  nand
  g2239
  (
    n2275,
    n1559,
    n1839,
    n2237,
    n2070
  );


  nand
  g2240
  (
    n2259,
    n2125,
    n1964,
    n1491,
    n1644
  );


  nor
  g2241
  (
    n2331,
    n2171,
    n1613,
    n1729,
    n2164
  );


  xor
  g2242
  (
    n2269,
    n1682,
    n2234,
    n2094,
    n1676
  );


  or
  g2243
  (
    n2349,
    n2165,
    n2076,
    n2221,
    n1740
  );


  nand
  g2244
  (
    n2397,
    n1918,
    n1447,
    n1938,
    n1739
  );


  nand
  g2245
  (
    n2403,
    n1632,
    n1574,
    n1624,
    n2032
  );


  or
  g2246
  (
    n2367,
    n2188,
    n1670,
    n2000,
    n1971
  );


  xor
  g2247
  (
    n2408,
    n1609,
    n2063,
    n1791,
    n1529
  );


  nor
  g2248
  (
    n2267,
    n2112,
    n1755,
    n2123,
    n1636
  );


  and
  g2249
  (
    n2308,
    n1566,
    n1823,
    n1954,
    n1833
  );


  or
  g2250
  (
    n2299,
    n1419,
    n1463,
    n2052,
    n2025
  );


  nor
  g2251
  (
    n2373,
    n2008,
    n1418,
    n1597,
    n2095
  );


  and
  g2252
  (
    n2292,
    n1786,
    n2046,
    n1553,
    n1503
  );


  xnor
  g2253
  (
    n2326,
    n1832,
    n1958,
    n1874,
    n1878
  );


  nor
  g2254
  (
    n2336,
    n1673,
    n1625,
    n1805,
    n1487
  );


  nor
  g2255
  (
    n2430,
    n1831,
    n2044,
    n1445,
    n1828
  );


  nor
  g2256
  (
    n2426,
    n1486,
    n2051,
    n2213,
    n1858
  );


  and
  g2257
  (
    n2333,
    n2131,
    n1662,
    n2086,
    n1523
  );


  xnor
  g2258
  (
    n2453,
    n1552,
    n1668,
    n1993,
    n1746
  );


  nor
  g2259
  (
    n2354,
    n2097,
    n2077,
    n1822,
    n2017
  );


  xnor
  g2260
  (
    n2450,
    n1836,
    n2007,
    n1431,
    n1745
  );


  and
  g2261
  (
    n2363,
    n2079,
    n1984,
    n1810,
    n1462
  );


  nand
  g2262
  (
    n2274,
    n2218,
    n1968,
    n2231,
    n1738
  );


  and
  g2263
  (
    n2346,
    n1801,
    n1960,
    n1873,
    n1758
  );


  xor
  g2264
  (
    n2378,
    n1542,
    n2181,
    n1998,
    n1944
  );


  nand
  g2265
  (
    n2328,
    n1666,
    n1556,
    n1942,
    n1816
  );


  or
  g2266
  (
    n2413,
    n2029,
    n1443,
    n2121,
    n2105
  );


  nand
  g2267
  (
    n2360,
    n1837,
    n1627,
    n1584,
    n1427
  );


  nand
  g2268
  (
    n2446,
    n1485,
    n2050,
    n1776,
    n1808
  );


  nor
  g2269
  (
    n2417,
    n1508,
    n2156,
    n1517,
    n2127
  );


  and
  g2270
  (
    n2284,
    n1880,
    n1453,
    n1907,
    n1647
  );


  xor
  g2271
  (
    n2422,
    n2238,
    n2116,
    n1896,
    n2130
  );


  xor
  g2272
  (
    n2303,
    n2190,
    n2219,
    n1886,
    n2096
  );


  or
  g2273
  (
    n2352,
    n1985,
    n1527,
    n2136,
    n1685
  );


  and
  g2274
  (
    n2401,
    n1558,
    n1561,
    n1737,
    n1425
  );


  and
  g2275
  (
    n2437,
    n2144,
    n1965,
    n2193,
    n1466
  );


  xor
  g2276
  (
    n2270,
    n1782,
    n2223,
    n1641,
    n1573
  );


  xnor
  g2277
  (
    n2390,
    n1712,
    n1921,
    n1765,
    n2151
  );


  nand
  g2278
  (
    n2278,
    n1688,
    n1638,
    n1847,
    n2011
  );


  nand
  g2279
  (
    n2432,
    n1507,
    n2147,
    n1477,
    n2005
  );


  nor
  g2280
  (
    n2258,
    n1877,
    n2245,
    n1988,
    n2220
  );


  xnor
  g2281
  (
    n2264,
    n2137,
    n1777,
    n1892,
    n1720
  );


  or
  g2282
  (
    n2280,
    n2192,
    n1975,
    n1820,
    n1580
  );


  xnor
  g2283
  (
    n2364,
    n2191,
    n1596,
    n2009,
    n1934
  );


  xnor
  g2284
  (
    n2348,
    n2014,
    n1494,
    n1920,
    n2159
  );


  nor
  g2285
  (
    n2254,
    n1577,
    n1623,
    n2196,
    n1626
  );


  and
  g2286
  (
    n2402,
    n1854,
    n2073,
    n1793,
    n2236
  );


  nor
  g2287
  (
    n2418,
    n1915,
    n2047,
    n1935,
    n1840
  );


  and
  g2288
  (
    n2307,
    n1595,
    n2207,
    n2224,
    n1518
  );


  and
  g2289
  (
    n2314,
    n1994,
    n1715,
    n2113,
    n1535
  );


  nor
  g2290
  (
    n2263,
    n1562,
    n1949,
    n1483,
    n1769
  );


  xor
  g2291
  (
    n2392,
    n2111,
    n1730,
    n1452,
    n2152
  );


  or
  g2292
  (
    n2250,
    n1812,
    n1498,
    n1774,
    n2026
  );


  nor
  g2293
  (
    n2358,
    n2182,
    n2067,
    n2118,
    n2027
  );


  xnor
  g2294
  (
    n2294,
    n1589,
    n1611,
    n1952,
    n2035
  );


  xnor
  g2295
  (
    n2375,
    n2078,
    n1894,
    n1783,
    n2200
  );


  nand
  g2296
  (
    n2290,
    n2226,
    n1570,
    n1744,
    n2179
  );


  and
  g2297
  (
    n2329,
    n2101,
    n1701,
    n1827,
    n1983
  );


  xnor
  g2298
  (
    n2411,
    n1862,
    n2064,
    n1931,
    n1937
  );


  and
  g2299
  (
    n2286,
    n2176,
    n2146,
    n1456,
    n2128
  );


  or
  g2300
  (
    n2345,
    n2021,
    n1864,
    n1591,
    n2040
  );


  xnor
  g2301
  (
    n2406,
    n2235,
    n2169,
    n1824,
    n1478
  );


  nand
  g2302
  (
    n2257,
    n1978,
    n2010,
    n1721,
    n1696
  );


  xnor
  g2303
  (
    n2289,
    n1586,
    n2054,
    n2177,
    n1665
  );


  xor
  g2304
  (
    n2381,
    n1629,
    n1593,
    n1619,
    n1516
  );


  and
  g2305
  (
    n2293,
    n1674,
    n2170,
    n2060,
    n1515
  );


  xor
  g2306
  (
    n2305,
    n1520,
    n1995,
    n1926,
    n2114
  );


  or
  g2307
  (
    n2441,
    n1587,
    n2003,
    n1564,
    n2175
  );


  or
  g2308
  (
    n2315,
    n1510,
    n1754,
    n1502,
    n2098
  );


  or
  g2309
  (
    n2319,
    n1505,
    n1449,
    n2041,
    n1655
  );


  nand
  g2310
  (
    n2320,
    n1480,
    n1764,
    n2015,
    n2155
  );


  nand
  g2311
  (
    n2423,
    n1557,
    n2115,
    n2085,
    n1440
  );


  xor
  g2312
  (
    n2276,
    n1699,
    n1605,
    n2173,
    n2088
  );


  xor
  g2313
  (
    n2266,
    n2199,
    n2001,
    n2216,
    n1635
  );


  and
  g2314
  (
    n2419,
    n1467,
    n2106,
    n1690,
    n2194
  );


  nor
  g2315
  (
    n2273,
    n2195,
    n2133,
    n1594,
    n1677
  );


  nor
  g2316
  (
    n2447,
    n1536,
    n1775,
    n1992,
    n1790
  );


  and
  g2317
  (
    n2252,
    n2172,
    n1436,
    n2150,
    n1838
  );


  or
  g2318
  (
    n2282,
    n1772,
    n1683,
    n1945,
    n1731
  );


  nand
  g2319
  (
    n2310,
    n1818,
    n1526,
    n2023,
    n1599
  );


  nand
  g2320
  (
    n2435,
    n1617,
    n1756,
    n1785,
    n1853
  );


  and
  g2321
  (
    n2454,
    n1702,
    n1809,
    n1667,
    n1490
  );


  xor
  g2322
  (
    n2316,
    n1807,
    n2024,
    n2187,
    n1735
  );


  and
  g2323
  (
    n2428,
    n1555,
    n1469,
    n2208,
    n1689
  );


  and
  g2324
  (
    n2251,
    n1612,
    n1637,
    n1863,
    n1439
  );


  and
  g2325
  (
    n2366,
    n1465,
    n2004,
    n1645,
    n1879
  );


  nand
  g2326
  (
    n2353,
    n2198,
    n1725,
    n1575,
    n1567
  );


  or
  g2327
  (
    n2404,
    n1770,
    n1496,
    n1967,
    n2048
  );


  and
  g2328
  (
    n2372,
    n1524,
    n2163,
    n1796,
    n1622
  );


  and
  g2329
  (
    n2379,
    n1590,
    n1541,
    n1663,
    n1424
  );


  xor
  g2330
  (
    n2265,
    n2006,
    n2240,
    n2033,
    n2074
  );


  xnor
  g2331
  (
    n2439,
    n1426,
    n1779,
    n1458,
    n1472
  );


  xnor
  g2332
  (
    n2433,
    n1976,
    n1800,
    n1766,
    n1819
  );


  xor
  g2333
  (
    n2261,
    n2056,
    n1870,
    n1885,
    n1813
  );


  and
  g2334
  (
    n2285,
    n2092,
    n1522,
    n1961,
    n1927
  );


  nand
  g2335
  (
    n2442,
    n1530,
    n1716,
    n1930,
    n1642
  );


  or
  g2336
  (
    n2304,
    n1649,
    n2142,
    n1719,
    n1736
  );


  xnor
  g2337
  (
    n2322,
    n2158,
    n1455,
    n1859,
    n1488
  );


  and
  g2338
  (
    n2389,
    n2117,
    n2202,
    n1946,
    n1955
  );


  xnor
  g2339
  (
    n2416,
    n1887,
    n1454,
    n1576,
    n1653
  );


  and
  g2340
  (
    n2271,
    n1545,
    n1759,
    n1763,
    n1817
  );


  xnor
  g2341
  (
    n2420,
    n1551,
    n1788,
    n1648,
    n1534
  );


  or
  g2342
  (
    n2339,
    n2089,
    n1861,
    n2055,
    n2167
  );


  nor
  g2343
  (
    n2384,
    n2135,
    n1694,
    n1750,
    n2038
  );


  nand
  g2344
  (
    n2391,
    n1607,
    n1728,
    n1875,
    n1658
  );


  and
  g2345
  (
    n2309,
    n1592,
    n1657,
    n2211,
    n2039
  );


  xor
  g2346
  (
    n2409,
    n1671,
    n1844,
    n1434,
    n1933
  );


  xor
  g2347
  (
    n2277,
    n1511,
    n1743,
    n1432,
    n1514
  );


  nor
  g2348
  (
    n2393,
    n1789,
    n1714,
    n1923,
    n2068
  );


  xor
  g2349
  (
    n2296,
    n1568,
    n1849,
    n1482,
    n1640
  );


  or
  g2350
  (
    n2287,
    n1428,
    n1856,
    n1459,
    n2072
  );


  or
  g2351
  (
    n2351,
    n1996,
    n1416,
    n1493,
    n1601
  );


  xor
  g2352
  (
    n2387,
    n1571,
    n1913,
    n1734,
    n1908
  );


  xor
  g2353
  (
    n2256,
    n1794,
    n2184,
    n2083,
    n2100
  );


  and
  g2354
  (
    n2395,
    n1684,
    n1980,
    n1940,
    n1604
  );


  nand
  g2355
  (
    n2410,
    n2087,
    n2036,
    n2197,
    n1916
  );


  and
  g2356
  (
    n2369,
    n1500,
    n2204,
    n1540,
    n1799
  );


  nor
  g2357
  (
    n2443,
    n1539,
    n1474,
    n2178,
    n1928
  );


  and
  g2358
  (
    n2449,
    n1829,
    n1634,
    n1437,
    n1977
  );


  xor
  g2359
  (
    n2248,
    n1479,
    n1811,
    n1563,
    n1509
  );


  xnor
  g2360
  (
    n2396,
    n1943,
    n1513,
    n2145,
    n1708
  );


  xnor
  g2361
  (
    n2376,
    n2108,
    n1646,
    n1948,
    n1780
  );


  xor
  g2362
  (
    n2444,
    n1792,
    n1962,
    n1504,
    n1546
  );


  xor
  g2363
  (
    n2400,
    n1585,
    n2162,
    n1565,
    n2102
  );


  nor
  g2364
  (
    n2337,
    n1707,
    n1986,
    n1578,
    n1969
  );


  xnor
  g2365
  (
    n2342,
    n1470,
    n2042,
    n1687,
    n1679
  );


  nand
  g2366
  (
    n2362,
    n2210,
    n2174,
    n2019,
    n2246
  );


  or
  g2367
  (
    n2262,
    n1990,
    n2122,
    n1722,
    n1767
  );


  nor
  g2368
  (
    n2359,
    n2206,
    n1497,
    n1956,
    n1651
  );


  and
  g2369
  (
    n2300,
    n1695,
    n1848,
    n2229,
    n1872
  );


  or
  g2370
  (
    n2436,
    n1554,
    n1845,
    n2043,
    n2228
  );


  or
  g2371
  (
    n2370,
    n2082,
    n2138,
    n1803,
    n2160
  );


  or
  g2372
  (
    n2302,
    n1987,
    n1989,
    n1429,
    n1741
  );


  xor
  g2373
  (
    n2297,
    n2140,
    n1981,
    n1678,
    n1492
  );


  and
  g2374
  (
    n2452,
    n1999,
    n1929,
    n1932,
    n1798
  );


  or
  g2375
  (
    n2330,
    n1826,
    n1675,
    n1686,
    n1691
  );


  and
  g2376
  (
    n2249,
    n1435,
    n1700,
    n2093,
    n1710
  );


  xor
  g2377
  (
    n2424,
    n2225,
    n1481,
    n2215,
    n1851
  );


  nand
  g2378
  (
    n2368,
    n2057,
    n1974,
    n2183,
    n1899
  );


  nor
  g2379
  (
    n2295,
    n1441,
    n1614,
    n2107,
    n1692
  );


  xor
  g2380
  (
    n2383,
    n1925,
    n1628,
    n2090,
    n2030
  );


  and
  g2381
  (
    n2361,
    n2053,
    n1888,
    n1543,
    n1753
  );


  or
  g2382
  (
    n2431,
    n1698,
    n1778,
    n1784,
    n1857
  );


  xor
  g2383
  (
    n2283,
    n1732,
    n1871,
    n2244,
    n1970
  );


  xnor
  g2384
  (
    n2405,
    n2241,
    n1583,
    n2186,
    n1855
  );


  xnor
  g2385
  (
    n2255,
    n2119,
    n2157,
    n1633,
    n1781
  );


  and
  g2386
  (
    n2312,
    n1953,
    n1475,
    n2065,
    n1902
  );


  xor
  g2387
  (
    n2347,
    n1901,
    n1834,
    n1537,
    n2075
  );


  and
  g2388
  (
    n2448,
    n2059,
    n1752,
    n1762,
    n1751
  );


  xnor
  g2389
  (
    n2371,
    n2124,
    n1868,
    n1664,
    n1650
  );


  nand
  g2390
  (
    n2281,
    n2031,
    n2209,
    n1444,
    n1717
  );


  and
  g2391
  (
    n2313,
    n1420,
    n2020,
    n1660,
    n1643
  );


  nand
  g2392
  (
    n2388,
    n1602,
    n1630,
    n1924,
    n1656
  );


  or
  g2393
  (
    n2445,
    n2189,
    n2103,
    n1771,
    n1904
  );


  nand
  g2394
  (
    n2355,
    n1603,
    n1821,
    n2212,
    n2132
  );


  xnor
  g2395
  (
    n2279,
    n1893,
    n1610,
    n1582,
    n2016
  );


  or
  g2396
  (
    n2398,
    n1941,
    n1866,
    n1423,
    n2058
  );


  nand
  g2397
  (
    n2344,
    n2045,
    n1713,
    n1917,
    n1489
  );


  nand
  g2398
  (
    n2385,
    n2069,
    n1865,
    n1903,
    n1814
  );


  or
  g2399
  (
    n2438,
    n1471,
    n1802,
    n1544,
    n1869
  );


  or
  g2400
  (
    n2382,
    n2126,
    n1841,
    n1900,
    n1600
  );


  and
  g2401
  (
    n2407,
    n1512,
    n1446,
    n2217,
    n1815
  );


  nand
  g2402
  (
    n2272,
    n1963,
    n1652,
    n1615,
    n2243
  );


  or
  g2403
  (
    n2429,
    n2022,
    n1706,
    n1897,
    n1438
  );


  nor
  g2404
  (
    n2321,
    n2203,
    n1835,
    n1538,
    n1620
  );


  nor
  g2405
  (
    n2332,
    n2166,
    n2002,
    n1906,
    n1889
  );


  nand
  g2406
  (
    n2412,
    n1982,
    n1608,
    n1912,
    n1951
  );


  nand
  g2407
  (
    n2425,
    n1867,
    n1547,
    n1416,
    n1499
  );


  nand
  g2408
  (
    n2323,
    n1616,
    n1890,
    n1884,
    n2154
  );


  or
  g2409
  (
    n2325,
    n1748,
    n2129,
    n1654,
    n1588
  );


  and
  g2410
  (
    n2327,
    n2013,
    n1606,
    n2018,
    n2214
  );


  xnor
  g2411
  (
    n2463,
    n2430,
    n2384,
    n2453,
    n2390
  );


  xnor
  g2412
  (
    n2464,
    n2334,
    n2447,
    n2364,
    n2427
  );


  xnor
  g2413
  (
    n2470,
    n2389,
    n2416,
    n2325,
    n2284
  );


  xor
  g2414
  (
    n2491,
    n2265,
    n2396,
    n2286,
    n2315
  );


  nand
  g2415
  (
    n2468,
    n2436,
    n2412,
    n2339,
    n2332
  );


  xor
  g2416
  (
    n2504,
    n2279,
    n2318,
    n2363,
    n2402
  );


  xor
  g2417
  (
    n2494,
    n2357,
    n2401,
    n2276,
    n2314
  );


  or
  g2418
  (
    n2493,
    n2309,
    n2285,
    n2330,
    n2264
  );


  xor
  g2419
  (
    n2473,
    n2410,
    n2373,
    n2277,
    n2352
  );


  nor
  g2420
  (
    n2476,
    n2391,
    n2441,
    n2261,
    n2299
  );


  xnor
  g2421
  (
    n2498,
    n2429,
    n2421,
    n2405,
    n2249
  );


  and
  g2422
  (
    n2455,
    n2298,
    n2404,
    n2392,
    n2250
  );


  xor
  g2423
  (
    n2474,
    n2440,
    n2452,
    n2362,
    n2375
  );


  nand
  g2424
  (
    n2502,
    n2344,
    n2377,
    n2259,
    n2293
  );


  xor
  g2425
  (
    n2503,
    n2247,
    n2454,
    n2303,
    n2443
  );


  or
  g2426
  (
    n2456,
    n2327,
    n2371,
    n2345,
    n2413
  );


  or
  g2427
  (
    n2469,
    n2423,
    n2320,
    n2350,
    n2400
  );


  nand
  g2428
  (
    n2489,
    n2358,
    n2305,
    n2346,
    n2267
  );


  nand
  g2429
  (
    n2495,
    n2269,
    n2317,
    n2349,
    n2343
  );


  xor
  g2430
  (
    n2465,
    n2354,
    n2415,
    n2382,
    n2256
  );


  xor
  g2431
  (
    n2457,
    n2433,
    n2395,
    n2383,
    n2329
  );


  nand
  g2432
  (
    n2461,
    n2281,
    n2380,
    n2434,
    n2424
  );


  or
  g2433
  (
    n2482,
    n2272,
    n2426,
    n2310,
    n2355
  );


  or
  g2434
  (
    n2462,
    n2356,
    n2406,
    n2294,
    n2425
  );


  nand
  g2435
  (
    n2505,
    n2291,
    n2365,
    n2326,
    n2445
  );


  nor
  g2436
  (
    n2501,
    n2278,
    n2268,
    n2372,
    n2283
  );


  nand
  g2437
  (
    n2497,
    n2255,
    n2311,
    n2258,
    n2398
  );


  nand
  g2438
  (
    n2478,
    n2342,
    n2446,
    n2316,
    n2409
  );


  nand
  g2439
  (
    n2466,
    n2335,
    n2351,
    n2399,
    n2312
  );


  and
  g2440
  (
    n2458,
    n2451,
    n2386,
    n2417,
    n2428
  );


  and
  g2441
  (
    KeyWire_0_31,
    n2266,
    n2324,
    n2381,
    n2275
  );


  xnor
  g2442
  (
    n2506,
    n2308,
    n2388,
    n2418,
    n2397
  );


  or
  g2443
  (
    n2479,
    n2302,
    n2360,
    n2270,
    n2288
  );


  xnor
  g2444
  (
    n2481,
    n2439,
    n2422,
    n2368,
    n2376
  );


  nand
  g2445
  (
    n2477,
    n2257,
    n2338,
    n2319,
    n2271
  );


  nand
  g2446
  (
    n2471,
    n2251,
    n2419,
    n2379,
    n2292
  );


  and
  g2447
  (
    KeyWire_0_18,
    n2378,
    n2273,
    n2297,
    n2304
  );


  or
  g2448
  (
    n2459,
    n2359,
    n2387,
    n2313,
    n2322
  );


  nor
  g2449
  (
    n2487,
    n2323,
    n2274,
    n2337,
    n2254
  );


  xor
  g2450
  (
    n2483,
    n2393,
    n2248,
    n2448,
    n2262
  );


  or
  g2451
  (
    n2499,
    n2385,
    n2403,
    n2260,
    n2321
  );


  xnor
  g2452
  (
    n2492,
    n2301,
    n2366,
    n2300,
    n2253
  );


  nand
  g2453
  (
    n2480,
    n2289,
    n2328,
    n2374,
    n2336
  );


  xnor
  g2454
  (
    n2496,
    n2414,
    n2367,
    n2408,
    n2280
  );


  xor
  g2455
  (
    n2475,
    n2435,
    n2407,
    n2290,
    n2394
  );


  nor
  g2456
  (
    n2486,
    n2444,
    n2361,
    n2370,
    n2411
  );


  xor
  g2457
  (
    n2467,
    n2287,
    n2442,
    n2449,
    n2340
  );


  xnor
  g2458
  (
    n2484,
    n2295,
    n2307,
    n2282,
    n2306
  );


  or
  g2459
  (
    n2490,
    n2347,
    n2353,
    n2431,
    n2450
  );


  or
  g2460
  (
    KeyWire_0_19,
    n2420,
    n2296,
    n2331,
    n2263
  );


  and
  g2461
  (
    n2500,
    n2333,
    n2432,
    n2348,
    n2252
  );


  xor
  g2462
  (
    n2460,
    n2437,
    n2341,
    n2369,
    n2438
  );


  nor
  g2463
  (
    n2518,
    n2505,
    n2501,
    n2485,
    n2484
  );


  nor
  g2464
  (
    KeyWire_0_2,
    n2466,
    n2486,
    n2456,
    n2477
  );


  nor
  g2465
  (
    n2516,
    n2494,
    n2504,
    n2461,
    n2503
  );


  or
  g2466
  (
    n2507,
    n2462,
    n2467,
    n2495,
    n2460
  );


  xnor
  g2467
  (
    n2511,
    n2488,
    n2491,
    n2500,
    n2468
  );


  nand
  g2468
  (
    n2513,
    n2465,
    n2472,
    n2497,
    n2499
  );


  nand
  g2469
  (
    n2514,
    n2469,
    n2459,
    n2481,
    n2483
  );


  nor
  g2470
  (
    n2512,
    n2458,
    n2478,
    n2463,
    n2476
  );


  nor
  g2471
  (
    n2509,
    n2480,
    n2490,
    n2464,
    n2489
  );


  xor
  g2472
  (
    n2510,
    n2496,
    n2457,
    n2502,
    n2493
  );


  or
  g2473
  (
    n2515,
    n2471,
    n2487,
    n2498,
    n2475
  );


  xnor
  g2474
  (
    n2508,
    n2482,
    n2506,
    n2470,
    n2492
  );


  or
  g2475
  (
    n2517,
    n2479,
    n2474,
    n2473,
    n2455
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n786,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n310,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n2519,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1966,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1648,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n225,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n2062,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1550,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1975,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n654,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n802,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n691,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n50,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n356,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1881,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n1342,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n829,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1620,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n2472,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n2488,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1655,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1090,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1272,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1029,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n382,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n2078,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n2142,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1424,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n2126,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n68,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1906,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n2485,
    KeyNOTWire_0_31
  );


endmodule

