// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_410 written by SynthGen on 2021/04/05 11:08:36
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_410 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n111, n106, n124, n110, n104, n132, n129, n125,
 n118, n119, n121, n108, n102, n109, n115, n112,
 n130, n123, n128, n101, n120, n131, n107, n103,
 n113, n117, n122, n126, n116, n105, n114, n127);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n111, n106, n124, n110, n104, n132, n129, n125,
 n118, n119, n121, n108, n102, n109, n115, n112,
 n130, n123, n128, n101, n120, n131, n107, n103,
 n113, n117, n122, n126, n116, n105, n114, n127;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

buf  g0 (n37, n1);
buf  g1 (n34, n2);
buf  g2 (n35, n2);
buf  g3 (n33, n1);
buf  g4 (n36, n1);
buf  g5 (n40, n34);
not  g6 (n56, n37);
buf  g7 (n49, n34);
buf  g8 (n50, n34);
buf  g9 (n53, n35);
not  g10 (n46, n33);
not  g11 (n55, n36);
buf  g12 (n44, n35);
not  g13 (n52, n35);
buf  g14 (n42, n33);
buf  g15 (n48, n37);
buf  g16 (n54, n36);
buf  g17 (n45, n36);
not  g18 (n41, n36);
buf  g19 (n39, n34);
not  g20 (n51, n37);
buf  g21 (n38, n35);
buf  g22 (n43, n33);
buf  g23 (n47, n37);
buf  g24 (n96, n54);
buf  g25 (n94, n40);
not  g26 (n93, n54);
not  g27 (n72, n45);
buf  g28 (n85, n9);
buf  g29 (n60, n26);
xnor g30 (n61, n31, n47, n48);
nor  g31 (n79, n28, n31, n18, n4);
xor  g32 (n88, n28, n38, n16, n48);
xnor g33 (n98, n53, n29, n14, n25);
xor  g34 (n92, n16, n5, n28, n43);
or   g35 (n82, n22, n19, n6, n21);
xnor g36 (n57, n52, n10, n7, n18);
xor  g37 (n71, n22, n9, n42, n26);
xnor g38 (n63, n44, n6, n32, n55);
nor  g39 (n64, n38, n25, n4, n41);
xnor g40 (n70, n39, n46, n49, n13);
nor  g41 (n95, n27, n27, n21, n46);
and  g42 (n99, n25, n47, n23, n3);
nor  g43 (n78, n46, n23, n49, n19);
and  g44 (n58, n43, n13, n53, n2);
or   g45 (n87, n5, n12, n25, n56);
and  g46 (n69, n50, n55, n40, n29);
nand g47 (n89, n7, n13, n39, n52);
nand g48 (n80, n17, n32, n30);
nor  g49 (n81, n18, n51, n45, n12);
nand g50 (n67, n6, n24, n30, n28);
nand g51 (n86, n24, n49, n27, n56);
nand g52 (n76, n14, n11, n3, n26);
and  g53 (n83, n17, n27, n9, n41);
nand g54 (n59, n12, n41, n3, n8);
and  g55 (n84, n53, n47, n51, n44);
and  g56 (n100, n8, n44, n56, n24);
nor  g57 (n77, n19, n17, n15, n31);
and  g58 (n68, n14, n15, n30, n20);
xor  g59 (n90, n23, n32, n8, n20);
or   g60 (n91, n31, n43, n42, n10);
and  g61 (n74, n38, n51, n55, n11);
xnor g62 (n62, n29, n54, n50, n52);
nor  g63 (n73, n26, n16, n5, n15);
or   g64 (n65, n40, n39, n7, n10);
xnor g65 (n75, n32, n24, n22, n48);
xnor g66 (n66, n50, n21, n29, n4);
nand g67 (n97, n20, n42, n11, n45);
xnor g68 (n104, n72, n78, n92, n59);
nor  g69 (n117, n81, n93, n80, n85);
or   g70 (n115, n59, n74, n65, n93);
xor  g71 (n106, n80, n95, n67, n97);
xor  g72 (n118, n100, n84, n76, n71);
nor  g73 (n124, n86, n62, n90, n59);
and  g74 (n131, n77, n72, n70, n63);
nor  g75 (n116, n97, n83, n95);
or   g76 (n105, n76, n64, n80, n96);
xnor g77 (n103, n91, n66, n58, n98);
or   g78 (n129, n70, n69, n62, n81);
xnor g79 (n101, n98, n60, n100, n78);
xnor g80 (n109, n99, n70, n85, n87);
xnor g81 (n121, n88, n61, n65, n77);
and  g82 (n102, n73, n67, n89, n63);
and  g83 (n111, n90, n73, n78, n72);
and  g84 (n127, n87, n92, n68, n79);
xor  g85 (n119, n94, n75, n74, n91);
xor  g86 (n113, n87, n96, n92, n71);
xnor g87 (n110, n67, n75, n94, n73);
nor  g88 (n114, n64, n71, n89, n79);
or   g89 (n107, n63, n83, n85, n65);
xnor g90 (n112, n77, n74, n88, n68);
nor  g91 (n120, n99, n60, n86, n75);
nand g92 (n128, n99, n86, n95, n66);
nand g93 (n123, n96, n81, n57, n62);
nor  g94 (n132, n82, n84, n88, n91);
xnor g95 (n122, n61, n98, n90, n69);
and  g96 (n125, n64, n61, n66, n84);
xnor g97 (n130, n60, n69, n76, n68);
xnor g98 (n126, n93, n79, n97, n82);
xor  g99 (n108, n89, n100, n82, n94);
endmodule
