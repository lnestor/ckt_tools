

module Stat_1000_109
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n912,
  n812,
  n867,
  n866,
  n806,
  n807,
  n833,
  n800,
  n906,
  n893,
  n860,
  n887,
  n909,
  n868,
  n848,
  n897,
  n853,
  n877,
  n904,
  n841,
  n811,
  n819,
  n832,
  n842,
  n875,
  n850,
  n1029,
  n1027,
  n1032,
  n1030,
  n1028,
  n1031
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n912;output n812;output n867;output n866;output n806;output n807;output n833;output n800;output n906;output n893;output n860;output n887;output n909;output n868;output n848;output n897;output n853;output n877;output n904;output n841;output n811;output n819;output n832;output n842;output n875;output n850;output n1029;output n1027;output n1032;output n1030;output n1028;output n1031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n801;wire n802;wire n803;wire n804;wire n805;wire n808;wire n809;wire n810;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n843;wire n844;wire n845;wire n846;wire n847;wire n849;wire n851;wire n852;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n861;wire n862;wire n863;wire n864;wire n865;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n876;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n888;wire n889;wire n890;wire n891;wire n892;wire n894;wire n895;wire n896;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n905;wire n907;wire n908;wire n910;wire n911;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n66,
    n13
  );


  not
  g1
  (
    n97,
    n3
  );


  not
  g2
  (
    n149,
    n5
  );


  buf
  g3
  (
    n130,
    n30
  );


  buf
  g4
  (
    KeyWire_0_15,
    n19
  );


  buf
  g5
  (
    n132,
    n30
  );


  not
  g6
  (
    n71,
    n7
  );


  not
  g7
  (
    n39,
    n28
  );


  not
  g8
  (
    n138,
    n32
  );


  not
  g9
  (
    n95,
    n18
  );


  not
  g10
  (
    n154,
    n6
  );


  not
  g11
  (
    KeyWire_0_12,
    n1
  );


  buf
  g12
  (
    n107,
    n9
  );


  not
  g13
  (
    n134,
    n8
  );


  buf
  g14
  (
    n68,
    n26
  );


  buf
  g15
  (
    n106,
    n4
  );


  buf
  g16
  (
    n114,
    n22
  );


  not
  g17
  (
    n135,
    n1
  );


  not
  g18
  (
    n113,
    n15
  );


  not
  g19
  (
    n99,
    n23
  );


  buf
  g20
  (
    n53,
    n20
  );


  not
  g21
  (
    n117,
    n9
  );


  buf
  g22
  (
    n96,
    n13
  );


  not
  g23
  (
    n159,
    n4
  );


  buf
  g24
  (
    n65,
    n5
  );


  buf
  g25
  (
    n62,
    n6
  );


  buf
  g26
  (
    n119,
    n20
  );


  buf
  g27
  (
    n120,
    n19
  );


  not
  g28
  (
    n72,
    n26
  );


  not
  g29
  (
    n157,
    n32
  );


  buf
  g30
  (
    n56,
    n2
  );


  not
  g31
  (
    n75,
    n12
  );


  not
  g32
  (
    n36,
    n9
  );


  buf
  g33
  (
    n102,
    n14
  );


  buf
  g34
  (
    n142,
    n21
  );


  not
  g35
  (
    n43,
    n24
  );


  not
  g36
  (
    n158,
    n20
  );


  not
  g37
  (
    n131,
    n25
  );


  not
  g38
  (
    n155,
    n10
  );


  buf
  g39
  (
    n55,
    n7
  );


  buf
  g40
  (
    n112,
    n11
  );


  not
  g41
  (
    n58,
    n2
  );


  buf
  g42
  (
    n45,
    n6
  );


  not
  g43
  (
    n145,
    n22
  );


  not
  g44
  (
    n81,
    n11
  );


  not
  g45
  (
    n70,
    n30
  );


  not
  g46
  (
    n49,
    n29
  );


  buf
  g47
  (
    n101,
    n18
  );


  not
  g48
  (
    n127,
    n29
  );


  not
  g49
  (
    n74,
    n29
  );


  not
  g50
  (
    n73,
    n3
  );


  not
  g51
  (
    n94,
    n30
  );


  buf
  g52
  (
    n33,
    n8
  );


  buf
  g53
  (
    n37,
    n28
  );


  not
  g54
  (
    n82,
    n8
  );


  not
  g55
  (
    n42,
    n23
  );


  buf
  g56
  (
    n148,
    n19
  );


  buf
  g57
  (
    n110,
    n16
  );


  buf
  g58
  (
    n115,
    n10
  );


  not
  g59
  (
    n76,
    n14
  );


  not
  g60
  (
    n80,
    n22
  );


  buf
  g61
  (
    n60,
    n25
  );


  buf
  g62
  (
    n103,
    n20
  );


  not
  g63
  (
    n153,
    n31
  );


  buf
  g64
  (
    n83,
    n5
  );


  buf
  g65
  (
    n116,
    n1
  );


  not
  g66
  (
    n123,
    n28
  );


  not
  g67
  (
    n84,
    n16
  );


  not
  g68
  (
    n124,
    n31
  );


  buf
  g69
  (
    n54,
    n12
  );


  not
  g70
  (
    n100,
    n27
  );


  buf
  g71
  (
    n89,
    n11
  );


  buf
  g72
  (
    n111,
    n13
  );


  not
  g73
  (
    n34,
    n32
  );


  buf
  g74
  (
    n78,
    n6
  );


  not
  g75
  (
    n87,
    n8
  );


  buf
  g76
  (
    n143,
    n28
  );


  buf
  g77
  (
    n69,
    n16
  );


  buf
  g78
  (
    n85,
    n2
  );


  buf
  g79
  (
    n152,
    n15
  );


  buf
  g80
  (
    n108,
    n26
  );


  buf
  g81
  (
    n146,
    n12
  );


  not
  g82
  (
    n46,
    n5
  );


  not
  g83
  (
    n150,
    n15
  );


  buf
  g84
  (
    n77,
    n10
  );


  buf
  g85
  (
    n61,
    n4
  );


  not
  g86
  (
    n160,
    n31
  );


  not
  g87
  (
    n90,
    n24
  );


  buf
  g88
  (
    n126,
    n17
  );


  not
  g89
  (
    n48,
    n4
  );


  buf
  g90
  (
    n140,
    n3
  );


  not
  g91
  (
    n151,
    n22
  );


  not
  g92
  (
    n51,
    n16
  );


  not
  g93
  (
    n104,
    n27
  );


  buf
  g94
  (
    n57,
    n21
  );


  buf
  g95
  (
    n50,
    n3
  );


  buf
  g96
  (
    n91,
    n17
  );


  not
  g97
  (
    n88,
    n27
  );


  not
  g98
  (
    n128,
    n14
  );


  buf
  g99
  (
    n136,
    n21
  );


  not
  g100
  (
    KeyWire_0_29,
    n15
  );


  buf
  g101
  (
    n144,
    n24
  );


  not
  g102
  (
    n139,
    n25
  );


  not
  g103
  (
    n63,
    n23
  );


  not
  g104
  (
    n52,
    n10
  );


  buf
  g105
  (
    n105,
    n26
  );


  buf
  g106
  (
    n86,
    n11
  );


  not
  g107
  (
    n109,
    n31
  );


  not
  g108
  (
    n133,
    n21
  );


  buf
  g109
  (
    n38,
    n29
  );


  not
  g110
  (
    n41,
    n19
  );


  buf
  g111
  (
    n125,
    n2
  );


  buf
  g112
  (
    n47,
    n9
  );


  not
  g113
  (
    n92,
    n12
  );


  buf
  g114
  (
    n137,
    n27
  );


  buf
  g115
  (
    n129,
    n1
  );


  buf
  g116
  (
    n156,
    n23
  );


  buf
  g117
  (
    KeyWire_0_23,
    n7
  );


  not
  g118
  (
    n35,
    n17
  );


  not
  g119
  (
    KeyWire_0_22,
    n24
  );


  not
  g120
  (
    n59,
    n25
  );


  buf
  g121
  (
    n98,
    n14
  );


  buf
  g122
  (
    n93,
    n13
  );


  not
  g123
  (
    n44,
    n17
  );


  buf
  g124
  (
    n121,
    n7
  );


  buf
  g125
  (
    n67,
    n18
  );


  buf
  g126
  (
    n141,
    n18
  );


  not
  g127
  (
    n64,
    n32
  );


  or
  g128
  (
    n266,
    n129,
    n42
  );


  xor
  g129
  (
    n250,
    n48,
    n138
  );


  nand
  g130
  (
    n304,
    n81,
    n142
  );


  nor
  g131
  (
    n277,
    n33,
    n127
  );


  xnor
  g132
  (
    n248,
    n45,
    n150
  );


  nand
  g133
  (
    n279,
    n46,
    n82
  );


  or
  g134
  (
    n296,
    n120,
    n132
  );


  xor
  g135
  (
    n303,
    n130,
    n111
  );


  or
  g136
  (
    n225,
    n96,
    n102
  );


  xor
  g137
  (
    n283,
    n47,
    n51
  );


  xor
  g138
  (
    n352,
    n65,
    n120
  );


  xnor
  g139
  (
    n344,
    n56,
    n137
  );


  nor
  g140
  (
    n251,
    n62,
    n159
  );


  or
  g141
  (
    n280,
    n43,
    n112
  );


  xnor
  g142
  (
    n342,
    n105,
    n71
  );


  nor
  g143
  (
    n325,
    n59,
    n124
  );


  xnor
  g144
  (
    n182,
    n58,
    n70
  );


  and
  g145
  (
    n346,
    n64,
    n83
  );


  xor
  g146
  (
    n338,
    n79,
    n154
  );


  nor
  g147
  (
    n215,
    n60,
    n123
  );


  nor
  g148
  (
    n244,
    n44,
    n35
  );


  and
  g149
  (
    n247,
    n120,
    n88
  );


  nand
  g150
  (
    n227,
    n148,
    n72
  );


  or
  g151
  (
    n276,
    n133,
    n113
  );


  nand
  g152
  (
    n230,
    n103,
    n71
  );


  xor
  g153
  (
    n191,
    n123,
    n43
  );


  and
  g154
  (
    n187,
    n63,
    n43
  );


  xnor
  g155
  (
    n184,
    n140,
    n41
  );


  nand
  g156
  (
    n299,
    n109,
    n123
  );


  and
  g157
  (
    n223,
    n36,
    n141
  );


  xnor
  g158
  (
    n188,
    n93,
    n138
  );


  and
  g159
  (
    n316,
    n100,
    n143
  );


  or
  g160
  (
    n246,
    n59,
    n156
  );


  xor
  g161
  (
    n336,
    n92,
    n134
  );


  xnor
  g162
  (
    n179,
    n71,
    n150
  );


  or
  g163
  (
    n337,
    n35,
    n60
  );


  and
  g164
  (
    n307,
    n91,
    n84
  );


  and
  g165
  (
    n309,
    n96,
    n61
  );


  and
  g166
  (
    n318,
    n68,
    n105
  );


  nand
  g167
  (
    n214,
    n102,
    n86
  );


  xor
  g168
  (
    n238,
    n101,
    n115
  );


  and
  g169
  (
    n270,
    n159,
    n112
  );


  or
  g170
  (
    n261,
    n50,
    n45
  );


  nand
  g171
  (
    n168,
    n90,
    n64
  );


  or
  g172
  (
    n190,
    n70,
    n146
  );


  not
  g173
  (
    n331,
    n34
  );


  and
  g174
  (
    n282,
    n35,
    n86
  );


  nor
  g175
  (
    n284,
    n132,
    n64
  );


  xor
  g176
  (
    n305,
    n126,
    n97
  );


  xor
  g177
  (
    n170,
    n57,
    n119
  );


  xor
  g178
  (
    n226,
    n117,
    n152
  );


  xor
  g179
  (
    n205,
    n125,
    n33
  );


  xor
  g180
  (
    n328,
    n149,
    n91
  );


  xor
  g181
  (
    n176,
    n124,
    n117
  );


  and
  g182
  (
    n294,
    n83,
    n122
  );


  nor
  g183
  (
    n194,
    n122,
    n79
  );


  xor
  g184
  (
    n163,
    n85,
    n133
  );


  and
  g185
  (
    n224,
    n59,
    n63
  );


  and
  g186
  (
    n203,
    n147,
    n129
  );


  or
  g187
  (
    n169,
    n126,
    n112
  );


  and
  g188
  (
    n197,
    n135,
    n68
  );


  or
  g189
  (
    n245,
    n148,
    n109
  );


  xor
  g190
  (
    n351,
    n100,
    n76
  );


  nand
  g191
  (
    n265,
    n131,
    n118
  );


  nand
  g192
  (
    n252,
    n97,
    n74
  );


  xnor
  g193
  (
    n240,
    n72,
    n94
  );


  and
  g194
  (
    n183,
    n106,
    n66
  );


  or
  g195
  (
    n171,
    n89,
    n153
  );


  xor
  g196
  (
    n285,
    n69,
    n138
  );


  xnor
  g197
  (
    n235,
    n92,
    n103
  );


  nand
  g198
  (
    n302,
    n155,
    n78
  );


  and
  g199
  (
    n345,
    n145,
    n124
  );


  nand
  g200
  (
    n311,
    n104,
    n132
  );


  and
  g201
  (
    n236,
    n47,
    n105
  );


  or
  g202
  (
    n249,
    n90,
    n154
  );


  and
  g203
  (
    n242,
    n89,
    n75
  );


  and
  g204
  (
    n233,
    n34,
    n71
  );


  and
  g205
  (
    n257,
    n134,
    n130
  );


  xnor
  g206
  (
    n339,
    n135,
    n98
  );


  or
  g207
  (
    n237,
    n53,
    n142
  );


  or
  g208
  (
    n263,
    n70,
    n100
  );


  nand
  g209
  (
    n216,
    n78,
    n160
  );


  xor
  g210
  (
    n269,
    n111,
    n156
  );


  xor
  g211
  (
    n241,
    n146,
    n115
  );


  and
  g212
  (
    n343,
    n81,
    n137
  );


  or
  g213
  (
    n255,
    n38,
    n58
  );


  nand
  g214
  (
    n254,
    n154,
    n133
  );


  or
  g215
  (
    n198,
    n87,
    n117
  );


  and
  g216
  (
    n165,
    n93,
    n51
  );


  nand
  g217
  (
    n330,
    n85,
    n77
  );


  or
  g218
  (
    n189,
    n86,
    n41
  );


  xor
  g219
  (
    n167,
    n44,
    n152
  );


  xnor
  g220
  (
    n239,
    n55,
    n150
  );


  xnor
  g221
  (
    KeyWire_0_9,
    n134,
    n94
  );


  xor
  g222
  (
    n295,
    n99,
    n138
  );


  and
  g223
  (
    n310,
    n160,
    n144
  );


  or
  g224
  (
    n210,
    n137,
    n40
  );


  nor
  g225
  (
    n232,
    n61,
    n102
  );


  and
  g226
  (
    n178,
    n139,
    n101
  );


  nand
  g227
  (
    n200,
    n98,
    n85
  );


  nor
  g228
  (
    n181,
    n108,
    n79
  );


  and
  g229
  (
    n334,
    n108,
    n95
  );


  nor
  g230
  (
    n208,
    n148,
    n155
  );


  nand
  g231
  (
    n287,
    n131,
    n118
  );


  or
  g232
  (
    n274,
    n49,
    n147
  );


  xnor
  g233
  (
    n297,
    n74,
    n77
  );


  and
  g234
  (
    n350,
    n155,
    n73
  );


  nand
  g235
  (
    n206,
    n63,
    n149
  );


  nor
  g236
  (
    n288,
    n113,
    n153
  );


  and
  g237
  (
    n207,
    n74,
    n130
  );


  or
  g238
  (
    n186,
    n42,
    n143
  );


  nand
  g239
  (
    n259,
    n90,
    n60
  );


  nand
  g240
  (
    n321,
    n141,
    n145
  );


  or
  g241
  (
    n175,
    n146,
    n128
  );


  xor
  g242
  (
    n260,
    n127,
    n51
  );


  xnor
  g243
  (
    n199,
    n37,
    n129
  );


  xor
  g244
  (
    KeyWire_0_19,
    n126,
    n156
  );


  and
  g245
  (
    n329,
    n86,
    n125
  );


  or
  g246
  (
    n315,
    n52,
    n54
  );


  nand
  g247
  (
    n243,
    n39,
    n61
  );


  nand
  g248
  (
    n192,
    n40,
    n82
  );


  nor
  g249
  (
    n217,
    n35,
    n160
  );


  or
  g250
  (
    n327,
    n70,
    n47
  );


  nand
  g251
  (
    n211,
    n104,
    n119
  );


  nand
  g252
  (
    n335,
    n140,
    n159
  );


  and
  g253
  (
    n173,
    n75,
    n69
  );


  xor
  g254
  (
    n209,
    n42,
    n151
  );


  nor
  g255
  (
    n272,
    n76,
    n82
  );


  or
  g256
  (
    n332,
    n89,
    n99
  );


  nor
  g257
  (
    n193,
    n90,
    n91
  );


  and
  g258
  (
    n317,
    n151,
    n87,
    n158,
    n111
  );


  nand
  g259
  (
    n220,
    n97,
    n154,
    n145,
    n127
  );


  xor
  g260
  (
    n319,
    n96,
    n121,
    n63
  );


  xnor
  g261
  (
    n196,
    n120,
    n157,
    n155,
    n68
  );


  nor
  g262
  (
    n323,
    n139,
    n139,
    n101,
    n50
  );


  nand
  g263
  (
    n278,
    n144,
    n61,
    n114,
    n57
  );


  and
  g264
  (
    n219,
    n116,
    n159,
    n57,
    n129
  );


  or
  g265
  (
    n161,
    n139,
    n80,
    n97,
    n49
  );


  or
  g266
  (
    n341,
    n157,
    n69,
    n55,
    n36
  );


  xor
  g267
  (
    n180,
    n143,
    n46,
    n145,
    n115
  );


  and
  g268
  (
    n322,
    n123,
    n72,
    n36,
    n113
  );


  or
  g269
  (
    n262,
    n54,
    n75,
    n135,
    n106
  );


  or
  g270
  (
    n218,
    n109,
    n39,
    n88
  );


  nand
  g271
  (
    n273,
    n39,
    n51,
    n110,
    n104
  );


  nand
  g272
  (
    n264,
    n80,
    n106,
    n94,
    n116
  );


  and
  g273
  (
    n271,
    n111,
    n37,
    n101,
    n89
  );


  xnor
  g274
  (
    n292,
    n49,
    n49,
    n135,
    n55
  );


  and
  g275
  (
    n301,
    n68,
    n48,
    n87,
    n92
  );


  xnor
  g276
  (
    n177,
    n110,
    n57,
    n131,
    n108
  );


  nand
  g277
  (
    n258,
    n94,
    n64,
    n55,
    n65
  );


  nand
  g278
  (
    n281,
    n99,
    n122,
    n67,
    n114
  );


  xor
  g279
  (
    n275,
    n110,
    n88,
    n85,
    n116
  );


  or
  g280
  (
    n222,
    n77,
    n77,
    n144,
    n93
  );


  and
  g281
  (
    n164,
    n124,
    n140,
    n48,
    n79
  );


  and
  g282
  (
    n312,
    n41,
    n122,
    n152,
    n93
  );


  or
  g283
  (
    n253,
    n73,
    n52,
    n107,
    n115
  );


  and
  g284
  (
    n204,
    n133,
    n40,
    n34,
    n73
  );


  xnor
  g285
  (
    n348,
    n128,
    n46,
    n106,
    n54
  );


  xor
  g286
  (
    n166,
    n67,
    n78,
    n141,
    n95
  );


  nand
  g287
  (
    n308,
    n98,
    n103,
    n134,
    n52
  );


  nand
  g288
  (
    n212,
    n118,
    n127,
    n80,
    n158
  );


  or
  g289
  (
    n286,
    n52,
    n160,
    n158,
    n45
  );


  nand
  g290
  (
    n353,
    n41,
    n144,
    n84,
    n156
  );


  and
  g291
  (
    n267,
    n146,
    n62,
    n98,
    n113
  );


  nor
  g292
  (
    n349,
    n92,
    n48,
    n132,
    n37
  );


  nor
  g293
  (
    n324,
    n69,
    n108,
    n42,
    n149
  );


  xor
  g294
  (
    n300,
    n152,
    n116,
    n136,
    n114
  );


  nor
  g295
  (
    n290,
    n117,
    n44,
    n136,
    n103
  );


  nand
  g296
  (
    n289,
    n78,
    n95,
    n99,
    n66
  );


  and
  g297
  (
    n333,
    n62,
    n33,
    n104,
    n59
  );


  nor
  g298
  (
    n202,
    n56,
    n66,
    n157,
    n141
  );


  xor
  g299
  (
    n201,
    n150,
    n112,
    n107,
    n102
  );


  xor
  g300
  (
    n298,
    n50,
    n137,
    n105,
    n45
  );


  nand
  g301
  (
    n174,
    n66,
    n131,
    n62,
    n142
  );


  or
  g302
  (
    n347,
    n53,
    n158,
    n73,
    n60
  );


  and
  g303
  (
    n313,
    n119,
    n67,
    n43,
    n83
  );


  nor
  g304
  (
    n306,
    n53,
    n36,
    n151,
    n121
  );


  nand
  g305
  (
    n256,
    n84,
    n67,
    n58,
    n126
  );


  or
  g306
  (
    n185,
    n118,
    n143,
    n153,
    n128
  );


  or
  g307
  (
    n229,
    n147,
    n147,
    n38,
    n40
  );


  xnor
  g308
  (
    n228,
    n65,
    n100,
    n140,
    n149
  );


  xor
  g309
  (
    n268,
    n37,
    n130,
    n136,
    n88
  );


  nor
  g310
  (
    n291,
    n125,
    n50,
    n56,
    n72
  );


  nand
  g311
  (
    n213,
    n54,
    n91,
    n107,
    n96
  );


  nand
  g312
  (
    n221,
    n95,
    n142,
    n56,
    n82
  );


  nor
  g313
  (
    n320,
    n121,
    n76,
    n119,
    n153
  );


  and
  g314
  (
    n234,
    n38,
    n87,
    n157,
    n136
  );


  or
  g315
  (
    n314,
    n53,
    n128,
    n151,
    n84
  );


  nor
  g316
  (
    n162,
    n38,
    n125,
    n47,
    n76
  );


  nand
  g317
  (
    KeyWire_0_13,
    n33,
    n148,
    n81,
    n75
  );


  nor
  g318
  (
    n340,
    n80,
    n83,
    n107,
    n46
  );


  or
  g319
  (
    n195,
    n74,
    n81,
    n109,
    n65
  );


  nor
  g320
  (
    n231,
    n44,
    n110,
    n58,
    n114
  );


  xor
  g321
  (
    n398,
    n317,
    n287,
    n236,
    n301
  );


  nand
  g322
  (
    n386,
    n162,
    n202,
    n205,
    n262
  );


  nand
  g323
  (
    n399,
    n206,
    n260,
    n229,
    n293
  );


  and
  g324
  (
    n429,
    n299,
    n287,
    n177,
    n310
  );


  xnor
  g325
  (
    n537,
    n231,
    n231,
    n336,
    n183
  );


  or
  g326
  (
    n454,
    n248,
    n308,
    n258,
    n254
  );


  nand
  g327
  (
    n495,
    n324,
    n176,
    n341,
    n200
  );


  nor
  g328
  (
    KeyWire_0_11,
    n184,
    n289,
    n288,
    n295
  );


  nand
  g329
  (
    n491,
    n301,
    n338,
    n276,
    n187
  );


  nor
  g330
  (
    n363,
    n292,
    n284,
    n318,
    n323
  );


  xnor
  g331
  (
    n376,
    n246,
    n178,
    n166,
    n278
  );


  and
  g332
  (
    n503,
    n263,
    n204,
    n163,
    n282
  );


  xnor
  g333
  (
    n360,
    n215,
    n261,
    n164,
    n240
  );


  xnor
  g334
  (
    n414,
    n277,
    n324,
    n225,
    n233
  );


  xnor
  g335
  (
    n524,
    n207,
    n304,
    n299,
    n315
  );


  xor
  g336
  (
    n387,
    n298,
    n236,
    n330,
    n211
  );


  and
  g337
  (
    n526,
    n313,
    n301,
    n325,
    n182
  );


  nand
  g338
  (
    n479,
    n172,
    n181,
    n334,
    n247
  );


  xor
  g339
  (
    n388,
    n328,
    n226,
    n284,
    n212
  );


  and
  g340
  (
    n416,
    n337,
    n270,
    n292,
    n216
  );


  nand
  g341
  (
    n518,
    n280,
    n322,
    n287,
    n249
  );


  xor
  g342
  (
    n474,
    n302,
    n173,
    n186,
    n252
  );


  nand
  g343
  (
    n478,
    n339,
    n193,
    n293,
    n281
  );


  nand
  g344
  (
    n447,
    n326,
    n210,
    n265,
    n298
  );


  xnor
  g345
  (
    n511,
    n250,
    n243,
    n216,
    n228
  );


  xor
  g346
  (
    n506,
    n248,
    n180,
    n221,
    n218
  );


  xor
  g347
  (
    n452,
    n213,
    n327,
    n172,
    n183
  );


  or
  g348
  (
    n505,
    n257,
    n205,
    n211,
    n307
  );


  nor
  g349
  (
    n497,
    n331,
    n243,
    n298,
    n165
  );


  or
  g350
  (
    n499,
    n321,
    n337,
    n269,
    n256
  );


  xor
  g351
  (
    n469,
    n213,
    n228,
    n238,
    n262
  );


  xnor
  g352
  (
    n400,
    n183,
    n222,
    n327,
    n170
  );


  xor
  g353
  (
    n451,
    n234,
    n307,
    n167,
    n293
  );


  and
  g354
  (
    n379,
    n246,
    n227,
    n204,
    n300
  );


  xor
  g355
  (
    n383,
    n195,
    n285,
    n310,
    n305
  );


  xnor
  g356
  (
    n409,
    n171,
    n191,
    n210,
    n267
  );


  nor
  g357
  (
    n514,
    n267,
    n290,
    n249,
    n198
  );


  nand
  g358
  (
    n446,
    n326,
    n223,
    n328,
    n190
  );


  xnor
  g359
  (
    n512,
    n193,
    n327,
    n272,
    n188
  );


  and
  g360
  (
    n397,
    n215,
    n297,
    n291,
    n175
  );


  xor
  g361
  (
    n445,
    n312,
    n198,
    n313,
    n176
  );


  nor
  g362
  (
    n450,
    n319,
    n248,
    n186
  );


  xnor
  g363
  (
    n507,
    n343,
    n202,
    n298,
    n329
  );


  xnor
  g364
  (
    n430,
    n252,
    n272,
    n340,
    n188
  );


  and
  g365
  (
    n457,
    n251,
    n270,
    n295,
    n313
  );


  or
  g366
  (
    n417,
    n247,
    n230,
    n292,
    n205
  );


  or
  g367
  (
    KeyWire_0_10,
    n220,
    n303,
    n215,
    n234
  );


  or
  g368
  (
    n465,
    n264,
    n175,
    n224,
    n302
  );


  nor
  g369
  (
    n408,
    n308,
    n273,
    n254,
    n203
  );


  nand
  g370
  (
    n401,
    n180,
    n200,
    n286,
    n182
  );


  nor
  g371
  (
    n356,
    n286,
    n337,
    n340,
    n276
  );


  and
  g372
  (
    n392,
    n324,
    n260,
    n278,
    n186
  );


  nand
  g373
  (
    n496,
    n313,
    n195,
    n266,
    n314
  );


  xor
  g374
  (
    n393,
    n344,
    n205,
    n333,
    n302
  );


  nand
  g375
  (
    n484,
    n296,
    n256,
    n230,
    n203
  );


  nor
  g376
  (
    n406,
    n306,
    n311,
    n241,
    n197
  );


  or
  g377
  (
    n536,
    n262,
    n227,
    n213,
    n261
  );


  or
  g378
  (
    n494,
    n176,
    n181,
    n224,
    n332
  );


  nor
  g379
  (
    n378,
    n254,
    n335,
    n344,
    n283
  );


  nor
  g380
  (
    n470,
    n239,
    n285,
    n168,
    n220
  );


  xor
  g381
  (
    n502,
    n291,
    n258,
    n262,
    n301
  );


  xor
  g382
  (
    n519,
    n243,
    n207,
    n172,
    n306
  );


  and
  g383
  (
    n382,
    n296,
    n321,
    n256,
    n227
  );


  nand
  g384
  (
    n528,
    n345,
    n319,
    n252,
    n299
  );


  xor
  g385
  (
    n355,
    n182,
    n200,
    n238,
    n187
  );


  nand
  g386
  (
    n443,
    n336,
    n241,
    n184,
    n204
  );


  nand
  g387
  (
    n373,
    n171,
    n271,
    n281,
    n286
  );


  nand
  g388
  (
    n438,
    n323,
    n236,
    n201,
    n237
  );


  or
  g389
  (
    n440,
    n188,
    n198,
    n161,
    n251
  );


  nand
  g390
  (
    n508,
    n318,
    n311,
    n202,
    n213
  );


  xnor
  g391
  (
    n531,
    n309,
    n290,
    n239,
    n173
  );


  or
  g392
  (
    n427,
    n339,
    n272,
    n271,
    n316
  );


  nor
  g393
  (
    n402,
    n335,
    n249,
    n242,
    n189
  );


  nor
  g394
  (
    n413,
    n274,
    n297,
    n327,
    n218
  );


  nor
  g395
  (
    n428,
    n210,
    n259,
    n277,
    n275
  );


  nor
  g396
  (
    KeyWire_0_31,
    n280,
    n314,
    n193,
    n212
  );


  xnor
  g397
  (
    n407,
    n260,
    n290,
    n294,
    n242
  );


  or
  g398
  (
    n359,
    n232,
    n315,
    n192,
    n199
  );


  nor
  g399
  (
    n492,
    n283,
    n294,
    n197,
    n185
  );


  xnor
  g400
  (
    n482,
    n328,
    n247,
    n161,
    n214
  );


  or
  g401
  (
    n405,
    n209,
    n253,
    n323,
    n245
  );


  or
  g402
  (
    n433,
    n259,
    n260,
    n322,
    n295
  );


  and
  g403
  (
    n442,
    n237,
    n261,
    n196
  );


  xor
  g404
  (
    n435,
    n230,
    n338,
    n203,
    n217
  );


  nand
  g405
  (
    n377,
    n169,
    n201,
    n219,
    n265
  );


  xor
  g406
  (
    n364,
    n268,
    n267,
    n339,
    n284
  );


  nor
  g407
  (
    n522,
    n333,
    n320,
    n342,
    n245
  );


  xnor
  g408
  (
    n432,
    n214,
    n182,
    n163,
    n255
  );


  nor
  g409
  (
    n426,
    n300,
    n171,
    n161,
    n256
  );


  and
  g410
  (
    n367,
    n181,
    n168,
    n273,
    n329
  );


  nand
  g411
  (
    n473,
    n274,
    n341,
    n216,
    n217
  );


  or
  g412
  (
    n501,
    n270,
    n324,
    n218,
    n185
  );


  or
  g413
  (
    n487,
    n167,
    n320,
    n305,
    n304
  );


  nand
  g414
  (
    n436,
    n217,
    n199,
    n292,
    n222
  );


  or
  g415
  (
    n418,
    n269,
    n248,
    n322,
    n170
  );


  nor
  g416
  (
    n460,
    n310,
    n331,
    n194,
    n295
  );


  and
  g417
  (
    n483,
    n193,
    n329,
    n238,
    n204
  );


  or
  g418
  (
    n381,
    n280,
    n237,
    n330,
    n225
  );


  xnor
  g419
  (
    n370,
    n183,
    n191,
    n209,
    n221
  );


  xor
  g420
  (
    n422,
    n291,
    n274,
    n264,
    n197
  );


  nor
  g421
  (
    n498,
    n244,
    n290,
    n272,
    n229
  );


  nor
  g422
  (
    n533,
    n163,
    n320,
    n276,
    n266
  );


  xor
  g423
  (
    n415,
    n253,
    n330,
    n333,
    n318
  );


  xor
  g424
  (
    n463,
    n164,
    n258,
    n266,
    n287
  );


  nor
  g425
  (
    n358,
    n214,
    n166,
    n232,
    n176
  );


  or
  g426
  (
    n372,
    n200,
    n267,
    n319,
    n343
  );


  nor
  g427
  (
    n410,
    n179,
    n206,
    n284,
    n252
  );


  and
  g428
  (
    n538,
    n293,
    n243,
    n217,
    n334
  );


  and
  g429
  (
    n365,
    n337,
    n181,
    n196,
    n187
  );


  xnor
  g430
  (
    n466,
    n194,
    n222,
    n236
  );


  xnor
  g431
  (
    n510,
    n227,
    n228,
    n199,
    n321
  );


  xor
  g432
  (
    n403,
    n226,
    n165,
    n309,
    n291
  );


  xnor
  g433
  (
    n455,
    n189,
    n338,
    n294,
    n178
  );


  xor
  g434
  (
    n419,
    n174,
    n259,
    n332,
    n286
  );


  and
  g435
  (
    n369,
    n208,
    n342,
    n237,
    n277
  );


  and
  g436
  (
    n412,
    n253,
    n233,
    n192,
    n338
  );


  and
  g437
  (
    n516,
    n224,
    n278,
    n315,
    n235
  );


  xor
  g438
  (
    n421,
    n162,
    n326,
    n253,
    n246
  );


  xnor
  g439
  (
    n384,
    n345,
    n274,
    n332,
    n179
  );


  xor
  g440
  (
    n481,
    n329,
    n164,
    n223,
    n273
  );


  or
  g441
  (
    n437,
    n315,
    n220,
    n234,
    n229
  );


  nand
  g442
  (
    n530,
    n328,
    n336,
    n317,
    n228
  );


  xnor
  g443
  (
    n488,
    n194,
    n206,
    n221,
    n174
  );


  xnor
  g444
  (
    n354,
    n190,
    n173,
    n196,
    n219
  );


  nor
  g445
  (
    n448,
    n178,
    n257,
    n189,
    n280
  );


  xor
  g446
  (
    n391,
    n164,
    n250,
    n178,
    n340
  );


  nand
  g447
  (
    n480,
    n245,
    n219,
    n254,
    n216
  );


  and
  g448
  (
    n424,
    n309,
    n316,
    n169,
    n321
  );


  nand
  g449
  (
    n509,
    n282,
    n331,
    n344,
    n245
  );


  nor
  g450
  (
    n423,
    n318,
    n308,
    n214,
    n180
  );


  xnor
  g451
  (
    n459,
    n282,
    n184,
    n275,
    n165
  );


  nor
  g452
  (
    n368,
    n255,
    n163,
    n302,
    n316
  );


  nor
  g453
  (
    n444,
    n219,
    n289,
    n206,
    n233
  );


  nor
  g454
  (
    n472,
    n322,
    n334,
    n317,
    n191
  );


  xor
  g455
  (
    n525,
    n263,
    n297,
    n304,
    n330
  );


  xor
  g456
  (
    n375,
    n196,
    n212,
    n190,
    n300
  );


  nand
  g457
  (
    n434,
    n273,
    n270,
    n317,
    n336
  );


  nor
  g458
  (
    n441,
    n251,
    n165,
    n312,
    n340
  );


  nor
  g459
  (
    n513,
    n172,
    n226,
    n307,
    n326
  );


  and
  g460
  (
    n504,
    n209,
    n265,
    n190,
    n294
  );


  and
  g461
  (
    n535,
    n188,
    n202,
    n185,
    n278
  );


  and
  g462
  (
    n449,
    n220,
    n345,
    n184,
    n223
  );


  nor
  g463
  (
    n490,
    n211,
    n296,
    n192,
    n283
  );


  and
  g464
  (
    n464,
    n225,
    n235,
    n195,
    n208
  );


  and
  g465
  (
    n489,
    n339,
    n224,
    n226,
    n275
  );


  nor
  g466
  (
    n357,
    n233,
    n232,
    n174,
    n279
  );


  nand
  g467
  (
    n527,
    n175,
    n189,
    n235,
    n168
  );


  nand
  g468
  (
    n523,
    n198,
    n335,
    n268,
    n207
  );


  or
  g469
  (
    n456,
    n269,
    n170,
    n215,
    n281
  );


  xor
  g470
  (
    n500,
    n276,
    n247,
    n212,
    n229
  );


  xor
  g471
  (
    n395,
    n288,
    n209,
    n266,
    n314
  );


  or
  g472
  (
    KeyWire_0_20,
    n242,
    n299,
    n325,
    n289
  );


  xnor
  g473
  (
    n486,
    n173,
    n208,
    n241,
    n283
  );


  xnor
  g474
  (
    n471,
    n296,
    n305,
    n171,
    n175
  );


  xor
  g475
  (
    n468,
    n179,
    n345,
    n210,
    n250
  );


  nand
  g476
  (
    n515,
    n238,
    n281,
    n334,
    n325
  );


  and
  g477
  (
    n467,
    n304,
    n241,
    n282,
    n167
  );


  nand
  g478
  (
    n361,
    n195,
    n255,
    n161,
    n170
  );


  xor
  g479
  (
    n458,
    n246,
    n314,
    n221,
    n192
  );


  or
  g480
  (
    n362,
    n180,
    n279,
    n342,
    n300
  );


  and
  g481
  (
    n371,
    n268,
    n307,
    n239,
    n207
  );


  xor
  g482
  (
    n532,
    n257,
    n341,
    n306,
    n265
  );


  nand
  g483
  (
    n420,
    n316,
    n303,
    n305,
    n263
  );


  xnor
  g484
  (
    KeyWire_0_14,
    n285,
    n342,
    n268,
    n232
  );


  nand
  g485
  (
    n475,
    n259,
    n311,
    n271,
    n162
  );


  xnor
  g486
  (
    n374,
    n303,
    n177,
    n279
  );


  and
  g487
  (
    n380,
    n312,
    n250,
    n306,
    n303
  );


  xnor
  g488
  (
    n485,
    n218,
    n201,
    n203,
    n308
  );


  xor
  g489
  (
    n476,
    n257,
    n288,
    n179,
    n166
  );


  nand
  g490
  (
    n411,
    n168,
    n194,
    n343,
    n325
  );


  or
  g491
  (
    n534,
    n211,
    n320,
    n174,
    n263
  );


  xor
  g492
  (
    n396,
    n244,
    n239,
    n223,
    n231
  );


  nor
  g493
  (
    n529,
    n230,
    n323,
    n331,
    n310
  );


  nand
  g494
  (
    n453,
    n277,
    n240,
    n271,
    n185
  );


  xnor
  g495
  (
    n366,
    n319,
    n162,
    n197,
    n244
  );


  xnor
  g496
  (
    n404,
    n269,
    n332,
    n258,
    n201
  );


  and
  g497
  (
    n425,
    n177,
    n231,
    n333,
    n244
  );


  xor
  g498
  (
    n493,
    n169,
    n309,
    n225,
    n208
  );


  xnor
  g499
  (
    n431,
    n169,
    n187,
    n240,
    n289
  );


  and
  g500
  (
    n521,
    n240,
    n199,
    n264,
    n341
  );


  xnor
  g501
  (
    n517,
    n288,
    n255,
    n312,
    n335
  );


  nor
  g502
  (
    n477,
    n191,
    n311,
    n166,
    n234
  );


  nor
  g503
  (
    n462,
    n285,
    n344,
    n279,
    n251
  );


  nand
  g504
  (
    n394,
    n249,
    n275,
    n343,
    n264
  );


  xor
  g505
  (
    n461,
    n297,
    n167,
    n235,
    n242
  );


  xor
  g506
  (
    n559,
    n365,
    n407,
    n414,
    n420
  );


  or
  g507
  (
    n546,
    n415,
    n440,
    n390,
    n423
  );


  and
  g508
  (
    n606,
    n443,
    n449,
    n434,
    n445
  );


  xor
  g509
  (
    n620,
    n395,
    n394,
    n413,
    n415
  );


  nand
  g510
  (
    n576,
    n467,
    n393,
    n398,
    n399
  );


  xnor
  g511
  (
    n543,
    n356,
    n452,
    n437,
    n449
  );


  xnor
  g512
  (
    n618,
    n358,
    n416,
    n461,
    n401
  );


  xnor
  g513
  (
    n579,
    n446,
    n436,
    n463,
    n382
  );


  or
  g514
  (
    n590,
    n406,
    n460,
    n450,
    n432
  );


  nor
  g515
  (
    n551,
    n385,
    n412,
    n399,
    n408
  );


  xor
  g516
  (
    n599,
    n397,
    n394,
    n425,
    n376
  );


  xnor
  g517
  (
    n541,
    n398,
    n357,
    n443,
    n435
  );


  nor
  g518
  (
    n561,
    n406,
    n405,
    n429,
    n459
  );


  nor
  g519
  (
    n603,
    n397,
    n463,
    n362,
    n450
  );


  xnor
  g520
  (
    n614,
    n426,
    n452,
    n466,
    n376
  );


  and
  g521
  (
    KeyWire_0_4,
    n410,
    n389,
    n460,
    n416
  );


  xor
  g522
  (
    n582,
    n378,
    n425,
    n457,
    n398
  );


  and
  g523
  (
    n597,
    n396,
    n396,
    n440,
    n392
  );


  xor
  g524
  (
    n548,
    n451,
    n377,
    n412
  );


  xnor
  g525
  (
    n595,
    n391,
    n359,
    n430,
    n415
  );


  nand
  g526
  (
    n564,
    n390,
    n424,
    n446,
    n417
  );


  xor
  g527
  (
    n568,
    n452,
    n430,
    n433,
    n409
  );


  xor
  g528
  (
    n593,
    n429,
    n437,
    n382,
    n461
  );


  nand
  g529
  (
    n550,
    n400,
    n468,
    n450,
    n458
  );


  and
  g530
  (
    n626,
    n397,
    n453,
    n444,
    n414
  );


  or
  g531
  (
    n633,
    n448,
    n431,
    n437,
    n408
  );


  and
  g532
  (
    n567,
    n419,
    n427,
    n440,
    n435
  );


  xor
  g533
  (
    n631,
    n465,
    n375,
    n384,
    n364
  );


  or
  g534
  (
    n585,
    n380,
    n427,
    n402,
    n435
  );


  xor
  g535
  (
    n557,
    n468,
    n417,
    n437,
    n389
  );


  xnor
  g536
  (
    n609,
    n411,
    n462,
    n389,
    n386
  );


  xor
  g537
  (
    n632,
    n401,
    n426,
    n444,
    n411
  );


  nand
  g538
  (
    KeyWire_0_24,
    n466,
    n421,
    n402,
    n400
  );


  xnor
  g539
  (
    n629,
    n433,
    n452,
    n409,
    n422
  );


  nor
  g540
  (
    n628,
    n378,
    n433,
    n403,
    n394
  );


  xor
  g541
  (
    n542,
    n418,
    n433,
    n424,
    n380
  );


  or
  g542
  (
    n560,
    n438,
    n405,
    n439
  );


  nand
  g543
  (
    n575,
    n413,
    n393,
    n448,
    n417
  );


  nand
  g544
  (
    n549,
    n455,
    n431,
    n385,
    n412
  );


  or
  g545
  (
    n547,
    n439,
    n401,
    n463,
    n384
  );


  and
  g546
  (
    n592,
    n429,
    n442,
    n413,
    n454
  );


  nand
  g547
  (
    KeyWire_0_30,
    n457,
    n392,
    n361
  );


  and
  g548
  (
    n581,
    n468,
    n453,
    n455,
    n419
  );


  or
  g549
  (
    n544,
    n368,
    n464,
    n442,
    n414
  );


  or
  g550
  (
    n552,
    n459,
    n354,
    n444,
    n456
  );


  xnor
  g551
  (
    n555,
    n448,
    n439,
    n363,
    n406
  );


  nand
  g552
  (
    n602,
    n379,
    n412,
    n366,
    n467
  );


  nor
  g553
  (
    n584,
    n436,
    n419,
    n383,
    n430
  );


  xor
  g554
  (
    KeyWire_0_28,
    n424,
    n465,
    n463,
    n399
  );


  nand
  g555
  (
    n587,
    n428,
    n424,
    n436,
    n418
  );


  xor
  g556
  (
    n625,
    n436,
    n385,
    n447,
    n425
  );


  or
  g557
  (
    n556,
    n360,
    n390,
    n456,
    n410
  );


  xor
  g558
  (
    n627,
    n355,
    n402,
    n371,
    n409
  );


  xor
  g559
  (
    n623,
    n403,
    n457,
    n445,
    n447
  );


  nor
  g560
  (
    n607,
    n398,
    n451,
    n445,
    n453
  );


  or
  g561
  (
    n613,
    n461,
    n380,
    n422,
    n441
  );


  xnor
  g562
  (
    n589,
    n378,
    n404,
    n431,
    n447
  );


  nor
  g563
  (
    n591,
    n465,
    n386,
    n407,
    n443
  );


  nor
  g564
  (
    n571,
    n399,
    n446,
    n455,
    n434
  );


  xnor
  g565
  (
    n563,
    n383,
    n428,
    n465,
    n418
  );


  xor
  g566
  (
    n594,
    n428,
    n420,
    n426,
    n448
  );


  nor
  g567
  (
    KeyWire_0_8,
    n408,
    n395,
    n375,
    n427
  );


  nor
  g568
  (
    n611,
    n458,
    n464,
    n441,
    n383
  );


  or
  g569
  (
    n583,
    n454,
    n432,
    n442,
    n459
  );


  xor
  g570
  (
    n600,
    n392,
    n391,
    n367,
    n420
  );


  xor
  g571
  (
    n598,
    n415,
    n382,
    n405,
    n443
  );


  or
  g572
  (
    n630,
    n467,
    n386,
    n426,
    n460
  );


  nor
  g573
  (
    n624,
    n391,
    n464,
    n440,
    n421
  );


  nor
  g574
  (
    n539,
    n373,
    n410,
    n369,
    n454
  );


  and
  g575
  (
    n588,
    n459,
    n429,
    n439,
    n403
  );


  and
  g576
  (
    n619,
    n396,
    n461,
    n387,
    n388
  );


  and
  g577
  (
    n574,
    n422,
    n441,
    n416,
    n404
  );


  nor
  g578
  (
    n615,
    n450,
    n441,
    n462,
    n414
  );


  or
  g579
  (
    n553,
    n393,
    n435,
    n456,
    n449
  );


  xor
  g580
  (
    n605,
    n402,
    n416,
    n431,
    n462
  );


  nand
  g581
  (
    n604,
    n451,
    n421,
    n454,
    n417
  );


  xnor
  g582
  (
    n570,
    n420,
    n395,
    n418,
    n466
  );


  nor
  g583
  (
    n580,
    n404,
    n464,
    n423,
    n422
  );


  xor
  g584
  (
    n577,
    n388,
    n466,
    n394,
    n376
  );


  xor
  g585
  (
    n569,
    n407,
    n397,
    n410,
    n423
  );


  nand
  g586
  (
    n616,
    n438,
    n430,
    n442,
    n421
  );


  or
  g587
  (
    n558,
    n400,
    n446,
    n445,
    n413
  );


  xor
  g588
  (
    n617,
    n411,
    n458,
    n396,
    n434
  );


  nand
  g589
  (
    n621,
    n375,
    n381,
    n468,
    n387
  );


  xnor
  g590
  (
    n610,
    n438,
    n404,
    n395,
    n428
  );


  or
  g591
  (
    n608,
    n388,
    n444,
    n377,
    n370
  );


  nand
  g592
  (
    n601,
    n411,
    n401,
    n447,
    n457
  );


  nand
  g593
  (
    n562,
    n453,
    n419,
    n374,
    n427
  );


  xnor
  g594
  (
    n586,
    n408,
    n460,
    n400,
    n432
  );


  xnor
  g595
  (
    n596,
    n393,
    n451,
    n381
  );


  or
  g596
  (
    n554,
    n434,
    n403,
    n455,
    n384
  );


  and
  g597
  (
    n566,
    n456,
    n438,
    n372,
    n406
  );


  nand
  g598
  (
    n573,
    n449,
    n432,
    n458,
    n379
  );


  xor
  g599
  (
    n578,
    n462,
    n387,
    n407,
    n467
  );


  xor
  g600
  (
    n572,
    n423,
    n379,
    n409,
    n425
  );


  or
  g601
  (
    n651,
    n544,
    n545,
    n556,
    n546
  );


  nand
  g602
  (
    n669,
    n552,
    n573,
    n574,
    n547
  );


  nand
  g603
  (
    n658,
    n568,
    n572,
    n566,
    n540
  );


  xor
  g604
  (
    n646,
    n566,
    n549,
    n583,
    n584
  );


  xnor
  g605
  (
    n647,
    n561,
    n576,
    n559,
    n572
  );


  nand
  g606
  (
    n644,
    n571,
    n562,
    n578
  );


  nand
  g607
  (
    n639,
    n557,
    n544,
    n581,
    n576
  );


  nor
  g608
  (
    n673,
    n573,
    n583,
    n542
  );


  xnor
  g609
  (
    n635,
    n578,
    n547,
    n554,
    n551
  );


  nand
  g610
  (
    n637,
    n555,
    n554,
    n552,
    n543
  );


  xor
  g611
  (
    n642,
    n544,
    n567,
    n580,
    n543
  );


  and
  g612
  (
    n660,
    n581,
    n550,
    n579,
    n573
  );


  xnor
  g613
  (
    n667,
    n583,
    n546,
    n584,
    n575
  );


  xnor
  g614
  (
    KeyWire_0_1,
    n577,
    n545,
    n547,
    n578
  );


  nand
  g615
  (
    n643,
    n568,
    n580,
    n574,
    n586
  );


  and
  g616
  (
    n656,
    n566,
    n586,
    n559,
    n553
  );


  and
  g617
  (
    n671,
    n576,
    n552,
    n574,
    n577
  );


  or
  g618
  (
    n655,
    n560,
    n545,
    n576,
    n567
  );


  xor
  g619
  (
    n670,
    n584,
    n542,
    n565,
    n548
  );


  and
  g620
  (
    n638,
    n554,
    n540,
    n568,
    n569
  );


  nor
  g621
  (
    n679,
    n557,
    n560,
    n564
  );


  and
  g622
  (
    n654,
    n541,
    n548,
    n562,
    n570
  );


  xor
  g623
  (
    n645,
    n556,
    n563,
    n555,
    n566
  );


  and
  g624
  (
    n650,
    n559,
    n561,
    n545,
    n579
  );


  xor
  g625
  (
    n652,
    n563,
    n577,
    n582,
    n550
  );


  and
  g626
  (
    n675,
    n549,
    n574,
    n560,
    n550
  );


  and
  g627
  (
    n636,
    n540,
    n549,
    n557,
    n555
  );


  nand
  g628
  (
    n663,
    n558,
    n584,
    n569
  );


  nor
  g629
  (
    n668,
    n565,
    n585,
    n553
  );


  nand
  g630
  (
    n648,
    n586,
    n585,
    n570,
    n563
  );


  xnor
  g631
  (
    n672,
    n552,
    n565,
    n579,
    n562
  );


  nand
  g632
  (
    n666,
    n544,
    n551,
    n582,
    n564
  );


  nand
  g633
  (
    n657,
    n577,
    n541,
    n580
  );


  nor
  g634
  (
    n662,
    n580,
    n571,
    n561,
    n582
  );


  and
  g635
  (
    n665,
    n543,
    n575,
    n583,
    n547
  );


  xnor
  g636
  (
    n674,
    n560,
    n567,
    n541,
    n571
  );


  xor
  g637
  (
    n659,
    n558,
    n558,
    n546,
    n553
  );


  and
  g638
  (
    n680,
    n570,
    n585,
    n553,
    n548
  );


  nor
  g639
  (
    n676,
    n581,
    n570,
    n565,
    n572
  );


  xnor
  g640
  (
    n678,
    n572,
    n575,
    n567,
    n586
  );


  or
  g641
  (
    KeyWire_0_17,
    n549,
    n579,
    n578,
    n581
  );


  nor
  g642
  (
    n641,
    n561,
    n551,
    n563,
    n556
  );


  and
  g643
  (
    n677,
    n551,
    n569,
    n542,
    n558
  );


  nand
  g644
  (
    n661,
    n557,
    n582,
    n556,
    n550
  );


  and
  g645
  (
    n649,
    n564,
    n539,
    n554,
    n546
  );


  and
  g646
  (
    n664,
    n568,
    n548,
    n559,
    n575
  );


  and
  g647
  (
    n640,
    n555,
    n543,
    n571,
    n573
  );


  and
  g648
  (
    n736,
    n346,
    n510,
    n485
  );


  xnor
  g649
  (
    n745,
    n522,
    n644,
    n654
  );


  nand
  g650
  (
    n694,
    n483,
    n651,
    n674
  );


  xor
  g651
  (
    n724,
    n488,
    n510,
    n346
  );


  nand
  g652
  (
    n689,
    n640,
    n492
  );


  xnor
  g653
  (
    n771,
    n641,
    n643,
    n501
  );


  and
  g654
  (
    n703,
    n512,
    n523,
    n661
  );


  nor
  g655
  (
    n684,
    n509,
    n672,
    n513
  );


  nor
  g656
  (
    n787,
    n491,
    n653,
    n517
  );


  xnor
  g657
  (
    n722,
    n472,
    n673,
    n667
  );


  nand
  g658
  (
    n710,
    n348,
    n641,
    n665
  );


  xnor
  g659
  (
    n693,
    n522,
    n657,
    n348
  );


  nand
  g660
  (
    n698,
    n646,
    n504,
    n353
  );


  and
  g661
  (
    n696,
    n514,
    n491,
    n653
  );


  and
  g662
  (
    n768,
    n649,
    n496,
    n350
  );


  nor
  g663
  (
    n761,
    n349,
    n659,
    n483
  );


  nor
  g664
  (
    n730,
    n508,
    n498,
    n470
  );


  and
  g665
  (
    n692,
    n472,
    n484,
    n518
  );


  nor
  g666
  (
    n723,
    n480,
    n486,
    n471
  );


  xor
  g667
  (
    n741,
    n475,
    n498,
    n645
  );


  nor
  g668
  (
    n720,
    n511,
    n646,
    n489
  );


  nor
  g669
  (
    n794,
    n657,
    n505,
    n635
  );


  nand
  g670
  (
    n721,
    n640,
    n509,
    n661
  );


  nand
  g671
  (
    n731,
    n639,
    n485,
    n664
  );


  xnor
  g672
  (
    n773,
    n347,
    n511,
    n642
  );


  nor
  g673
  (
    n712,
    n478,
    n668,
    n649
  );


  or
  g674
  (
    n789,
    n658,
    n666,
    n522
  );


  nand
  g675
  (
    n738,
    n668,
    n636,
    n671
  );


  or
  g676
  (
    n701,
    n667,
    n480,
    n657
  );


  xnor
  g677
  (
    n708,
    n476,
    n507,
    n349
  );


  and
  g678
  (
    n718,
    n654,
    n656,
    n653
  );


  or
  g679
  (
    n681,
    n474,
    n520,
    n501
  );


  nand
  g680
  (
    n779,
    n524,
    n646,
    n676
  );


  and
  g681
  (
    n759,
    n666,
    n668,
    n523
  );


  xnor
  g682
  (
    n733,
    n490,
    n651,
    n493
  );


  and
  g683
  (
    n797,
    n650,
    n525,
    n469
  );


  or
  g684
  (
    n739,
    n505,
    n651,
    n473
  );


  nor
  g685
  (
    n780,
    n472,
    n658,
    n521
  );


  xor
  g686
  (
    n749,
    n511,
    n643
  );


  or
  g687
  (
    n735,
    n519,
    n495,
    n507
  );


  xor
  g688
  (
    n752,
    n513,
    n525,
    n669
  );


  and
  g689
  (
    n753,
    n523,
    n346,
    n512
  );


  nand
  g690
  (
    n782,
    n352,
    n638,
    n487
  );


  or
  g691
  (
    n763,
    n519,
    n492,
    n472
  );


  and
  g692
  (
    n747,
    n483,
    n347,
    n644,
    n351
  );


  nand
  g693
  (
    KeyWire_0_21,
    n639,
    n641,
    n507,
    n636
  );


  or
  g694
  (
    n740,
    n497,
    n479,
    n635,
    n511
  );


  xor
  g695
  (
    n772,
    n481,
    n482,
    n515,
    n649
  );


  nor
  g696
  (
    n695,
    n496,
    n642,
    n500,
    n659
  );


  nor
  g697
  (
    n777,
    n510,
    n503,
    n516,
    n660
  );


  xor
  g698
  (
    n713,
    n508,
    n493,
    n495,
    n350
  );


  nand
  g699
  (
    n778,
    n665,
    n504,
    n674,
    n643
  );


  nor
  g700
  (
    n767,
    n666,
    n647,
    n508,
    n481
  );


  xor
  g701
  (
    n742,
    n352,
    n474,
    n644,
    n673
  );


  xor
  g702
  (
    n748,
    n659,
    n673,
    n674,
    n657
  );


  or
  g703
  (
    n715,
    n491,
    n656,
    n349,
    n676
  );


  or
  g704
  (
    n783,
    n637,
    n514,
    n485,
    n500
  );


  xnor
  g705
  (
    n727,
    n489,
    n669,
    n524,
    n508
  );


  nor
  g706
  (
    n691,
    n675,
    n524,
    n638,
    n351
  );


  and
  g707
  (
    n683,
    n498,
    n654,
    n471,
    n487
  );


  nand
  g708
  (
    n682,
    n479,
    n475,
    n353,
    n658
  );


  xnor
  g709
  (
    n756,
    n488,
    n493,
    n518,
    n523
  );


  xor
  g710
  (
    n781,
    n499,
    n501,
    n513,
    n662
  );


  and
  g711
  (
    n769,
    n512,
    n487,
    n503,
    n496
  );


  nand
  g712
  (
    n757,
    n514,
    n652,
    n478,
    n672
  );


  nand
  g713
  (
    n786,
    n647,
    n485,
    n634,
    n348
  );


  xnor
  g714
  (
    n766,
    n667,
    n670,
    n473,
    n502
  );


  xnor
  g715
  (
    n776,
    n503,
    n479,
    n667,
    n639
  );


  or
  g716
  (
    n743,
    n517,
    n350,
    n656,
    n484
  );


  xor
  g717
  (
    n704,
    n494,
    n671,
    n473,
    n652
  );


  nand
  g718
  (
    n798,
    n517,
    n655,
    n651,
    n514
  );


  nor
  g719
  (
    n716,
    n486,
    n491,
    n506,
    n672
  );


  nor
  g720
  (
    n788,
    n663,
    n650,
    n635,
    n470
  );


  nand
  g721
  (
    n726,
    n521,
    n647,
    n645,
    n493
  );


  nand
  g722
  (
    n750,
    n655,
    n471,
    n496,
    n671
  );


  and
  g723
  (
    n754,
    n637,
    n500,
    n478,
    n513
  );


  nand
  g724
  (
    n728,
    n640,
    n469,
    n516,
    n490
  );


  nor
  g725
  (
    n795,
    n645,
    n636,
    n515,
    n646
  );


  xnor
  g726
  (
    n758,
    n518,
    n478,
    n648,
    n504
  );


  nand
  g727
  (
    n770,
    n515,
    n637,
    n502,
    n505
  );


  or
  g728
  (
    n793,
    n494,
    n510,
    n353,
    n675
  );


  xnor
  g729
  (
    n717,
    n495,
    n642,
    n351,
    n669
  );


  and
  g730
  (
    n792,
    n661,
    n518,
    n477,
    n673
  );


  nor
  g731
  (
    n706,
    n660,
    n473,
    n500,
    n509
  );


  nand
  g732
  (
    n732,
    n494,
    n480,
    n484,
    n671
  );


  and
  g733
  (
    n765,
    n658,
    n346,
    n664,
    n353
  );


  nand
  g734
  (
    n790,
    n489,
    n504,
    n497,
    n498
  );


  nor
  g735
  (
    KeyWire_0_26,
    n652,
    n519,
    n672,
    n488
  );


  xor
  g736
  (
    n737,
    n664,
    n674,
    n648,
    n470
  );


  nor
  g737
  (
    n744,
    n469,
    n477,
    n634,
    n675
  );


  xor
  g738
  (
    n725,
    n642,
    n635,
    n668,
    n502
  );


  nand
  g739
  (
    n686,
    n516,
    n486,
    n499,
    n347
  );


  nor
  g740
  (
    KeyWire_0_18,
    n497,
    n664,
    n638,
    n506
  );


  or
  g741
  (
    n709,
    n516,
    n479,
    n512,
    n524
  );


  xnor
  g742
  (
    n702,
    n515,
    n475,
    n520,
    n650
  );


  xnor
  g743
  (
    n687,
    n525,
    n499,
    n648,
    n475
  );


  nor
  g744
  (
    n760,
    n640,
    n495,
    n351,
    n492
  );


  xnor
  g745
  (
    n719,
    n645,
    n347,
    n644,
    n655
  );


  nor
  g746
  (
    n746,
    n637,
    n648,
    n647,
    n476
  );


  xor
  g747
  (
    n711,
    n497,
    n670,
    n639,
    n654
  );


  xor
  g748
  (
    n799,
    n675,
    n525,
    n474,
    n521
  );


  nand
  g749
  (
    n688,
    n503,
    n663,
    n659,
    n483
  );


  xor
  g750
  (
    n796,
    n476,
    n676,
    n477,
    n470
  );


  or
  g751
  (
    n774,
    n490,
    n480,
    n506,
    n469
  );


  nor
  g752
  (
    n762,
    n522,
    n352,
    n666,
    n482
  );


  and
  g753
  (
    n755,
    n520,
    n526,
    n349,
    n655
  );


  nand
  g754
  (
    n791,
    n519,
    n490,
    n517,
    n499
  );


  and
  g755
  (
    n697,
    n638,
    n484,
    n634,
    n482
  );


  xor
  g756
  (
    KeyWire_0_6,
    n650,
    n476,
    n348,
    n663
  );


  nand
  g757
  (
    n784,
    n507,
    n660,
    n501,
    n481
  );


  and
  g758
  (
    n700,
    n636,
    n488,
    n481,
    n661
  );


  xnor
  g759
  (
    n775,
    n489,
    n474,
    n653,
    n662
  );


  or
  g760
  (
    n705,
    n486,
    n665,
    n471,
    n502
  );


  or
  g761
  (
    n764,
    n663,
    n521,
    n641,
    n669
  );


  xor
  g762
  (
    n685,
    n487,
    n652,
    n665,
    n352
  );


  nor
  g763
  (
    n729,
    n350,
    n662,
    n649,
    n656
  );


  nor
  g764
  (
    n699,
    n505,
    n506,
    n662,
    n494
  );


  xnor
  g765
  (
    n707,
    n509,
    n634,
    n482,
    n660
  );


  xnor
  g766
  (
    n785,
    n520,
    n670,
    n477
  );


  nor
  g767
  (
    n829,
    n716,
    n771,
    n762,
    n759
  );


  or
  g768
  (
    n922,
    n591,
    n799,
    n796,
    n721
  );


  and
  g769
  (
    n859,
    n526,
    n692,
    n734,
    n713
  );


  or
  g770
  (
    n824,
    n753,
    n745,
    n714,
    n699
  );


  or
  g771
  (
    n813,
    n742,
    n754,
    n769,
    n770
  );


  xor
  g772
  (
    n814,
    n792,
    n776,
    n781,
    n590
  );


  or
  g773
  (
    n907,
    n769,
    n692,
    n771,
    n763
  );


  nor
  g774
  (
    n877,
    n690,
    n756,
    n783,
    n781
  );


  xor
  g775
  (
    n863,
    n776,
    n719,
    n731,
    n779
  );


  or
  g776
  (
    n856,
    n726,
    n744,
    n716,
    n697
  );


  nand
  g777
  (
    n895,
    n796,
    n730,
    n702,
    n729
  );


  and
  g778
  (
    n812,
    n703,
    n774,
    n732,
    n765
  );


  nand
  g779
  (
    n850,
    n775,
    n798,
    n765,
    n723
  );


  xor
  g780
  (
    n888,
    n685,
    n715,
    n745,
    n728
  );


  or
  g781
  (
    n876,
    n757,
    n784,
    n690,
    n791
  );


  nor
  g782
  (
    n900,
    n768,
    n775,
    n697,
    n705
  );


  nor
  g783
  (
    n828,
    n736,
    n743,
    n778,
    n691
  );


  nand
  g784
  (
    n887,
    n590,
    n723,
    n693,
    n772
  );


  xor
  g785
  (
    n866,
    n771,
    n698,
    n735,
    n711
  );


  or
  g786
  (
    n896,
    n747,
    n725,
    n683,
    n778
  );


  xnor
  g787
  (
    KeyWire_0_0,
    n682,
    n724,
    n733,
    n720
  );


  and
  g788
  (
    n830,
    n789,
    n717,
    n792,
    n767
  );


  nor
  g789
  (
    n911,
    n737,
    n730,
    n715,
    n718
  );


  xnor
  g790
  (
    n847,
    n588,
    n588,
    n750,
    n741
  );


  xor
  g791
  (
    n878,
    n720,
    n789,
    n793,
    n698
  );


  xnor
  g792
  (
    n848,
    n791,
    n716,
    n711,
    n794
  );


  nor
  g793
  (
    n916,
    n695,
    n712,
    n691,
    n749
  );


  nor
  g794
  (
    n890,
    n693,
    n779,
    n721,
    n689
  );


  nand
  g795
  (
    n831,
    n762,
    n738,
    n708,
    n683
  );


  nand
  g796
  (
    n919,
    n706,
    n755,
    n780,
    n784
  );


  nand
  g797
  (
    n827,
    n757,
    n752,
    n713,
    n731
  );


  nor
  g798
  (
    n899,
    n710,
    n691,
    n762,
    n780
  );


  nor
  g799
  (
    n864,
    n698,
    n721,
    n780,
    n797
  );


  xor
  g800
  (
    n903,
    n715,
    n777,
    n687,
    n765
  );


  nor
  g801
  (
    n879,
    n728,
    n681,
    n785
  );


  nor
  g802
  (
    n815,
    n751,
    n735,
    n684,
    n700
  );


  xor
  g803
  (
    n811,
    n682,
    n728,
    n782,
    n711
  );


  xnor
  g804
  (
    n868,
    n716,
    n776,
    n789,
    n689
  );


  or
  g805
  (
    n867,
    n737,
    n776,
    n784,
    n704
  );


  xor
  g806
  (
    n817,
    n752,
    n732,
    n714,
    n760
  );


  nor
  g807
  (
    n897,
    n692,
    n686,
    n694,
    n741
  );


  nor
  g808
  (
    n885,
    n591,
    n722,
    n745,
    n730
  );


  and
  g809
  (
    n825,
    n717,
    n708,
    n782,
    n684
  );


  nand
  g810
  (
    n838,
    n686,
    n790,
    n729,
    n783
  );


  nor
  g811
  (
    n915,
    n709,
    n587,
    n727,
    n769
  );


  xnor
  g812
  (
    n912,
    n727,
    n589,
    n777,
    n791
  );


  or
  g813
  (
    n892,
    n785,
    n703,
    n701,
    n794
  );


  nand
  g814
  (
    n803,
    n701,
    n722,
    n699,
    n760
  );


  xnor
  g815
  (
    n883,
    n591,
    n736,
    n749,
    n696
  );


  xnor
  g816
  (
    n834,
    n755,
    n739,
    n693,
    n698
  );


  xnor
  g817
  (
    n906,
    n713,
    n787,
    n797,
    n757
  );


  xnor
  g818
  (
    n875,
    n685,
    n759,
    n739,
    n756
  );


  and
  g819
  (
    n881,
    n704,
    n745,
    n701,
    n736
  );


  xnor
  g820
  (
    n886,
    n795,
    n686,
    n765,
    n699
  );


  and
  g821
  (
    n901,
    n734,
    n767,
    n792,
    n756
  );


  nor
  g822
  (
    n893,
    n681,
    n687,
    n706,
    n742
  );


  xor
  g823
  (
    n839,
    n761,
    n799,
    n712,
    n749
  );


  nand
  g824
  (
    n820,
    n696,
    n744,
    n782,
    n682
  );


  nor
  g825
  (
    n874,
    n683,
    n718,
    n743,
    n703
  );


  nand
  g826
  (
    n908,
    n707,
    n683,
    n783,
    n794
  );


  xnor
  g827
  (
    n869,
    n795,
    n690,
    n694,
    n793
  );


  or
  g828
  (
    n894,
    n709,
    n587,
    n733,
    n722
  );


  or
  g829
  (
    n823,
    n751,
    n732,
    n777,
    n747
  );


  and
  g830
  (
    n826,
    n748,
    n694,
    n749,
    n781
  );


  or
  g831
  (
    n855,
    n748,
    n798,
    n782,
    n723
  );


  xnor
  g832
  (
    n843,
    n724,
    n739,
    n710,
    n753
  );


  and
  g833
  (
    n810,
    n763,
    n705,
    n797,
    n790
  );


  nor
  g834
  (
    n818,
    n748,
    n688,
    n589,
    n744
  );


  xnor
  g835
  (
    n909,
    n708,
    n777,
    n718,
    n692
  );


  nor
  g836
  (
    n821,
    n739,
    n705,
    n707,
    n715
  );


  and
  g837
  (
    n905,
    n706,
    n689,
    n774,
    n755
  );


  nand
  g838
  (
    n918,
    n773,
    n734,
    n766,
    n763
  );


  xor
  g839
  (
    n805,
    n746,
    n751,
    n720,
    n772
  );


  or
  g840
  (
    n802,
    n704,
    n588,
    n685,
    n725
  );


  or
  g841
  (
    n872,
    n697,
    n733,
    n767,
    n787
  );


  or
  g842
  (
    n837,
    n766,
    n778,
    n725,
    n729
  );


  xor
  g843
  (
    n920,
    n740,
    n769,
    n795,
    n731
  );


  xnor
  g844
  (
    n889,
    n695,
    n710,
    n719,
    n721
  );


  nor
  g845
  (
    n832,
    n790,
    n764,
    n714,
    n768
  );


  or
  g846
  (
    n854,
    n746,
    n772,
    n751,
    n754
  );


  nor
  g847
  (
    n845,
    n726,
    n790,
    n740,
    n701
  );


  xor
  g848
  (
    n853,
    n796,
    n735,
    n788,
    n741
  );


  or
  g849
  (
    n914,
    n699,
    n743,
    n727,
    n738
  );


  nor
  g850
  (
    n835,
    n794,
    n770,
    n757,
    n696
  );


  or
  g851
  (
    n870,
    n737,
    n764,
    n717,
    n693
  );


  nor
  g852
  (
    n816,
    n742,
    n750,
    n746,
    n768
  );


  and
  g853
  (
    n884,
    n764,
    n732,
    n587,
    n754
  );


  xnor
  g854
  (
    KeyWire_0_27,
    n785,
    n711,
    n799,
    n725
  );


  nor
  g855
  (
    n923,
    n727,
    n728,
    n773,
    n755
  );


  nand
  g856
  (
    n860,
    n707,
    n710,
    n696,
    n752
  );


  xor
  g857
  (
    n822,
    n761,
    n722,
    n589,
    n774
  );


  nand
  g858
  (
    n902,
    n750,
    n781,
    n686,
    n738
  );


  nand
  g859
  (
    n851,
    n759,
    n775,
    n724,
    n700
  );


  xor
  g860
  (
    n891,
    n799,
    n786,
    n759,
    n590
  );


  nand
  g861
  (
    n836,
    n753,
    n719,
    n736,
    n587
  );


  xor
  g862
  (
    n801,
    n787,
    n787,
    n720,
    n797
  );


  xor
  g863
  (
    n800,
    n754,
    n793,
    n764,
    n791
  );


  and
  g864
  (
    n804,
    n752,
    n684,
    n767,
    n798
  );


  xnor
  g865
  (
    n833,
    n700,
    n702,
    n712,
    n766
  );


  nor
  g866
  (
    n844,
    n763,
    n703,
    n775,
    n688
  );


  and
  g867
  (
    n857,
    n729,
    n695,
    n774,
    n684
  );


  or
  g868
  (
    n898,
    n713,
    n706,
    n768,
    n770
  );


  and
  g869
  (
    n840,
    n718,
    n786,
    n726,
    n734
  );


  nor
  g870
  (
    n904,
    n730,
    n760,
    n779,
    n788
  );


  and
  g871
  (
    n852,
    n771,
    n694,
    n750,
    n762
  );


  xnor
  g872
  (
    n862,
    n695,
    n687,
    n778,
    n784
  );


  or
  g873
  (
    n849,
    n786,
    n795,
    n743,
    n773
  );


  nor
  g874
  (
    n807,
    n588,
    n702,
    n697,
    n753
  );


  nor
  g875
  (
    n913,
    n798,
    n591,
    n758,
    n726
  );


  or
  g876
  (
    n917,
    n772,
    n773,
    n779,
    n761
  );


  or
  g877
  (
    KeyWire_0_7,
    n780,
    n789,
    n760,
    n758
  );


  xor
  g878
  (
    n808,
    n788,
    n682,
    n738,
    n761
  );


  xor
  g879
  (
    n842,
    n724,
    n704,
    n756,
    n681
  );


  nand
  g880
  (
    n880,
    n709,
    n709,
    n714,
    n689
  );


  xnor
  g881
  (
    n819,
    n758,
    n712,
    n733,
    n691
  );


  xnor
  g882
  (
    n865,
    n705,
    n740,
    n793,
    n685
  );


  xor
  g883
  (
    n809,
    n747,
    n702,
    n700,
    n687
  );


  nand
  g884
  (
    n861,
    n792,
    n719,
    n688,
    n747
  );


  or
  g885
  (
    n910,
    n707,
    n589,
    n748,
    n590
  );


  nor
  g886
  (
    n858,
    n723,
    n766,
    n688,
    n731
  );


  and
  g887
  (
    n873,
    n741,
    n740,
    n735,
    n770
  );


  xor
  g888
  (
    n871,
    n788,
    n717,
    n708,
    n783
  );


  nor
  g889
  (
    n882,
    n690,
    n746,
    n742,
    n796
  );


  nor
  g890
  (
    n806,
    n744,
    n737,
    n758,
    n786
  );


  nor
  g891
  (
    n975,
    n677,
    n529,
    n906,
    n624
  );


  xnor
  g892
  (
    n1002,
    n921,
    n838,
    n828,
    n678
  );


  or
  g893
  (
    n989,
    n916,
    n887,
    n629,
    n530
  );


  xnor
  g894
  (
    n965,
    n678,
    n619,
    n532,
    n898
  );


  and
  g895
  (
    n958,
    n604,
    n537,
    n530,
    n593
  );


  and
  g896
  (
    n941,
    n592,
    n532,
    n835,
    n537
  );


  xor
  g897
  (
    n940,
    n830,
    n619,
    n892,
    n596
  );


  or
  g898
  (
    n932,
    n533,
    n883,
    n536,
    n623
  );


  xnor
  g899
  (
    n972,
    n615,
    n620,
    n902,
    n531
  );


  or
  g900
  (
    n938,
    n613,
    n864,
    n604,
    n600
  );


  or
  g901
  (
    n935,
    n538,
    n856,
    n615,
    n891
  );


  nand
  g902
  (
    n939,
    n629,
    n612,
    n628,
    n602
  );


  nor
  g903
  (
    n1001,
    n923,
    n908,
    n530,
    n831
  );


  and
  g904
  (
    n998,
    n594,
    n848,
    n592,
    n536
  );


  nand
  g905
  (
    n980,
    n603,
    n617,
    n911,
    n600
  );


  or
  g906
  (
    n931,
    n599,
    n615,
    n626,
    n608
  );


  nor
  g907
  (
    n990,
    n619,
    n622,
    n530,
    n534
  );


  or
  g908
  (
    n1000,
    n623,
    n592,
    n910,
    n622
  );


  or
  g909
  (
    n945,
    n875,
    n836,
    n536,
    n680
  );


  xor
  g910
  (
    n952,
    n531,
    n612,
    n877,
    n619
  );


  xor
  g911
  (
    n963,
    n867,
    n609,
    n597,
    n919
  );


  xor
  g912
  (
    n971,
    n628,
    n605,
    n617,
    n595
  );


  xor
  g913
  (
    KeyWire_0_3,
    n533,
    n628,
    n529,
    n535
  );


  nor
  g914
  (
    n930,
    n680,
    n677,
    n839,
    n593
  );


  xnor
  g915
  (
    n992,
    n614,
    n608,
    n625,
    n872
  );


  and
  g916
  (
    n997,
    n677,
    n621,
    n600,
    n611
  );


  or
  g917
  (
    n984,
    n614,
    n598,
    n677,
    n844
  );


  and
  g918
  (
    n981,
    n869,
    n881,
    n534,
    n625
  );


  xor
  g919
  (
    n996,
    n676,
    n596,
    n901,
    n595
  );


  nand
  g920
  (
    n955,
    n611,
    n832,
    n890,
    n871
  );


  xnor
  g921
  (
    KeyWire_0_5,
    n618,
    n527,
    n626,
    n627
  );


  nand
  g922
  (
    n927,
    n538,
    n620,
    n629
  );


  or
  g923
  (
    KeyWire_0_2,
    n873,
    n907,
    n616,
    n678
  );


  xnor
  g924
  (
    n926,
    n857,
    n528,
    n598,
    n601
  );


  and
  g925
  (
    n994,
    n526,
    n605,
    n528,
    n603
  );


  or
  g926
  (
    n951,
    n594,
    n847,
    n621,
    n897
  );


  nor
  g927
  (
    n979,
    n599,
    n863,
    n886,
    n879
  );


  nor
  g928
  (
    n960,
    n833,
    n614,
    n628,
    n920
  );


  xnor
  g929
  (
    n943,
    n613,
    n528,
    n837,
    n827
  );


  xnor
  g930
  (
    n973,
    n840,
    n882,
    n531,
    n870
  );


  and
  g931
  (
    n999,
    n611,
    n621,
    n627,
    n603
  );


  nor
  g932
  (
    n933,
    n533,
    n680,
    n889,
    n878
  );


  xor
  g933
  (
    n956,
    n626,
    n826,
    n627,
    n594
  );


  or
  g934
  (
    n928,
    n915,
    n612,
    n845,
    n617
  );


  nor
  g935
  (
    n924,
    n606,
    n605,
    n842,
    n527
  );


  and
  g936
  (
    n944,
    n623,
    n593,
    n609,
    n884
  );


  xor
  g937
  (
    n957,
    n903,
    n853,
    n599,
    n593
  );


  nor
  g938
  (
    n986,
    n528,
    n529,
    n874,
    n535
  );


  xor
  g939
  (
    n966,
    n606,
    n904,
    n625,
    n607
  );


  nand
  g940
  (
    n953,
    n860,
    n538,
    n855
  );


  or
  g941
  (
    n947,
    n598,
    n913,
    n834,
    n613
  );


  nor
  g942
  (
    n976,
    n829,
    n602,
    n532,
    n599
  );


  xnor
  g943
  (
    n969,
    n606,
    n597,
    n533,
    n680
  );


  or
  g944
  (
    n946,
    n598,
    n620,
    n885,
    n527
  );


  xor
  g945
  (
    n978,
    n609,
    n601,
    n862,
    n597
  );


  xor
  g946
  (
    n983,
    n917,
    n621,
    n529,
    n608
  );


  or
  g947
  (
    KeyWire_0_25,
    n880,
    n678,
    n909,
    n622
  );


  xnor
  g948
  (
    KeyWire_0_16,
    n859,
    n535,
    n613,
    n861
  );


  xnor
  g949
  (
    n954,
    n900,
    n618,
    n604,
    n610
  );


  or
  g950
  (
    n991,
    n914,
    n600,
    n624,
    n618
  );


  or
  g951
  (
    n948,
    n609,
    n602,
    n597,
    n624
  );


  xnor
  g952
  (
    n942,
    n602,
    n679,
    n868,
    n858
  );


  and
  g953
  (
    n949,
    n627,
    n626,
    n596,
    n866
  );


  nand
  g954
  (
    n937,
    n604,
    n607,
    n851,
    n537
  );


  nand
  g955
  (
    n968,
    n592,
    n854,
    n679,
    n618
  );


  and
  g956
  (
    n934,
    n625,
    n624,
    n610,
    n536
  );


  nor
  g957
  (
    n995,
    n623,
    n531,
    n841,
    n899
  );


  xnor
  g958
  (
    n985,
    n534,
    n876,
    n679,
    n526
  );


  nor
  g959
  (
    n961,
    n606,
    n616,
    n605,
    n595
  );


  and
  g960
  (
    n925,
    n601,
    n603,
    n615,
    n895
  );


  nand
  g961
  (
    n950,
    n527,
    n614,
    n610
  );


  nand
  g962
  (
    n970,
    n893,
    n532,
    n607,
    n918
  );


  and
  g963
  (
    n967,
    n846,
    n535,
    n894,
    n617
  );


  nand
  g964
  (
    n929,
    n608,
    n534,
    n888,
    n595
  );


  nor
  g965
  (
    n974,
    n905,
    n843,
    n611,
    n616
  );


  nand
  g966
  (
    n962,
    n896,
    n612,
    n537,
    n616
  );


  and
  g967
  (
    n936,
    n849,
    n865,
    n922,
    n594
  );


  or
  g968
  (
    n987,
    n601,
    n850,
    n679,
    n596
  );


  and
  g969
  (
    n977,
    n607,
    n912,
    n852,
    n622
  );


  or
  g970
  (
    n1005,
    n961,
    n994,
    n969,
    n633
  );


  xnor
  g971
  (
    n1022,
    n632,
    n938,
    n987,
    n976
  );


  or
  g972
  (
    n1018,
    n630,
    n956,
    n943,
    n989
  );


  nand
  g973
  (
    n1015,
    n930,
    n629,
    n931,
    n940
  );


  xnor
  g974
  (
    n1020,
    n632,
    n949,
    n925,
    n966
  );


  nand
  g975
  (
    n1004,
    n937,
    n630,
    n983,
    n953
  );


  xor
  g976
  (
    n1025,
    n960,
    n996,
    n947,
    n995
  );


  and
  g977
  (
    n1003,
    n979,
    n941,
    n984,
    n993
  );


  xor
  g978
  (
    n1023,
    n973,
    n1002,
    n992,
    n928
  );


  nand
  g979
  (
    n1008,
    n630,
    n952,
    n631,
    n632
  );


  or
  g980
  (
    n1013,
    n967,
    n939,
    n998,
    n631
  );


  or
  g981
  (
    n1026,
    n942,
    n997,
    n633,
    n946
  );


  xor
  g982
  (
    n1024,
    n929,
    n968,
    n631,
    n999
  );


  nor
  g983
  (
    n1014,
    n633,
    n932,
    n927,
    n632
  );


  nand
  g984
  (
    n1012,
    n965,
    n990,
    n1000,
    n958
  );


  or
  g985
  (
    n1017,
    n954,
    n944,
    n948,
    n991
  );


  nand
  g986
  (
    n1019,
    n631,
    n972,
    n977,
    n936
  );


  nand
  g987
  (
    n1016,
    n955,
    n935,
    n951,
    n982
  );


  xnor
  g988
  (
    n1007,
    n959,
    n981,
    n986,
    n950
  );


  or
  g989
  (
    n1009,
    n988,
    n926,
    n974,
    n985
  );


  xnor
  g990
  (
    n1006,
    n633,
    n934,
    n933,
    n971
  );


  xor
  g991
  (
    n1011,
    n1001,
    n945,
    n964,
    n978
  );


  nor
  g992
  (
    n1021,
    n962,
    n975,
    n980,
    n957
  );


  and
  g993
  (
    n1010,
    n970,
    n924,
    n963,
    n630
  );


  xnor
  g994
  (
    n1028,
    n1018,
    n1026,
    n1008,
    n1024
  );


  nor
  g995
  (
    n1030,
    n1012,
    n1016,
    n1005,
    n1019
  );


  xor
  g996
  (
    n1032,
    n1021,
    n1009,
    n1017,
    n1004
  );


  xor
  g997
  (
    n1027,
    n1025,
    n1003,
    n1006,
    n1010
  );


  and
  g998
  (
    n1031,
    n1015,
    n1022,
    n1011,
    n1014
  );


  and
  g999
  (
    n1029,
    n1023,
    n1020,
    n1007,
    n1013
  );


  xnor
  KeyGate_0_0
  (
    n846,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n653,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n959,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n988,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n540,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n993,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n734,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n841,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n545,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n293,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n390,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n520,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n79,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n326,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n389,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n147,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n982,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n634,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n751,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n172,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n385,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n690,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n122,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n40,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n565,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n964,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n714,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n921,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n622,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n118,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n612,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n439,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


