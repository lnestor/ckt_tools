// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_55 written by SynthGen on 2021/04/05 11:22:31
module Stat_100_55( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n98, n103, n107, n109, n104, n112, n131, n117,
 n113, n126, n116, n120, n114, n115, n132, n108,
 n127, n121, n122, n128, n111, n106, n125, n123,
 n102, n118, n105, n129, n110, n119, n130, n124);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n98, n103, n107, n109, n104, n112, n131, n117,
 n113, n126, n116, n120, n114, n115, n132, n108,
 n127, n121, n122, n128, n111, n106, n125, n123,
 n102, n118, n105, n129, n110, n119, n130, n124;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n99, n100, n101;

not  g0 (n33, n9);
buf  g1 (n37, n4);
buf  g2 (n42, n6);
buf  g3 (n41, n10);
buf  g4 (n38, n3);
buf  g5 (n36, n2);
buf  g6 (n34, n5);
buf  g7 (n39, n1);
buf  g8 (n40, n8);
not  g9 (n35, n7);
buf  g10 (n74, n36);
not  g11 (n46, n35);
not  g12 (n59, n36);
not  g13 (n61, n34);
buf  g14 (n44, n38);
buf  g15 (n57, n12);
not  g16 (n62, n37);
buf  g17 (n52, n38);
buf  g18 (n67, n37);
not  g19 (n49, n40);
not  g20 (n69, n35);
not  g21 (n77, n38);
buf  g22 (n60, n11);
buf  g23 (n50, n38);
buf  g24 (n63, n34);
buf  g25 (n70, n37);
buf  g26 (n47, n39);
not  g27 (n65, n40);
not  g28 (n76, n13);
not  g29 (n68, n39);
buf  g30 (n56, n33);
not  g31 (n64, n36);
not  g32 (n58, n33);
buf  g33 (n53, n41);
not  g34 (n54, n35);
not  g35 (n43, n33);
buf  g36 (n71, n34);
not  g37 (n66, n35);
buf  g38 (n45, n33);
not  g39 (n55, n37);
buf  g40 (n75, n39);
not  g41 (n73, n40);
buf  g42 (n72, n39);
buf  g43 (n51, n36);
or   g44 (n48, n40, n34, n41);
nor  g45 (n78, n22, n46, n24, n32);
nor  g46 (n80, n32, n32, n16, n31);
nand g47 (n81, n43, n29, n47, n23);
and  g48 (n79, n18, n45, n20, n21);
nand g49 (n82, n30, n30, n44, n14);
or   g50 (n85, n28, n19, n25, n50);
or   g51 (n83, n51, n49, n17, n27);
nor  g52 (n84, n26, n31, n48, n15);
buf  g53 (n92, n80);
not  g54 (n97, n83);
not  g55 (n86, n53);
not  g56 (n100, n42);
not  g57 (n94, n42);
not  g58 (n91, n83);
buf  g59 (n88, n32);
buf  g60 (n87, n55);
buf  g61 (n99, n55);
buf  g62 (n101, n83);
xor  g63 (n89, n54, n82);
and  g64 (n96, n79, n85, n41, n84);
or   g65 (n90, n52, n84, n82);
and  g66 (n93, n82, n54, n42);
and  g67 (n95, n84, n53, n54, n83);
xor  g68 (n98, n84, n42, n81, n78);
and  g69 (n132, n58, n73, n65, n62);
or   g70 (n115, n68, n70, n61, n69);
nand g71 (n106, n59, n61, n56, n100);
or   g72 (n128, n74, n66, n72, n62);
xnor g73 (n108, n55, n70, n63, n92);
xnor g74 (n123, n87, n56, n64, n95);
nor  g75 (n104, n67, n88, n61, n60);
xor  g76 (n114, n68, n77, n74, n64);
nor  g77 (n110, n75, n101, n55, n67);
or   g78 (n125, n65, n97, n71, n60);
xor  g79 (n120, n56, n62, n99, n100);
xor  g80 (n111, n100, n62, n74, n91);
xnor g81 (n126, n96, n58, n67, n90);
nand g82 (n121, n57, n66, n99, n69);
nor  g83 (n116, n75, n69, n59, n94);
xnor g84 (n118, n72, n97, n61, n98);
nand g85 (n112, n75, n59, n57, n100);
and  g86 (n107, n64, n85, n58, n77);
and  g87 (n103, n69, n98, n65);
xnor g88 (n102, n56, n76, n73);
xnor g89 (n130, n89, n59, n97, n74);
nand g90 (n109, n101, n66, n71);
nor  g91 (n122, n76, n97, n71, n86);
xnor g92 (n124, n63, n63, n99, n75);
xnor g93 (n113, n60, n76, n85, n101);
and  g94 (n105, n77, n73, n72, n68);
and  g95 (n127, n57, n70, n66, n85);
xor  g96 (n117, n99, n68, n73, n58);
nand g97 (n119, n64, n98, n101, n70);
nand g98 (n129, n93, n63, n65, n67);
and  g99 (n131, n72, n57, n60, n77);
endmodule
