

module Stat_3000_307
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1840,
  n1835,
  n1829,
  n1833,
  n1843,
  n1841,
  n1837,
  n1834,
  n1839,
  n1831,
  n1832,
  n1846,
  n1836,
  n1842,
  n1867,
  n1866,
  n3024,
  n3020,
  n3029,
  n3023,
  n3019,
  n3017,
  n3032,
  n3030,
  n3025,
  n3022,
  n3028,
  n3021,
  n3031,
  n3027,
  n3026,
  n3018,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1840;
  output n1835;
  output n1829;
  output n1833;
  output n1843;
  output n1841;
  output n1837;
  output n1834;
  output n1839;
  output n1831;
  output n1832;
  output n1846;
  output n1836;
  output n1842;
  output n1867;
  output n1866;
  output n3024;
  output n3020;
  output n3029;
  output n3023;
  output n3019;
  output n3017;
  output n3032;
  output n3030;
  output n3025;
  output n3022;
  output n3028;
  output n3021;
  output n3031;
  output n3027;
  output n3026;
  output n3018;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1830;
  wire n1838;
  wire n1844;
  wire n1845;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n113,
    n31
  );


  buf
  g1
  (
    n86,
    n25
  );


  buf
  g2
  (
    n126,
    n8
  );


  not
  g3
  (
    n69,
    n32
  );


  buf
  g4
  (
    n49,
    n30
  );


  not
  g5
  (
    n150,
    n23
  );


  buf
  g6
  (
    n71,
    n25
  );


  not
  g7
  (
    n144,
    n19
  );


  not
  g8
  (
    n134,
    n28
  );


  not
  g9
  (
    n37,
    n26
  );


  not
  g10
  (
    n55,
    n9
  );


  buf
  g11
  (
    n63,
    n32
  );


  not
  g12
  (
    n114,
    n4
  );


  not
  g13
  (
    n156,
    n6
  );


  buf
  g14
  (
    n56,
    n11
  );


  buf
  g15
  (
    n92,
    n16
  );


  buf
  g16
  (
    n98,
    n4
  );


  buf
  g17
  (
    n72,
    n31
  );


  not
  g18
  (
    n50,
    n29
  );


  not
  g19
  (
    n103,
    n14
  );


  not
  g20
  (
    n66,
    n2
  );


  buf
  g21
  (
    n127,
    n9
  );


  buf
  g22
  (
    n73,
    n29
  );


  not
  g23
  (
    n94,
    n17
  );


  buf
  g24
  (
    n80,
    n11
  );


  buf
  g25
  (
    n135,
    n31
  );


  not
  g26
  (
    n88,
    n6
  );


  buf
  g27
  (
    n87,
    n16
  );


  not
  g28
  (
    n99,
    n3
  );


  buf
  g29
  (
    n35,
    n27
  );


  buf
  g30
  (
    n138,
    n24
  );


  not
  g31
  (
    n136,
    n14
  );


  buf
  g32
  (
    n137,
    n21
  );


  buf
  g33
  (
    n102,
    n18
  );


  not
  g34
  (
    n128,
    n20
  );


  buf
  g35
  (
    n154,
    n5
  );


  not
  g36
  (
    n120,
    n7
  );


  buf
  g37
  (
    n81,
    n25
  );


  buf
  g38
  (
    n96,
    n22
  );


  not
  g39
  (
    n97,
    n5
  );


  not
  g40
  (
    n34,
    n15
  );


  buf
  g41
  (
    n83,
    n32
  );


  buf
  g42
  (
    n57,
    n2
  );


  not
  g43
  (
    n116,
    n11
  );


  not
  g44
  (
    n39,
    n1
  );


  buf
  g45
  (
    n54,
    n17
  );


  buf
  g46
  (
    n90,
    n12
  );


  not
  g47
  (
    n142,
    n31
  );


  not
  g48
  (
    n115,
    n13
  );


  buf
  g49
  (
    n124,
    n16
  );


  not
  g50
  (
    n132,
    n32
  );


  not
  g51
  (
    n157,
    n10
  );


  buf
  g52
  (
    n67,
    n2
  );


  not
  g53
  (
    n59,
    n26
  );


  not
  g54
  (
    n61,
    n23
  );


  not
  g55
  (
    n111,
    n4
  );


  not
  g56
  (
    n38,
    n3
  );


  not
  g57
  (
    n82,
    n13
  );


  not
  g58
  (
    n143,
    n27
  );


  buf
  g59
  (
    n147,
    n5
  );


  buf
  g60
  (
    n101,
    n14
  );


  not
  g61
  (
    n42,
    n19
  );


  buf
  g62
  (
    n40,
    n15
  );


  not
  g63
  (
    n130,
    n6
  );


  buf
  g64
  (
    n107,
    n7
  );


  not
  g65
  (
    n43,
    n20
  );


  buf
  g66
  (
    n74,
    n22
  );


  not
  g67
  (
    n119,
    n28
  );


  buf
  g68
  (
    n75,
    n24
  );


  buf
  g69
  (
    n117,
    n9
  );


  buf
  g70
  (
    n79,
    n29
  );


  buf
  g71
  (
    n46,
    n28
  );


  not
  g72
  (
    n100,
    n22
  );


  buf
  g73
  (
    n151,
    n12
  );


  not
  g74
  (
    n145,
    n12
  );


  buf
  g75
  (
    n158,
    n23
  );


  not
  g76
  (
    n62,
    n19
  );


  buf
  g77
  (
    n121,
    n19
  );


  buf
  g78
  (
    n122,
    n24
  );


  not
  g79
  (
    n95,
    n28
  );


  buf
  g80
  (
    n33,
    n9
  );


  buf
  g81
  (
    n110,
    n8
  );


  not
  g82
  (
    n84,
    n1
  );


  buf
  g83
  (
    n108,
    n10
  );


  buf
  g84
  (
    n104,
    n18
  );


  buf
  g85
  (
    n139,
    n8
  );


  buf
  g86
  (
    n125,
    n4
  );


  not
  g87
  (
    n133,
    n10
  );


  buf
  g88
  (
    n91,
    n2
  );


  buf
  g89
  (
    n45,
    n29
  );


  buf
  g90
  (
    n155,
    n23
  );


  buf
  g91
  (
    n36,
    n15
  );


  buf
  g92
  (
    n70,
    n7
  );


  not
  g93
  (
    n78,
    n14
  );


  not
  g94
  (
    n106,
    n30
  );


  buf
  g95
  (
    n148,
    n26
  );


  buf
  g96
  (
    n109,
    n13
  );


  buf
  g97
  (
    n123,
    n30
  );


  buf
  g98
  (
    n160,
    n18
  );


  not
  g99
  (
    n141,
    n13
  );


  not
  g100
  (
    n89,
    n27
  );


  not
  g101
  (
    n68,
    n21
  );


  buf
  g102
  (
    n77,
    n5
  );


  buf
  g103
  (
    n129,
    n20
  );


  not
  g104
  (
    n52,
    n11
  );


  buf
  g105
  (
    n93,
    n20
  );


  buf
  g106
  (
    n58,
    n30
  );


  not
  g107
  (
    n76,
    n25
  );


  buf
  g108
  (
    n153,
    n1
  );


  buf
  g109
  (
    n149,
    n7
  );


  not
  g110
  (
    n65,
    n22
  );


  buf
  g111
  (
    n47,
    n8
  );


  not
  g112
  (
    n146,
    n21
  );


  not
  g113
  (
    n140,
    n17
  );


  buf
  g114
  (
    n41,
    n16
  );


  buf
  g115
  (
    n48,
    n10
  );


  buf
  g116
  (
    n118,
    n12
  );


  buf
  g117
  (
    n131,
    n6
  );


  buf
  g118
  (
    n64,
    n1
  );


  not
  g119
  (
    n53,
    n17
  );


  not
  g120
  (
    n159,
    n3
  );


  not
  g121
  (
    n44,
    n21
  );


  buf
  g122
  (
    n85,
    n24
  );


  buf
  g123
  (
    n51,
    n26
  );


  buf
  g124
  (
    n112,
    n27
  );


  not
  g125
  (
    n105,
    n3
  );


  buf
  g126
  (
    n60,
    n18
  );


  not
  g127
  (
    n152,
    n15
  );


  buf
  g128
  (
    n654,
    n134
  );


  buf
  g129
  (
    n345,
    n43
  );


  not
  g130
  (
    n606,
    n130
  );


  buf
  g131
  (
    n635,
    n118
  );


  not
  g132
  (
    n233,
    n84
  );


  buf
  g133
  (
    n627,
    n140
  );


  not
  g134
  (
    n652,
    n152
  );


  buf
  g135
  (
    n413,
    n78
  );


  not
  g136
  (
    n380,
    n37
  );


  not
  g137
  (
    n261,
    n83
  );


  not
  g138
  (
    n375,
    n33
  );


  buf
  g139
  (
    n499,
    n133
  );


  not
  g140
  (
    n318,
    n86
  );


  not
  g141
  (
    n523,
    n82
  );


  buf
  g142
  (
    n300,
    n58
  );


  buf
  g143
  (
    n636,
    n133
  );


  buf
  g144
  (
    n554,
    n153
  );


  not
  g145
  (
    n368,
    n55
  );


  buf
  g146
  (
    n540,
    n158
  );


  buf
  g147
  (
    n632,
    n82
  );


  buf
  g148
  (
    n476,
    n132
  );


  not
  g149
  (
    n537,
    n103
  );


  not
  g150
  (
    n195,
    n140
  );


  not
  g151
  (
    n197,
    n138
  );


  buf
  g152
  (
    n250,
    n89
  );


  buf
  g153
  (
    n641,
    n126
  );


  buf
  g154
  (
    n623,
    n65
  );


  not
  g155
  (
    n462,
    n41
  );


  not
  g156
  (
    n452,
    n100
  );


  buf
  g157
  (
    n517,
    n67
  );


  buf
  g158
  (
    n604,
    n48
  );


  not
  g159
  (
    n385,
    n142
  );


  buf
  g160
  (
    n486,
    n135
  );


  not
  g161
  (
    n474,
    n102
  );


  not
  g162
  (
    n498,
    n136
  );


  not
  g163
  (
    n613,
    n59
  );


  buf
  g164
  (
    n576,
    n74
  );


  buf
  g165
  (
    n320,
    n123
  );


  not
  g166
  (
    n362,
    n125
  );


  buf
  g167
  (
    n524,
    n93
  );


  buf
  g168
  (
    n629,
    n52
  );


  buf
  g169
  (
    n198,
    n84
  );


  not
  g170
  (
    n400,
    n110
  );


  buf
  g171
  (
    n553,
    n152
  );


  buf
  g172
  (
    n428,
    n46
  );


  buf
  g173
  (
    n242,
    n122
  );


  not
  g174
  (
    n188,
    n57
  );


  not
  g175
  (
    n263,
    n85
  );


  not
  g176
  (
    n401,
    n109
  );


  buf
  g177
  (
    n256,
    n108
  );


  buf
  g178
  (
    n522,
    n122
  );


  buf
  g179
  (
    n642,
    n98
  );


  not
  g180
  (
    n186,
    n38
  );


  not
  g181
  (
    n218,
    n41
  );


  buf
  g182
  (
    n502,
    n93
  );


  buf
  g183
  (
    n459,
    n156
  );


  not
  g184
  (
    n232,
    n127
  );


  buf
  g185
  (
    n526,
    n158
  );


  buf
  g186
  (
    n311,
    n85
  );


  buf
  g187
  (
    n442,
    n124
  );


  buf
  g188
  (
    n396,
    n60
  );


  buf
  g189
  (
    n237,
    n103
  );


  buf
  g190
  (
    n620,
    n40
  );


  not
  g191
  (
    n663,
    n131
  );


  buf
  g192
  (
    n568,
    n60
  );


  not
  g193
  (
    n253,
    n118
  );


  buf
  g194
  (
    n203,
    n61
  );


  not
  g195
  (
    n411,
    n108
  );


  not
  g196
  (
    n225,
    n135
  );


  buf
  g197
  (
    n190,
    n92
  );


  buf
  g198
  (
    n588,
    n145
  );


  not
  g199
  (
    n319,
    n64
  );


  not
  g200
  (
    n231,
    n117
  );


  not
  g201
  (
    n162,
    n109
  );


  not
  g202
  (
    n390,
    n39
  );


  not
  g203
  (
    n166,
    n47
  );


  buf
  g204
  (
    n520,
    n130
  );


  buf
  g205
  (
    n355,
    n119
  );


  buf
  g206
  (
    n182,
    n58
  );


  buf
  g207
  (
    n591,
    n35
  );


  buf
  g208
  (
    n359,
    n76
  );


  not
  g209
  (
    n449,
    n106
  );


  buf
  g210
  (
    n445,
    n68
  );


  buf
  g211
  (
    n471,
    n114
  );


  not
  g212
  (
    n614,
    n150
  );


  not
  g213
  (
    n421,
    n51
  );


  not
  g214
  (
    n434,
    n143
  );


  buf
  g215
  (
    n496,
    n64
  );


  buf
  g216
  (
    n647,
    n39
  );


  not
  g217
  (
    n608,
    n146
  );


  not
  g218
  (
    n532,
    n57
  );


  not
  g219
  (
    n451,
    n144
  );


  buf
  g220
  (
    n293,
    n56
  );


  not
  g221
  (
    n335,
    n135
  );


  buf
  g222
  (
    n597,
    n116
  );


  not
  g223
  (
    n333,
    n47
  );


  not
  g224
  (
    n201,
    n92
  );


  buf
  g225
  (
    n603,
    n96
  );


  not
  g226
  (
    n339,
    n153
  );


  buf
  g227
  (
    n668,
    n79
  );


  not
  g228
  (
    n251,
    n87
  );


  not
  g229
  (
    n189,
    n100
  );


  not
  g230
  (
    n356,
    n60
  );


  buf
  g231
  (
    n179,
    n157
  );


  not
  g232
  (
    n582,
    n42
  );


  buf
  g233
  (
    n220,
    n154
  );


  buf
  g234
  (
    n301,
    n106
  );


  not
  g235
  (
    n316,
    n36
  );


  not
  g236
  (
    n450,
    n139
  );


  not
  g237
  (
    n408,
    n95
  );


  not
  g238
  (
    n351,
    n107
  );


  not
  g239
  (
    n460,
    n70
  );


  buf
  g240
  (
    n264,
    n55
  );


  not
  g241
  (
    n625,
    n150
  );


  not
  g242
  (
    n489,
    n97
  );


  not
  g243
  (
    n260,
    n141
  );


  not
  g244
  (
    n639,
    n73
  );


  buf
  g245
  (
    n247,
    n99
  );


  not
  g246
  (
    n653,
    n69
  );


  not
  g247
  (
    n399,
    n120
  );


  buf
  g248
  (
    n270,
    n59
  );


  not
  g249
  (
    n432,
    n46
  );


  not
  g250
  (
    n555,
    n129
  );


  buf
  g251
  (
    n516,
    n39
  );


  not
  g252
  (
    n172,
    n142
  );


  not
  g253
  (
    n202,
    n138
  );


  buf
  g254
  (
    n626,
    n105
  );


  not
  g255
  (
    n384,
    n38
  );


  buf
  g256
  (
    n191,
    n50
  );


  not
  g257
  (
    n545,
    n38
  );


  not
  g258
  (
    n181,
    n76
  );


  not
  g259
  (
    n170,
    n67
  );


  buf
  g260
  (
    n376,
    n114
  );


  not
  g261
  (
    n306,
    n97
  );


  buf
  g262
  (
    n477,
    n128
  );


  buf
  g263
  (
    n238,
    n125
  );


  buf
  g264
  (
    n531,
    n98
  );


  buf
  g265
  (
    n328,
    n145
  );


  buf
  g266
  (
    n577,
    n82
  );


  not
  g267
  (
    n248,
    n105
  );


  not
  g268
  (
    n276,
    n87
  );


  not
  g269
  (
    n495,
    n86
  );


  buf
  g270
  (
    n561,
    n54
  );


  buf
  g271
  (
    n404,
    n102
  );


  buf
  g272
  (
    n364,
    n61
  );


  buf
  g273
  (
    n363,
    n137
  );


  buf
  g274
  (
    n464,
    n68
  );


  buf
  g275
  (
    n317,
    n91
  );


  not
  g276
  (
    n277,
    n160
  );


  not
  g277
  (
    n571,
    n94
  );


  not
  g278
  (
    n479,
    n136
  );


  buf
  g279
  (
    n552,
    n130
  );


  not
  g280
  (
    n574,
    n56
  );


  not
  g281
  (
    n533,
    n121
  );


  not
  g282
  (
    n650,
    n112
  );


  not
  g283
  (
    n511,
    n94
  );


  buf
  g284
  (
    n426,
    n68
  );


  not
  g285
  (
    n525,
    n114
  );


  buf
  g286
  (
    n584,
    n74
  );


  buf
  g287
  (
    n192,
    n43
  );


  buf
  g288
  (
    n558,
    n37
  );


  buf
  g289
  (
    n267,
    n141
  );


  buf
  g290
  (
    n453,
    n125
  );


  buf
  g291
  (
    n633,
    n51
  );


  not
  g292
  (
    n587,
    n93
  );


  not
  g293
  (
    n176,
    n127
  );


  not
  g294
  (
    n435,
    n148
  );


  not
  g295
  (
    n550,
    n140
  );


  not
  g296
  (
    n329,
    n147
  );


  not
  g297
  (
    n235,
    n128
  );


  buf
  g298
  (
    n560,
    n41
  );


  buf
  g299
  (
    n485,
    n89
  );


  buf
  g300
  (
    n472,
    n160
  );


  buf
  g301
  (
    n337,
    n49
  );


  not
  g302
  (
    n322,
    n52
  );


  not
  g303
  (
    n430,
    n132
  );


  not
  g304
  (
    n619,
    n115
  );


  not
  g305
  (
    n341,
    n88
  );


  buf
  g306
  (
    n559,
    n79
  );


  not
  g307
  (
    n634,
    n103
  );


  buf
  g308
  (
    n374,
    n107
  );


  buf
  g309
  (
    n425,
    n95
  );


  not
  g310
  (
    n163,
    n116
  );


  not
  g311
  (
    n503,
    n46
  );


  not
  g312
  (
    n478,
    n72
  );


  buf
  g313
  (
    n269,
    n58
  );


  not
  g314
  (
    n278,
    n85
  );


  buf
  g315
  (
    n416,
    n61
  );


  buf
  g316
  (
    n482,
    n96
  );


  buf
  g317
  (
    n229,
    n143
  );


  buf
  g318
  (
    n284,
    n44
  );


  buf
  g319
  (
    n296,
    n75
  );


  buf
  g320
  (
    n648,
    n149
  );


  not
  g321
  (
    n392,
    n87
  );


  buf
  g322
  (
    n444,
    n154
  );


  not
  g323
  (
    n466,
    n101
  );


  buf
  g324
  (
    n423,
    n76
  );


  not
  g325
  (
    n395,
    n63
  );


  not
  g326
  (
    n222,
    n159
  );


  not
  g327
  (
    n369,
    n54
  );


  not
  g328
  (
    n657,
    n65
  );


  not
  g329
  (
    n378,
    n157
  );


  buf
  g330
  (
    n564,
    n132
  );


  not
  g331
  (
    n327,
    n40
  );


  not
  g332
  (
    n325,
    n150
  );


  buf
  g333
  (
    n655,
    n111
  );


  buf
  g334
  (
    n212,
    n51
  );


  not
  g335
  (
    n507,
    n42
  );


  not
  g336
  (
    n406,
    n45
  );


  not
  g337
  (
    n309,
    n73
  );


  not
  g338
  (
    n565,
    n97
  );


  buf
  g339
  (
    n349,
    n128
  );


  not
  g340
  (
    n615,
    n75
  );


  not
  g341
  (
    n468,
    n78
  );


  buf
  g342
  (
    n446,
    n123
  );


  buf
  g343
  (
    n539,
    n117
  );


  buf
  g344
  (
    n630,
    n121
  );


  not
  g345
  (
    n656,
    n43
  );


  not
  g346
  (
    n410,
    n35
  );


  not
  g347
  (
    n458,
    n67
  );


  not
  g348
  (
    n649,
    n119
  );


  buf
  g349
  (
    n169,
    n77
  );


  buf
  g350
  (
    n204,
    n76
  );


  not
  g351
  (
    n433,
    n131
  );


  buf
  g352
  (
    n470,
    n127
  );


  not
  g353
  (
    n262,
    n44
  );


  not
  g354
  (
    n481,
    n62
  );


  not
  g355
  (
    n310,
    n40
  );


  buf
  g356
  (
    n493,
    n149
  );


  not
  g357
  (
    n455,
    n42
  );


  buf
  g358
  (
    n535,
    n63
  );


  not
  g359
  (
    n377,
    n83
  );


  not
  g360
  (
    n226,
    n144
  );


  not
  g361
  (
    n196,
    n104
  );


  buf
  g362
  (
    n213,
    n109
  );


  buf
  g363
  (
    n618,
    n62
  );


  buf
  g364
  (
    n346,
    n49
  );


  buf
  g365
  (
    n504,
    n154
  );


  not
  g366
  (
    n415,
    n43
  );


  not
  g367
  (
    n424,
    n69
  );


  buf
  g368
  (
    n440,
    n91
  );


  buf
  g369
  (
    n272,
    n80
  );


  not
  g370
  (
    n330,
    n91
  );


  not
  g371
  (
    n326,
    n146
  );


  buf
  g372
  (
    n287,
    n149
  );


  not
  g373
  (
    n572,
    n66
  );


  buf
  g374
  (
    n372,
    n53
  );


  buf
  g375
  (
    n397,
    n148
  );


  not
  g376
  (
    n500,
    n39
  );


  buf
  g377
  (
    n549,
    n141
  );


  not
  g378
  (
    n244,
    n133
  );


  not
  g379
  (
    n383,
    n156
  );


  buf
  g380
  (
    n230,
    n152
  );


  buf
  g381
  (
    n427,
    n95
  );


  buf
  g382
  (
    n417,
    n95
  );


  not
  g383
  (
    n402,
    n116
  );


  buf
  g384
  (
    n193,
    n36
  );


  not
  g385
  (
    n484,
    n101
  );


  buf
  g386
  (
    n366,
    n49
  );


  not
  g387
  (
    n598,
    n104
  );


  buf
  g388
  (
    n360,
    n157
  );


  buf
  g389
  (
    n586,
    n81
  );


  buf
  g390
  (
    n601,
    n65
  );


  not
  g391
  (
    n557,
    n120
  );


  not
  g392
  (
    n505,
    n47
  );


  not
  g393
  (
    n469,
    n137
  );


  not
  g394
  (
    n543,
    n118
  );


  not
  g395
  (
    n611,
    n148
  );


  buf
  g396
  (
    n671,
    n104
  );


  not
  g397
  (
    n542,
    n72
  );


  not
  g398
  (
    n285,
    n158
  );


  not
  g399
  (
    n570,
    n136
  );


  buf
  g400
  (
    n596,
    n160
  );


  not
  g401
  (
    n666,
    n123
  );


  not
  g402
  (
    n518,
    n45
  );


  buf
  g403
  (
    n297,
    n52
  );


  not
  g404
  (
    n334,
    n138
  );


  not
  g405
  (
    n578,
    n54
  );


  not
  g406
  (
    n536,
    n131
  );


  not
  g407
  (
    n185,
    n136
  );


  buf
  g408
  (
    n646,
    n151
  );


  buf
  g409
  (
    n447,
    n53
  );


  buf
  g410
  (
    n438,
    n96
  );


  not
  g411
  (
    n483,
    n105
  );


  not
  g412
  (
    n461,
    n93
  );


  buf
  g413
  (
    n254,
    n108
  );


  not
  g414
  (
    n344,
    n144
  );


  buf
  g415
  (
    n640,
    n98
  );


  buf
  g416
  (
    n294,
    n73
  );


  buf
  g417
  (
    n209,
    n59
  );


  buf
  g418
  (
    n579,
    n142
  );


  buf
  g419
  (
    n609,
    n156
  );


  not
  g420
  (
    n658,
    n49
  );


  not
  g421
  (
    n631,
    n69
  );


  buf
  g422
  (
    n506,
    n53
  );


  not
  g423
  (
    n279,
    n72
  );


  buf
  g424
  (
    n224,
    n34
  );


  buf
  g425
  (
    n194,
    n52
  );


  not
  g426
  (
    n422,
    n149
  );


  not
  g427
  (
    n580,
    n44
  );


  not
  g428
  (
    n480,
    n102
  );


  buf
  g429
  (
    n645,
    n151
  );


  not
  g430
  (
    n307,
    n85
  );


  not
  g431
  (
    n295,
    n34
  );


  not
  g432
  (
    n281,
    n33
  );


  buf
  g433
  (
    n527,
    n57
  );


  buf
  g434
  (
    n575,
    n153
  );


  buf
  g435
  (
    n605,
    n143
  );


  not
  g436
  (
    n274,
    n104
  );


  not
  g437
  (
    n431,
    n150
  );


  buf
  g438
  (
    n407,
    n156
  );


  not
  g439
  (
    n405,
    n82
  );


  buf
  g440
  (
    n381,
    n115
  );


  buf
  g441
  (
    n566,
    n107
  );


  not
  g442
  (
    n239,
    n146
  );


  buf
  g443
  (
    n534,
    n112
  );


  buf
  g444
  (
    n429,
    n56
  );


  not
  g445
  (
    n314,
    n46
  );


  not
  g446
  (
    n454,
    n88
  );


  not
  g447
  (
    n547,
    n86
  );


  not
  g448
  (
    n236,
    n48
  );


  not
  g449
  (
    n210,
    n48
  );


  buf
  g450
  (
    n227,
    n159
  );


  not
  g451
  (
    n273,
    n90
  );


  not
  g452
  (
    n621,
    n37
  );


  buf
  g453
  (
    n252,
    n63
  );


  not
  g454
  (
    n669,
    n124
  );


  not
  g455
  (
    n388,
    n113
  );


  buf
  g456
  (
    n289,
    n50
  );


  buf
  g457
  (
    n266,
    n138
  );


  buf
  g458
  (
    n573,
    n51
  );


  not
  g459
  (
    n513,
    n119
  );


  buf
  g460
  (
    n569,
    n74
  );


  not
  g461
  (
    n662,
    n74
  );


  not
  g462
  (
    n528,
    n78
  );


  buf
  g463
  (
    n398,
    n101
  );


  buf
  g464
  (
    n286,
    n86
  );


  buf
  g465
  (
    n304,
    n134
  );


  buf
  g466
  (
    n412,
    n58
  );


  buf
  g467
  (
    n643,
    n34
  );


  not
  g468
  (
    n556,
    n45
  );


  buf
  g469
  (
    n409,
    n122
  );


  not
  g470
  (
    n177,
    n71
  );


  not
  g471
  (
    n443,
    n90
  );


  buf
  g472
  (
    n538,
    n100
  );


  not
  g473
  (
    n245,
    n102
  );


  buf
  g474
  (
    n303,
    n145
  );


  not
  g475
  (
    n206,
    n115
  );


  buf
  g476
  (
    n241,
    n77
  );


  not
  g477
  (
    n665,
    n80
  );


  buf
  g478
  (
    n208,
    n110
  );


  buf
  g479
  (
    n187,
    n62
  );


  not
  g480
  (
    n246,
    n99
  );


  not
  g481
  (
    n288,
    n99
  );


  buf
  g482
  (
    n324,
    n50
  );


  not
  g483
  (
    n667,
    n112
  );


  buf
  g484
  (
    n389,
    n105
  );


  not
  g485
  (
    n200,
    n100
  );


  buf
  g486
  (
    n331,
    n126
  );


  not
  g487
  (
    n420,
    n84
  );


  buf
  g488
  (
    n265,
    n63
  );


  buf
  g489
  (
    n298,
    n37
  );


  not
  g490
  (
    n161,
    n120
  );


  not
  g491
  (
    n371,
    n81
  );


  not
  g492
  (
    n216,
    n137
  );


  not
  g493
  (
    n271,
    n88
  );


  not
  g494
  (
    n219,
    n142
  );


  buf
  g495
  (
    n541,
    n147
  );


  not
  g496
  (
    n299,
    n155
  );


  not
  g497
  (
    n592,
    n70
  );


  buf
  g498
  (
    n521,
    n65
  );


  buf
  g499
  (
    n174,
    n115
  );


  buf
  g500
  (
    n168,
    n107
  );


  not
  g501
  (
    n211,
    n123
  );


  buf
  g502
  (
    n215,
    n126
  );


  not
  g503
  (
    n628,
    n68
  );


  buf
  g504
  (
    n361,
    n114
  );


  buf
  g505
  (
    n180,
    n47
  );


  buf
  g506
  (
    n512,
    n124
  );


  not
  g507
  (
    n456,
    n112
  );


  buf
  g508
  (
    n487,
    n144
  );


  not
  g509
  (
    n544,
    n117
  );


  buf
  g510
  (
    n457,
    n154
  );


  not
  g511
  (
    n313,
    n134
  );


  not
  g512
  (
    n228,
    n134
  );


  buf
  g513
  (
    n332,
    n98
  );


  buf
  g514
  (
    n370,
    n80
  );


  buf
  g515
  (
    n367,
    n159
  );


  buf
  g516
  (
    n217,
    n137
  );


  not
  g517
  (
    n546,
    n34
  );


  buf
  g518
  (
    n515,
    n111
  );


  not
  g519
  (
    n638,
    n35
  );


  not
  g520
  (
    n593,
    n81
  );


  buf
  g521
  (
    n491,
    n64
  );


  not
  g522
  (
    n467,
    n126
  );


  not
  g523
  (
    n519,
    n66
  );


  not
  g524
  (
    n350,
    n79
  );


  buf
  g525
  (
    n321,
    n129
  );


  buf
  g526
  (
    n386,
    n54
  );


  not
  g527
  (
    n514,
    n59
  );


  not
  g528
  (
    n664,
    n69
  );


  not
  g529
  (
    n165,
    n67
  );


  buf
  g530
  (
    n353,
    n35
  );


  buf
  g531
  (
    n599,
    n83
  );


  buf
  g532
  (
    n488,
    n55
  );


  buf
  g533
  (
    KeyWire_0_6,
    n91
  );


  not
  g534
  (
    n268,
    n75
  );


  not
  g535
  (
    n205,
    n128
  );


  not
  g536
  (
    n583,
    n89
  );


  buf
  g537
  (
    n403,
    n90
  );


  buf
  g538
  (
    n548,
    n73
  );


  not
  g539
  (
    n336,
    n72
  );


  not
  g540
  (
    n617,
    n147
  );


  not
  g541
  (
    n373,
    n155
  );


  buf
  g542
  (
    n275,
    n152
  );


  not
  g543
  (
    n595,
    n118
  );


  buf
  g544
  (
    n465,
    n94
  );


  buf
  g545
  (
    n234,
    n124
  );


  not
  g546
  (
    n610,
    n117
  );


  buf
  g547
  (
    n624,
    n80
  );


  buf
  g548
  (
    n567,
    n33
  );


  buf
  g549
  (
    n291,
    n77
  );


  not
  g550
  (
    n183,
    n110
  );


  buf
  g551
  (
    n441,
    n64
  );


  not
  g552
  (
    n473,
    n33
  );


  not
  g553
  (
    n660,
    n88
  );


  not
  g554
  (
    n240,
    n145
  );


  not
  g555
  (
    n382,
    n55
  );


  buf
  g556
  (
    n302,
    n146
  );


  buf
  g557
  (
    n659,
    n89
  );


  not
  g558
  (
    n616,
    n120
  );


  not
  g559
  (
    n207,
    n56
  );


  not
  g560
  (
    n651,
    n135
  );


  not
  g561
  (
    n342,
    n121
  );


  not
  g562
  (
    n199,
    n97
  );


  not
  g563
  (
    n258,
    n141
  );


  buf
  g564
  (
    n221,
    n77
  );


  not
  g565
  (
    n637,
    n40
  );


  buf
  g566
  (
    n347,
    n62
  );


  buf
  g567
  (
    n255,
    n157
  );


  buf
  g568
  (
    n510,
    n53
  );


  buf
  g569
  (
    n292,
    n101
  );


  buf
  g570
  (
    n340,
    n158
  );


  buf
  g571
  (
    n352,
    n94
  );


  buf
  g572
  (
    n354,
    n147
  );


  buf
  g573
  (
    n600,
    n139
  );


  buf
  g574
  (
    n670,
    n84
  );


  not
  g575
  (
    n393,
    n71
  );


  not
  g576
  (
    n508,
    n127
  );


  buf
  g577
  (
    n563,
    n125
  );


  buf
  g578
  (
    n607,
    n111
  );


  not
  g579
  (
    n358,
    n109
  );


  buf
  g580
  (
    n494,
    n103
  );


  buf
  g581
  (
    n497,
    n45
  );


  not
  g582
  (
    n391,
    n42
  );


  buf
  g583
  (
    n283,
    n48
  );


  buf
  g584
  (
    n581,
    n70
  );


  not
  g585
  (
    n280,
    n130
  );


  not
  g586
  (
    n529,
    n83
  );


  buf
  g587
  (
    n164,
    n44
  );


  not
  g588
  (
    n439,
    n79
  );


  buf
  g589
  (
    n348,
    n70
  );


  not
  g590
  (
    n562,
    n132
  );


  not
  g591
  (
    n463,
    n108
  );


  not
  g592
  (
    n448,
    n116
  );


  buf
  g593
  (
    n612,
    n151
  );


  buf
  g594
  (
    n644,
    n110
  );


  not
  g595
  (
    n418,
    n50
  );


  buf
  g596
  (
    n585,
    n38
  );


  not
  g597
  (
    n622,
    n113
  );


  buf
  g598
  (
    n323,
    n155
  );


  not
  g599
  (
    n509,
    n36
  );


  not
  g600
  (
    n437,
    n155
  );


  not
  g601
  (
    n305,
    n41
  );


  buf
  g602
  (
    n387,
    n36
  );


  not
  g603
  (
    n184,
    n106
  );


  not
  g604
  (
    n315,
    n148
  );


  buf
  g605
  (
    n223,
    n131
  );


  not
  g606
  (
    n589,
    n129
  );


  buf
  g607
  (
    n290,
    n66
  );


  not
  g608
  (
    n343,
    n140
  );


  not
  g609
  (
    n243,
    n78
  );


  not
  g610
  (
    n175,
    n99
  );


  buf
  g611
  (
    n178,
    n113
  );


  not
  g612
  (
    n501,
    n133
  );


  buf
  g613
  (
    n173,
    n122
  );


  not
  g614
  (
    n492,
    n106
  );


  buf
  g615
  (
    n365,
    n90
  );


  buf
  g616
  (
    n214,
    n121
  );


  buf
  g617
  (
    n249,
    n66
  );


  not
  g618
  (
    n436,
    n87
  );


  not
  g619
  (
    n259,
    n60
  );


  not
  g620
  (
    n590,
    n71
  );


  buf
  g621
  (
    n282,
    n111
  );


  not
  g622
  (
    n312,
    n153
  );


  buf
  g623
  (
    n257,
    n139
  );


  not
  g624
  (
    n171,
    n119
  );


  buf
  g625
  (
    n419,
    n113
  );


  buf
  g626
  (
    n602,
    n139
  );


  buf
  g627
  (
    n551,
    n129
  );


  not
  g628
  (
    n379,
    n71
  );


  buf
  g629
  (
    n167,
    n159
  );


  buf
  g630
  (
    n357,
    n92
  );


  buf
  g631
  (
    n490,
    n92
  );


  buf
  g632
  (
    n338,
    n143
  );


  not
  g633
  (
    n530,
    n96
  );


  not
  g634
  (
    n594,
    n75
  );


  buf
  g635
  (
    n414,
    n61
  );


  not
  g636
  (
    n661,
    n57
  );


  not
  g637
  (
    n394,
    n81
  );


  buf
  g638
  (
    n308,
    n151
  );


  buf
  g639
  (
    n807,
    n526
  );


  buf
  g640
  (
    n938,
    n569
  );


  not
  g641
  (
    n1055,
    n431
  );


  not
  g642
  (
    n1100,
    n505
  );


  buf
  g643
  (
    n1197,
    n407
  );


  buf
  g644
  (
    n881,
    n323
  );


  not
  g645
  (
    n1126,
    n503
  );


  not
  g646
  (
    n745,
    n210
  );


  buf
  g647
  (
    n1178,
    n564
  );


  buf
  g648
  (
    n1158,
    n233
  );


  not
  g649
  (
    n997,
    n333
  );


  not
  g650
  (
    n1038,
    n365
  );


  not
  g651
  (
    n761,
    n430
  );


  buf
  g652
  (
    n974,
    n472
  );


  not
  g653
  (
    n1106,
    n221
  );


  not
  g654
  (
    n894,
    n557
  );


  buf
  g655
  (
    n1184,
    n301
  );


  not
  g656
  (
    n1410,
    n368
  );


  buf
  g657
  (
    n846,
    n484
  );


  buf
  g658
  (
    n792,
    n386
  );


  not
  g659
  (
    n944,
    n205
  );


  buf
  g660
  (
    n879,
    n461
  );


  not
  g661
  (
    n1185,
    n412
  );


  not
  g662
  (
    n1044,
    n465
  );


  buf
  g663
  (
    n1059,
    n224
  );


  buf
  g664
  (
    n697,
    n487
  );


  buf
  g665
  (
    n1395,
    n175
  );


  not
  g666
  (
    n1367,
    n559
  );


  not
  g667
  (
    n773,
    n294
  );


  not
  g668
  (
    n1135,
    n298
  );


  buf
  g669
  (
    n758,
    n560
  );


  buf
  g670
  (
    n805,
    n538
  );


  buf
  g671
  (
    n1161,
    n549
  );


  not
  g672
  (
    n1407,
    n395
  );


  buf
  g673
  (
    n836,
    n186
  );


  not
  g674
  (
    n977,
    n252
  );


  buf
  g675
  (
    n1130,
    n440
  );


  not
  g676
  (
    n853,
    n265
  );


  not
  g677
  (
    n714,
    n333
  );


  buf
  g678
  (
    n1193,
    n482
  );


  buf
  g679
  (
    n1369,
    n174
  );


  not
  g680
  (
    n987,
    n164
  );


  not
  g681
  (
    n771,
    n417
  );


  buf
  g682
  (
    n1203,
    n409
  );


  buf
  g683
  (
    n1334,
    n486
  );


  not
  g684
  (
    n871,
    n242
  );


  not
  g685
  (
    n1314,
    n465
  );


  not
  g686
  (
    n810,
    n334
  );


  not
  g687
  (
    n812,
    n199
  );


  buf
  g688
  (
    n1436,
    n514
  );


  not
  g689
  (
    n1311,
    n489
  );


  buf
  g690
  (
    n1413,
    n450
  );


  not
  g691
  (
    n1182,
    n555
  );


  not
  g692
  (
    n715,
    n421
  );


  not
  g693
  (
    n953,
    n334
  );


  buf
  g694
  (
    n728,
    n264
  );


  buf
  g695
  (
    n1264,
    n534
  );


  not
  g696
  (
    n1062,
    n249
  );


  buf
  g697
  (
    n1388,
    n407
  );


  buf
  g698
  (
    n719,
    n350
  );


  buf
  g699
  (
    KeyWire_0_4,
    n420
  );


  buf
  g700
  (
    n1363,
    n210
  );


  buf
  g701
  (
    n850,
    n549
  );


  not
  g702
  (
    n1120,
    n518
  );


  buf
  g703
  (
    n907,
    n231
  );


  buf
  g704
  (
    n1128,
    n413
  );


  buf
  g705
  (
    KeyWire_0_8,
    n262
  );


  buf
  g706
  (
    n884,
    n308
  );


  buf
  g707
  (
    n1332,
    n177
  );


  not
  g708
  (
    n718,
    n268
  );


  buf
  g709
  (
    n901,
    n561
  );


  not
  g710
  (
    n1076,
    n179
  );


  not
  g711
  (
    n1049,
    n298
  );


  not
  g712
  (
    n949,
    n195
  );


  buf
  g713
  (
    n683,
    n361
  );


  buf
  g714
  (
    n932,
    n428
  );


  not
  g715
  (
    n916,
    n203
  );


  buf
  g716
  (
    n1122,
    n486
  );


  not
  g717
  (
    n769,
    n552
  );


  not
  g718
  (
    n1352,
    n349
  );


  not
  g719
  (
    n1090,
    n527
  );


  buf
  g720
  (
    n1426,
    n389
  );


  not
  g721
  (
    n1226,
    n241
  );


  buf
  g722
  (
    n1181,
    n457
  );


  not
  g723
  (
    n694,
    n431
  );


  not
  g724
  (
    n1249,
    n562
  );


  buf
  g725
  (
    n1392,
    n437
  );


  not
  g726
  (
    n1280,
    n178
  );


  not
  g727
  (
    n724,
    n215
  );


  buf
  g728
  (
    n1269,
    n192
  );


  buf
  g729
  (
    n1299,
    n317
  );


  not
  g730
  (
    n896,
    n545
  );


  buf
  g731
  (
    n1419,
    n258
  );


  not
  g732
  (
    n1208,
    n462
  );


  buf
  g733
  (
    n1134,
    n235
  );


  not
  g734
  (
    n1321,
    n187
  );


  buf
  g735
  (
    n927,
    n472
  );


  not
  g736
  (
    n1375,
    n321
  );


  not
  g737
  (
    n1254,
    n432
  );


  not
  g738
  (
    n1276,
    n229
  );


  not
  g739
  (
    n1348,
    n179
  );


  not
  g740
  (
    n1333,
    n418
  );


  not
  g741
  (
    n795,
    n264
  );


  not
  g742
  (
    n1089,
    n368
  );


  not
  g743
  (
    n1032,
    n318
  );


  buf
  g744
  (
    n851,
    n428
  );


  buf
  g745
  (
    n1206,
    n361
  );


  not
  g746
  (
    n1060,
    n176
  );


  buf
  g747
  (
    n1157,
    n533
  );


  buf
  g748
  (
    n1180,
    n474
  );


  not
  g749
  (
    n804,
    n268
  );


  buf
  g750
  (
    n1317,
    n358
  );


  buf
  g751
  (
    n1361,
    n452
  );


  buf
  g752
  (
    n1042,
    n351
  );


  buf
  g753
  (
    n999,
    n226
  );


  not
  g754
  (
    n1217,
    n419
  );


  not
  g755
  (
    n972,
    n403
  );


  not
  g756
  (
    n931,
    n505
  );


  not
  g757
  (
    n736,
    n199
  );


  not
  g758
  (
    n1406,
    n391
  );


  not
  g759
  (
    n847,
    n348
  );


  buf
  g760
  (
    n917,
    n331
  );


  buf
  g761
  (
    n1286,
    n511
  );


  not
  g762
  (
    n754,
    n457
  );


  not
  g763
  (
    n891,
    n220
  );


  not
  g764
  (
    n906,
    n494
  );


  buf
  g765
  (
    n1414,
    n209
  );


  not
  g766
  (
    n1095,
    n423
  );


  not
  g767
  (
    n1043,
    n225
  );


  not
  g768
  (
    n994,
    n389
  );


  not
  g769
  (
    n698,
    n386
  );


  buf
  g770
  (
    n1313,
    n399
  );


  buf
  g771
  (
    n965,
    n347
  );


  buf
  g772
  (
    n760,
    n383
  );


  buf
  g773
  (
    n1343,
    n529
  );


  not
  g774
  (
    n1019,
    n233
  );


  buf
  g775
  (
    n834,
    n255
  );


  not
  g776
  (
    n1296,
    n543
  );


  buf
  g777
  (
    n845,
    n485
  );


  not
  g778
  (
    n740,
    n195
  );


  not
  g779
  (
    n1131,
    n434
  );


  not
  g780
  (
    n1405,
    n341
  );


  not
  g781
  (
    n722,
    n180
  );


  not
  g782
  (
    n682,
    n192
  );


  not
  g783
  (
    n1191,
    n462
  );


  buf
  g784
  (
    n969,
    n393
  );


  buf
  g785
  (
    n1210,
    n239
  );


  not
  g786
  (
    n674,
    n459
  );


  not
  g787
  (
    n854,
    n246
  );


  buf
  g788
  (
    n1243,
    n208
  );


  buf
  g789
  (
    n877,
    n330
  );


  not
  g790
  (
    n1379,
    n260
  );


  buf
  g791
  (
    n744,
    n449
  );


  buf
  g792
  (
    n756,
    n167
  );


  not
  g793
  (
    n898,
    n196
  );


  not
  g794
  (
    n1347,
    n252
  );


  buf
  g795
  (
    n1329,
    n464
  );


  buf
  g796
  (
    n1036,
    n550
  );


  not
  g797
  (
    n904,
    n249
  );


  buf
  g798
  (
    KeyWire_0_13,
    n180
  );


  buf
  g799
  (
    n1002,
    n520
  );


  not
  g800
  (
    n741,
    n457
  );


  buf
  g801
  (
    n1295,
    n174
  );


  not
  g802
  (
    n1279,
    n285
  );


  buf
  g803
  (
    n873,
    n258
  );


  buf
  g804
  (
    n1201,
    n548
  );


  buf
  g805
  (
    n1417,
    n253
  );


  buf
  g806
  (
    n1171,
    n427
  );


  not
  g807
  (
    n1058,
    n345
  );


  buf
  g808
  (
    n1163,
    n428
  );


  not
  g809
  (
    n779,
    n257
  );


  not
  g810
  (
    n940,
    n513
  );


  buf
  g811
  (
    n1451,
    n369
  );


  not
  g812
  (
    n1053,
    n231
  );


  buf
  g813
  (
    n1097,
    n383
  );


  not
  g814
  (
    n1111,
    n480
  );


  buf
  g815
  (
    n1415,
    n462
  );


  buf
  g816
  (
    n685,
    n272
  );


  not
  g817
  (
    n1235,
    n189
  );


  not
  g818
  (
    n919,
    n448
  );


  not
  g819
  (
    n1165,
    n247
  );


  buf
  g820
  (
    n1270,
    n476
  );


  not
  g821
  (
    n713,
    n352
  );


  not
  g822
  (
    n1285,
    n281
  );


  not
  g823
  (
    n785,
    n303
  );


  buf
  g824
  (
    n1207,
    n399
  );


  not
  g825
  (
    n1104,
    n198
  );


  not
  g826
  (
    n1001,
    n541
  );


  buf
  g827
  (
    n1113,
    n473
  );


  not
  g828
  (
    n1288,
    n515
  );


  buf
  g829
  (
    n1428,
    n320
  );


  not
  g830
  (
    n1302,
    n470
  );


  buf
  g831
  (
    n1213,
    n202
  );


  not
  g832
  (
    n833,
    n287
  );


  buf
  g833
  (
    n1219,
    n476
  );


  not
  g834
  (
    n1354,
    n481
  );


  buf
  g835
  (
    n895,
    n527
  );


  not
  g836
  (
    n1025,
    n191
  );


  buf
  g837
  (
    n1046,
    n331
  );


  buf
  g838
  (
    n1237,
    n343
  );


  buf
  g839
  (
    n930,
    n310
  );


  not
  g840
  (
    n702,
    n268
  );


  not
  g841
  (
    n1227,
    n333
  );


  not
  g842
  (
    n1422,
    n499
  );


  not
  g843
  (
    n1433,
    n288
  );


  not
  g844
  (
    n1374,
    n504
  );


  buf
  g845
  (
    n686,
    n429
  );


  not
  g846
  (
    n1127,
    n190
  );


  not
  g847
  (
    n1246,
    n379
  );


  buf
  g848
  (
    n1256,
    n562
  );


  buf
  g849
  (
    n692,
    n451
  );


  not
  g850
  (
    n787,
    n535
  );


  not
  g851
  (
    n687,
    n263
  );


  buf
  g852
  (
    n1423,
    n357
  );


  buf
  g853
  (
    n1024,
    n435
  );


  buf
  g854
  (
    n1438,
    n236
  );


  not
  g855
  (
    n1109,
    n224
  );


  buf
  g856
  (
    n1045,
    n437
  );


  not
  g857
  (
    n1010,
    n250
  );


  buf
  g858
  (
    n908,
    n220
  );


  buf
  g859
  (
    n1092,
    n432
  );


  buf
  g860
  (
    n748,
    n294
  );


  buf
  g861
  (
    n1322,
    n243
  );


  buf
  g862
  (
    n1306,
    n302
  );


  buf
  g863
  (
    n1020,
    n237
  );


  not
  g864
  (
    n1265,
    n410
  );


  buf
  g865
  (
    n1396,
    n300
  );


  not
  g866
  (
    n902,
    n313
  );


  buf
  g867
  (
    n1102,
    n282
  );


  not
  g868
  (
    n1132,
    n222
  );


  not
  g869
  (
    n1139,
    n221
  );


  not
  g870
  (
    n1238,
    n393
  );


  not
  g871
  (
    n937,
    n262
  );


  buf
  g872
  (
    n696,
    n262
  );


  not
  g873
  (
    n1366,
    n542
  );


  not
  g874
  (
    n936,
    n266
  );


  not
  g875
  (
    n1124,
    n234
  );


  buf
  g876
  (
    n874,
    n570
  );


  not
  g877
  (
    n1224,
    n390
  );


  buf
  g878
  (
    n1205,
    n209
  );


  not
  g879
  (
    n684,
    n454
  );


  not
  g880
  (
    n943,
    n269
  );


  not
  g881
  (
    n984,
    n518
  );


  buf
  g882
  (
    n1026,
    n494
  );


  buf
  g883
  (
    n726,
    n254
  );


  buf
  g884
  (
    n1412,
    n539
  );


  not
  g885
  (
    n1117,
    n479
  );


  buf
  g886
  (
    n889,
    n217
  );


  buf
  g887
  (
    n1156,
    n227
  );


  buf
  g888
  (
    n1067,
    n458
  );


  not
  g889
  (
    n1373,
    n163
  );


  buf
  g890
  (
    n840,
    n531
  );


  not
  g891
  (
    n1284,
    n360
  );


  buf
  g892
  (
    n1051,
    n496
  );


  buf
  g893
  (
    n897,
    n246
  );


  buf
  g894
  (
    n738,
    n411
  );


  not
  g895
  (
    n680,
    n235
  );


  buf
  g896
  (
    n825,
    n563
  );


  not
  g897
  (
    n958,
    n321
  );


  not
  g898
  (
    n951,
    n293
  );


  buf
  g899
  (
    n811,
    n229
  );


  not
  g900
  (
    n1258,
    n240
  );


  buf
  g901
  (
    n732,
    n329
  );


  buf
  g902
  (
    n1389,
    n513
  );


  buf
  g903
  (
    n746,
    n344
  );


  buf
  g904
  (
    n727,
    n515
  );


  not
  g905
  (
    n842,
    n491
  );


  buf
  g906
  (
    n1027,
    n301
  );


  not
  g907
  (
    n878,
    n207
  );


  buf
  g908
  (
    n992,
    n248
  );


  buf
  g909
  (
    n1303,
    n461
  );


  not
  g910
  (
    n695,
    n188
  );


  buf
  g911
  (
    n1261,
    n373
  );


  buf
  g912
  (
    KeyWire_0_14,
    n314
  );


  not
  g913
  (
    n747,
    n522
  );


  buf
  g914
  (
    n1223,
    n459
  );


  buf
  g915
  (
    n869,
    n245
  );


  buf
  g916
  (
    n915,
    n547
  );


  buf
  g917
  (
    n1137,
    n497
  );


  not
  g918
  (
    n1175,
    n442
  );


  not
  g919
  (
    n776,
    n502
  );


  not
  g920
  (
    n913,
    n433
  );


  not
  g921
  (
    n1229,
    n359
  );


  buf
  g922
  (
    n971,
    n370
  );


  buf
  g923
  (
    n1228,
    n328
  );


  buf
  g924
  (
    n1315,
    n498
  );


  buf
  g925
  (
    n993,
    n546
  );


  not
  g926
  (
    n1272,
    n387
  );


  not
  g927
  (
    n1318,
    n213
  );


  buf
  g928
  (
    n1421,
    n165
  );


  not
  g929
  (
    n799,
    n305
  );


  buf
  g930
  (
    n1071,
    n569
  );


  not
  g931
  (
    n1119,
    n363
  );


  buf
  g932
  (
    n1431,
    n404
  );


  buf
  g933
  (
    n725,
    n404
  );


  not
  g934
  (
    n1084,
    n418
  );


  buf
  g935
  (
    n967,
    n430
  );


  not
  g936
  (
    n942,
    n425
  );


  buf
  g937
  (
    n988,
    n365
  );


  buf
  g938
  (
    n1103,
    n336
  );


  not
  g939
  (
    n1174,
    n319
  );


  not
  g940
  (
    n1023,
    n480
  );


  buf
  g941
  (
    n1337,
    n492
  );


  buf
  g942
  (
    n1003,
    n507
  );


  buf
  g943
  (
    n1344,
    n263
  );


  not
  g944
  (
    n996,
    n547
  );


  buf
  g945
  (
    n848,
    n517
  );


  buf
  g946
  (
    n1188,
    n516
  );


  buf
  g947
  (
    n768,
    n211
  );


  not
  g948
  (
    n1293,
    n163
  );


  not
  g949
  (
    n1064,
    n453
  );


  not
  g950
  (
    n843,
    n425
  );


  not
  g951
  (
    n690,
    n482
  );


  not
  g952
  (
    n1098,
    n491
  );


  buf
  g953
  (
    n925,
    n502
  );


  not
  g954
  (
    n1196,
    n531
  );


  buf
  g955
  (
    n794,
    n411
  );


  not
  g956
  (
    n826,
    n235
  );


  buf
  g957
  (
    n1186,
    n304
  );


  buf
  g958
  (
    n1241,
    n215
  );


  buf
  g959
  (
    n839,
    n284
  );


  buf
  g960
  (
    n1271,
    n426
  );


  buf
  g961
  (
    n1034,
    n294
  );


  buf
  g962
  (
    n887,
    n170
  );


  not
  g963
  (
    n1377,
    n343
  );


  not
  g964
  (
    n1247,
    n467
  );


  not
  g965
  (
    n1448,
    n292
  );


  not
  g966
  (
    n1006,
    n208
  );


  not
  g967
  (
    n1039,
    n477
  );


  buf
  g968
  (
    n1439,
    n182
  );


  not
  g969
  (
    n829,
    n422
  );


  not
  g970
  (
    n815,
    n486
  );


  buf
  g971
  (
    n1022,
    n325
  );


  buf
  g972
  (
    n1007,
    n478
  );


  buf
  g973
  (
    n1194,
    n309
  );


  not
  g974
  (
    n1147,
    n556
  );


  not
  g975
  (
    n716,
    n238
  );


  buf
  g976
  (
    n905,
    n546
  );


  buf
  g977
  (
    n966,
    n184
  );


  buf
  g978
  (
    n723,
    n187
  );


  not
  g979
  (
    n1121,
    n247
  );


  not
  g980
  (
    n1239,
    n237
  );


  buf
  g981
  (
    n1298,
    n228
  );


  buf
  g982
  (
    n1079,
    n180
  );


  buf
  g983
  (
    n1397,
    n414
  );


  not
  g984
  (
    n976,
    n338
  );


  not
  g985
  (
    n1250,
    n500
  );


  not
  g986
  (
    n1072,
    n326
  );


  not
  g987
  (
    n1140,
    n216
  );


  not
  g988
  (
    n1052,
    n342
  );


  buf
  g989
  (
    n712,
    n521
  );


  not
  g990
  (
    n918,
    n433
  );


  not
  g991
  (
    n1112,
    n439
  );


  buf
  g992
  (
    n1234,
    n185
  );


  not
  g993
  (
    n1364,
    n239
  );


  buf
  g994
  (
    n1088,
    n423
  );


  buf
  g995
  (
    n817,
    n346
  );


  buf
  g996
  (
    n1115,
    n249
  );


  not
  g997
  (
    n1325,
    n501
  );


  buf
  g998
  (
    n1091,
    n361
  );


  buf
  g999
  (
    n1014,
    n180
  );


  not
  g1000
  (
    n809,
    n319
  );


  not
  g1001
  (
    n990,
    n330
  );


  buf
  g1002
  (
    n1068,
    n266
  );


  buf
  g1003
  (
    n995,
    n501
  );


  not
  g1004
  (
    n998,
    n359
  );


  not
  g1005
  (
    n720,
    n475
  );


  not
  g1006
  (
    n1399,
    n181
  );


  not
  g1007
  (
    n1173,
    n293
  );


  buf
  g1008
  (
    n1409,
    n318
  );


  buf
  g1009
  (
    n1324,
    n391
  );


  buf
  g1010
  (
    n956,
    n506
  );


  buf
  g1011
  (
    n742,
    n170
  );


  buf
  g1012
  (
    n858,
    n521
  );


  not
  g1013
  (
    n946,
    n218
  );


  buf
  g1014
  (
    n1323,
    n492
  );


  not
  g1015
  (
    n1168,
    n257
  );


  buf
  g1016
  (
    n1394,
    n206
  );


  not
  g1017
  (
    n1376,
    n410
  );


  buf
  g1018
  (
    n1297,
    n316
  );


  not
  g1019
  (
    n1190,
    n331
  );


  not
  g1020
  (
    n1031,
    n465
  );


  not
  g1021
  (
    n920,
    n406
  );


  not
  g1022
  (
    n1080,
    n433
  );


  buf
  g1023
  (
    n893,
    n446
  );


  buf
  g1024
  (
    n1105,
    n391
  );


  buf
  g1025
  (
    n1030,
    n232
  );


  not
  g1026
  (
    n1304,
    n302
  );


  buf
  g1027
  (
    n1078,
    n209
  );


  not
  g1028
  (
    n861,
    n412
  );


  not
  g1029
  (
    n1093,
    n287
  );


  not
  g1030
  (
    n1177,
    n269
  );


  not
  g1031
  (
    n806,
    n199
  );


  buf
  g1032
  (
    n1434,
    n335
  );


  not
  g1033
  (
    n1145,
    n495
  );


  buf
  g1034
  (
    n767,
    n554
  );


  not
  g1035
  (
    n1274,
    n336
  );


  not
  g1036
  (
    n1259,
    n538
  );


  buf
  g1037
  (
    n1085,
    n468
  );


  buf
  g1038
  (
    n798,
    n335
  );


  not
  g1039
  (
    n816,
    n479
  );


  buf
  g1040
  (
    n678,
    n545
  );


  not
  g1041
  (
    n859,
    n302
  );


  not
  g1042
  (
    n672,
    n495
  );


  not
  g1043
  (
    n1440,
    n163
  );


  buf
  g1044
  (
    n753,
    n176
  );


  not
  g1045
  (
    n870,
    n372
  );


  not
  g1046
  (
    n1222,
    n475
  );


  not
  g1047
  (
    n764,
    n403
  );


  buf
  g1048
  (
    n790,
    n242
  );


  buf
  g1049
  (
    n935,
    n535
  );


  not
  g1050
  (
    n819,
    n207
  );


  not
  g1051
  (
    n1041,
    n368
  );


  buf
  g1052
  (
    n982,
    n564
  );


  buf
  g1053
  (
    n757,
    n269
  );


  not
  g1054
  (
    n1357,
    n273
  );


  not
  g1055
  (
    n783,
    n357
  );


  not
  g1056
  (
    n1360,
    n388
  );


  buf
  g1057
  (
    n820,
    n164
  );


  not
  g1058
  (
    n890,
    n453
  );


  buf
  g1059
  (
    n784,
    n336
  );


  buf
  g1060
  (
    n1096,
    n405
  );


  buf
  g1061
  (
    KeyWire_0_11,
    n311
  );


  buf
  g1062
  (
    n1164,
    n193
  );


  not
  g1063
  (
    n964,
    n385
  );


  not
  g1064
  (
    n703,
    n484
  );


  not
  g1065
  (
    n1035,
    n405
  );


  buf
  g1066
  (
    n1004,
    n309
  );


  buf
  g1067
  (
    n1262,
    n517
  );


  buf
  g1068
  (
    n1424,
    n320
  );


  buf
  g1069
  (
    n1075,
    n440
  );


  buf
  g1070
  (
    n1142,
    n201
  );


  not
  g1071
  (
    n1435,
    n470
  );


  buf
  g1072
  (
    n1442,
    n171
  );


  not
  g1073
  (
    n1443,
    n487
  );


  buf
  g1074
  (
    n1013,
    n401
  );


  buf
  g1075
  (
    n1266,
    n282
  );


  buf
  g1076
  (
    n1152,
    n174
  );


  buf
  g1077
  (
    n1048,
    n349
  );


  not
  g1078
  (
    n823,
    n193
  );


  not
  g1079
  (
    n963,
    n220
  );


  not
  g1080
  (
    n885,
    n269
  );


  not
  g1081
  (
    n911,
    n177
  );


  buf
  g1082
  (
    n1444,
    n568
  );


  not
  g1083
  (
    n1278,
    n402
  );


  not
  g1084
  (
    n955,
    n536
  );


  not
  g1085
  (
    n923,
    n308
  );


  not
  g1086
  (
    n1225,
    n360
  );


  not
  g1087
  (
    n1368,
    n524
  );


  not
  g1088
  (
    n948,
    n367
  );


  buf
  g1089
  (
    n699,
    n347
  );


  not
  g1090
  (
    n1170,
    n162
  );


  buf
  g1091
  (
    n1365,
    n563
  );


  buf
  g1092
  (
    n778,
    n453
  );


  buf
  g1093
  (
    n882,
    n464
  );


  not
  g1094
  (
    n926,
    n565
  );


  buf
  g1095
  (
    n1326,
    n274
  );


  buf
  g1096
  (
    n772,
    n260
  );


  not
  g1097
  (
    n1342,
    n537
  );


  buf
  g1098
  (
    n770,
    n394
  );


  not
  g1099
  (
    n888,
    n483
  );


  not
  g1100
  (
    n872,
    n287
  );


  buf
  g1101
  (
    n1403,
    n330
  );


  buf
  g1102
  (
    n835,
    n326
  );


  buf
  g1103
  (
    n1340,
    n285
  );


  buf
  g1104
  (
    n1328,
    n418
  );


  not
  g1105
  (
    n929,
    n512
  );


  buf
  g1106
  (
    n765,
    n532
  );


  not
  g1107
  (
    n1125,
    n234
  );


  buf
  g1108
  (
    n1404,
    n355
  );


  buf
  g1109
  (
    n1218,
    n532
  );


  not
  g1110
  (
    n857,
    n536
  );


  buf
  g1111
  (
    n1384,
    n516
  );


  not
  g1112
  (
    n774,
    n219
  );


  not
  g1113
  (
    n868,
    n395
  );


  not
  g1114
  (
    n751,
    n563
  );


  buf
  g1115
  (
    n1005,
    n204
  );


  buf
  g1116
  (
    n860,
    n381
  );


  buf
  g1117
  (
    n1446,
    n409
  );


  buf
  g1118
  (
    n970,
    n182
  );


  not
  g1119
  (
    n1065,
    n230
  );


  not
  g1120
  (
    n1211,
    n227
  );


  not
  g1121
  (
    n1385,
    n176
  );


  not
  g1122
  (
    n1154,
    n390
  );


  not
  g1123
  (
    n689,
    n338
  );


  buf
  g1124
  (
    n1146,
    n435
  );


  buf
  g1125
  (
    n864,
    n352
  );


  not
  g1126
  (
    n705,
    n297
  );


  not
  g1127
  (
    KeyWire_0_2,
    n408
  );


  not
  g1128
  (
    n1341,
    n280
  );


  not
  g1129
  (
    n679,
    n174
  );


  not
  g1130
  (
    n849,
    n282
  );


  buf
  g1131
  (
    n1275,
    n539
  );


  not
  g1132
  (
    n1202,
    n440
  );


  buf
  g1133
  (
    n1452,
    n358
  );


  not
  g1134
  (
    n1215,
    n188
  );


  buf
  g1135
  (
    n838,
    n441
  );


  not
  g1136
  (
    n1192,
    n177
  );


  not
  g1137
  (
    n677,
    n169
  );


  nand
  g1138
  (
    n681,
    n178,
    n443,
    n439,
    n197
  );


  xor
  g1139
  (
    n1012,
    n280,
    n544,
    n500,
    n243
  );


  xor
  g1140
  (
    n989,
    n519,
    n201,
    n404,
    n554
  );


  and
  g1141
  (
    n1320,
    n185,
    n505,
    n332,
    n445
  );


  xor
  g1142
  (
    n1214,
    n195,
    n173,
    n340,
    n237
  );


  xor
  g1143
  (
    n735,
    n498,
    n559,
    n534,
    n566
  );


  and
  g1144
  (
    n1350,
    n405,
    n389,
    n363,
    n456
  );


  and
  g1145
  (
    n1114,
    n343,
    n166,
    n414,
    n270
  );


  and
  g1146
  (
    n880,
    n528,
    n201,
    n163,
    n194
  );


  nand
  g1147
  (
    n1273,
    n378,
    n195,
    n175,
    n339
  );


  nor
  g1148
  (
    n968,
    n340,
    n481,
    n339,
    n405
  );


  or
  g1149
  (
    n1400,
    n168,
    n341,
    n375,
    n199
  );


  xnor
  g1150
  (
    n1390,
    n366,
    n566,
    n529,
    n324
  );


  xnor
  g1151
  (
    n1216,
    n533,
    n261,
    n309,
    n492
  );


  nor
  g1152
  (
    n1356,
    n550,
    n384,
    n567,
    n507
  );


  xor
  g1153
  (
    n1308,
    n403,
    n539,
    n322,
    n451
  );


  or
  g1154
  (
    n947,
    n223,
    n417,
    n212,
    n306
  );


  xnor
  g1155
  (
    n1429,
    n504,
    n426,
    n396,
    n462
  );


  xnor
  g1156
  (
    n844,
    n395,
    n493,
    n355,
    n290
  );


  xor
  g1157
  (
    n981,
    n340,
    n494,
    n480,
    n309
  );


  or
  g1158
  (
    n1172,
    n442,
    n366,
    n506,
    n380
  );


  and
  g1159
  (
    n1355,
    n311,
    n207,
    n266,
    n162
  );


  xnor
  g1160
  (
    n1252,
    n356,
    n528,
    n407,
    n511
  );


  and
  g1161
  (
    n831,
    n193,
    n303,
    n469,
    n291
  );


  and
  g1162
  (
    n1083,
    n184,
    n342,
    n419,
    n239
  );


  or
  g1163
  (
    n914,
    n277,
    n231,
    n166,
    n232
  );


  nor
  g1164
  (
    n1336,
    n557,
    n297,
    n295,
    n299
  );


  nand
  g1165
  (
    n1445,
    n522,
    n321,
    n350,
    n556
  );


  nor
  g1166
  (
    n1110,
    n275,
    n445,
    n283,
    n333
  );


  and
  g1167
  (
    n960,
    n290,
    n293,
    n300,
    n447
  );


  nand
  g1168
  (
    n952,
    n512,
    n218,
    n244,
    n438
  );


  and
  g1169
  (
    n1242,
    n423,
    n537,
    n259,
    n548
  );


  nand
  g1170
  (
    n1150,
    n419,
    n188,
    n459,
    n535
  );


  and
  g1171
  (
    n1441,
    n191,
    n339,
    n500,
    n356
  );


  xor
  g1172
  (
    n922,
    n221,
    n458,
    n475,
    n540
  );


  nor
  g1173
  (
    n1290,
    n493,
    n276,
    n194,
    n458
  );


  xnor
  g1174
  (
    n1330,
    n466,
    n499,
    n434,
    n490
  );


  xor
  g1175
  (
    n841,
    n461,
    n198,
    n305,
    n325
  );


  xnor
  g1176
  (
    n867,
    n447,
    n224,
    n466,
    n258
  );


  xnor
  g1177
  (
    n1263,
    n416,
    n337,
    n353,
    n275
  );


  xnor
  g1178
  (
    n781,
    n373,
    n415,
    n528,
    n183
  );


  or
  g1179
  (
    n1289,
    n353,
    n379,
    n342,
    n453
  );


  xor
  g1180
  (
    n763,
    n416,
    n285,
    n210,
    n272
  );


  or
  g1181
  (
    n912,
    n303,
    n499,
    n289,
    n390
  );


  or
  g1182
  (
    n1319,
    n471,
    n336,
    n460,
    n452
  );


  xnor
  g1183
  (
    n800,
    n364,
    n559,
    n310,
    n280
  );


  or
  g1184
  (
    n1416,
    n502,
    n378,
    n530,
    n510
  );


  xnor
  g1185
  (
    n941,
    n442,
    n417,
    n374,
    n392
  );


  xnor
  g1186
  (
    n1148,
    n236,
    n239,
    n184,
    n536
  );


  xnor
  g1187
  (
    n777,
    n378,
    n322,
    n430,
    n537
  );


  nand
  g1188
  (
    n730,
    n257,
    n448,
    n255,
    n488
  );


  or
  g1189
  (
    n1240,
    n169,
    n566,
    n335,
    n416
  );


  nand
  g1190
  (
    n750,
    n421,
    n449,
    n325,
    n553
  );


  xor
  g1191
  (
    n1144,
    n491,
    n278,
    n196,
    n466
  );


  xor
  g1192
  (
    n1420,
    n545,
    n178,
    n554,
    n212
  );


  nand
  g1193
  (
    n759,
    n519,
    n356,
    n396
  );


  nor
  g1194
  (
    n1050,
    n303,
    n413,
    n384,
    n421
  );


  xor
  g1195
  (
    n1040,
    n165,
    n426,
    n307,
    n502
  );


  nand
  g1196
  (
    n704,
    n305,
    n277,
    n247,
    n532
  );


  nor
  g1197
  (
    n1371,
    n509,
    n337,
    n463,
    n306
  );


  xnor
  g1198
  (
    n700,
    n277,
    n404,
    n223,
    n460
  );


  nor
  g1199
  (
    n1138,
    n176,
    n463,
    n181,
    n423
  );


  nor
  g1200
  (
    n675,
    n208,
    n200,
    n496,
    n503
  );


  or
  g1201
  (
    n1391,
    n474,
    n238,
    n540,
    n441
  );


  xnor
  g1202
  (
    n1449,
    n417,
    n433,
    n217,
    n347
  );


  or
  g1203
  (
    n1370,
    n541,
    n550,
    n523,
    n376
  );


  and
  g1204
  (
    n743,
    n491,
    n504,
    n379,
    n422
  );


  nor
  g1205
  (
    n1220,
    n532,
    n287,
    n486,
    n334
  );


  xnor
  g1206
  (
    n1346,
    n523,
    n527,
    n251,
    n265
  );


  nor
  g1207
  (
    n1437,
    n547,
    n534,
    n519,
    n445
  );


  and
  g1208
  (
    n762,
    n485,
    n399,
    n542,
    n365
  );


  nor
  g1209
  (
    n1008,
    n545,
    n367,
    n510,
    n363
  );


  xor
  g1210
  (
    n1310,
    n330,
    n429,
    n377,
    n354
  );


  xor
  g1211
  (
    n793,
    n224,
    n547,
    n390,
    n185
  );


  xnor
  g1212
  (
    n1453,
    n452,
    n544,
    n321,
    n197
  );


  and
  g1213
  (
    n1345,
    n442,
    n364,
    n345,
    n373
  );


  nand
  g1214
  (
    n802,
    n231,
    n521,
    n169,
    n381
  );


  and
  g1215
  (
    n892,
    n261,
    n523,
    n509,
    n544
  );


  nor
  g1216
  (
    n1017,
    n385,
    n503,
    n265,
    n472
  );


  xor
  g1217
  (
    n1300,
    n435,
    n286,
    n570,
    n171
  );


  or
  g1218
  (
    n1335,
    n243,
    n561,
    n520,
    n315
  );


  or
  g1219
  (
    n1454,
    n429,
    n273,
    n267,
    n395
  );


  nand
  g1220
  (
    n1047,
    n543,
    n296,
    n256,
    n517
  );


  nand
  g1221
  (
    n775,
    n191,
    n499,
    n421,
    n283
  );


  xor
  g1222
  (
    n979,
    n289,
    n489,
    n514,
    n387
  );


  or
  g1223
  (
    n1393,
    n457,
    n322,
    n313,
    n482
  );


  and
  g1224
  (
    n903,
    n177,
    n274,
    n172,
    n427
  );


  xnor
  g1225
  (
    n803,
    n567,
    n171,
    n346,
    n427
  );


  xor
  g1226
  (
    n1151,
    n444,
    n256,
    n249,
    n471
  );


  nand
  g1227
  (
    n1232,
    n394,
    n445,
    n376,
    n567
  );


  or
  g1228
  (
    n1099,
    n259,
    n295,
    n449,
    n291
  );


  xnor
  g1229
  (
    n986,
    n507,
    n381,
    n266,
    n478
  );


  xnor
  g1230
  (
    n813,
    n456,
    n512,
    n244,
    n508
  );


  nand
  g1231
  (
    n827,
    n250,
    n270,
    n275,
    n443
  );


  xor
  g1232
  (
    n1380,
    n564,
    n341,
    n415,
    n359
  );


  xnor
  g1233
  (
    n1267,
    n169,
    n362,
    n190,
    n204
  );


  nor
  g1234
  (
    n934,
    n506,
    n230,
    n233,
    n392
  );


  nand
  g1235
  (
    n1338,
    n485,
    n398,
    n268,
    n455
  );


  xor
  g1236
  (
    n862,
    n274,
    n437,
    n347,
    n228
  );


  xor
  g1237
  (
    n786,
    n299,
    n202,
    n253,
    n234
  );


  xor
  g1238
  (
    n1086,
    n202,
    n400,
    n272,
    n412
  );


  xor
  g1239
  (
    n1073,
    n289,
    n229,
    n264,
    n422
  );


  xor
  g1240
  (
    n978,
    n397,
    n271,
    n286,
    n340
  );


  and
  g1241
  (
    n1401,
    n497,
    n161,
    n304,
    n383
  );


  nand
  g1242
  (
    n789,
    n344,
    n189,
    n553,
    n406
  );


  or
  g1243
  (
    n1129,
    n494,
    n483,
    n296,
    n518
  );


  or
  g1244
  (
    n1312,
    n455,
    n288,
    n200,
    n248
  );


  nand
  g1245
  (
    n1070,
    n172,
    n207,
    n394,
    n222
  );


  and
  g1246
  (
    n1257,
    n391,
    n529,
    n200,
    n302
  );


  nand
  g1247
  (
    n962,
    n271,
    n393,
    n300,
    n186
  );


  nand
  g1248
  (
    n1309,
    n357,
    n541,
    n276,
    n482
  );


  and
  g1249
  (
    n1255,
    n387,
    n533,
    n346,
    n367
  );


  xnor
  g1250
  (
    n883,
    n375,
    n427,
    n490,
    n318
  );


  xor
  g1251
  (
    n1077,
    n290,
    n376,
    n382,
    n388
  );


  or
  g1252
  (
    n957,
    n407,
    n534,
    n498,
    n194
  );


  or
  g1253
  (
    n945,
    n211,
    n307,
    n558,
    n424
  );


  nor
  g1254
  (
    n1066,
    n162,
    n278,
    n173,
    n345
  );


  nor
  g1255
  (
    n818,
    n539,
    n288,
    n267,
    n524
  );


  nor
  g1256
  (
    n1141,
    n292,
    n335,
    n552,
    n476
  );


  or
  g1257
  (
    n991,
    n215,
    n470,
    n213,
    n327
  );


  xnor
  g1258
  (
    n1450,
    n196,
    n216,
    n444,
    n414
  );


  nand
  g1259
  (
    n1195,
    n510,
    n324,
    n167,
    n531
  );


  xnor
  g1260
  (
    n1349,
    n329,
    n254,
    n566,
    n443
  );


  xnor
  g1261
  (
    n1455,
    n527,
    n366,
    n446,
    n310
  );


  nor
  g1262
  (
    n1294,
    n505,
    n204,
    n409,
    n480
  );


  xnor
  g1263
  (
    n1169,
    n240,
    n468,
    n406,
    n460
  );


  xnor
  g1264
  (
    n1108,
    n316,
    n270,
    n454,
    n370
  );


  xor
  g1265
  (
    n1236,
    n206,
    n431,
    n565,
    n350
  );


  xor
  g1266
  (
    n1033,
    n522,
    n408,
    n278,
    n564
  );


  nand
  g1267
  (
    n1245,
    n323,
    n293,
    n238,
    n161
  );


  nand
  g1268
  (
    n830,
    n477,
    n229,
    n451,
    n489
  );


  xnor
  g1269
  (
    n673,
    n173,
    n338,
    n273,
    n447
  );


  nor
  g1270
  (
    n828,
    n450,
    n267,
    n362,
    n276
  );


  xor
  g1271
  (
    n801,
    n379,
    n464,
    n289,
    n260
  );


  nand
  g1272
  (
    n1233,
    n256,
    n471,
    n313,
    n197
  );


  and
  g1273
  (
    n852,
    n555,
    n488,
    n196,
    n251
  );


  or
  g1274
  (
    n856,
    n168,
    n219,
    n308,
    n428
  );


  and
  g1275
  (
    n1029,
    n400,
    n528,
    n183,
    n353
  );


  and
  g1276
  (
    n1143,
    n371,
    n246,
    n306,
    n463
  );


  and
  g1277
  (
    n1291,
    n307,
    n314,
    n219,
    n364
  );


  nor
  g1278
  (
    n1331,
    n175,
    n317,
    n284,
    n456
  );


  nor
  g1279
  (
    n737,
    n326,
    n346,
    n487,
    n179
  );


  and
  g1280
  (
    n1402,
    n220,
    n555,
    n479,
    n353
  );


  nand
  g1281
  (
    n1292,
    n468,
    n397,
    n473,
    n298
  );


  and
  g1282
  (
    n688,
    n166,
    n168,
    n396,
    n531
  );


  or
  g1283
  (
    n1362,
    n402,
    n173,
    n292,
    n242
  );


  xnor
  g1284
  (
    n1054,
    n374,
    n543,
    n398,
    n538
  );


  nand
  g1285
  (
    n755,
    n213,
    n225,
    n525,
    n203
  );


  nor
  g1286
  (
    n1069,
    n438,
    n294,
    n439,
    n372
  );


  nand
  g1287
  (
    n788,
    n568,
    n250,
    n569,
    n481
  );


  or
  g1288
  (
    n959,
    n202,
    n412,
    n214,
    n474
  );


  nor
  g1289
  (
    n980,
    n388,
    n444,
    n472,
    n467
  );


  and
  g1290
  (
    n1268,
    n323,
    n332,
    n230,
    n530
  );


  or
  g1291
  (
    n1425,
    n551,
    n299,
    n469,
    n556
  );


  or
  g1292
  (
    n1372,
    n410,
    n222,
    n469,
    n370
  );


  nor
  g1293
  (
    n729,
    n508,
    n257,
    n170,
    n232
  );


  and
  g1294
  (
    n1101,
    n312,
    n358,
    n386,
    n565
  );


  nand
  g1295
  (
    n921,
    n443,
    n385,
    n397,
    n216
  );


  xnor
  g1296
  (
    n1204,
    n515,
    n351,
    n256,
    n553
  );


  xor
  g1297
  (
    n983,
    n235,
    n178,
    n167,
    n562
  );


  xnor
  g1298
  (
    n1260,
    n504,
    n323,
    n225,
    n380
  );


  and
  g1299
  (
    n1094,
    n209,
    n497,
    n370,
    n381
  );


  xnor
  g1300
  (
    n1277,
    n317,
    n552,
    n459,
    n324
  );


  xor
  g1301
  (
    n1176,
    n349,
    n228,
    n369,
    n397
  );


  and
  g1302
  (
    n1305,
    n253,
    n446,
    n422,
    n314
  );


  xor
  g1303
  (
    n797,
    n533,
    n448,
    n230,
    n327
  );


  nor
  g1304
  (
    n876,
    n366,
    n282,
    n514,
    n351
  );


  xor
  g1305
  (
    KeyWire_0_7,
    n484,
    n365,
    n299,
    n467
  );


  nand
  g1306
  (
    n1082,
    n311,
    n286,
    n261,
    n560
  );


  nand
  g1307
  (
    n780,
    n411,
    n410,
    n217,
    n377
  );


  and
  g1308
  (
    KeyWire_0_10,
    n483,
    n319,
    n349,
    n329
  );


  nand
  g1309
  (
    n1382,
    n343,
    n219,
    n454,
    n455
  );


  xor
  g1310
  (
    n837,
    n255,
    n398,
    n436,
    n372
  );


  or
  g1311
  (
    n973,
    n312,
    n431,
    n279,
    n435
  );


  nor
  g1312
  (
    n950,
    n284,
    n312,
    n508,
    n255
  );


  and
  g1313
  (
    n1307,
    n489,
    n513,
    n495,
    n377
  );


  nand
  g1314
  (
    n822,
    n172,
    n424,
    n184,
    n450
  );


  xnor
  g1315
  (
    n1000,
    n473,
    n240,
    n456,
    n563
  );


  xnor
  g1316
  (
    n1087,
    n205,
    n521,
    n439,
    n408
  );


  xnor
  g1317
  (
    n821,
    n241,
    n212,
    n332,
    n389
  );


  xor
  g1318
  (
    n1011,
    n380,
    n198,
    n454,
    n460
  );


  nor
  g1319
  (
    n933,
    n408,
    n194,
    n285,
    n441
  );


  xor
  g1320
  (
    n1432,
    n481,
    n254,
    n187,
    n226
  );


  xor
  g1321
  (
    n1061,
    n413,
    n186,
    n436,
    n450
  );


  and
  g1322
  (
    n1358,
    n307,
    n265,
    n165,
    n204
  );


  or
  g1323
  (
    n985,
    n223,
    n337,
    n469,
    n384
  );


  xor
  g1324
  (
    n1378,
    n271,
    n236,
    n305,
    n328
  );


  xnor
  g1325
  (
    n875,
    n524,
    n306,
    n473,
    n440
  );


  xor
  g1326
  (
    n710,
    n483,
    n530,
    n315,
    n320
  );


  xnor
  g1327
  (
    n752,
    n279,
    n203,
    n301,
    n546
  );


  or
  g1328
  (
    n1123,
    n192,
    n167,
    n267,
    n217
  );


  nand
  g1329
  (
    n1037,
    n296,
    n198,
    n348,
    n316
  );


  xor
  g1330
  (
    n1359,
    n203,
    n226,
    n233,
    n540
  );


  xor
  g1331
  (
    n701,
    n236,
    n201,
    n315,
    n471
  );


  nor
  g1332
  (
    n1159,
    n296,
    n183,
    n298,
    n411
  );


  nor
  g1333
  (
    n928,
    n371,
    n182,
    n549,
    n331
  );


  or
  g1334
  (
    n1116,
    n490,
    n253,
    n488,
    n377
  );


  and
  g1335
  (
    n1386,
    n525,
    n429,
    n225,
    n247
  );


  xnor
  g1336
  (
    n766,
    n280,
    n222,
    n419,
    n214
  );


  xor
  g1337
  (
    n1287,
    n540,
    n441,
    n570,
    n378
  );


  nor
  g1338
  (
    n1056,
    n474,
    n258,
    n354,
    n328
  );


  nor
  g1339
  (
    n1153,
    n488,
    n344,
    n324,
    n218
  );


  or
  g1340
  (
    n706,
    n313,
    n283,
    n541,
    n434
  );


  nand
  g1341
  (
    n1447,
    n357,
    n496,
    n211,
    n387
  );


  or
  g1342
  (
    n711,
    n317,
    n250,
    n227,
    n558
  );


  or
  g1343
  (
    n749,
    n271,
    n291,
    n288,
    n186
  );


  or
  g1344
  (
    n1353,
    n360,
    n206,
    n273,
    n190
  );


  nand
  g1345
  (
    n1253,
    n374,
    n213,
    n400,
    n369
  );


  nor
  g1346
  (
    n1381,
    n318,
    n278,
    n542,
    n295
  );


  and
  g1347
  (
    n961,
    n212,
    n197,
    n512,
    n348
  );


  xnor
  g1348
  (
    n863,
    n561,
    n382,
    n270,
    n497
  );


  nand
  g1349
  (
    n717,
    n297,
    n308,
    n200,
    n479
  );


  and
  g1350
  (
    n1015,
    n424,
    n286,
    n358,
    n434
  );


  and
  g1351
  (
    n1383,
    n432,
    n161,
    n218,
    n501
  );


  xnor
  g1352
  (
    n1387,
    n314,
    n371,
    n300,
    n551
  );


  and
  g1353
  (
    n791,
    n251,
    n393,
    n511,
    n341
  );


  xnor
  g1354
  (
    n1351,
    n383,
    n264,
    n447,
    n511
  );


  xnor
  g1355
  (
    n1209,
    n339,
    n187,
    n487,
    n232
  );


  or
  g1356
  (
    n886,
    n466,
    n329,
    n507,
    n162
  );


  and
  g1357
  (
    n924,
    n364,
    n181,
    n355,
    n399
  );


  or
  g1358
  (
    n1411,
    n376,
    n241,
    n179,
    n524
  );


  xnor
  g1359
  (
    n796,
    n205,
    n477,
    n508,
    n560
  );


  xor
  g1360
  (
    n1136,
    n281,
    n520,
    n430,
    n555
  );


  nand
  g1361
  (
    n1408,
    n252,
    n215,
    n221,
    n425
  );


  nor
  g1362
  (
    n1231,
    n263,
    n530,
    n401,
    n192
  );


  xor
  g1363
  (
    n808,
    n245,
    n248,
    n535,
    n553
  );


  xor
  g1364
  (
    n899,
    n291,
    n506,
    n359,
    n557
  );


  xnor
  g1365
  (
    n1021,
    n242,
    n375,
    n223,
    n208
  );


  or
  g1366
  (
    n1212,
    n315,
    n476,
    n211,
    n327
  );


  xor
  g1367
  (
    n1316,
    n562,
    n363,
    n161,
    n354
  );


  nand
  g1368
  (
    n900,
    n401,
    n415,
    n382,
    n544
  );


  xor
  g1369
  (
    n1418,
    n561,
    n328,
    n384,
    n181
  );


  nor
  g1370
  (
    n731,
    n292,
    n360,
    n518,
    n325
  );


  nand
  g1371
  (
    n1166,
    n478,
    n168,
    n465,
    n373
  );


  and
  g1372
  (
    n939,
    n234,
    n170,
    n538,
    n311
  );


  xnor
  g1373
  (
    n1189,
    n189,
    n245,
    n259,
    n254
  );


  xor
  g1374
  (
    n1198,
    n171,
    n500,
    n380,
    n556
  );


  nand
  g1375
  (
    n1057,
    n352,
    n551,
    n426,
    n525
  );


  nand
  g1376
  (
    n866,
    n501,
    n388,
    n420,
    n164
  );


  nand
  g1377
  (
    n676,
    n546,
    n558,
    n467,
    n517
  );


  and
  g1378
  (
    n1282,
    n568,
    n560,
    n396,
    n351
  );


  nor
  g1379
  (
    n739,
    n526,
    n438,
    n263,
    n185
  );


  or
  g1380
  (
    n1081,
    n362,
    n227,
    n350,
    n543
  );


  nor
  g1381
  (
    n1327,
    n355,
    n554,
    n345,
    n392
  );


  nor
  g1382
  (
    n1183,
    n244,
    n228,
    n310,
    n542
  );


  xnor
  g1383
  (
    n824,
    n413,
    n344,
    n477,
    n274
  );


  and
  g1384
  (
    n1301,
    n243,
    n437,
    n334,
    n210
  );


  xnor
  g1385
  (
    n1248,
    n327,
    n206,
    n259,
    n240
  );


  nor
  g1386
  (
    n1063,
    n338,
    n183,
    n172,
    n478
  );


  and
  g1387
  (
    n1281,
    n495,
    n446,
    n526,
    n385
  );


  xor
  g1388
  (
    n832,
    n252,
    n272,
    n496,
    n414
  );


  and
  g1389
  (
    n1162,
    n295,
    n452,
    n559,
    n403
  );


  nor
  g1390
  (
    n1028,
    n342,
    n175,
    n337,
    n520
  );


  and
  g1391
  (
    n1230,
    n416,
    n444,
    n361,
    n362
  );


  nand
  g1392
  (
    n1187,
    n415,
    n375,
    n550,
    n283
  );


  nand
  g1393
  (
    n1251,
    n386,
    n238,
    n262,
    n322
  );


  nor
  g1394
  (
    n1167,
    n245,
    n537,
    n438,
    n392
  );


  xor
  g1395
  (
    n1244,
    n526,
    n493,
    n449,
    n515
  );


  nand
  g1396
  (
    n1200,
    n448,
    n425,
    n367,
    n522
  );


  xor
  g1397
  (
    n855,
    n394,
    n398,
    n569,
    n558
  );


  nand
  g1398
  (
    n708,
    n326,
    n368,
    n492,
    n189
  );


  nand
  g1399
  (
    n1133,
    n432,
    n464,
    n418,
    n319
  );


  and
  g1400
  (
    n909,
    n371,
    n348,
    n567,
    n509
  );


  and
  g1401
  (
    n1018,
    n277,
    n193,
    n458,
    n248
  );


  nor
  g1402
  (
    n1016,
    n372,
    n514,
    n216,
    n190
  );


  nand
  g1403
  (
    n733,
    n164,
    n513,
    n166,
    n191
  );


  nor
  g1404
  (
    n782,
    n402,
    n214,
    n551,
    n519
  );


  nor
  g1405
  (
    n1398,
    n297,
    n165,
    n468,
    n301
  );


  nand
  g1406
  (
    n1074,
    n276,
    n568,
    n548,
    n523
  );


  or
  g1407
  (
    n1221,
    n525,
    n493,
    n246,
    n455
  );


  nand
  g1408
  (
    n814,
    n279,
    n332,
    n275,
    n557
  );


  and
  g1409
  (
    n975,
    n382,
    n463,
    n529,
    n237
  );


  xnor
  g1410
  (
    n1430,
    n436,
    n241,
    n475,
    n214
  );


  nor
  g1411
  (
    n707,
    n281,
    n420,
    n316,
    n516
  );


  nand
  g1412
  (
    n1149,
    n470,
    n354,
    n516,
    n260
  );


  or
  g1413
  (
    n1118,
    n484,
    n536,
    n304,
    n312
  );


  xor
  g1414
  (
    n1179,
    n420,
    n290,
    n188,
    n436
  );


  xor
  g1415
  (
    n721,
    n510,
    n320,
    n281,
    n485
  );


  nor
  g1416
  (
    n1427,
    n284,
    n503,
    n498,
    n549
  );


  nor
  g1417
  (
    n734,
    n352,
    n182,
    n279,
    n261
  );


  and
  g1418
  (
    n1283,
    n226,
    n424,
    n451,
    n409
  );


  or
  g1419
  (
    n1199,
    n461,
    n509,
    n251,
    n369
  );


  and
  g1420
  (
    n1339,
    n304,
    n548,
    n490,
    n552
  );


  xnor
  g1421
  (
    n910,
    n244,
    n401,
    n565,
    n374
  );


  nand
  g1422
  (
    n1160,
    n406,
    n205,
    n402,
    n400
  );


  nand
  g1423
  (
    n1723,
    n729,
    n1240,
    n1305,
    n1038
  );


  nand
  g1424
  (
    n1604,
    n1164,
    n1172,
    n852,
    n731
  );


  or
  g1425
  (
    n1661,
    n789,
    n1296,
    n753,
    n1239
  );


  and
  g1426
  (
    n1539,
    n966,
    n1117,
    n1081,
    n1263
  );


  xor
  g1427
  (
    n1496,
    n810,
    n1259,
    n1277,
    n1110
  );


  nor
  g1428
  (
    n1501,
    n774,
    n926,
    n1248,
    n855
  );


  nand
  g1429
  (
    n1636,
    n1207,
    n898,
    n725,
    n1205
  );


  nand
  g1430
  (
    n1738,
    n936,
    n1048,
    n1220,
    n835
  );


  and
  g1431
  (
    n1813,
    n746,
    n1094,
    n1168,
    n1133
  );


  or
  g1432
  (
    n1789,
    n1112,
    n799,
    n1078,
    n683
  );


  xnor
  g1433
  (
    n1671,
    n1069,
    n1174,
    n1054,
    n1204
  );


  and
  g1434
  (
    n1668,
    n1149,
    n1287,
    n1265,
    n1218
  );


  and
  g1435
  (
    n1515,
    n1082,
    n1205,
    n798,
    n1308
  );


  xor
  g1436
  (
    n1649,
    n717,
    n1052,
    n791,
    n1106
  );


  and
  g1437
  (
    n1602,
    n1178,
    n1140,
    n1046
  );


  nor
  g1438
  (
    n1729,
    n730,
    n1048,
    n1279
  );


  xnor
  g1439
  (
    n1489,
    n1134,
    n1103,
    n946,
    n1127
  );


  and
  g1440
  (
    n1562,
    n887,
    n1301,
    n865,
    n991
  );


  xor
  g1441
  (
    n1590,
    n733,
    n1301,
    n739,
    n1112
  );


  xor
  g1442
  (
    n1566,
    n1174,
    n1280,
    n1022,
    n1100
  );


  and
  g1443
  (
    n1804,
    n1214,
    n924,
    n1030,
    n1213
  );


  or
  g1444
  (
    n1462,
    n1216,
    n1195,
    n1047,
    n1222
  );


  or
  g1445
  (
    n1619,
    n1045,
    n1160,
    n1251,
    n1199
  );


  nand
  g1446
  (
    n1548,
    n1198,
    n689,
    n1295,
    n876
  );


  xnor
  g1447
  (
    n1537,
    n1146,
    n1209,
    n1155,
    n1285
  );


  or
  g1448
  (
    n1512,
    n932,
    n947,
    n1200,
    n823
  );


  nor
  g1449
  (
    n1825,
    n1193,
    n1200,
    n1154,
    n1134
  );


  and
  g1450
  (
    n1513,
    n1230,
    n883,
    n1152,
    n1225
  );


  nand
  g1451
  (
    n1497,
    n1209,
    n1245,
    n1111,
    n1083
  );


  and
  g1452
  (
    n1592,
    n812,
    n716,
    n1267,
    n856
  );


  or
  g1453
  (
    n1805,
    n1053,
    n1101,
    n1288,
    n1208
  );


  xnor
  g1454
  (
    n1646,
    n1027,
    n1109,
    n1262,
    n1308
  );


  nand
  g1455
  (
    n1568,
    n1049,
    n1121,
    n727,
    n864
  );


  nor
  g1456
  (
    n1586,
    n1174,
    n1125,
    n1141,
    n1309
  );


  or
  g1457
  (
    n1521,
    n1069,
    n1252,
    n1180,
    n1102
  );


  nand
  g1458
  (
    n1616,
    n1208,
    n1002,
    n1050,
    n901
  );


  and
  g1459
  (
    n1612,
    n1109,
    n1235,
    n1124,
    n1188
  );


  xor
  g1460
  (
    n1480,
    n1272,
    n1029,
    n1010,
    n1211
  );


  nor
  g1461
  (
    n1570,
    n1226,
    n1208,
    n684,
    n1266
  );


  or
  g1462
  (
    n1599,
    n1213,
    n1200,
    n1286,
    n1235
  );


  xor
  g1463
  (
    n1818,
    n1021,
    n760,
    n766,
    n1018
  );


  nor
  g1464
  (
    n1740,
    n1218,
    n1217,
    n944,
    n826
  );


  nor
  g1465
  (
    n1719,
    n1086,
    n1019,
    n1263,
    n1203
  );


  and
  g1466
  (
    n1603,
    n1236,
    n1280,
    n1127,
    n1257
  );


  xor
  g1467
  (
    n1531,
    n1004,
    n1078,
    n1143,
    n1067
  );


  nand
  g1468
  (
    n1808,
    n912,
    n1241,
    n1159,
    n1118
  );


  xnor
  g1469
  (
    n1508,
    n1117,
    n1251,
    n1104,
    n1160
  );


  xnor
  g1470
  (
    n1494,
    n1236,
    n1258,
    n1132,
    n1268
  );


  and
  g1471
  (
    n1742,
    n1210,
    n1006,
    n1255,
    n1039
  );


  xnor
  g1472
  (
    n1575,
    n1124,
    n1304,
    n1261,
    n1169
  );


  nor
  g1473
  (
    n1609,
    n1186,
    n986,
    n1241,
    n1057
  );


  nor
  g1474
  (
    n1734,
    n1249,
    n1149,
    n906,
    n719
  );


  xnor
  g1475
  (
    n1682,
    n1150,
    n1233,
    n1193,
    n1194
  );


  xor
  g1476
  (
    n1736,
    n880,
    n763,
    n1081,
    n1192
  );


  nand
  g1477
  (
    n1746,
    n801,
    n1222,
    n1149,
    n1025
  );


  xor
  g1478
  (
    n1544,
    n1310,
    n1304,
    n1262,
    n1011
  );


  nor
  g1479
  (
    n1666,
    n1210,
    n1277,
    n1087,
    n1004
  );


  nand
  g1480
  (
    n1563,
    n1119,
    n1098,
    n896,
    n1230
  );


  xor
  g1481
  (
    n1755,
    n1015,
    n1275,
    n1163,
    n1059
  );


  xor
  g1482
  (
    n1553,
    n1009,
    n1154,
    n679,
    n879
  );


  nor
  g1483
  (
    n1510,
    n831,
    n1108,
    n1196,
    n1071
  );


  xor
  g1484
  (
    n1696,
    n1100,
    n802,
    n1308,
    n1085
  );


  xor
  g1485
  (
    n1713,
    n903,
    n1063,
    n1033,
    n1043
  );


  xor
  g1486
  (
    n1468,
    n1192,
    n1196,
    n1287,
    n1303
  );


  xor
  g1487
  (
    n1632,
    n1247,
    n1305,
    n1185,
    n829
  );


  xor
  g1488
  (
    n1624,
    n1147,
    n803,
    n1202,
    n960
  );


  nand
  g1489
  (
    n1556,
    n1092,
    n1228,
    n1276,
    n1160
  );


  or
  g1490
  (
    n1662,
    n1050,
    n680,
    n745,
    n1238
  );


  or
  g1491
  (
    n1795,
    n1169,
    n1221,
    n1222,
    n1255
  );


  nor
  g1492
  (
    n1718,
    n1309,
    n1135,
    n1261,
    n1102
  );


  xnor
  g1493
  (
    n1467,
    n1270,
    n1073,
    n1256,
    n1120
  );


  and
  g1494
  (
    n1552,
    n1232,
    n1151,
    n1063,
    n1041
  );


  xnor
  g1495
  (
    n1518,
    n1290,
    n1013,
    n1075,
    n976
  );


  nor
  g1496
  (
    n1773,
    n1179,
    n1121,
    n1262,
    n1096
  );


  xor
  g1497
  (
    n1584,
    n1154,
    n1300,
    n853,
    n1189
  );


  or
  g1498
  (
    n1765,
    n703,
    n917,
    n1255,
    n1259
  );


  nand
  g1499
  (
    n1461,
    n1270,
    n1145,
    n1168,
    n1272
  );


  xor
  g1500
  (
    n1703,
    n1019,
    n1127,
    n952,
    n1179
  );


  nor
  g1501
  (
    n1727,
    n1045,
    n1268,
    n1060,
    n712
  );


  xor
  g1502
  (
    n1751,
    n1076,
    n1212,
    n1203,
    n1066
  );


  or
  g1503
  (
    n1546,
    n1193,
    n1122,
    n1079,
    n1247
  );


  nand
  g1504
  (
    n1793,
    n941,
    n1269,
    n1036,
    n1206
  );


  or
  g1505
  (
    n1485,
    n1294,
    n1077,
    n1153,
    n764
  );


  nand
  g1506
  (
    n1761,
    n1032,
    n893,
    n1055,
    n889
  );


  xnor
  g1507
  (
    n1634,
    n1260,
    n1091,
    n697,
    n1070
  );


  or
  g1508
  (
    n1655,
    n685,
    n985,
    n1298,
    n1049
  );


  nand
  g1509
  (
    n1557,
    n1054,
    n1111,
    n817,
    n1151
  );


  xor
  g1510
  (
    n1694,
    n1290,
    n1204,
    n1098,
    n1310
  );


  and
  g1511
  (
    n1763,
    n1264,
    n1168,
    n1069,
    n1061
  );


  and
  g1512
  (
    n1555,
    n1119,
    n1071,
    n1307,
    n1123
  );


  and
  g1513
  (
    n1684,
    n845,
    n1075,
    n827,
    n1224
  );


  xor
  g1514
  (
    n1564,
    n1025,
    n1290,
    n1162,
    n1229
  );


  nand
  g1515
  (
    n1611,
    n1006,
    n776,
    n869,
    n1050
  );


  nor
  g1516
  (
    n1675,
    n1087,
    n850,
    n1090,
    n1170
  );


  nor
  g1517
  (
    n1528,
    n1113,
    n1214,
    n1107,
    n1161
  );


  or
  g1518
  (
    n1486,
    n1113,
    n1285,
    n1132,
    n1159
  );


  and
  g1519
  (
    n1645,
    n1074,
    n1052,
    n1123,
    n1136
  );


  xor
  g1520
  (
    n1629,
    n874,
    n1103,
    n1086,
    n1012
  );


  nand
  g1521
  (
    n1520,
    n1055,
    n1214,
    n1292,
    n1269
  );


  nand
  g1522
  (
    n1756,
    n1087,
    n1045,
    n1060,
    n1079
  );


  or
  g1523
  (
    n1667,
    n1061,
    n1176,
    n743,
    n1197
  );


  and
  g1524
  (
    n1591,
    n1084,
    n772,
    n1284,
    n1148
  );


  xnor
  g1525
  (
    n1759,
    n1166,
    n690,
    n1129,
    n822
  );


  xnor
  g1526
  (
    n1673,
    n1141,
    n1169,
    n1296,
    n1131
  );


  nand
  g1527
  (
    n1743,
    n1223,
    n1262,
    n1284,
    n1084
  );


  nand
  g1528
  (
    n1705,
    n1095,
    n934,
    n1131,
    n1159
  );


  and
  g1529
  (
    n1571,
    n1138,
    n1210,
    n1112,
    n1139
  );


  or
  g1530
  (
    n1551,
    n1306,
    n1020,
    n672,
    n1231
  );


  and
  g1531
  (
    n1504,
    n1081,
    n1232,
    n1046,
    n1093
  );


  xor
  g1532
  (
    n1782,
    n701,
    n940,
    n1097,
    n1104
  );


  xor
  g1533
  (
    n1500,
    n811,
    n1195,
    n1238,
    n1158
  );


  xor
  g1534
  (
    n1690,
    n1257,
    n1085,
    n1278,
    n841
  );


  nand
  g1535
  (
    n1472,
    n1137,
    n1281,
    n1167,
    n1258
  );


  xnor
  g1536
  (
    n1550,
    n1057,
    n1195,
    n965,
    n982
  );


  nand
  g1537
  (
    n1643,
    n935,
    n1066,
    n1142,
    n1289
  );


  nand
  g1538
  (
    n1752,
    n714,
    n752,
    n1169,
    n1274
  );


  nor
  g1539
  (
    n1771,
    n868,
    n771,
    n1056,
    n1234
  );


  xor
  g1540
  (
    n1683,
    n878,
    n735,
    n1212,
    n1098
  );


  and
  g1541
  (
    n1698,
    n1086,
    n1107,
    n709,
    n1226
  );


  xnor
  g1542
  (
    n1822,
    n1225,
    n700,
    n1122,
    n1106
  );


  nand
  g1543
  (
    n1583,
    n1260,
    n1295,
    n1201,
    n1182
  );


  nor
  g1544
  (
    n1790,
    n1283,
    n1303,
    n1156,
    n1204
  );


  xnor
  g1545
  (
    n1511,
    n1159,
    n1053,
    n1177,
    n1270
  );


  and
  g1546
  (
    n1498,
    n1094,
    n1275,
    n1183,
    n1135
  );


  xnor
  g1547
  (
    n1823,
    n1231,
    n870,
    n1267,
    n1105
  );


  xor
  g1548
  (
    n1796,
    n920,
    n1062,
    n1068,
    n1080
  );


  nand
  g1549
  (
    n1588,
    n1103,
    n1161,
    n1082,
    n1254
  );


  nor
  g1550
  (
    n1710,
    n828,
    n1000,
    n1176,
    n877
  );


  xor
  g1551
  (
    n1691,
    n972,
    n1292,
    n1265,
    n1099
  );


  and
  g1552
  (
    n1768,
    n1220,
    n1190,
    n1205,
    n796
  );


  or
  g1553
  (
    n1600,
    n820,
    n1071,
    n1161,
    n1075
  );


  or
  g1554
  (
    n1760,
    n854,
    n1059,
    n1147,
    n711
  );


  xor
  g1555
  (
    n1711,
    n998,
    n1283,
    n1093,
    n1246
  );


  and
  g1556
  (
    n1466,
    n1095,
    n968,
    n1298,
    n1224
  );


  nor
  g1557
  (
    n1799,
    n1176,
    n902,
    n1120,
    n1066
  );


  nand
  g1558
  (
    n1596,
    n925,
    n1252,
    n1306,
    n1085
  );


  nand
  g1559
  (
    n1493,
    n1181,
    n1168,
    n904,
    n1177
  );


  nor
  g1560
  (
    n1597,
    n1069,
    n1080,
    n967,
    n1229
  );


  or
  g1561
  (
    n1741,
    n1096,
    n1286,
    n698,
    n989
  );


  and
  g1562
  (
    n1569,
    n1104,
    n1215,
    n1023,
    n1034
  );


  xor
  g1563
  (
    n1465,
    n955,
    n1089,
    n1183,
    n1235
  );


  nand
  g1564
  (
    n1777,
    n1206,
    n1292,
    n995,
    n1080
  );


  xnor
  g1565
  (
    n1614,
    n1188,
    n1225,
    n1116,
    n1299
  );


  or
  g1566
  (
    n1639,
    n1138,
    n1049,
    n1181,
    n1219
  );


  nand
  g1567
  (
    n1700,
    n786,
    n1129,
    n702,
    n866
  );


  nor
  g1568
  (
    n1502,
    n1252,
    n1074,
    n1266,
    n1227
  );


  xnor
  g1569
  (
    n1664,
    n1225,
    n778,
    n1256,
    n1246
  );


  nor
  g1570
  (
    n1582,
    n1297,
    n958,
    n1288,
    n1250
  );


  and
  g1571
  (
    n1744,
    n1009,
    n1198,
    n814,
    n1083
  );


  and
  g1572
  (
    n1627,
    n1017,
    n1194,
    n1244,
    n805
  );


  nand
  g1573
  (
    n1618,
    n675,
    n1269,
    n1148,
    n734
  );


  and
  g1574
  (
    n1784,
    n1062,
    n994,
    n1104,
    n1046
  );


  xor
  g1575
  (
    n1826,
    n1220,
    n694,
    n833,
    n1035
  );


  nor
  g1576
  (
    n1473,
    n930,
    n678,
    n1137,
    n1053
  );


  and
  g1577
  (
    n1471,
    n886,
    n1089,
    n1179,
    n1007
  );


  xnor
  g1578
  (
    n1476,
    n1088,
    n882,
    n1126,
    n1091
  );


  and
  g1579
  (
    n1686,
    n1166,
    n1281,
    n1044,
    n1273
  );


  xor
  g1580
  (
    n1687,
    n964,
    n728,
    n1117,
    n1191
  );


  xnor
  g1581
  (
    n1534,
    n1067,
    n1073,
    n1131,
    n1283
  );


  xor
  g1582
  (
    n1491,
    n688,
    n1133,
    n1181,
    n1166
  );


  nor
  g1583
  (
    n1764,
    n1120,
    n1178,
    n806,
    n1227
  );


  nand
  g1584
  (
    n1578,
    n1081,
    n1274,
    n1094,
    n1213
  );


  and
  g1585
  (
    n1716,
    n1133,
    n1198,
    n1308,
    n867
  );


  nand
  g1586
  (
    n1469,
    n1289,
    n1157,
    n1036,
    n1300
  );


  or
  g1587
  (
    n1697,
    n1061,
    n1250,
    n1087,
    n1129
  );


  xnor
  g1588
  (
    n1458,
    n1146,
    n1171,
    n1038,
    n830
  );


  or
  g1589
  (
    n1625,
    n1183,
    n1248,
    n1190,
    n1088
  );


  xnor
  g1590
  (
    n1692,
    n1040,
    n1037,
    n1010,
    n809
  );


  xnor
  g1591
  (
    n1540,
    n1302,
    n1259,
    n1311,
    n1143
  );


  nand
  g1592
  (
    n1483,
    n1049,
    n1141,
    n1042,
    n1139
  );


  xor
  g1593
  (
    n1785,
    n1071,
    n1216,
    n978,
    n1101
  );


  and
  g1594
  (
    n1487,
    n1128,
    n1175,
    n1130,
    n1020
  );


  nor
  g1595
  (
    n1554,
    n1170,
    n1206,
    n1300,
    n1240
  );


  xor
  g1596
  (
    n1580,
    n1121,
    n1241,
    n1164,
    n758
  );


  nor
  g1597
  (
    n1622,
    n1116,
    n1279,
    n1229,
    n1129
  );


  nand
  g1598
  (
    n1648,
    n1301,
    n1068,
    n1195,
    n1001
  );


  xnor
  g1599
  (
    n1613,
    n1136,
    n1187,
    n1297,
    n1130
  );


  and
  g1600
  (
    n1620,
    n1239,
    n1022,
    n1097,
    n1131
  );


  xor
  g1601
  (
    n1728,
    n1086,
    n1028,
    n927,
    n718
  );


  xnor
  g1602
  (
    n1689,
    n1105,
    n1080,
    n1045,
    n1089
  );


  and
  g1603
  (
    n1748,
    n858,
    n1306,
    n1044,
    n1224
  );


  and
  g1604
  (
    n1474,
    n732,
    n983,
    n1164,
    n1217
  );


  and
  g1605
  (
    n1561,
    n816,
    n1051,
    n1196,
    n1249
  );


  xnor
  g1606
  (
    n1670,
    n1024,
    n1200,
    n1165,
    n1135
  );


  xor
  g1607
  (
    n1730,
    n909,
    n1109,
    n1167,
    n1037
  );


  xor
  g1608
  (
    n1617,
    n1302,
    n1046,
    n1124,
    n1294
  );


  or
  g1609
  (
    n1798,
    n1152,
    n1163,
    n1291,
    n687
  );


  or
  g1610
  (
    n1519,
    n1207,
    n1092,
    n1171,
    n1218
  );


  and
  g1611
  (
    n1786,
    n1243,
    n1078,
    n1271,
    n1109
  );


  and
  g1612
  (
    n1516,
    n1030,
    n1288,
    n1052,
    n705
  );


  nand
  g1613
  (
    n1635,
    n1170,
    n1058,
    n1060,
    n1072
  );


  and
  g1614
  (
    n1753,
    n1106,
    n1153,
    n1296,
    n720
  );


  xnor
  g1615
  (
    n1573,
    n937,
    n769,
    n1226,
    n1222
  );


  nand
  g1616
  (
    n1749,
    n736,
    n1298,
    n1066,
    n1085
  );


  nor
  g1617
  (
    n1638,
    n933,
    n1220,
    n1003,
    n1140
  );


  xnor
  g1618
  (
    n1601,
    n1244,
    n1134,
    n1291,
    n1175
  );


  xor
  g1619
  (
    n1810,
    n993,
    n1241,
    n1148,
    n1243
  );


  xnor
  g1620
  (
    n1637,
    n1056,
    n1047,
    n1219,
    n1210
  );


  and
  g1621
  (
    n1669,
    n832,
    n1215,
    n928,
    n1260
  );


  and
  g1622
  (
    n1776,
    n1144,
    n1281,
    n1258,
    n1097
  );


  xor
  g1623
  (
    n1607,
    n1167,
    n1110,
    n808,
    n1185
  );


  nand
  g1624
  (
    n1576,
    n1290,
    n1072,
    n692,
    n1255
  );


  or
  g1625
  (
    n1802,
    n1047,
    n1078,
    n1265,
    n1024
  );


  and
  g1626
  (
    n1674,
    n1192,
    n1031,
    n840,
    n1296
  );


  xnor
  g1627
  (
    n1470,
    n1145,
    n945,
    n740,
    n1079
  );


  or
  g1628
  (
    n1526,
    n923,
    n1122,
    n996,
    n862
  );


  nand
  g1629
  (
    n1457,
    n1256,
    n686,
    n1221,
    n794
  );


  and
  g1630
  (
    n1820,
    n915,
    n1128,
    n781,
    n1029
  );


  or
  g1631
  (
    n1581,
    n1065,
    n1152,
    n1105,
    n1063
  );


  xnor
  g1632
  (
    n1701,
    n1221,
    n969,
    n1216,
    n1305
  );


  or
  g1633
  (
    n1817,
    n1098,
    n875,
    n1253,
    n1276
  );


  xor
  g1634
  (
    n1572,
    n1287,
    n957,
    n1145,
    n1207
  );


  xor
  g1635
  (
    n1814,
    n1180,
    n779,
    n1077,
    n1282
  );


  nor
  g1636
  (
    n1788,
    n1128,
    n1148,
    n1043,
    n782
  );


  nor
  g1637
  (
    n1647,
    n1289,
    n1005,
    n1102,
    n1191
  );


  or
  g1638
  (
    n1652,
    n1115,
    n1246,
    n1055,
    n1174
  );


  nand
  g1639
  (
    n1787,
    n1126,
    n1120,
    n1186,
    n848
  );


  or
  g1640
  (
    n1704,
    n1075,
    n1014,
    n1035,
    n860
  );


  and
  g1641
  (
    n1589,
    n1242,
    n1233,
    n834,
    n894
  );


  and
  g1642
  (
    n1606,
    n1186,
    n1108,
    n1183,
    n1311
  );


  xnor
  g1643
  (
    n1815,
    n842,
    n1297,
    n1309,
    n837
  );


  and
  g1644
  (
    n1482,
    n777,
    n1306,
    n761,
    n1157
  );


  and
  g1645
  (
    n1712,
    n1212,
    n962,
    n1201,
    n1084
  );


  or
  g1646
  (
    n1809,
    n1088,
    n813,
    n1001,
    n1229
  );


  and
  g1647
  (
    n1812,
    n1053,
    n1261,
    n1052,
    n1211
  );


  or
  g1648
  (
    n1523,
    n1211,
    n1123,
    n1122,
    n1042
  );


  nand
  g1649
  (
    n1714,
    n943,
    n1090,
    n1175,
    n1242
  );


  nand
  g1650
  (
    n1679,
    n1013,
    n1260,
    n916,
    n1155
  );


  nor
  g1651
  (
    n1792,
    n1271,
    n1252,
    n1125,
    n1212
  );


  xor
  g1652
  (
    n1681,
    n1016,
    n961,
    n1272,
    n1043
  );


  nand
  g1653
  (
    n1766,
    n1011,
    n1307,
    n1099,
    n857
  );


  nand
  g1654
  (
    n1747,
    n1207,
    n744,
    n1163,
    n1278
  );


  nor
  g1655
  (
    n1806,
    n1248,
    n708,
    n1043,
    n1251
  );


  nor
  g1656
  (
    n1505,
    n1270,
    n1056,
    n1003,
    n1047
  );


  nand
  g1657
  (
    n1492,
    n1064,
    n1108,
    n1057,
    n885
  );


  xnor
  g1658
  (
    n1598,
    n1238,
    n1188,
    n748,
    n873
  );


  xor
  g1659
  (
    n1463,
    n1067,
    n1180,
    n1193,
    n1197
  );


  xor
  g1660
  (
    n1524,
    n1279,
    n1156,
    n959,
    n1187
  );


  xnor
  g1661
  (
    n1651,
    n676,
    n1230,
    n755,
    n1272
  );


  xor
  g1662
  (
    n1783,
    n1279,
    n1082,
    n1055,
    n981
  );


  and
  g1663
  (
    n1680,
    n767,
    n843,
    n1311,
    n1056
  );


  and
  g1664
  (
    n1720,
    n1105,
    n1079,
    n1301,
    n1150
  );


  nand
  g1665
  (
    n1781,
    n987,
    n1018,
    n1147,
    n1282
  );


  xnor
  g1666
  (
    n1538,
    n1136,
    n1032,
    n1249,
    n1189
  );


  nor
  g1667
  (
    n1517,
    n1215,
    n1100,
    n1092,
    n1263
  );


  and
  g1668
  (
    n1685,
    n999,
    n1201,
    n890,
    n1155
  );


  xnor
  g1669
  (
    n1800,
    n1135,
    n1254,
    n1305,
    n1095
  );


  nor
  g1670
  (
    n1610,
    n1162,
    n1114,
    n1058,
    n1184
  );


  and
  g1671
  (
    n1565,
    n888,
    n1160,
    n1293,
    n1203
  );


  xnor
  g1672
  (
    n1656,
    n765,
    n1253,
    n1299,
    n1283
  );


  or
  g1673
  (
    n1535,
    n724,
    n1194,
    n1118,
    n884
  );


  and
  g1674
  (
    n1642,
    n1286,
    n1238,
    n913,
    n1116
  );


  nor
  g1675
  (
    n1641,
    n1108,
    n1138,
    n1291,
    n1233
  );


  or
  g1676
  (
    n1536,
    n1132,
    n836,
    n1133,
    n1017
  );


  xnor
  g1677
  (
    n1542,
    n1202,
    n1070,
    n999,
    n1126
  );


  xnor
  g1678
  (
    n1456,
    n1237,
    n1227,
    n1278,
    n1154
  );


  xor
  g1679
  (
    n1791,
    n1138,
    n1033,
    n1248,
    n804
  );


  xnor
  g1680
  (
    n1595,
    n1065,
    n751,
    n1170,
    n1057
  );


  xnor
  g1681
  (
    n1762,
    n1267,
    n1147,
    n762,
    n1064
  );


  and
  g1682
  (
    n1507,
    n1224,
    n1092,
    n914,
    n1274
  );


  and
  g1683
  (
    n1631,
    n1125,
    n1254,
    n1294,
    n1008
  );


  xnor
  g1684
  (
    n1827,
    n1280,
    n1236,
    n797,
    n825
  );


  nor
  g1685
  (
    n1626,
    n707,
    n1072,
    n1249,
    n1099
  );


  nor
  g1686
  (
    n1478,
    n1101,
    n1005,
    n815,
    n1068
  );


  nor
  g1687
  (
    n1658,
    n1076,
    n975,
    n1041,
    n1269
  );


  nor
  g1688
  (
    n1794,
    n1221,
    n984,
    n1008,
    n1295
  );


  and
  g1689
  (
    n1549,
    n1012,
    n742,
    n750,
    n1153
  );


  and
  g1690
  (
    n1770,
    n783,
    n1171,
    n1130,
    n1064
  );


  xnor
  g1691
  (
    n1732,
    n1285,
    n1307,
    n780,
    n1251
  );


  or
  g1692
  (
    n1758,
    n1250,
    n1172,
    n1285,
    n1074
  );


  xnor
  g1693
  (
    n1750,
    n1062,
    n1244,
    n1146,
    n1058
  );


  and
  g1694
  (
    n1663,
    n1149,
    n1197,
    n1259,
    n1114
  );


  xor
  g1695
  (
    n1533,
    n1058,
    n948,
    n921,
    n1172
  );


  or
  g1696
  (
    n1717,
    n721,
    n1060,
    n775,
    n1026
  );


  nand
  g1697
  (
    n1811,
    n695,
    n911,
    n1311,
    n773
  );


  xor
  g1698
  (
    n1731,
    n696,
    n1118,
    n1217,
    n1236
  );


  nor
  g1699
  (
    n1816,
    n1051,
    n1194,
    n1178,
    n1208
  );


  or
  g1700
  (
    n1541,
    n1143,
    n1239,
    n1115,
    n1177
  );


  and
  g1701
  (
    n1522,
    n1067,
    n1287,
    n1309,
    n1093
  );


  xor
  g1702
  (
    n1779,
    n929,
    n1162,
    n1111,
    n970
  );


  and
  g1703
  (
    n1543,
    n1209,
    n1076,
    n1261,
    n1121
  );


  xnor
  g1704
  (
    n1585,
    n1099,
    n1276,
    n1277,
    n1299
  );


  or
  g1705
  (
    n1567,
    n1281,
    n1185,
    n1107,
    n1139
  );


  xnor
  g1706
  (
    n1699,
    n1114,
    n1039,
    n1117,
    n1091
  );


  xnor
  g1707
  (
    n1678,
    n1264,
    n1097,
    n1288,
    n807
  );


  and
  g1708
  (
    n1650,
    n785,
    n954,
    n1275,
    n1190
  );


  or
  g1709
  (
    n1488,
    n792,
    n1218,
    n1034,
    n1184
  );


  nor
  g1710
  (
    n1628,
    n1083,
    n1167,
    n997,
    n949
  );


  xnor
  g1711
  (
    n1460,
    n1116,
    n1192,
    n824,
    n938
  );


  nand
  g1712
  (
    n1514,
    n1188,
    n726,
    n1295,
    n1070
  );


  nor
  g1713
  (
    n1653,
    n1090,
    n1143,
    n1257,
    n1196
  );


  nor
  g1714
  (
    n1615,
    n1090,
    n1044,
    n1273,
    n1063
  );


  nand
  g1715
  (
    n1545,
    n1231,
    n682,
    n1158,
    n1021
  );


  nand
  g1716
  (
    n1722,
    n851,
    n1302,
    n1245,
    n1119
  );


  nor
  g1717
  (
    n1702,
    n723,
    n922,
    n1095,
    n1082
  );


  and
  g1718
  (
    n1693,
    n1165,
    n1216,
    n1271,
    n1294
  );


  xor
  g1719
  (
    n1660,
    n677,
    n1102,
    n1186,
    n839
  );


  or
  g1720
  (
    n1527,
    n1227,
    n1000,
    n881,
    n1083
  );


  or
  g1721
  (
    n1828,
    n1184,
    n1051,
    n1134,
    n1266
  );


  xnor
  g1722
  (
    n1824,
    n715,
    n1123,
    n1280,
    n1182
  );


  or
  g1723
  (
    n1757,
    n1074,
    n1164,
    n795,
    n977
  );


  xor
  g1724
  (
    n1803,
    n988,
    n1158,
    n1065,
    n1189
  );


  or
  g1725
  (
    n1706,
    n800,
    n1165,
    n1219,
    n908
  );


  nor
  g1726
  (
    n1640,
    n1264,
    n1303,
    n1150,
    n950
  );


  xor
  g1727
  (
    n1780,
    n1094,
    n1158,
    n838,
    n1191
  );


  and
  g1728
  (
    n1506,
    n1153,
    n1234,
    n872,
    n1050
  );


  or
  g1729
  (
    n1774,
    n1237,
    n1059,
    n741,
    n1219
  );


  nor
  g1730
  (
    n1547,
    n1031,
    n861,
    n1084,
    n1258
  );


  xnor
  g1731
  (
    n1745,
    n1127,
    n1278,
    n1243,
    n1291
  );


  or
  g1732
  (
    n1475,
    n1115,
    n1237,
    n951,
    n1211
  );


  xnor
  g1733
  (
    n1724,
    n1275,
    n1293,
    n1051,
    n1040
  );


  nor
  g1734
  (
    n1688,
    n770,
    n1146,
    n1292,
    n1177
  );


  nor
  g1735
  (
    n1577,
    n1245,
    n790,
    n1172,
    n1256
  );


  nor
  g1736
  (
    n1587,
    n1124,
    n1187,
    n821,
    n1199
  );


  and
  g1737
  (
    n1594,
    n1054,
    n1273,
    n1093,
    n1228
  );


  nand
  g1738
  (
    n1797,
    n1232,
    n891,
    n1298,
    n1110
  );


  nor
  g1739
  (
    n1560,
    n1198,
    n859,
    n1226,
    n1233
  );


  nor
  g1740
  (
    n1726,
    n1070,
    n1304,
    n1182,
    n1268
  );


  xnor
  g1741
  (
    n1659,
    n1101,
    n1163,
    n1171,
    n1115
  );


  nor
  g1742
  (
    n1676,
    n942,
    n974,
    n899,
    n863
  );


  xor
  g1743
  (
    n1737,
    n1293,
    n971,
    n847,
    n1214
  );


  nand
  g1744
  (
    n1665,
    n990,
    n1023,
    n1182,
    n749
  );


  nand
  g1745
  (
    n1769,
    n1299,
    n1077,
    n738,
    n1223
  );


  nor
  g1746
  (
    n1530,
    n681,
    n1235,
    n1231,
    n787
  );


  xnor
  g1747
  (
    n1529,
    n1273,
    n1203,
    n1199,
    n1062
  );


  or
  g1748
  (
    n1821,
    n1088,
    n1156,
    n956,
    n1113
  );


  xor
  g1749
  (
    n1707,
    n1184,
    n1173,
    n1282,
    n691
  );


  nor
  g1750
  (
    n1630,
    n699,
    n784,
    n895,
    n1173
  );


  nor
  g1751
  (
    n1644,
    n1197,
    n1059,
    n1137,
    n1271
  );


  or
  g1752
  (
    n1767,
    n1042,
    n892,
    n1180,
    n953
  );


  or
  g1753
  (
    n1819,
    n693,
    n900,
    n1243,
    n722
  );


  or
  g1754
  (
    n1479,
    n1199,
    n1130,
    n673,
    n1027
  );


  nand
  g1755
  (
    n1754,
    n1072,
    n818,
    n1119,
    n747
  );


  nand
  g1756
  (
    n1708,
    n1254,
    n1155,
    n1282,
    n704
  );


  or
  g1757
  (
    n1509,
    n1026,
    n844,
    n1247,
    n1242
  );


  nor
  g1758
  (
    n1525,
    n710,
    n1178,
    n1150,
    n1205
  );


  xor
  g1759
  (
    n1477,
    n1297,
    n1202,
    n1002,
    n939
  );


  xnor
  g1760
  (
    n1621,
    n1215,
    n1106,
    n1310,
    n1136
  );


  or
  g1761
  (
    n1481,
    n1204,
    n910,
    n1103,
    n846
  );


  or
  g1762
  (
    n1579,
    n1228,
    n1113,
    n1165,
    n1175
  );


  and
  g1763
  (
    n1605,
    n793,
    n706,
    n1144,
    n1028
  );


  xor
  g1764
  (
    n1459,
    n1065,
    n713,
    n1276,
    n1114
  );


  xor
  g1765
  (
    n1733,
    n1213,
    n1176,
    n1107,
    n1244
  );


  xor
  g1766
  (
    n1558,
    n1289,
    n1016,
    n1187,
    n1077
  );


  or
  g1767
  (
    n1593,
    n1179,
    n1277,
    n905,
    n1157
  );


  xor
  g1768
  (
    n1715,
    n737,
    n1304,
    n1144,
    n1142
  );


  xor
  g1769
  (
    n1559,
    n1015,
    n1310,
    n1173,
    n1247
  );


  nor
  g1770
  (
    n1503,
    n1230,
    n1217,
    n759,
    n1206
  );


  or
  g1771
  (
    n1721,
    n1162,
    n1267,
    n1125,
    n1173
  );


  nor
  g1772
  (
    n1464,
    n674,
    n979,
    n1302,
    n1151
  );


  xnor
  g1773
  (
    n1695,
    n897,
    n1142,
    n1253,
    n918
  );


  xnor
  g1774
  (
    n1490,
    n1189,
    n1303,
    n1048,
    n1064
  );


  xnor
  g1775
  (
    n1725,
    n1242,
    n1307,
    n1181,
    n1234
  );


  or
  g1776
  (
    n1657,
    n1257,
    n1112,
    n1228,
    n1073
  );


  and
  g1777
  (
    n1709,
    n1091,
    n819,
    n1007,
    n1089
  );


  or
  g1778
  (
    n1807,
    n1240,
    n1161,
    n1054,
    n1263
  );


  or
  g1779
  (
    n1677,
    n1061,
    n1096,
    n980,
    n1073
  );


  nand
  g1780
  (
    n1772,
    n1284,
    n907,
    n1190,
    n1152
  );


  nor
  g1781
  (
    n1633,
    n1157,
    n1293,
    n1253,
    n1156
  );


  nor
  g1782
  (
    n1654,
    n1145,
    n1266,
    n1201,
    n1284
  );


  or
  g1783
  (
    n1775,
    n849,
    n1286,
    n1191,
    n1118
  );


  nor
  g1784
  (
    n1608,
    n756,
    n1300,
    n788,
    n1139
  );


  nand
  g1785
  (
    n1801,
    n1223,
    n1202,
    n1014,
    n919
  );


  xor
  g1786
  (
    n1574,
    n1264,
    n1111,
    n1237,
    n973
  );


  xor
  g1787
  (
    n1484,
    n1128,
    n1246,
    n1240,
    n1144
  );


  or
  g1788
  (
    n1623,
    n1141,
    n1209,
    n1044,
    n1137
  );


  or
  g1789
  (
    n1739,
    n931,
    n1068,
    n1110,
    n1265
  );


  xnor
  g1790
  (
    n1532,
    n1274,
    n1142,
    n1166,
    n1245
  );


  xor
  g1791
  (
    n1495,
    n768,
    n1076,
    n1232,
    n1100
  );


  or
  g1792
  (
    n1778,
    n1250,
    n1223,
    n1126,
    n1151
  );


  nand
  g1793
  (
    n1735,
    n1132,
    n1234,
    n754,
    n963
  );


  nand
  g1794
  (
    n1499,
    n757,
    n1239,
    n992,
    n1096
  );


  xor
  g1795
  (
    n1672,
    n1268,
    n1140,
    n1185,
    n871
  );


  or
  g1796
  (
    n1831,
    n1481,
    n1456,
    n1464,
    n1513
  );


  nor
  g1797
  (
    n1844,
    n1502,
    n1465,
    n1463,
    n1477
  );


  and
  g1798
  (
    n1840,
    n1526,
    n1462,
    n1493,
    n1519
  );


  and
  g1799
  (
    n1843,
    n1486,
    n1479,
    n1527,
    n1499
  );


  nor
  g1800
  (
    n1839,
    n1483,
    n1488,
    n1517,
    n1498
  );


  nand
  g1801
  (
    n1830,
    n1470,
    n1492,
    n1478,
    n1487
  );


  xor
  g1802
  (
    n1838,
    n1500,
    n1522,
    n1518,
    n1459
  );


  xnor
  g1803
  (
    n1833,
    n1495,
    n1521,
    n1480,
    n1476
  );


  nor
  g1804
  (
    n1834,
    n1503,
    n1523,
    n1515,
    n1510
  );


  or
  g1805
  (
    n1846,
    n1472,
    n1496,
    n1511,
    n1512
  );


  nand
  g1806
  (
    n1835,
    n1507,
    n1473,
    n1460,
    n1467
  );


  or
  g1807
  (
    n1832,
    n1497,
    n1525,
    n1506,
    n1491
  );


  nand
  g1808
  (
    n1829,
    n1469,
    n1514,
    n1457,
    n1461
  );


  xor
  g1809
  (
    n1845,
    n1505,
    n1482,
    n1485,
    n1494
  );


  xnor
  g1810
  (
    n1842,
    n1504,
    n1484,
    n1509,
    n1489
  );


  or
  g1811
  (
    n1836,
    n1508,
    n1475,
    n1471,
    n1524
  );


  nor
  g1812
  (
    n1841,
    n1490,
    n1501,
    n1516,
    n1520
  );


  and
  g1813
  (
    n1837,
    n1458,
    n1474,
    n1468,
    n1466
  );


  buf
  g1814
  (
    n1849,
    n1844
  );


  not
  g1815
  (
    n1848,
    n1843
  );


  buf
  g1816
  (
    n1847,
    n1845
  );


  nand
  g1817
  (
    n1855,
    n575,
    n575,
    n571,
    n573
  );


  xnor
  g1818
  (
    n1853,
    n575,
    n1847
  );


  nor
  g1819
  (
    n1852,
    n573,
    n1848,
    n571,
    n1849
  );


  or
  g1820
  (
    n1858,
    n572,
    n576,
    n574
  );


  xor
  g1821
  (
    n1850,
    n1848,
    n576,
    n1849
  );


  nand
  g1822
  (
    n1857,
    n577,
    n573,
    n576,
    n578
  );


  nand
  g1823
  (
    n1859,
    n577,
    n571,
    n576
  );


  or
  g1824
  (
    n1854,
    n575,
    n572,
    n570
  );


  nand
  g1825
  (
    n1851,
    n577,
    n572,
    n1849,
    n1848
  );


  xnor
  g1826
  (
    n1856,
    n573,
    n577,
    n574
  );


  not
  g1827
  (
    n1862,
    n1312
  );


  buf
  g1828
  (
    n1860,
    n1851
  );


  not
  g1829
  (
    n1863,
    n1853
  );


  nand
  g1830
  (
    n1861,
    n1852,
    n1312
  );


  xor
  g1831
  (
    n1864,
    n1850,
    n1312,
    n1854
  );


  buf
  g1832
  (
    n1865,
    n1860
  );


  or
  g1833
  (
    n1869,
    n1315,
    n1313
  );


  and
  g1834
  (
    n1866,
    n1865,
    n1315,
    n1314
  );


  and
  g1835
  (
    n1867,
    n1865,
    n1314
  );


  and
  g1836
  (
    n1868,
    n1865,
    n1313,
    n1315
  );


  or
  g1837
  (
    n1870,
    n1529,
    n1530,
    n1528,
    n1868
  );


  buf
  g1838
  (
    n1872,
    n1870
  );


  not
  g1839
  (
    n1871,
    n1870
  );


  xnor
  g1840
  (
    n1874,
    n579,
    n1871,
    n580,
    n581
  );


  or
  g1841
  (
    n1879,
    n581,
    n582,
    n579
  );


  nand
  g1842
  (
    n1880,
    n583,
    n579,
    n1871,
    n582
  );


  xor
  g1843
  (
    n1877,
    n1871,
    n581,
    n1872,
    n583
  );


  or
  g1844
  (
    n1875,
    n578,
    n1872
  );


  nor
  g1845
  (
    n1876,
    n580,
    n582,
    n583
  );


  and
  g1846
  (
    n1873,
    n580,
    n578,
    n579,
    n584
  );


  nor
  g1847
  (
    n1878,
    n578,
    n580,
    n581,
    n1871
  );


  xnor
  g1848
  (
    n1881,
    n1876,
    n1318,
    n1316
  );


  nor
  g1849
  (
    n1882,
    n1874,
    n1320,
    n1319
  );


  nand
  g1850
  (
    n1885,
    n1318,
    n1316
  );


  and
  g1851
  (
    n1884,
    n1317,
    n1319,
    n1873,
    n1875
  );


  or
  g1852
  (
    n1886,
    n1319,
    n1878,
    n1317
  );


  and
  g1853
  (
    n1883,
    n1877,
    n1316,
    n1320,
    n1317
  );


  or
  g1854
  (
    n1889,
    n1536,
    n1533,
    n1539,
    n1535
  );


  or
  g1855
  (
    n1890,
    n1534,
    n1884,
    n1537,
    n1532
  );


  or
  g1856
  (
    n1888,
    n1881,
    n1540,
    n1542,
    n1538
  );


  xnor
  g1857
  (
    n1887,
    n1541,
    n1882,
    n1531,
    n1883
  );


  not
  g1858
  (
    n1893,
    n1888
  );


  buf
  g1859
  (
    n1894,
    n1889
  );


  buf
  g1860
  (
    n1898,
    n1889
  );


  buf
  g1861
  (
    n1896,
    n1887
  );


  buf
  g1862
  (
    n1897,
    n1890
  );


  buf
  g1863
  (
    n1895,
    n1543
  );


  buf
  g1864
  (
    n1891,
    n1890
  );


  or
  g1865
  (
    n1892,
    n1889,
    n1890,
    n1846
  );


  not
  g1866
  (
    n1901,
    n1891
  );


  not
  g1867
  (
    n1899,
    n1891
  );


  buf
  g1868
  (
    n1900,
    n1891
  );


  not
  g1869
  (
    n1902,
    n1892
  );


  buf
  g1870
  (
    n1909,
    n1900
  );


  not
  g1871
  (
    n1908,
    n1899
  );


  not
  g1872
  (
    n1910,
    n1901
  );


  not
  g1873
  (
    n1911,
    n1900
  );


  buf
  g1874
  (
    n1912,
    n1899
  );


  buf
  g1875
  (
    n1904,
    n1900
  );


  buf
  g1876
  (
    n1907,
    n1900
  );


  not
  g1877
  (
    n1906,
    n1901
  );


  buf
  g1878
  (
    n1903,
    n1899
  );


  not
  g1879
  (
    n1905,
    n1899
  );


  buf
  g1880
  (
    n1931,
    n1910
  );


  buf
  g1881
  (
    n1921,
    n1908
  );


  not
  g1882
  (
    n1938,
    n1909
  );


  buf
  g1883
  (
    n1913,
    n1906
  );


  buf
  g1884
  (
    n1930,
    n1908
  );


  not
  g1885
  (
    n1915,
    n1910
  );


  not
  g1886
  (
    n1920,
    n1910
  );


  not
  g1887
  (
    n1927,
    n1907
  );


  buf
  g1888
  (
    n1939,
    n1905
  );


  buf
  g1889
  (
    n1933,
    n1908
  );


  buf
  g1890
  (
    n1937,
    n1904
  );


  not
  g1891
  (
    n1924,
    n1904
  );


  buf
  g1892
  (
    n1934,
    n1909
  );


  not
  g1893
  (
    n1926,
    n1903
  );


  not
  g1894
  (
    n1917,
    n1906
  );


  buf
  g1895
  (
    n1932,
    n1907
  );


  buf
  g1896
  (
    n1928,
    n1904
  );


  buf
  g1897
  (
    n1944,
    n1904
  );


  buf
  g1898
  (
    n1918,
    n1909
  );


  not
  g1899
  (
    n1925,
    n1910
  );


  not
  g1900
  (
    n1919,
    n1905
  );


  not
  g1901
  (
    n1929,
    n1908
  );


  not
  g1902
  (
    n1936,
    n1907
  );


  buf
  g1903
  (
    n1935,
    n1905
  );


  not
  g1904
  (
    n1943,
    n1906
  );


  not
  g1905
  (
    n1941,
    n1903
  );


  not
  g1906
  (
    n1942,
    n1903
  );


  not
  g1907
  (
    n1916,
    n1909
  );


  buf
  g1908
  (
    n1923,
    n1903
  );


  buf
  g1909
  (
    n1940,
    n1905
  );


  not
  g1910
  (
    n1914,
    n1906
  );


  buf
  g1911
  (
    n1922,
    n1907
  );


  xnor
  g1912
  (
    n2006,
    n1595,
    n1943,
    n1599
  );


  nor
  g1913
  (
    n2032,
    n1698,
    n1563,
    n1940
  );


  xor
  g1914
  (
    n1997,
    n1570,
    n1864,
    n1944
  );


  or
  g1915
  (
    n2030,
    n1800,
    n1714,
    n1324
  );


  or
  g1916
  (
    n1945,
    n1778,
    n1940,
    n1937
  );


  xor
  g1917
  (
    n2027,
    n1929,
    n1600,
    n1928
  );


  nor
  g1918
  (
    n1960,
    n1717,
    n1721,
    n1547
  );


  nor
  g1919
  (
    n1995,
    n1933,
    n1786,
    n1742
  );


  xnor
  g1920
  (
    n1987,
    n1793,
    n1747,
    n1933
  );


  nand
  g1921
  (
    n2047,
    n1649,
    n1914,
    n1779
  );


  xnor
  g1922
  (
    n1974,
    n1918,
    n1709,
    n584
  );


  or
  g1923
  (
    n1975,
    n1325,
    n1612,
    n1680
  );


  and
  g1924
  (
    n2041,
    n1713,
    n1770,
    n1691
  );


  nor
  g1925
  (
    n1999,
    n1806,
    n1648,
    n1798
  );


  xor
  g1926
  (
    n2038,
    n1663,
    n1555,
    n1936
  );


  xor
  g1927
  (
    KeyWire_0_9,
    n1864,
    n584,
    n1584
  );


  or
  g1928
  (
    n1958,
    n1619,
    n1930,
    n1936
  );


  nor
  g1929
  (
    n2010,
    n1753,
    n1692,
    n1926
  );


  or
  g1930
  (
    n1982,
    n1723,
    n1931,
    n1935
  );


  nand
  g1931
  (
    n2005,
    n1607,
    n1322,
    n1735
  );


  xor
  g1932
  (
    n2066,
    n1924,
    n1758,
    n1637
  );


  nand
  g1933
  (
    n1986,
    n1771,
    n1681,
    n586
  );


  or
  g1934
  (
    n2034,
    n1931,
    n1938,
    n1792
  );


  nor
  g1935
  (
    n2043,
    n1575,
    n1922,
    n1919
  );


  xor
  g1936
  (
    n2029,
    n1939,
    n1630,
    n1716
  );


  xor
  g1937
  (
    n2042,
    n1775,
    n1554,
    n1917
  );


  xnor
  g1938
  (
    n1947,
    n1659,
    n1914,
    n1743
  );


  nor
  g1939
  (
    n1959,
    n1578,
    n1810,
    n1777
  );


  and
  g1940
  (
    n2053,
    n1928,
    n1924,
    n1785
  );


  xor
  g1941
  (
    n2001,
    n1918,
    n1320,
    n1923
  );


  xnor
  g1942
  (
    n1985,
    n1622,
    n1605,
    n1802
  );


  and
  g1943
  (
    n1971,
    n1935,
    n1568,
    n1751
  );


  nor
  g1944
  (
    n2011,
    n1321,
    n1926,
    n1572
  );


  nand
  g1945
  (
    n2060,
    n1323,
    n1737,
    n1664
  );


  nor
  g1946
  (
    n2046,
    n1789,
    n1860,
    n1934
  );


  xnor
  g1947
  (
    n2002,
    n1682,
    n1734,
    n1585
  );


  xnor
  g1948
  (
    n2065,
    n1557,
    n1638,
    n1641
  );


  or
  g1949
  (
    n2048,
    n1624,
    n1918,
    n1941
  );


  nor
  g1950
  (
    n2003,
    n1566,
    n1803,
    n1586
  );


  xnor
  g1951
  (
    n2063,
    n1929,
    n1863,
    n1614
  );


  xor
  g1952
  (
    n1957,
    n1725,
    n1610,
    n1322
  );


  or
  g1953
  (
    n1994,
    n1632,
    n585,
    n1577
  );


  xnor
  g1954
  (
    n2068,
    n1732,
    n1921,
    n1658
  );


  or
  g1955
  (
    n2023,
    n1929,
    n1784,
    n1943
  );


  and
  g1956
  (
    n2051,
    n1923,
    n1915,
    n1927
  );


  xnor
  g1957
  (
    n2031,
    n1643,
    n1712,
    n1808
  );


  xnor
  g1958
  (
    n2013,
    n1931,
    n1756,
    n1932
  );


  or
  g1959
  (
    n1980,
    n1863,
    n1677,
    n1799
  );


  nand
  g1960
  (
    n2017,
    n1769,
    n1601,
    n1938
  );


  and
  g1961
  (
    n2040,
    n1809,
    n1918,
    n1683
  );


  nand
  g1962
  (
    n2057,
    n1938,
    n1930,
    n1913
  );


  nand
  g1963
  (
    n1993,
    n1767,
    n1937,
    n1327
  );


  nand
  g1964
  (
    n1984,
    n1939,
    n1944,
    n1774
  );


  nand
  g1965
  (
    n2033,
    n1323,
    n1917,
    n1724
  );


  or
  g1966
  (
    n1953,
    n1764,
    n1588,
    n1760
  );


  xnor
  g1967
  (
    n1981,
    n1679,
    n1629,
    n1943
  );


  xor
  g1968
  (
    n1962,
    n1564,
    n1860,
    n1687
  );


  nand
  g1969
  (
    n1964,
    n1720,
    n1551,
    n1780
  );


  xor
  g1970
  (
    n2059,
    n1589,
    n1695,
    n1730
  );


  xnor
  g1971
  (
    n1948,
    n1604,
    n1927,
    n1916
  );


  xnor
  g1972
  (
    n1963,
    n1791,
    n1736,
    n1662
  );


  or
  g1973
  (
    n2028,
    n1913,
    n1321,
    n1917
  );


  and
  g1974
  (
    n2070,
    n1699,
    n1921,
    n1688
  );


  nand
  g1975
  (
    n2045,
    n1703,
    n1652,
    n1707,
    n1548
  );


  and
  g1976
  (
    n2008,
    n1773,
    n1561,
    n1602,
    n1558
  );


  nor
  g1977
  (
    n2020,
    n1861,
    n1796,
    n1696,
    n1934
  );


  or
  g1978
  (
    n1967,
    n1651,
    n1863,
    n1325,
    n1794
  );


  xor
  g1979
  (
    n1989,
    n1657,
    n1940,
    n1569,
    n1325
  );


  nand
  g1980
  (
    n2064,
    n1766,
    n1623,
    n1722,
    n1655
  );


  nor
  g1981
  (
    n1990,
    n1581,
    n1921,
    n1801,
    n1693
  );


  nand
  g1982
  (
    n1946,
    n1861,
    n585,
    n1740,
    n1749
  );


  nand
  g1983
  (
    n1992,
    n1923,
    n1697,
    n1625,
    n1782
  );


  or
  g1984
  (
    n1949,
    n1689,
    n1705,
    n1861,
    n1567
  );


  xnor
  g1985
  (
    n2019,
    n1661,
    n1924,
    n1320,
    n1583
  );


  xor
  g1986
  (
    n1956,
    n1938,
    n1762,
    n1748,
    n1606
  );


  or
  g1987
  (
    n1961,
    n1765,
    n1653,
    n1931,
    n1744
  );


  nor
  g1988
  (
    n1998,
    n1615,
    n585,
    n1731,
    n1324
  );


  xnor
  g1989
  (
    n2022,
    n1710,
    n1711,
    n1942
  );


  xnor
  g1990
  (
    n2025,
    n1934,
    n1862,
    n1939,
    n1666
  );


  xor
  g1991
  (
    n1983,
    n1805,
    n1923,
    n1728,
    n1613
  );


  and
  g1992
  (
    n2009,
    n1862,
    n1660,
    n1326,
    n1807
  );


  or
  g1993
  (
    n1951,
    n1565,
    n1919,
    n1694,
    n1933
  );


  xnor
  g1994
  (
    n2015,
    n1916,
    n1700,
    n1592,
    n1635
  );


  xnor
  g1995
  (
    n2061,
    n1325,
    n1627,
    n1914,
    n1915
  );


  xnor
  g1996
  (
    n2007,
    n1591,
    n1864,
    n1783,
    n1776
  );


  nand
  g1997
  (
    n2049,
    n1560,
    n1644,
    n1579,
    n1940
  );


  or
  g1998
  (
    n1952,
    n1324,
    n1795,
    n1628,
    n1936
  );


  or
  g1999
  (
    n2021,
    n1676,
    n1944,
    n1935,
    n1757
  );


  or
  g2000
  (
    n2012,
    n1690,
    n1929,
    n1754,
    n1544
  );


  nor
  g2001
  (
    n2072,
    n1925,
    n1633,
    n1675,
    n1686
  );


  and
  g2002
  (
    n1988,
    n1322,
    n1597,
    n1708,
    n1603
  );


  and
  g2003
  (
    n1950,
    n1667,
    n1671,
    n586,
    n1553
  );


  and
  g2004
  (
    n1972,
    n1943,
    n1930,
    n1768,
    n1741
  );


  xor
  g2005
  (
    n1973,
    n1919,
    n1718,
    n1932,
    n1552
  );


  xor
  g2006
  (
    n2062,
    n1941,
    n1922,
    n1913,
    n1862
  );


  xnor
  g2007
  (
    n2000,
    n1590,
    n1608,
    n1704,
    n1587
  );


  xnor
  g2008
  (
    n2024,
    n1788,
    n1321,
    n1787,
    n1670
  );


  or
  g2009
  (
    n2058,
    n1656,
    n1915,
    n1642,
    n1942
  );


  or
  g2010
  (
    n2044,
    n1739,
    n1936,
    n1634,
    n1729
  );


  nor
  g2011
  (
    n2016,
    n584,
    n1727,
    n1752,
    n1559
  );


  xor
  g2012
  (
    n1996,
    n1925,
    n1862,
    n1546,
    n1920
  );


  or
  g2013
  (
    n2050,
    n1755,
    n1935,
    n1631,
    n1326
  );


  nand
  g2014
  (
    n2069,
    n585,
    n1647,
    n1750,
    n1594
  );


  nor
  g2015
  (
    n2036,
    n1738,
    n1763,
    n1869,
    n1678
  );


  nand
  g2016
  (
    n1977,
    n1915,
    n1930,
    n1611,
    n1942
  );


  or
  g2017
  (
    n1976,
    n1562,
    n1937,
    n1927,
    n1733
  );


  xor
  g2018
  (
    n1979,
    n1715,
    n1616,
    n1934,
    n1321
  );


  xnor
  g2019
  (
    n1955,
    n1326,
    n1618,
    n1323,
    n1927
  );


  or
  g2020
  (
    n1970,
    n1545,
    n1933,
    n1719,
    n1609
  );


  nor
  g2021
  (
    n2035,
    n1916,
    n1582,
    n1672,
    n1549
  );


  nor
  g2022
  (
    n2014,
    n1922,
    n1645,
    n1925,
    n1550
  );


  or
  g2023
  (
    n2067,
    n1684,
    n1668,
    n1790,
    n1673
  );


  nand
  g2024
  (
    n1968,
    n1924,
    n1639,
    n1928,
    n1617
  );


  nand
  g2025
  (
    n2026,
    n1804,
    n1925,
    n1941,
    n1571
  );


  and
  g2026
  (
    n1965,
    n1621,
    n1654,
    n1797,
    n1916
  );


  xnor
  g2027
  (
    n1966,
    n1702,
    n1646,
    n1920,
    n1939
  );


  or
  g2028
  (
    n2056,
    n1922,
    n1598,
    n1926,
    n1928
  );


  xnor
  g2029
  (
    n2054,
    n1920,
    n1650,
    n1759,
    n1932
  );


  xor
  g2030
  (
    n1978,
    n1913,
    n1573,
    n1640,
    n1937
  );


  or
  g2031
  (
    n1969,
    n1920,
    n1669,
    n1745,
    n1580
  );


  and
  g2032
  (
    n1954,
    n1636,
    n1944,
    n1665,
    n1917
  );


  nor
  g2033
  (
    n2055,
    n1701,
    n1781,
    n1746,
    n1921
  );


  nor
  g2034
  (
    n2039,
    n1726,
    n1685,
    n1326,
    n1863
  );


  or
  g2035
  (
    n1991,
    n1706,
    n1761,
    n1626,
    n1574
  );


  nand
  g2036
  (
    n2018,
    n1576,
    n1914,
    n1941,
    n1926
  );


  or
  g2037
  (
    n2037,
    n1919,
    n1556,
    n1596,
    n1323
  );


  nand
  g2038
  (
    n2052,
    n1932,
    n1772,
    n1324,
    n1593
  );


  or
  g2039
  (
    n2071,
    n1811,
    n1674,
    n1322,
    n1620
  );


  buf
  g2040
  (
    n2075,
    n1947
  );


  buf
  g2041
  (
    n2078,
    n1947
  );


  buf
  g2042
  (
    n2079,
    n1946
  );


  not
  g2043
  (
    n2086,
    n1946
  );


  not
  g2044
  (
    n2080,
    n1948
  );


  buf
  g2045
  (
    n2083,
    n1945
  );


  not
  g2046
  (
    n2074,
    n1945
  );


  not
  g2047
  (
    n2073,
    n1946
  );


  buf
  g2048
  (
    n2077,
    n1948
  );


  not
  g2049
  (
    n2084,
    n1948
  );


  buf
  g2050
  (
    n2085,
    n1947
  );


  not
  g2051
  (
    n2081,
    n1947
  );


  buf
  g2052
  (
    n2088,
    n1948
  );


  buf
  g2053
  (
    n2087,
    n1945
  );


  buf
  g2054
  (
    n2082,
    n1946
  );


  buf
  g2055
  (
    n2076,
    n1945
  );


  not
  g2056
  (
    n2092,
    n2075
  );


  not
  g2057
  (
    n2108,
    n2079
  );


  not
  g2058
  (
    n2096,
    n2078
  );


  buf
  g2059
  (
    n2109,
    n2073
  );


  not
  g2060
  (
    n2114,
    n2073
  );


  not
  g2061
  (
    n2099,
    n2080
  );


  not
  g2062
  (
    n2095,
    n2073
  );


  not
  g2063
  (
    n2104,
    n2076
  );


  not
  g2064
  (
    n2103,
    n2077
  );


  not
  g2065
  (
    n2117,
    n2076
  );


  buf
  g2066
  (
    n2116,
    n2078
  );


  not
  g2067
  (
    n2101,
    n2076
  );


  not
  g2068
  (
    n2113,
    n2079
  );


  buf
  g2069
  (
    n2089,
    n2074
  );


  not
  g2070
  (
    n2111,
    n2074
  );


  not
  g2071
  (
    n2102,
    n2077
  );


  buf
  g2072
  (
    KeyWire_0_15,
    n2077
  );


  not
  g2073
  (
    n2112,
    n2075
  );


  not
  g2074
  (
    n2093,
    n2073
  );


  not
  g2075
  (
    n2100,
    n2080
  );


  buf
  g2076
  (
    n2094,
    n2077
  );


  not
  g2077
  (
    n2098,
    n2079
  );


  buf
  g2078
  (
    n2118,
    n2075
  );


  not
  g2079
  (
    n2091,
    n2076
  );


  not
  g2080
  (
    n2105,
    n2079
  );


  buf
  g2081
  (
    n2090,
    n2078
  );


  buf
  g2082
  (
    n2110,
    n2075
  );


  not
  g2083
  (
    n2107,
    n2078
  );


  buf
  g2084
  (
    n2115,
    n2074
  );


  buf
  g2085
  (
    n2097,
    n2074
  );


  not
  g2086
  (
    n2122,
    n1348
  );


  buf
  g2087
  (
    n2164,
    n2109
  );


  buf
  g2088
  (
    n2149,
    n1858
  );


  buf
  g2089
  (
    n2219,
    n1334
  );


  not
  g2090
  (
    n2236,
    n1346
  );


  buf
  g2091
  (
    n2157,
    n2111
  );


  buf
  g2092
  (
    n2142,
    n1812
  );


  buf
  g2093
  (
    n2233,
    n1813
  );


  buf
  g2094
  (
    n2174,
    n1332
  );


  buf
  g2095
  (
    n2146,
    n1949
  );


  not
  g2096
  (
    n2159,
    n2114
  );


  buf
  g2097
  (
    n2185,
    n2106
  );


  not
  g2098
  (
    n2193,
    n2115
  );


  buf
  g2099
  (
    n2161,
    n2094
  );


  buf
  g2100
  (
    n2134,
    n2116
  );


  not
  g2101
  (
    n2204,
    n2118
  );


  not
  g2102
  (
    n2133,
    n2108
  );


  not
  g2103
  (
    n2148,
    n1856
  );


  buf
  g2104
  (
    n2163,
    n1827
  );


  not
  g2105
  (
    n2129,
    n2098
  );


  buf
  g2106
  (
    n2184,
    n1333
  );


  buf
  g2107
  (
    n2169,
    n2103
  );


  not
  g2108
  (
    n2173,
    n1332
  );


  not
  g2109
  (
    n2198,
    n1815
  );


  not
  g2110
  (
    n2192,
    n2095
  );


  buf
  g2111
  (
    n2183,
    n1335
  );


  not
  g2112
  (
    n2124,
    n1347
  );


  not
  g2113
  (
    n2227,
    n2091
  );


  buf
  g2114
  (
    n2152,
    n2094
  );


  not
  g2115
  (
    n2225,
    n2101
  );


  not
  g2116
  (
    n2143,
    n1331
  );


  buf
  g2117
  (
    n2162,
    n1341
  );


  buf
  g2118
  (
    n2190,
    n2106
  );


  not
  g2119
  (
    n2232,
    n2101
  );


  not
  g2120
  (
    n2207,
    n2092
  );


  buf
  g2121
  (
    n2121,
    n2099
  );


  not
  g2122
  (
    n2166,
    n1349
  );


  not
  g2123
  (
    n2195,
    n2099
  );


  not
  g2124
  (
    n2135,
    n1338
  );


  not
  g2125
  (
    n2139,
    n2100
  );


  buf
  g2126
  (
    n2217,
    n1327
  );


  not
  g2127
  (
    n2226,
    n1347
  );


  not
  g2128
  (
    n2201,
    n2101
  );


  not
  g2129
  (
    n2186,
    n2093
  );


  buf
  g2130
  (
    n2130,
    n2111
  );


  not
  g2131
  (
    n2213,
    n1329
  );


  buf
  g2132
  (
    n2200,
    n2115
  );


  buf
  g2133
  (
    n2228,
    n1327
  );


  not
  g2134
  (
    n2177,
    n1338
  );


  not
  g2135
  (
    n2223,
    n2101
  );


  not
  g2136
  (
    n2231,
    n1327
  );


  buf
  g2137
  (
    n2238,
    n2102
  );


  buf
  g2138
  (
    n2120,
    n1822
  );


  buf
  g2139
  (
    n2176,
    n2110
  );


  not
  g2140
  (
    n2153,
    n1333
  );


  buf
  g2141
  (
    n2214,
    n2113
  );


  buf
  g2142
  (
    n2119,
    n2112
  );


  not
  g2143
  (
    n2189,
    n2117
  );


  buf
  g2144
  (
    n2222,
    n1346
  );


  not
  g2145
  (
    n2125,
    n1339
  );


  buf
  g2146
  (
    n2132,
    n2115
  );


  not
  g2147
  (
    n2151,
    n1344
  );


  not
  g2148
  (
    n2137,
    n1330
  );


  not
  g2149
  (
    n2203,
    n1329
  );


  buf
  g2150
  (
    n2179,
    n1329
  );


  not
  g2151
  (
    n2224,
    n1816
  );


  buf
  g2152
  (
    n2175,
    n1341
  );


  buf
  g2153
  (
    n2235,
    n1340
  );


  buf
  g2154
  (
    n2220,
    n1350
  );


  buf
  g2155
  (
    n2215,
    n1818
  );


  buf
  g2156
  (
    n2178,
    n2110
  );


  buf
  g2157
  (
    n2155,
    n1855
  );


  not
  g2158
  (
    n2216,
    n1826
  );


  not
  g2159
  (
    n2229,
    n2097
  );


  buf
  g2160
  (
    n2123,
    n1343
  );


  buf
  g2161
  (
    n2156,
    n2099
  );


  not
  g2162
  (
    n2188,
    n2114
  );


  buf
  g2163
  (
    n2210,
    n1339
  );


  not
  g2164
  (
    n2230,
    n2117
  );


  not
  g2165
  (
    n2167,
    n1336
  );


  buf
  g2166
  (
    n2165,
    n1348
  );


  nand
  g2167
  (
    n2206,
    n1825,
    n1336,
    n2116,
    n1348
  );


  nand
  g2168
  (
    n2202,
    n2113,
    n1817,
    n2097,
    n1335
  );


  or
  g2169
  (
    n2194,
    n1328,
    n2102,
    n1346,
    n2104
  );


  xor
  g2170
  (
    n2208,
    n1349,
    n2096,
    n1345,
    n1344
  );


  xor
  g2171
  (
    n2145,
    n2111,
    n1819,
    n1341,
    n2100
  );


  nand
  g2172
  (
    n2172,
    n1335,
    n2118,
    n2092,
    n2115
  );


  or
  g2173
  (
    n2171,
    n1334,
    n2114,
    n2107,
    n2089
  );


  nor
  g2174
  (
    KeyWire_0_3,
    n1334,
    n1348,
    n2112,
    n2114
  );


  xnor
  g2175
  (
    n2211,
    n2118,
    n2091,
    n1334,
    n2102
  );


  or
  g2176
  (
    n2237,
    n2110,
    n1345,
    n1344,
    n2090
  );


  xor
  g2177
  (
    n2144,
    n1328,
    n1864,
    n2091,
    n2112
  );


  xnor
  g2178
  (
    n2147,
    n1347,
    n2110,
    n2095,
    n1345
  );


  nand
  g2179
  (
    n2199,
    n1343,
    n2100,
    n1336,
    n2106
  );


  and
  g2180
  (
    n2136,
    n1338,
    n1340,
    n2118,
    n2113
  );


  xnor
  g2181
  (
    n2154,
    n1337,
    n1341,
    n2107,
    n2095
  );


  nand
  g2182
  (
    n2205,
    n1330,
    n2105,
    n2089,
    n1338
  );


  or
  g2183
  (
    n2140,
    n2117,
    n2098,
    n2093,
    n2108
  );


  nand
  g2184
  (
    n2181,
    n2104,
    n1332,
    n2105,
    n1337
  );


  nand
  g2185
  (
    n2170,
    n2090,
    n1337,
    n2095,
    n1340
  );


  xor
  g2186
  (
    n2187,
    n2103,
    n2097,
    n2093,
    n1342
  );


  xnor
  g2187
  (
    n2196,
    n1331,
    n1337,
    n2099,
    n2109
  );


  and
  g2188
  (
    n2126,
    n1824,
    n2117,
    n1330,
    n1342
  );


  or
  g2189
  (
    n2158,
    n2090,
    n1823,
    n1342,
    n1349
  );


  and
  g2190
  (
    n2127,
    n2090,
    n2098,
    n2107,
    n1331
  );


  xor
  g2191
  (
    n2150,
    n2091,
    n2092,
    n2103,
    n1814
  );


  and
  g2192
  (
    n2131,
    n1347,
    n2096,
    n1340,
    n1828
  );


  nor
  g2193
  (
    n2182,
    n1344,
    n2089,
    n1335,
    n2104
  );


  xnor
  g2194
  (
    n2221,
    n2111,
    n1820,
    n1857,
    n1330
  );


  xnor
  g2195
  (
    n2197,
    n2092,
    n1331,
    n2094,
    n2112
  );


  xnor
  g2196
  (
    n2212,
    n1859,
    n2116,
    n2109,
    n2105
  );


  nand
  g2197
  (
    n2209,
    n1329,
    n2094,
    n1349,
    n1343
  );


  or
  g2198
  (
    n2168,
    n1333,
    n1345,
    n1332,
    n2097
  );


  xnor
  g2199
  (
    n2180,
    n1821,
    n2089,
    n1339,
    n2103
  );


  nand
  g2200
  (
    n2128,
    n1336,
    n2093,
    n2102,
    n1333
  );


  nor
  g2201
  (
    n2141,
    n2113,
    n1339,
    n2106,
    n1343
  );


  xnor
  g2202
  (
    n2218,
    n2105,
    n1328,
    n2108,
    n2096
  );


  xnor
  g2203
  (
    n2191,
    n2108,
    n1342,
    n2100,
    n2080
  );


  nand
  g2204
  (
    n2234,
    n2104,
    n2107,
    n2098,
    n2116
  );


  or
  g2205
  (
    n2160,
    n1328,
    n1346,
    n2109,
    n2096
  );


  not
  g2206
  (
    n2601,
    n1952
  );


  not
  g2207
  (
    n2298,
    n2043
  );


  buf
  g2208
  (
    n2455,
    n2005
  );


  buf
  g2209
  (
    n2550,
    n2084
  );


  not
  g2210
  (
    n2549,
    n596
  );


  not
  g2211
  (
    n2371,
    n652
  );


  not
  g2212
  (
    n2573,
    n2009
  );


  not
  g2213
  (
    n2566,
    n666
  );


  buf
  g2214
  (
    n2400,
    n1975
  );


  not
  g2215
  (
    n2249,
    n2220
  );


  not
  g2216
  (
    n2410,
    n596
  );


  not
  g2217
  (
    n2284,
    n1957
  );


  not
  g2218
  (
    n2470,
    n669
  );


  buf
  g2219
  (
    n2457,
    n647
  );


  not
  g2220
  (
    n2534,
    n2127
  );


  buf
  g2221
  (
    n2345,
    n667
  );


  not
  g2222
  (
    n2598,
    n1949
  );


  buf
  g2223
  (
    n2610,
    n1994
  );


  buf
  g2224
  (
    n2522,
    n2022
  );


  not
  g2225
  (
    n2579,
    n2130
  );


  not
  g2226
  (
    n2502,
    n617
  );


  not
  g2227
  (
    n2423,
    n2043
  );


  buf
  g2228
  (
    n2537,
    n1978
  );


  buf
  g2229
  (
    n2270,
    n2063
  );


  buf
  g2230
  (
    n2321,
    n2063
  );


  buf
  g2231
  (
    n2446,
    n1985
  );


  not
  g2232
  (
    n2367,
    n2017
  );


  buf
  g2233
  (
    n2278,
    n2197
  );


  buf
  g2234
  (
    n2543,
    n658
  );


  not
  g2235
  (
    n2370,
    n2162
  );


  not
  g2236
  (
    n2616,
    n2135
  );


  not
  g2237
  (
    n2487,
    n2131
  );


  not
  g2238
  (
    n2529,
    n2129
  );


  buf
  g2239
  (
    n2327,
    n1953
  );


  buf
  g2240
  (
    n2299,
    n2027
  );


  buf
  g2241
  (
    n2331,
    n645
  );


  buf
  g2242
  (
    n2514,
    n2124
  );


  buf
  g2243
  (
    n2356,
    n2017
  );


  buf
  g2244
  (
    n2464,
    n2061
  );


  buf
  g2245
  (
    n2336,
    n2231
  );


  not
  g2246
  (
    n2448,
    n2067
  );


  buf
  g2247
  (
    n2332,
    n1970
  );


  buf
  g2248
  (
    n2561,
    n650
  );


  not
  g2249
  (
    n2435,
    n2132
  );


  not
  g2250
  (
    n2396,
    n2206
  );


  not
  g2251
  (
    n2281,
    n631
  );


  buf
  g2252
  (
    n2294,
    n2146
  );


  buf
  g2253
  (
    n2468,
    n2190
  );


  buf
  g2254
  (
    n2243,
    n2129
  );


  not
  g2255
  (
    n2337,
    n2016
  );


  buf
  g2256
  (
    n2307,
    n2145
  );


  not
  g2257
  (
    n2443,
    n2221
  );


  buf
  g2258
  (
    n2256,
    n2185
  );


  buf
  g2259
  (
    n2578,
    n650
  );


  not
  g2260
  (
    n2295,
    n2222
  );


  not
  g2261
  (
    n2260,
    n1993
  );


  nor
  g2262
  (
    n2300,
    n2083,
    n2140,
    n612,
    n2188
  );


  or
  g2263
  (
    n2605,
    n600,
    n2163,
    n2173,
    n2154
  );


  or
  g2264
  (
    n2389,
    n2064,
    n2139,
    n2132,
    n2004
  );


  xnor
  g2265
  (
    n2449,
    n635,
    n2208,
    n2155,
    n2031
  );


  xnor
  g2266
  (
    n2528,
    n2156,
    n2030,
    n668,
    n2131
  );


  and
  g2267
  (
    n2374,
    n2010,
    n2161,
    n2048,
    n2151
  );


  xor
  g2268
  (
    n2597,
    n2122,
    n1985,
    n1972,
    n635
  );


  or
  g2269
  (
    n2413,
    n2152,
    n2014,
    n1951,
    n2009
  );


  nand
  g2270
  (
    n2556,
    n1965,
    n2214,
    n2082,
    n2050
  );


  and
  g2271
  (
    n2612,
    n2124,
    n599,
    n601,
    n2055
  );


  or
  g2272
  (
    n2335,
    n2136,
    n626,
    n2199,
    n1958
  );


  nor
  g2273
  (
    n2465,
    n623,
    n2161,
    n624,
    n2037
  );


  or
  g2274
  (
    n2290,
    n592,
    n2181,
    n2054,
    n2174
  );


  xor
  g2275
  (
    n2359,
    n2002,
    n598,
    n2126,
    n2231
  );


  and
  g2276
  (
    n2478,
    n591,
    n1996,
    n603,
    n2193
  );


  xnor
  g2277
  (
    n2599,
    n2147,
    n2165,
    n2151,
    n603
  );


  and
  g2278
  (
    n2461,
    n2148,
    n2209,
    n631,
    n1999
  );


  or
  g2279
  (
    n2607,
    n629,
    n1969,
    n2139,
    n2212
  );


  nor
  g2280
  (
    n2267,
    n2180,
    n2141,
    n1987,
    n668
  );


  nor
  g2281
  (
    n2554,
    n2150,
    n2217,
    n2051
  );


  or
  g2282
  (
    n2254,
    n2055,
    n1961,
    n2086,
    n2020
  );


  nor
  g2283
  (
    n2242,
    n2207,
    n2222,
    n2150,
    n632
  );


  or
  g2284
  (
    n2386,
    n2167,
    n2187,
    n2224,
    n1969
  );


  nand
  g2285
  (
    n2262,
    n2003,
    n657,
    n2231,
    n1977
  );


  nand
  g2286
  (
    n2585,
    n2047,
    n650,
    n2029,
    n622
  );


  xor
  g2287
  (
    n2593,
    n2068,
    n2175,
    n590,
    n622
  );


  xnor
  g2288
  (
    n2521,
    n645,
    n618,
    n2120,
    n1955
  );


  and
  g2289
  (
    n2445,
    n2051,
    n1972,
    n642,
    n2027
  );


  nand
  g2290
  (
    n2481,
    n2199,
    n2127,
    n2201,
    n610
  );


  and
  g2291
  (
    n2407,
    n2138,
    n2181,
    n671,
    n2018
  );


  nand
  g2292
  (
    n2434,
    n2130,
    n2225,
    n2173,
    n1959
  );


  nor
  g2293
  (
    n2474,
    n1977,
    n2085,
    n622,
    n2032
  );


  and
  g2294
  (
    n2546,
    n613,
    n633,
    n1974,
    n2213
  );


  nand
  g2295
  (
    n2248,
    n657,
    n2203,
    n2214,
    n2012
  );


  and
  g2296
  (
    n2308,
    n2223,
    n2173,
    n643,
    n599
  );


  xnor
  g2297
  (
    n2325,
    n2065,
    n2211,
    n2143,
    n2149
  );


  and
  g2298
  (
    n2568,
    n599,
    n636,
    n2043,
    n1992
  );


  xor
  g2299
  (
    n2313,
    n1985,
    n593,
    n1960,
    n611
  );


  nand
  g2300
  (
    n2343,
    n2123,
    n2171,
    n1956,
    n1989
  );


  and
  g2301
  (
    n2338,
    n2205,
    n2200,
    n2161,
    n1979
  );


  xor
  g2302
  (
    n2426,
    n2153,
    n602,
    n2135,
    n2032
  );


  xor
  g2303
  (
    n2419,
    n2210,
    n2208,
    n609,
    n2212
  );


  xnor
  g2304
  (
    n2286,
    n2207,
    n2194,
    n2036,
    n636
  );


  xor
  g2305
  (
    n2437,
    n2222,
    n2052,
    n2000,
    n615
  );


  and
  g2306
  (
    n2586,
    n604,
    n2149,
    n2003,
    n1988
  );


  xor
  g2307
  (
    n2490,
    n2197,
    n2158,
    n640,
    n2050
  );


  xor
  g2308
  (
    n2259,
    n2158,
    n2206,
    n618,
    n2085
  );


  nand
  g2309
  (
    n2329,
    n2156,
    n2122,
    n2057,
    n2087
  );


  nand
  g2310
  (
    n2440,
    n2035,
    n2232,
    n660,
    n2179
  );


  nor
  g2311
  (
    n2408,
    n2159,
    n640,
    n657,
    n2060
  );


  or
  g2312
  (
    n2289,
    n1879,
    n1971,
    n2082,
    n1880
  );


  and
  g2313
  (
    n2314,
    n1963,
    n604,
    n1990,
    n2003
  );


  xor
  g2314
  (
    n2342,
    n2151,
    n2162,
    n2229,
    n1969
  );


  and
  g2315
  (
    n2240,
    n659,
    n2009,
    n1975,
    n641
  );


  and
  g2316
  (
    n2392,
    n2227,
    n2067,
    n2023,
    n648
  );


  nand
  g2317
  (
    n2344,
    n2035,
    n651,
    n2024,
    n2048
  );


  xnor
  g2318
  (
    n2297,
    n1974,
    n2221,
    n2125,
    n627
  );


  nor
  g2319
  (
    n2312,
    n1879,
    n653,
    n632,
    n2083
  );


  and
  g2320
  (
    n2526,
    n1999,
    n592,
    n2170,
    n2123
  );


  xor
  g2321
  (
    n2358,
    n2051,
    n2040,
    n2020,
    n2201
  );


  xnor
  g2322
  (
    n2296,
    n2126,
    n1991,
    n628,
    n2004
  );


  and
  g2323
  (
    n2536,
    n638,
    n2219,
    n2152,
    n610
  );


  and
  g2324
  (
    n2339,
    n2008,
    n2229,
    n614,
    n2178
  );


  or
  g2325
  (
    n2424,
    n2233,
    n2164,
    n2191,
    n1952
  );


  and
  g2326
  (
    n2603,
    n651,
    n1991,
    n2006,
    n2032
  );


  nor
  g2327
  (
    n2504,
    n2177,
    n654,
    n2146,
    n1960
  );


  xor
  g2328
  (
    n2614,
    n2210,
    n664,
    n2038,
    n643
  );


  and
  g2329
  (
    n2495,
    n2191,
    n2194,
    n2230,
    n590
  );


  and
  g2330
  (
    n2466,
    n2033,
    n2007,
    n2164,
    n2176
  );


  and
  g2331
  (
    n2430,
    n1953,
    n2157,
    n1964,
    n607
  );


  xor
  g2332
  (
    n2282,
    n1980,
    n597,
    n1976,
    n2064
  );


  and
  g2333
  (
    n2483,
    n1350,
    n650,
    n611,
    n2180
  );


  xnor
  g2334
  (
    n2600,
    n2037,
    n2050,
    n1982,
    n1989
  );


  or
  g2335
  (
    n2571,
    n2010,
    n625,
    n609,
    n669
  );


  nor
  g2336
  (
    n2456,
    n1964,
    n2202,
    n2199,
    n2149
  );


  xnor
  g2337
  (
    n2606,
    n2211,
    n2063,
    n616,
    n2042
  );


  and
  g2338
  (
    n2244,
    n2038,
    n1976,
    n2041,
    n1351
  );


  nor
  g2339
  (
    n2401,
    n2184,
    n637,
    n2030,
    n667
  );


  nor
  g2340
  (
    n2469,
    n2142,
    n1955,
    n2192,
    n648
  );


  nand
  g2341
  (
    n2569,
    n2063,
    n2037,
    n1966,
    n2158
  );


  nand
  g2342
  (
    n2372,
    n2199,
    n1987,
    n2142,
    n1954
  );


  or
  g2343
  (
    n2283,
    n2213,
    n2235,
    n2171,
    n1968
  );


  and
  g2344
  (
    n2247,
    n2227,
    n667,
    n2042,
    n1998
  );


  or
  g2345
  (
    n2444,
    n2143,
    n2176,
    n608,
    n2155
  );


  nand
  g2346
  (
    n2503,
    n660,
    n607,
    n663,
    n619
  );


  and
  g2347
  (
    n2263,
    n591,
    n2166,
    n2219,
    n1999
  );


  or
  g2348
  (
    n2275,
    n666,
    n1950,
    n1987,
    n2059
  );


  nand
  g2349
  (
    n2428,
    n2219,
    n2152,
    n2146,
    n2065
  );


  and
  g2350
  (
    n2375,
    n586,
    n2234,
    n1949,
    n2024
  );


  or
  g2351
  (
    n2274,
    n1993,
    n2119,
    n1997,
    n2040
  );


  nand
  g2352
  (
    n2398,
    n2000,
    n2133,
    n1978,
    n2233
  );


  xnor
  g2353
  (
    n2508,
    n640,
    n1998,
    n2224,
    n2015
  );


  xnor
  g2354
  (
    n2551,
    n2068,
    n2088,
    n646,
    n2229
  );


  and
  g2355
  (
    n2391,
    n612,
    n2038,
    n2085,
    n2169
  );


  nor
  g2356
  (
    n2513,
    n2087,
    n2131,
    n2210,
    n2157
  );


  or
  g2357
  (
    n2330,
    n2120,
    n2125,
    n2182,
    n648
  );


  or
  g2358
  (
    n2277,
    n2225,
    n2046,
    n641,
    n598
  );


  nand
  g2359
  (
    n2500,
    n2014,
    n589,
    n591,
    n1989
  );


  or
  g2360
  (
    n2480,
    n644,
    n2165,
    n2059,
    n1880
  );


  xor
  g2361
  (
    n2378,
    n2046,
    n1951,
    n587,
    n2198
  );


  xnor
  g2362
  (
    n2390,
    n2049,
    n1995,
    n588,
    n2216
  );


  xnor
  g2363
  (
    n2559,
    n2031,
    n2082,
    n2189,
    n2149
  );


  and
  g2364
  (
    n2509,
    n2182,
    n1973,
    n597,
    n2119
  );


  xnor
  g2365
  (
    n2454,
    n2159,
    n2126,
    n2137,
    n647
  );


  nor
  g2366
  (
    n2575,
    n2168,
    n2030,
    n2213,
    n665
  );


  nand
  g2367
  (
    n2310,
    n2224,
    n2041,
    n2186,
    n2167
  );


  xnor
  g2368
  (
    n2591,
    n617,
    n1973,
    n1994,
    n621
  );


  nand
  g2369
  (
    n2420,
    n2203,
    n1965,
    n2019,
    n2029
  );


  xnor
  g2370
  (
    n2531,
    n662,
    n1997,
    n610,
    n2227
  );


  nand
  g2371
  (
    n2590,
    n594,
    n2047,
    n2136,
    n2172
  );


  xor
  g2372
  (
    n2524,
    n2195,
    n2012,
    n2161,
    n2197
  );


  xnor
  g2373
  (
    n2475,
    n588,
    n651,
    n661,
    n2235
  );


  or
  g2374
  (
    n2304,
    n1988,
    n2184,
    n623,
    n661
  );


  nand
  g2375
  (
    n2280,
    n2230,
    n2138,
    n2168,
    n634
  );


  nor
  g2376
  (
    n2518,
    n2025,
    n1999,
    n605,
    n2160
  );


  nor
  g2377
  (
    n2511,
    n2175,
    n2142,
    n2224,
    n662
  );


  xor
  g2378
  (
    n2562,
    n614,
    n1954,
    n1979,
    n2154
  );


  xor
  g2379
  (
    n2293,
    n2155,
    n2186,
    n2020,
    n2041
  );


  nor
  g2380
  (
    n2517,
    n663,
    n1957,
    n613,
    n2206
  );


  xnor
  g2381
  (
    n2496,
    n1983,
    n2028,
    n595,
    n2015
  );


  xor
  g2382
  (
    n2364,
    n2029,
    n2197,
    n2140,
    n656
  );


  and
  g2383
  (
    n2403,
    n1971,
    n1962,
    n1979,
    n635
  );


  xor
  g2384
  (
    n2324,
    n2171,
    n607,
    n649,
    n1981
  );


  xor
  g2385
  (
    n2276,
    n1995,
    n2140,
    n1961,
    n2009
  );


  or
  g2386
  (
    n2552,
    n611,
    n619,
    n628,
    n2213
  );


  nor
  g2387
  (
    n2576,
    n607,
    n2054,
    n2012,
    n2209
  );


  xor
  g2388
  (
    n2425,
    n1981,
    n2060,
    n601,
    n592
  );


  xor
  g2389
  (
    n2501,
    n644,
    n2233,
    n635,
    n2058
  );


  nor
  g2390
  (
    n2602,
    n1986,
    n2121,
    n2024,
    n2037
  );


  or
  g2391
  (
    n2587,
    n1967,
    n2140,
    n2232,
    n2062
  );


  or
  g2392
  (
    n2458,
    n2200,
    n2179,
    n1978,
    n2182
  );


  or
  g2393
  (
    n2473,
    n1878,
    n1950,
    n1965,
    n2189
  );


  or
  g2394
  (
    n2472,
    n2218,
    n2188,
    n630,
    n649
  );


  xor
  g2395
  (
    n2318,
    n2084,
    n662,
    n2024,
    n2228
  );


  xnor
  g2396
  (
    n2442,
    n2012,
    n2026,
    n2022,
    n609
  );


  xor
  g2397
  (
    n2380,
    n620,
    n2204,
    n1968,
    n663
  );


  nor
  g2398
  (
    n2432,
    n2230,
    n630,
    n2234,
    n1962
  );


  and
  g2399
  (
    n2545,
    n2162,
    n1985,
    n2014,
    n2221
  );


  nand
  g2400
  (
    n2351,
    n2200,
    n2016,
    n2046,
    n619
  );


  or
  g2401
  (
    n2476,
    n2128,
    n599,
    n2144,
    n2029
  );


  nand
  g2402
  (
    n2608,
    n2017,
    n2055,
    n594,
    n2023
  );


  xnor
  g2403
  (
    n2451,
    n2172,
    n2121,
    n2205,
    n656
  );


  nor
  g2404
  (
    n2394,
    n2201,
    n2217,
    n2087,
    n2145
  );


  nor
  g2405
  (
    n2431,
    n2129,
    n2015,
    n2027,
    n1954
  );


  nand
  g2406
  (
    n2258,
    n2141,
    n1967,
    n2144,
    n2039
  );


  xor
  g2407
  (
    n2405,
    n2163,
    n2160,
    n1989,
    n1976
  );


  xnor
  g2408
  (
    n2592,
    n1970,
    n2021,
    n2051,
    n2058
  );


  and
  g2409
  (
    n2581,
    n2136,
    n2205,
    n2150,
    n616
  );


  nand
  g2410
  (
    n2497,
    n2220,
    n2163,
    n2013,
    n594
  );


  or
  g2411
  (
    n2346,
    n593,
    n1992,
    n2057,
    n2221
  );


  xnor
  g2412
  (
    n2527,
    n2148,
    n2226,
    n633,
    n637
  );


  or
  g2413
  (
    n2273,
    n1951,
    n2026,
    n2021,
    n2086
  );


  and
  g2414
  (
    n2540,
    n642,
    n2204,
    n2231,
    n2081
  );


  xnor
  g2415
  (
    n2309,
    n587,
    n2068,
    n2008,
    n634
  );


  and
  g2416
  (
    n2357,
    n2178,
    n2030,
    n2173,
    n2185
  );


  and
  g2417
  (
    n2557,
    n2069,
    n2196,
    n2068,
    n1996
  );


  nor
  g2418
  (
    n2530,
    n2191,
    n2223,
    n2083,
    n1980
  );


  and
  g2419
  (
    n2565,
    n2121,
    n639,
    n2061,
    n2232
  );


  and
  g2420
  (
    n2311,
    n646,
    n2025,
    n2160,
    n2036
  );


  xor
  g2421
  (
    n2572,
    n1998,
    n629,
    n2180,
    n637
  );


  xnor
  g2422
  (
    n2538,
    n601,
    n2081,
    n2045,
    n588
  );


  and
  g2423
  (
    n2411,
    n1975,
    n1954,
    n2137,
    n2040
  );


  xor
  g2424
  (
    n2609,
    n2223,
    n631,
    n2062,
    n2011
  );


  and
  g2425
  (
    n2305,
    n2202,
    n1994,
    n2192,
    n1960
  );


  and
  g2426
  (
    n2422,
    n670,
    n654,
    n2054,
    n623
  );


  nand
  g2427
  (
    n2441,
    n2187,
    n666,
    n644,
    n2169
  );


  and
  g2428
  (
    n2547,
    n2081,
    n2216,
    n2055,
    n1964
  );


  nand
  g2429
  (
    n2488,
    n2060,
    n2004,
    n2136,
    n643
  );


  xnor
  g2430
  (
    n2373,
    n1953,
    n2045,
    n600,
    n1964
  );


  xnor
  g2431
  (
    n2381,
    n2011,
    n2052,
    n1350,
    n2219
  );


  xor
  g2432
  (
    n2253,
    n2058,
    n2167,
    n669,
    n1993
  );


  nor
  g2433
  (
    n2594,
    n2206,
    n659,
    n2122,
    n637
  );


  and
  g2434
  (
    n2489,
    n2170,
    n2028,
    n2008,
    n2122
  );


  xnor
  g2435
  (
    n2515,
    n2201,
    n2124,
    n1994,
    n2016
  );


  nor
  g2436
  (
    n2560,
    n2204,
    n2202,
    n2141,
    n2134
  );


  or
  g2437
  (
    n2414,
    n2017,
    n2066,
    n602,
    n2083
  );


  or
  g2438
  (
    n2264,
    n1963,
    n2194,
    n2048,
    n2059
  );


  xor
  g2439
  (
    n2302,
    n587,
    n2134,
    n2195,
    n2192
  );


  and
  g2440
  (
    n2417,
    n2165,
    n592,
    n653,
    n2172
  );


  or
  g2441
  (
    n2519,
    n2190,
    n2176,
    n1978,
    n2142
  );


  nor
  g2442
  (
    n2499,
    n2125,
    n2148,
    n2181,
    n2207
  );


  xor
  g2443
  (
    n2584,
    n2021,
    n2002,
    n1879,
    n2044
  );


  or
  g2444
  (
    n2418,
    n1955,
    n1983,
    n2031,
    n2157
  );


  nor
  g2445
  (
    n2412,
    n2132,
    n2005,
    n2168,
    n1878
  );


  xor
  g2446
  (
    n2317,
    n2042,
    n2057,
    n2234,
    n606
  );


  xnor
  g2447
  (
    n2341,
    n1982,
    n1950,
    n669,
    n617
  );


  nand
  g2448
  (
    n2319,
    n638,
    n2025,
    n606,
    n2189
  );


  or
  g2449
  (
    n2382,
    n2034,
    n631,
    n655,
    n660
  );


  nand
  g2450
  (
    n2520,
    n593,
    n642,
    n2088,
    n2139
  );


  nand
  g2451
  (
    n2363,
    n2194,
    n2053,
    n2159,
    n626
  );


  xor
  g2452
  (
    n2246,
    n608,
    n1986,
    n627,
    n657
  );


  and
  g2453
  (
    n2485,
    n2177,
    n664,
    n2033,
    n2195
  );


  xor
  g2454
  (
    n2506,
    n2000,
    n595,
    n656,
    n2156
  );


  nor
  g2455
  (
    n2388,
    n2209,
    n655,
    n2036,
    n2013
  );


  nand
  g2456
  (
    n2429,
    n594,
    n2163,
    n639,
    n2196
  );


  nor
  g2457
  (
    n2368,
    n2067,
    n2156,
    n1955,
    n2178
  );


  nor
  g2458
  (
    n2493,
    n2175,
    n2204,
    n608,
    n659
  );


  nor
  g2459
  (
    n2596,
    n2016,
    n2133,
    n2044,
    n2159
  );


  and
  g2460
  (
    n2399,
    n589,
    n2025,
    n2137,
    n2184
  );


  xnor
  g2461
  (
    n2553,
    n2044,
    n2234,
    n1971,
    n1988
  );


  xor
  g2462
  (
    n2523,
    n664,
    n1966,
    n2128,
    n2069
  );


  nand
  g2463
  (
    n2482,
    n2035,
    n2215,
    n2200,
    n2046
  );


  nor
  g2464
  (
    n2484,
    n654,
    n668,
    n2137,
    n1972
  );


  and
  g2465
  (
    n2334,
    n2154,
    n615,
    n2225,
    n2147
  );


  xnor
  g2466
  (
    n2404,
    n1968,
    n652,
    n671,
    n2082
  );


  or
  g2467
  (
    n2257,
    n2220,
    n2171,
    n2048,
    n2157
  );


  or
  g2468
  (
    n2326,
    n2170,
    n618,
    n2052,
    n2139
  );


  xnor
  g2469
  (
    n2548,
    n2177,
    n2162,
    n656,
    n2028
  );


  xnor
  g2470
  (
    n2416,
    n2147,
    n2223,
    n2208,
    n2119
  );


  xnor
  g2471
  (
    n2486,
    n1351,
    n1980,
    n623,
    n1959
  );


  xnor
  g2472
  (
    n2510,
    n626,
    n2166,
    n587,
    n621
  );


  or
  g2473
  (
    n2383,
    n612,
    n589,
    n643,
    n2210
  );


  nand
  g2474
  (
    n2409,
    n2138,
    n2198,
    n2034,
    n586
  );


  nand
  g2475
  (
    n2265,
    n2215,
    n647,
    n1984,
    n2062
  );


  nand
  g2476
  (
    n2369,
    n2135,
    n2047,
    n2121,
    n645
  );


  xor
  g2477
  (
    n2491,
    n2128,
    n667,
    n2067,
    n2179
  );


  nor
  g2478
  (
    n2479,
    n663,
    n2002,
    n1961,
    n1984
  );


  xor
  g2479
  (
    n2555,
    n2143,
    n1974,
    n632,
    n2188
  );


  or
  g2480
  (
    n2362,
    n1970,
    n603,
    n2229,
    n1951
  );


  nand
  g2481
  (
    n2376,
    n2123,
    n2165,
    n2228,
    n2064
  );


  or
  g2482
  (
    n2245,
    n621,
    n2144,
    n2155,
    n2177
  );


  nor
  g2483
  (
    n2406,
    n2007,
    n2033,
    n670,
    n2196
  );


  nor
  g2484
  (
    n2463,
    n1984,
    n2023,
    n2195,
    n664
  );


  xnor
  g2485
  (
    n2462,
    n1979,
    n2039,
    n615,
    n2026
  );


  xor
  g2486
  (
    n2415,
    n1976,
    n1990,
    n2185,
    n597
  );


  nor
  g2487
  (
    n2507,
    n2129,
    n606,
    n2036,
    n2010
  );


  nor
  g2488
  (
    n2361,
    n2125,
    n621,
    n2087,
    n660
  );


  nand
  g2489
  (
    n2349,
    n2023,
    n608,
    n2066,
    n2169
  );


  xor
  g2490
  (
    n2558,
    n645,
    n609,
    n2027,
    n2003
  );


  and
  g2491
  (
    n2533,
    n2226,
    n595,
    n1880,
    n2054
  );


  and
  g2492
  (
    n2563,
    n1990,
    n618,
    n2081,
    n1986
  );


  and
  g2493
  (
    n2241,
    n2203,
    n2128,
    n598,
    n2022
  );


  or
  g2494
  (
    n2255,
    n2232,
    n2052,
    n602,
    n2178
  );


  and
  g2495
  (
    n2516,
    n1879,
    n2119,
    n1991,
    n1973
  );


  or
  g2496
  (
    n2393,
    n2154,
    n2146,
    n2225,
    n1960
  );


  xor
  g2497
  (
    n2301,
    n665,
    n661,
    n2174,
    n2183
  );


  xor
  g2498
  (
    n2542,
    n596,
    n2228,
    n670,
    n633
  );


  and
  g2499
  (
    n2285,
    n2187,
    n2193,
    n2214,
    n622
  );


  xor
  g2500
  (
    n2397,
    n2222,
    n2209,
    n2132,
    n2179
  );


  or
  g2501
  (
    n2272,
    n2011,
    n2064,
    n597,
    n2032
  );


  or
  g2502
  (
    n2452,
    n641,
    n2191,
    n603,
    n2193
  );


  xnor
  g2503
  (
    n2604,
    n2035,
    n2186,
    n628,
    n601
  );


  nor
  g2504
  (
    n2567,
    n2062,
    n2022,
    n1987,
    n615
  );


  xor
  g2505
  (
    n2268,
    n1352,
    n641,
    n2175,
    n2039
  );


  xnor
  g2506
  (
    n2271,
    n1984,
    n1995,
    n1982,
    n636
  );


  xnor
  g2507
  (
    n2589,
    n625,
    n606,
    n596,
    n642
  );


  xnor
  g2508
  (
    n2365,
    n590,
    n2141,
    n1983,
    n613
  );


  xnor
  g2509
  (
    n2251,
    n2170,
    n1958,
    n624,
    n2226
  );


  nand
  g2510
  (
    n2316,
    n2145,
    n2230,
    n2026,
    n613
  );


  nor
  g2511
  (
    n2328,
    n2019,
    n1969,
    n2020,
    n617
  );


  nand
  g2512
  (
    n2377,
    n1959,
    n616,
    n654,
    n2031
  );


  and
  g2513
  (
    n2544,
    n1968,
    n2007,
    n2164,
    n2034
  );


  or
  g2514
  (
    n2494,
    n2053,
    n2152,
    n1967,
    n2001
  );


  xor
  g2515
  (
    n2291,
    n1351,
    n2181,
    n2217,
    n2056
  );


  nor
  g2516
  (
    n2347,
    n2059,
    n2047,
    n2144,
    n2045
  );


  xnor
  g2517
  (
    n2615,
    n1949,
    n646,
    n1966,
    n2211
  );


  and
  g2518
  (
    n2570,
    n602,
    n633,
    n1996,
    n2188
  );


  and
  g2519
  (
    n2577,
    n2127,
    n593,
    n2190,
    n2005
  );


  xor
  g2520
  (
    n2323,
    n611,
    n1992,
    n1352,
    n2034
  );


  nor
  g2521
  (
    n2261,
    n1950,
    n1962,
    n2061,
    n589
  );


  or
  g2522
  (
    n2535,
    n619,
    n2057,
    n1970,
    n2056
  );


  xor
  g2523
  (
    KeyWire_0_5,
    n2066,
    n2124,
    n639,
    n2043
  );


  and
  g2524
  (
    n2395,
    n588,
    n2056,
    n1958,
    n2018
  );


  nand
  g2525
  (
    n2315,
    n2205,
    n2151,
    n2214,
    n2187
  );


  and
  g2526
  (
    n2427,
    n2218,
    n1352,
    n2053,
    n2021
  );


  xor
  g2527
  (
    n2402,
    n2131,
    n634,
    n2084,
    n2007
  );


  and
  g2528
  (
    n2505,
    n2014,
    n2180,
    n2123,
    n2065
  );


  xor
  g2529
  (
    n2580,
    n2018,
    n1350,
    n2120,
    n638
  );


  xor
  g2530
  (
    n2453,
    n620,
    n1957,
    n2049,
    n2174
  );


  or
  g2531
  (
    n2574,
    n2153,
    n2019,
    n1973,
    n2198
  );


  or
  g2532
  (
    n2303,
    n1972,
    n2000,
    n2186,
    n616
  );


  or
  g2533
  (
    n2471,
    n591,
    n1977,
    n2228,
    n2189
  );


  and
  g2534
  (
    n2352,
    n2227,
    n2183,
    n2084
  );


  or
  g2535
  (
    n2340,
    n2166,
    n1880,
    n1980,
    n1974
  );


  xnor
  g2536
  (
    n2541,
    n2167,
    n640,
    n610,
    n2008
  );


  nor
  g2537
  (
    n2525,
    n2182,
    n628,
    n2039,
    n620
  );


  nor
  g2538
  (
    n2583,
    n2183,
    n2001,
    n2019
  );


  xor
  g2539
  (
    n2582,
    n2065,
    n2086,
    n655,
    n2005
  );


  xnor
  g2540
  (
    n2492,
    n2134,
    n2015,
    n1997,
    n2001
  );


  nor
  g2541
  (
    n2354,
    n2135,
    n632,
    n2066,
    n604
  );


  xor
  g2542
  (
    n2279,
    n625,
    n658,
    n1986,
    n2088
  );


  nor
  g2543
  (
    n2512,
    n2049,
    n2006,
    n624,
    n1966
  );


  and
  g2544
  (
    n2460,
    n2233,
    n1995,
    n2045,
    n2058
  );


  xor
  g2545
  (
    n2287,
    n1963,
    n2050,
    n2053,
    n1982
  );


  nand
  g2546
  (
    n2360,
    n1993,
    n1959,
    n2198,
    n1990
  );


  and
  g2547
  (
    n2387,
    n1971,
    n1962,
    n2193,
    n595
  );


  xnor
  g2548
  (
    n2459,
    n612,
    n2218,
    n2127,
    n627
  );


  nor
  g2549
  (
    n2477,
    n624,
    n1981,
    n2011,
    n646
  );


  or
  g2550
  (
    n2348,
    n2060,
    n2148,
    n671
  );


  xor
  g2551
  (
    n2250,
    n600,
    n2138,
    n2147,
    n1952
  );


  nor
  g2552
  (
    n2333,
    n1988,
    n1956,
    n2044,
    n614
  );


  nand
  g2553
  (
    n2421,
    n600,
    n2207,
    n648,
    n630
  );


  or
  g2554
  (
    n2498,
    n653,
    n1963,
    n620,
    n2185
  );


  nor
  g2555
  (
    n2355,
    n2133,
    n2216,
    n653,
    n644
  );


  xnor
  g2556
  (
    n2439,
    n659,
    n1952,
    n665,
    n2042
  );


  nand
  g2557
  (
    n2239,
    n2013,
    n2216,
    n1983,
    n2158
  );


  nand
  g2558
  (
    n2532,
    n634,
    n2010,
    n590,
    n2226
  );


  nand
  g2559
  (
    n2433,
    n647,
    n2086,
    n1953,
    n2153
  );


  or
  g2560
  (
    n2611,
    n1961,
    n2169,
    n658,
    n1956
  );


  or
  g2561
  (
    n2322,
    n2013,
    n2033,
    n2080,
    n2150
  );


  and
  g2562
  (
    n2564,
    n1992,
    n1957,
    n2211,
    n2028
  );


  nand
  g2563
  (
    n2320,
    n2049,
    n1956,
    n2041,
    n2153
  );


  xor
  g2564
  (
    n2269,
    n605,
    n630,
    n668,
    n2220
  );


  nor
  g2565
  (
    n2588,
    n2069,
    n652,
    n626,
    n2203
  );


  xor
  g2566
  (
    n2350,
    n2212,
    n605,
    n1351,
    n2085
  );


  xnor
  g2567
  (
    n2366,
    n629,
    n2208,
    n2218,
    n2133
  );


  nor
  g2568
  (
    n2450,
    n2164,
    n649,
    n627,
    n2192
  );


  xnor
  g2569
  (
    n2447,
    n2215,
    n2184,
    n639,
    n2143
  );


  nor
  g2570
  (
    n2379,
    n666,
    n2168,
    n2145,
    n2040
  );


  nand
  g2571
  (
    n2353,
    n658,
    n2006,
    n2196,
    n1965
  );


  nor
  g2572
  (
    n2539,
    n2130,
    n2061,
    n638,
    n2174
  );


  nand
  g2573
  (
    n2288,
    n2038,
    n1997,
    n614,
    n1878
  );


  and
  g2574
  (
    n2306,
    n662,
    n605,
    n636,
    n1977
  );


  xnor
  g2575
  (
    n2438,
    n655,
    n2069,
    n649,
    n661
  );


  nand
  g2576
  (
    n2252,
    n2190,
    n604,
    n2130,
    n629
  );


  nor
  g2577
  (
    n2385,
    n625,
    n665,
    n2202,
    n2172
  );


  or
  g2578
  (
    n2595,
    n2018,
    n2215,
    n652,
    n2120
  );


  xor
  g2579
  (
    n2266,
    n1991,
    n1998,
    n598,
    n2212
  );


  or
  g2580
  (
    n2292,
    n2056,
    n2160,
    n2004,
    n2134
  );


  and
  g2581
  (
    n2613,
    n1981,
    n670,
    n1958,
    n2176
  );


  nand
  g2582
  (
    n2436,
    n1975,
    n1967,
    n1996,
    n2166
  );


  xor
  g2583
  (
    n2384,
    n2002,
    n651,
    n2126,
    n2006
  );


  and
  g2584
  (
    n2619,
    n2070,
    n2246
  );


  not
  g2585
  (
    n2624,
    n2070
  );


  and
  g2586
  (
    n2622,
    n2244,
    n2072
  );


  xor
  g2587
  (
    n2620,
    n2072,
    n2245
  );


  buf
  g2588
  (
    n2617,
    n2071
  );


  xor
  g2589
  (
    n2623,
    n2072,
    n2242,
    n2239,
    n2243
  );


  or
  g2590
  (
    n2621,
    n2071,
    n2070,
    n2240,
    n1886
  );


  xnor
  g2591
  (
    n2618,
    n1885,
    n2071,
    n2241,
    n1352
  );


  not
  g2592
  (
    n2631,
    n2621
  );


  buf
  g2593
  (
    n2628,
    n2619
  );


  buf
  g2594
  (
    n2629,
    n2617
  );


  not
  g2595
  (
    n2634,
    n2623
  );


  not
  g2596
  (
    n2625,
    n2622
  );


  buf
  g2597
  (
    n2636,
    n2624
  );


  not
  g2598
  (
    n2637,
    n2623
  );


  not
  g2599
  (
    n2638,
    n2623
  );


  buf
  g2600
  (
    n2627,
    n2622
  );


  buf
  g2601
  (
    n2632,
    n2620
  );


  buf
  g2602
  (
    n2640,
    n2624
  );


  buf
  g2603
  (
    n2630,
    n2624
  );


  not
  g2604
  (
    n2635,
    n2621
  );


  buf
  g2605
  (
    n2633,
    n2622
  );


  not
  g2606
  (
    n2639,
    n2618
  );


  buf
  g2607
  (
    n2626,
    n2621
  );


  buf
  g2608
  (
    n2691,
    n2626
  );


  not
  g2609
  (
    n2684,
    n1894
  );


  not
  g2610
  (
    n2651,
    n2254
  );


  buf
  g2611
  (
    n2678,
    n1893
  );


  buf
  g2612
  (
    n2660,
    n2286
  );


  not
  g2613
  (
    n2647,
    n2274
  );


  buf
  g2614
  (
    n2689,
    n2625
  );


  not
  g2615
  (
    n2659,
    n2628
  );


  not
  g2616
  (
    n2672,
    n2637
  );


  not
  g2617
  (
    n2683,
    n1892
  );


  buf
  g2618
  (
    n2667,
    n2640
  );


  not
  g2619
  (
    n2656,
    n2291
  );


  not
  g2620
  (
    n2670,
    n2278
  );


  not
  g2621
  (
    n2654,
    n2639
  );


  not
  g2622
  (
    n2664,
    n2264
  );


  not
  g2623
  (
    n2676,
    n2248
  );


  not
  g2624
  (
    n2657,
    n2304
  );


  buf
  g2625
  (
    n2641,
    n2297
  );


  buf
  g2626
  (
    n2685,
    n1898
  );


  buf
  g2627
  (
    n2699,
    n2625
  );


  not
  g2628
  (
    n2701,
    n2631
  );


  buf
  g2629
  (
    n2674,
    n1895
  );


  not
  g2630
  (
    n2661,
    n2632
  );


  not
  g2631
  (
    n2700,
    n2629
  );


  buf
  g2632
  (
    n2696,
    n2273
  );


  not
  g2633
  (
    n2694,
    n2628
  );


  not
  g2634
  (
    n2695,
    n1894
  );


  buf
  g2635
  (
    n2644,
    n2309
  );


  buf
  g2636
  (
    n2671,
    n1896
  );


  buf
  g2637
  (
    n2665,
    n2626
  );


  buf
  g2638
  (
    n2669,
    n2634
  );


  or
  g2639
  (
    n2687,
    n2279,
    n1895
  );


  xor
  g2640
  (
    n2703,
    n2631,
    n2280,
    n2247,
    n2268
  );


  xnor
  g2641
  (
    n2682,
    n2636,
    n2300,
    n2633,
    n2638
  );


  nand
  g2642
  (
    n2642,
    n2314,
    n2630,
    n2634,
    n1895
  );


  xnor
  g2643
  (
    n2652,
    n2629,
    n1894,
    n2630,
    n1893
  );


  xnor
  g2644
  (
    n2658,
    n2634,
    n2282,
    n2638,
    n1893
  );


  or
  g2645
  (
    n2648,
    n2271,
    n2635,
    n2250,
    n2276
  );


  and
  g2646
  (
    n2702,
    n2275,
    n2285,
    n2307,
    n2257
  );


  or
  g2647
  (
    n2679,
    n2295,
    n2632,
    n2293,
    n2289
  );


  nor
  g2648
  (
    n2697,
    n2261,
    n1896,
    n2302,
    n2252
  );


  nand
  g2649
  (
    n2688,
    n2249,
    n1896,
    n2633,
    n2631
  );


  and
  g2650
  (
    n2649,
    n1892,
    n2303,
    n2072,
    n2288
  );


  xor
  g2651
  (
    n2650,
    n2628,
    n2639,
    n2310,
    n2311
  );


  nor
  g2652
  (
    n2643,
    n1897,
    n2632,
    n2255,
    n2636
  );


  xnor
  g2653
  (
    n2663,
    n2632,
    n2635,
    n2639,
    n2284
  );


  nor
  g2654
  (
    n2686,
    n2627,
    n2637,
    n2263,
    n2251
  );


  nor
  g2655
  (
    n2655,
    n2637,
    n2633,
    n1893,
    n2629
  );


  and
  g2656
  (
    n2677,
    n2308,
    n2277,
    n2635,
    n2270
  );


  xor
  g2657
  (
    n2690,
    n1896,
    n1892,
    n2625,
    n2627
  );


  or
  g2658
  (
    n2704,
    n2287,
    n2633,
    n2634,
    n2306
  );


  and
  g2659
  (
    n2698,
    n2296,
    n2631,
    n2638,
    n2626
  );


  xor
  g2660
  (
    n2666,
    n2635,
    n2256,
    n1894,
    n2640
  );


  xor
  g2661
  (
    n2673,
    n1898,
    n2636,
    n2266,
    n2253
  );


  nor
  g2662
  (
    n2692,
    n2272,
    n2299,
    n2281,
    n2638
  );


  or
  g2663
  (
    n2681,
    n2088,
    n2283,
    n2625,
    n1895
  );


  nand
  g2664
  (
    n2668,
    n2630,
    n1898,
    n2627
  );


  xor
  g2665
  (
    n2653,
    n2301,
    n2640,
    n2630,
    n2629
  );


  or
  g2666
  (
    n2693,
    n2292,
    n2637,
    n2298,
    n2626
  );


  nand
  g2667
  (
    n2662,
    n2265,
    n2627,
    n2258,
    n1897
  );


  xnor
  g2668
  (
    n2675,
    n2269,
    n2639,
    n2305,
    n1897
  );


  or
  g2669
  (
    n2645,
    n2640,
    n2262,
    n2628,
    n2260
  );


  nor
  g2670
  (
    n2680,
    n2259,
    n1897,
    n2267,
    n2290
  );


  nand
  g2671
  (
    n2646,
    n2312,
    n2313,
    n2294,
    n2636
  );


  xnor
  g2672
  (
    n2794,
    n2691,
    n2592,
    n2465,
    n1408
  );


  and
  g2673
  (
    n2816,
    n1372,
    n1362,
    n2654,
    n2528
  );


  and
  g2674
  (
    n2744,
    n2517,
    n2481,
    n1419,
    n1354
  );


  or
  g2675
  (
    n2792,
    n2681,
    n2500,
    n2345,
    n1355
  );


  nor
  g2676
  (
    n2882,
    n1401,
    n2505,
    n1421,
    n2515
  );


  or
  g2677
  (
    n2837,
    n2565,
    n2573,
    n2319,
    n1405
  );


  or
  g2678
  (
    n2797,
    n1440,
    n2397,
    n2702,
    n2678
  );


  nor
  g2679
  (
    n2724,
    n1431,
    n1425,
    n2684,
    n1375
  );


  and
  g2680
  (
    n2860,
    n1369,
    n1449,
    n1444,
    n1387
  );


  nor
  g2681
  (
    n2745,
    n1447,
    n2661,
    n2413,
    n2673
  );


  nand
  g2682
  (
    n2734,
    n2696,
    n2686,
    n2486,
    n1448
  );


  xnor
  g2683
  (
    n2814,
    n1415,
    n1436,
    n1404,
    n2608
  );


  nand
  g2684
  (
    n2843,
    n2698,
    n1426,
    n1360,
    n1357
  );


  and
  g2685
  (
    n2866,
    n1437,
    n2688,
    n2480,
    n2694
  );


  xor
  g2686
  (
    n2854,
    n2359,
    n2683,
    n2494,
    n2375
  );


  xnor
  g2687
  (
    n2875,
    n2662,
    n2649,
    n2694,
    n2437
  );


  or
  g2688
  (
    n2772,
    n2464,
    n2453,
    n2337,
    n2490
  );


  xnor
  g2689
  (
    n2948,
    n1414,
    n1374,
    n2237,
    n1402
  );


  and
  g2690
  (
    n2751,
    n1427,
    n2419,
    n2661,
    n2540
  );


  xor
  g2691
  (
    n2940,
    n1424,
    n2410,
    n160,
    n2326
  );


  nand
  g2692
  (
    KeyWire_0_0,
    n1362,
    n2447,
    n2657,
    n1388
  );


  nand
  g2693
  (
    n2855,
    n1902,
    n1420,
    n2510,
    n1454
  );


  nand
  g2694
  (
    n2717,
    n1429,
    n2401,
    n2542,
    n1363
  );


  or
  g2695
  (
    n2914,
    n2651,
    n1901,
    n2699,
    n2332
  );


  or
  g2696
  (
    n2802,
    n2667,
    n2695,
    n1416,
    n1424
  );


  nand
  g2697
  (
    n2928,
    n2365,
    n1450,
    n2555,
    n2689
  );


  and
  g2698
  (
    n2881,
    n2439,
    n1357,
    n1417,
    n2700
  );


  and
  g2699
  (
    n2768,
    n1394,
    n2703,
    n1377,
    n2654
  );


  xor
  g2700
  (
    n2715,
    n2696,
    n2691,
    n1450,
    n2471
  );


  nor
  g2701
  (
    n2919,
    n2316,
    n2405,
    n1427,
    n1419
  );


  nor
  g2702
  (
    n2900,
    n1357,
    n1431,
    n2612,
    n1365
  );


  xnor
  g2703
  (
    n2818,
    n2660,
    n1412,
    n1365,
    n2701
  );


  or
  g2704
  (
    n2933,
    n2516,
    n2651,
    n1364,
    n2373
  );


  nand
  g2705
  (
    n2842,
    n2686,
    n1412,
    n1394,
    n2457
  );


  nor
  g2706
  (
    n2781,
    n2398,
    n2649,
    n2651,
    n1354
  );


  or
  g2707
  (
    n2722,
    n2522,
    n1404,
    n2646,
    n2655
  );


  nor
  g2708
  (
    n2812,
    n2421,
    n2320,
    n2686,
    n2534
  );


  nand
  g2709
  (
    n2851,
    n2446,
    n2520,
    n1405,
    n1384
  );


  nand
  g2710
  (
    n2924,
    n1437,
    n2660,
    n1407,
    n1383
  );


  nor
  g2711
  (
    n2813,
    n2689,
    n2390,
    n2645,
    n2695
  );


  or
  g2712
  (
    n2735,
    n1368,
    n2354,
    n1427,
    n1358
  );


  xnor
  g2713
  (
    n2801,
    n1354,
    n1362,
    n2647,
    n1371
  );


  and
  g2714
  (
    n2778,
    n2697,
    n2489,
    n1374,
    n1363
  );


  xnor
  g2715
  (
    n2757,
    n2677,
    n2323,
    n1406,
    n1385
  );


  xnor
  g2716
  (
    n2718,
    n1391,
    n2644,
    n2697,
    n2680
  );


  nand
  g2717
  (
    n2748,
    n2384,
    n2325,
    n2409,
    n2676
  );


  xnor
  g2718
  (
    n2936,
    n1365,
    n2435,
    n2581,
    n1435
  );


  and
  g2719
  (
    n2821,
    n2461,
    n1400,
    n1441,
    n1399
  );


  nor
  g2720
  (
    n2938,
    n2602,
    n1439,
    n2683,
    n1451
  );


  xnor
  g2721
  (
    n2926,
    n1391,
    n1420,
    n2535,
    n1400
  );


  xor
  g2722
  (
    n2798,
    n2669,
    n2681,
    n1412,
    n1455
  );


  xnor
  g2723
  (
    n2896,
    n1417,
    n2670,
    n2671,
    n2543
  );


  xor
  g2724
  (
    n2943,
    n1440,
    n2682,
    n2663,
    n2483
  );


  nor
  g2725
  (
    n2836,
    n2491,
    n2400,
    n2645,
    n1446
  );


  nand
  g2726
  (
    n2951,
    n1418,
    n2324,
    n2649,
    n1408
  );


  xor
  g2727
  (
    n2720,
    n2476,
    n2648,
    n2507,
    n2512
  );


  nor
  g2728
  (
    n2820,
    n2659,
    n1358,
    n2668,
    n2689
  );


  xor
  g2729
  (
    n2769,
    n1445,
    n1447,
    n2643
  );


  or
  g2730
  (
    n2915,
    n1441,
    n2653,
    n2467,
    n1438
  );


  xor
  g2731
  (
    n2890,
    n1359,
    n2395,
    n2680,
    n1382
  );


  nor
  g2732
  (
    n2927,
    n1409,
    n2366,
    n2697,
    n1386
  );


  xnor
  g2733
  (
    n2904,
    n2669,
    n2424,
    n1361,
    n2677
  );


  or
  g2734
  (
    n2796,
    n2562,
    n2646,
    n2672,
    n2474
  );


  and
  g2735
  (
    n2775,
    n1417,
    n2686,
    n2448,
    n1431
  );


  and
  g2736
  (
    n2749,
    n2650,
    n1388,
    n2652,
    n2473
  );


  nand
  g2737
  (
    n2947,
    n1356,
    n2702,
    n1373,
    n1405
  );


  xor
  g2738
  (
    n2844,
    n2315,
    n1403,
    n1435,
    n2683
  );


  or
  g2739
  (
    n2791,
    n1393,
    n2553,
    n2469,
    n2591
  );


  xnor
  g2740
  (
    n2771,
    n2429,
    n2442,
    n1444,
    n2586
  );


  xnor
  g2741
  (
    n2859,
    n1429,
    n2672,
    n1388,
    n2597
  );


  nand
  g2742
  (
    n2830,
    n2501,
    n2417,
    n2679,
    n2666
  );


  or
  g2743
  (
    n2780,
    n2704,
    n2470,
    n2668,
    n2703
  );


  xnor
  g2744
  (
    n2815,
    n1368,
    n2659,
    n2392,
    n1438
  );


  xor
  g2745
  (
    n2942,
    n2655,
    n2572,
    n2660,
    n1444
  );


  or
  g2746
  (
    n2767,
    n1445,
    n2466,
    n2545,
    n1387
  );


  and
  g2747
  (
    n2823,
    n2508,
    n1375,
    n2338,
    n2653
  );


  and
  g2748
  (
    n2764,
    n2647,
    n1354,
    n1443,
    n2674
  );


  xor
  g2749
  (
    n2827,
    n2689,
    n1398,
    n2699,
    n1386
  );


  or
  g2750
  (
    n2742,
    n2526,
    n1413,
    n2564,
    n2402
  );


  xor
  g2751
  (
    n2788,
    n2673,
    n2333,
    n2530,
    n2653
  );


  and
  g2752
  (
    n2723,
    n2541,
    n2687,
    n2664,
    n1360
  );


  xor
  g2753
  (
    n2874,
    n1392,
    n2654,
    n2361,
    n2682
  );


  xor
  g2754
  (
    n2833,
    n1381,
    n2646,
    n2607,
    n2680
  );


  xnor
  g2755
  (
    n2829,
    n1381,
    n2676,
    n1368,
    n1443
  );


  xor
  g2756
  (
    n2785,
    n2443,
    n1371,
    n2418,
    n2690
  );


  xnor
  g2757
  (
    n2863,
    n2692,
    n1394,
    n2355,
    n1356
  );


  and
  g2758
  (
    n2870,
    n2658,
    n1439,
    n2652,
    n2693
  );


  xnor
  g2759
  (
    n2872,
    n2647,
    n2667,
    n2423,
    n2645
  );


  and
  g2760
  (
    n2736,
    n2440,
    n2605,
    n1390,
    n1416
  );


  xnor
  g2761
  (
    n2714,
    n1409,
    n2680,
    n2677,
    n2657
  );


  or
  g2762
  (
    n2784,
    n2678,
    n1374,
    n1422,
    n2321
  );


  nand
  g2763
  (
    n2807,
    n1396,
    n1430,
    n2665,
    n1422
  );


  xor
  g2764
  (
    n2810,
    n1408,
    n1364,
    n1363,
    n2678
  );


  xor
  g2765
  (
    n2883,
    n2691,
    n2544,
    n1428,
    n2644
  );


  nand
  g2766
  (
    n2712,
    n1363,
    n2580,
    n2672,
    n2613
  );


  xnor
  g2767
  (
    n2732,
    n1384,
    n1392,
    n1418,
    n2648
  );


  or
  g2768
  (
    n2888,
    n1439,
    n1377,
    n2237,
    n1383
  );


  xor
  g2769
  (
    n2803,
    n2569,
    n1440,
    n2644,
    n1421
  );


  or
  g2770
  (
    n2941,
    n1378,
    n1445,
    n2650,
    n2682
  );


  and
  g2771
  (
    n2905,
    n1448,
    n2521,
    n1399,
    n2700
  );


  or
  g2772
  (
    n2728,
    n1358,
    n2644,
    n1353,
    n2403
  );


  xnor
  g2773
  (
    n2824,
    n2693,
    n2388,
    n1453,
    n2601
  );


  nor
  g2774
  (
    n2886,
    n2616,
    n1385,
    n1404,
    n2347
  );


  and
  g2775
  (
    n2822,
    n1402,
    n2381,
    n2391,
    n2687
  );


  nand
  g2776
  (
    n2952,
    n1411,
    n1376,
    n1423,
    n2344
  );


  and
  g2777
  (
    n2777,
    n2578,
    n1366,
    n1425,
    n2615
  );


  nor
  g2778
  (
    n2950,
    n2658,
    n1353,
    n1421,
    n1902
  );


  nand
  g2779
  (
    n2917,
    n2551,
    n2585,
    n2529,
    n2329
  );


  xnor
  g2780
  (
    KeyWire_0_12,
    n2660,
    n1440,
    n2666,
    n2674
  );


  xor
  g2781
  (
    n2795,
    n1392,
    n1369,
    n1370,
    n1401
  );


  nand
  g2782
  (
    n2897,
    n2451,
    n1413,
    n2379,
    n1383
  );


  nor
  g2783
  (
    n2727,
    n2690,
    n2422,
    n2679,
    n2380
  );


  nor
  g2784
  (
    n2920,
    n2695,
    n1373,
    n2702,
    n1449
  );


  xor
  g2785
  (
    n2770,
    n2694,
    n1372,
    n1435,
    n1396
  );


  and
  g2786
  (
    n2945,
    n1385,
    n2673,
    n2382,
    n2604
  );


  nor
  g2787
  (
    n2892,
    n1403,
    n2697,
    n1415,
    n1409
  );


  nand
  g2788
  (
    n2907,
    n1423,
    n2698,
    n2456,
    n2675
  );


  xor
  g2789
  (
    n2916,
    n1426,
    n1367,
    n2460,
    n1379
  );


  xor
  g2790
  (
    n2935,
    n2387,
    n2430,
    n2681,
    n2504
  );


  xor
  g2791
  (
    n2806,
    n1418,
    n2675,
    n2536,
    n1399
  );


  or
  g2792
  (
    n2865,
    n2584,
    n1415,
    n1361,
    n2598
  );


  xnor
  g2793
  (
    n2739,
    n2698,
    n1381,
    n1414,
    n1386
  );


  nand
  g2794
  (
    n2711,
    n2676,
    n2571,
    n1411,
    n1402
  );


  xnor
  g2795
  (
    n2853,
    n1359,
    n1368,
    n2575,
    n2236
  );


  or
  g2796
  (
    n2949,
    n2485,
    n1373,
    n2657,
    n2343
  );


  and
  g2797
  (
    n2709,
    n1404,
    n2463,
    n2554,
    n2236
  );


  nand
  g2798
  (
    n2759,
    n2568,
    n1418,
    n2548,
    n2561
  );


  or
  g2799
  (
    n2925,
    n1446,
    n1412,
    n2350,
    n2670
  );


  nand
  g2800
  (
    n2835,
    n1442,
    n2317,
    n2533,
    n1434
  );


  nand
  g2801
  (
    n2856,
    n2472,
    n2434,
    n2525,
    n2654
  );


  xor
  g2802
  (
    n2783,
    n2674,
    n2656,
    n1376,
    n1366
  );


  nand
  g2803
  (
    n2877,
    n2590,
    n1447,
    n2342,
    n2656
  );


  xnor
  g2804
  (
    n2809,
    n1380,
    n1380,
    n2649,
    n2643
  );


  and
  g2805
  (
    n2887,
    n2588,
    n1364,
    n1390,
    n2532
  );


  nand
  g2806
  (
    n2930,
    n1442,
    n1410,
    n2687,
    n2334
  );


  and
  g2807
  (
    n2755,
    n1375,
    n1396,
    n1455,
    n1453
  );


  or
  g2808
  (
    n2817,
    n2374,
    n1369,
    n2671,
    n2611
  );


  and
  g2809
  (
    n2903,
    n1371,
    n1454,
    n2701,
    n1390
  );


  nand
  g2810
  (
    n2901,
    n1392,
    n1393,
    n2537,
    n1378
  );


  nor
  g2811
  (
    n2869,
    n1376,
    n2664,
    n2527,
    n2331
  );


  or
  g2812
  (
    n2752,
    n2673,
    n1435,
    n2593,
    n2428
  );


  nand
  g2813
  (
    n2831,
    n1355,
    n1408,
    n1407,
    n2589
  );


  xor
  g2814
  (
    n2832,
    n1397,
    n2238,
    n2438,
    n2479
  );


  nor
  g2815
  (
    n2707,
    n1402,
    n1393,
    n1365,
    n1399
  );


  and
  g2816
  (
    n2811,
    n2596,
    n1382,
    n2523,
    n1902
  );


  or
  g2817
  (
    n2839,
    n2519,
    n1397,
    n1433,
    n2558
  );


  and
  g2818
  (
    n2850,
    n1361,
    n1366,
    n1406,
    n1430
  );


  xor
  g2819
  (
    n2804,
    n2679,
    n2692,
    n1434,
    n1389
  );


  xnor
  g2820
  (
    n2828,
    n1430,
    n2514,
    n1452,
    n2703
  );


  or
  g2821
  (
    n2846,
    n2546,
    n1367,
    n1452,
    n2661
  );


  and
  g2822
  (
    n2731,
    n2351,
    n1379,
    n1426,
    n2336
  );


  nor
  g2823
  (
    n2799,
    n2518,
    n2704,
    n1443,
    n2436
  );


  xor
  g2824
  (
    n2841,
    n1397,
    n2656,
    n2349,
    n2700
  );


  and
  g2825
  (
    n2884,
    n1359,
    n2455,
    n1353,
    n1384
  );


  nand
  g2826
  (
    n2932,
    n1436,
    n2549,
    n1401,
    n1409
  );


  nor
  g2827
  (
    n2922,
    n2511,
    n1410,
    n1432,
    n2687
  );


  or
  g2828
  (
    n2730,
    n2587,
    n2666,
    n1391,
    n2702
  );


  nor
  g2829
  (
    n2738,
    n2655,
    n2238,
    n1367,
    n2684
  );


  xnor
  g2830
  (
    n2871,
    n1387,
    n2356,
    n1355,
    n1451
  );


  xnor
  g2831
  (
    n2939,
    n2651,
    n2616,
    n2696,
    n2657
  );


  xnor
  g2832
  (
    n2852,
    n2704,
    n2369,
    n2371,
    n2559
  );


  nor
  g2833
  (
    n2847,
    n2652,
    n1449,
    n2404,
    n2478
  );


  xnor
  g2834
  (
    n2743,
    n2577,
    n1433,
    n1413,
    n1396
  );


  nor
  g2835
  (
    n2834,
    n2665,
    n2645,
    n1378,
    n2496
  );


  xor
  g2836
  (
    n2946,
    n1400,
    n2493,
    n2416,
    n2346
  );


  nand
  g2837
  (
    n2760,
    n2372,
    n1403,
    n2431,
    n2445
  );


  or
  g2838
  (
    n2782,
    n2450,
    n2676,
    n1425,
    n1379
  );


  nor
  g2839
  (
    n2895,
    n2412,
    n1403,
    n2433,
    n2368
  );


  or
  g2840
  (
    n2705,
    n1413,
    n2570,
    n2701,
    n2662
  );


  xor
  g2841
  (
    n2774,
    n1381,
    n1450,
    n2449,
    n2643
  );


  nand
  g2842
  (
    n2921,
    n2385,
    n1356,
    n2693,
    n2653
  );


  nand
  g2843
  (
    n2719,
    n2360,
    n2502,
    n1398,
    n1377
  );


  xor
  g2844
  (
    n2733,
    n1380,
    n1442,
    n2667,
    n1419
  );


  nor
  g2845
  (
    n2762,
    n2685,
    n2358,
    n1438,
    n2566
  );


  nor
  g2846
  (
    n2910,
    n2650,
    n1438,
    n2669
  );


  xnor
  g2847
  (
    n2912,
    n2609,
    n2671,
    n1446,
    n1420
  );


  and
  g2848
  (
    n2867,
    n1357,
    n1360,
    n2327,
    n2616
  );


  xor
  g2849
  (
    n2754,
    n1370,
    n2704,
    n1398,
    n2614
  );


  xor
  g2850
  (
    n2800,
    n2650,
    n2685,
    n1353,
    n1386
  );


  or
  g2851
  (
    n2885,
    n1395,
    n2394,
    n1394,
    n2698
  );


  nor
  g2852
  (
    n2765,
    n2497,
    n2667,
    n1446,
    n1416
  );


  and
  g2853
  (
    n2880,
    n2454,
    n2378,
    n2659,
    n2700
  );


  and
  g2854
  (
    n2741,
    n2503,
    n2475,
    n2642,
    n2363
  );


  and
  g2855
  (
    n2934,
    n2678,
    n1390,
    n1383,
    n1452
  );


  nand
  g2856
  (
    n2944,
    n2524,
    n1405,
    n1391,
    n2647
  );


  and
  g2857
  (
    n2848,
    n1406,
    n2663,
    n2681,
    n2665
  );


  or
  g2858
  (
    n2753,
    n1432,
    n2389,
    n1400,
    n2685
  );


  xor
  g2859
  (
    n2861,
    n2459,
    n1430,
    n1427,
    n1398
  );


  and
  g2860
  (
    n2766,
    n2642,
    n2236,
    n2600,
    n1355
  );


  and
  g2861
  (
    n2878,
    n1431,
    n2420,
    n1454
  );


  or
  g2862
  (
    n2894,
    n2238,
    n2642,
    n1449,
    n1372
  );


  xnor
  g2863
  (
    n2913,
    n2432,
    n2335,
    n1367,
    n1428
  );


  nor
  g2864
  (
    n2793,
    n1420,
    n2648,
    n1428,
    n2352
  );


  or
  g2865
  (
    n2849,
    n2701,
    n1385,
    n2487,
    n1417
  );


  nand
  g2866
  (
    n2906,
    n1429,
    n1424,
    n2560,
    n2672
  );


  xor
  g2867
  (
    n2789,
    n1447,
    n2426,
    n2610,
    n2663
  );


  nand
  g2868
  (
    n2746,
    n1361,
    n1437,
    n2237,
    n1434
  );


  nor
  g2869
  (
    n2790,
    n2661,
    n1425,
    n2699,
    n1377
  );


  or
  g2870
  (
    n2864,
    n2367,
    n2458,
    n2377,
    n2671
  );


  nor
  g2871
  (
    n2908,
    n2427,
    n2658,
    n2563,
    n1445
  );


  and
  g2872
  (
    n2761,
    n1432,
    n1901,
    n2462,
    n2322
  );


  and
  g2873
  (
    n2706,
    n1389,
    n2663,
    n2665,
    n2694
  );


  xnor
  g2874
  (
    n2729,
    n1360,
    n2576,
    n2509,
    n2238
  );


  xor
  g2875
  (
    n2929,
    n2668,
    n1395,
    n1370,
    n2690
  );


  xor
  g2876
  (
    n2825,
    n2574,
    n1407,
    n2582,
    n2691
  );


  xnor
  g2877
  (
    n2862,
    n2513,
    n1371,
    n2376,
    n2677
  );


  or
  g2878
  (
    n2891,
    n2383,
    n2641,
    n1407,
    n1411
  );


  nor
  g2879
  (
    n2819,
    n2646,
    n2393,
    n1397,
    n2557
  );


  or
  g2880
  (
    n2805,
    n2341,
    n1429,
    n2407,
    n2688
  );


  nor
  g2881
  (
    n2787,
    n1378,
    n1372,
    n2685,
    n2482
  );


  nand
  g2882
  (
    n2758,
    n1416,
    n1436,
    n2583,
    n2688
  );


  xor
  g2883
  (
    n2737,
    n2498,
    n2556,
    n1395,
    n2599
  );


  nand
  g2884
  (
    n2750,
    n2679,
    n2648,
    n2703,
    n2547
  );


  xnor
  g2885
  (
    n2713,
    n1422,
    n2330,
    n2506,
    n2658
  );


  nor
  g2886
  (
    n2899,
    n1382,
    n2531,
    n2370,
    n2579
  );


  or
  g2887
  (
    n2725,
    n2235,
    n2684,
    n1433
  );


  or
  g2888
  (
    n2776,
    n1362,
    n2688,
    n2656,
    n2675
  );


  xnor
  g2889
  (
    n2923,
    n1401,
    n2364,
    n1389,
    n1441
  );


  xnor
  g2890
  (
    n2876,
    n2693,
    n1374,
    n2237,
    n2495
  );


  nand
  g2891
  (
    n2808,
    n2484,
    n2664,
    n1393,
    n1373
  );


  xor
  g2892
  (
    n2937,
    n1902,
    n2670,
    n1451,
    n2452
  );


  nor
  g2893
  (
    n2858,
    n1388,
    n1414,
    n2603,
    n2683
  );


  nand
  g2894
  (
    n2779,
    n1441,
    n2662,
    n2499,
    n1415
  );


  xor
  g2895
  (
    n2826,
    n2668,
    n1451,
    n2477,
    n1424
  );


  nand
  g2896
  (
    n2911,
    n1434,
    n1444,
    n1423,
    n1369
  );


  nand
  g2897
  (
    n2909,
    n1442,
    n2595,
    n2690,
    n1384
  );


  xnor
  g2898
  (
    n2845,
    n2675,
    n2414,
    n2415,
    n2666
  );


  xnor
  g2899
  (
    n2902,
    n1406,
    n2386,
    n1422,
    n2659
  );


  or
  g2900
  (
    n2747,
    n1419,
    n1414,
    n2692,
    n1443
  );


  nor
  g2901
  (
    n2873,
    n1358,
    n1423,
    n2538,
    n2641
  );


  xor
  g2902
  (
    n2721,
    n1395,
    n2444,
    n2641,
    n2340
  );


  xor
  g2903
  (
    n2868,
    n1375,
    n2492,
    n1448,
    n2642
  );


  xnor
  g2904
  (
    n2716,
    n2552,
    n1389,
    n1359,
    n2339
  );


  or
  g2905
  (
    n2710,
    n1439,
    n1380,
    n2662,
    n1366
  );


  nand
  g2906
  (
    n2786,
    n2328,
    n1428,
    n1379,
    n2318
  );


  and
  g2907
  (
    n2740,
    n2699,
    n2652,
    n1433,
    n2664
  );


  xor
  g2908
  (
    n2773,
    n1410,
    n2408,
    n2696,
    n2441
  );


  and
  g2909
  (
    n2931,
    n2235,
    n1411,
    n2362,
    n2655
  );


  or
  g2910
  (
    n2898,
    n2682,
    n2488,
    n2674,
    n1436
  );


  xnor
  g2911
  (
    n2840,
    n2468,
    n2539,
    n1410,
    n2550
  );


  nand
  g2912
  (
    n2893,
    n1364,
    n1453,
    n2695,
    n1450
  );


  and
  g2913
  (
    n2838,
    n1432,
    n2357,
    n2567,
    n1426
  );


  nor
  g2914
  (
    n2889,
    n1452,
    n1455,
    n2399,
    n1448
  );


  nand
  g2915
  (
    n2918,
    n1387,
    n2236,
    n1437,
    n1455
  );


  or
  g2916
  (
    n2726,
    n2594,
    n2396,
    n1421,
    n2670
  );


  xnor
  g2917
  (
    n2708,
    n2606,
    n1356,
    n2692,
    n1382
  );


  nor
  g2918
  (
    n2879,
    n2406,
    n2411,
    n2353,
    n1453
  );


  xnor
  g2919
  (
    n2756,
    n1376,
    n2425,
    n2348,
    n1370
  );


  nor
  g2920
  (
    n2999,
    n2821,
    n2877,
    n2771,
    n1912
  );


  nand
  g2921
  (
    n2989,
    n2897,
    n2710,
    n2775,
    n2722
  );


  or
  g2922
  (
    n2995,
    n2876,
    n2875,
    n2943,
    n2840
  );


  xnor
  g2923
  (
    n3006,
    n2705,
    n2904,
    n2736,
    n2852
  );


  xnor
  g2924
  (
    n2979,
    n2865,
    n2822,
    n2874,
    n2930
  );


  xor
  g2925
  (
    n2977,
    n1911,
    n2887,
    n2913,
    n2939
  );


  xnor
  g2926
  (
    n3009,
    n2915,
    n2753,
    n2889,
    n2818
  );


  or
  g2927
  (
    n2975,
    n2933,
    n2867,
    n2751,
    n2756
  );


  nand
  g2928
  (
    n2998,
    n2895,
    n2906,
    n2911,
    n2839
  );


  nand
  g2929
  (
    n3016,
    n2814,
    n2725,
    n1911,
    n2836
  );


  nor
  g2930
  (
    n2984,
    n2755,
    n2908,
    n2944,
    n2860
  );


  xor
  g2931
  (
    n2992,
    n2924,
    n2805,
    n2768,
    n2949
  );


  nand
  g2932
  (
    n2969,
    n2918,
    n2824,
    n2901,
    n2729
  );


  xor
  g2933
  (
    n2976,
    n2873,
    n2782,
    n2929,
    n2932
  );


  xnor
  g2934
  (
    n3015,
    n2854,
    n2793,
    n1912,
    n2850
  );


  xnor
  g2935
  (
    n2997,
    n2721,
    n2816,
    n2749,
    n2763
  );


  nor
  g2936
  (
    n2981,
    n2807,
    n2893,
    n2886,
    n2864
  );


  nor
  g2937
  (
    n2967,
    n2902,
    n2828,
    n1911,
    n2734
  );


  or
  g2938
  (
    n2988,
    n1912,
    n2802,
    n2842,
    n2861
  );


  nand
  g2939
  (
    n2970,
    n2727,
    n2796,
    n2863,
    n2869
  );


  or
  g2940
  (
    n3005,
    n2896,
    n2898,
    n2788,
    n1911
  );


  nand
  g2941
  (
    n2961,
    n2937,
    n2928,
    n2952,
    n2765
  );


  xnor
  g2942
  (
    n2963,
    n2759,
    n2858,
    n2792,
    n2799
  );


  and
  g2943
  (
    n2994,
    n2733,
    n2879,
    n2740,
    n2833
  );


  and
  g2944
  (
    n3004,
    n2914,
    n2744,
    n2743,
    n2757
  );


  and
  g2945
  (
    n3010,
    n2856,
    n2794,
    n2945,
    n2724
  );


  xnor
  g2946
  (
    n2983,
    n2741,
    n2769,
    n2767,
    n2866
  );


  nand
  g2947
  (
    n2957,
    n2880,
    n2927,
    n2885,
    n2938
  );


  nor
  g2948
  (
    n2958,
    n2925,
    n2888,
    n2719,
    n2935
  );


  nand
  g2949
  (
    KeyWire_0_1,
    n2829,
    n2855,
    n2826,
    n2709
  );


  and
  g2950
  (
    n2953,
    n2832,
    n2778,
    n2789,
    n2909
  );


  nand
  g2951
  (
    n3003,
    n2810,
    n2786,
    n2857,
    n2730
  );


  and
  g2952
  (
    n2964,
    n2819,
    n2809,
    n2762,
    n2849
  );


  nor
  g2953
  (
    n2991,
    n2834,
    n2916,
    n2838,
    n2732
  );


  xnor
  g2954
  (
    n3002,
    n2817,
    n2776,
    n2712,
    n2899
  );


  nand
  g2955
  (
    n2959,
    n2714,
    n2773,
    n2890,
    n2770
  );


  xnor
  g2956
  (
    n2965,
    n2891,
    n2823,
    n2803,
    n2737
  );


  nand
  g2957
  (
    n2960,
    n2947,
    n2827,
    n2907,
    n2951
  );


  nand
  g2958
  (
    n3014,
    n2774,
    n2790,
    n2777,
    n2920
  );


  xor
  g2959
  (
    n2980,
    n2871,
    n2706,
    n2715,
    n2934
  );


  nor
  g2960
  (
    n2955,
    n2711,
    n2851,
    n2795,
    n2848
  );


  and
  g2961
  (
    n3011,
    n2830,
    n2812,
    n2844,
    n2742
  );


  xor
  g2962
  (
    n2971,
    n2784,
    n2806,
    n2931,
    n2881
  );


  nand
  g2963
  (
    n2978,
    n2707,
    n2798,
    n2738,
    n2859
  );


  nor
  g2964
  (
    n2993,
    n2811,
    n2720,
    n2900,
    n2716
  );


  nor
  g2965
  (
    n2968,
    n2797,
    n2785,
    n2841,
    n2750
  );


  nor
  g2966
  (
    n2982,
    n2870,
    n2772,
    n2921,
    n2800
  );


  xnor
  g2967
  (
    n3007,
    n2948,
    n2746,
    n2905,
    n2808
  );


  nor
  g2968
  (
    n3012,
    n2843,
    n2835,
    n2941,
    n2853
  );


  nand
  g2969
  (
    n2954,
    n2783,
    n2940,
    n2922,
    n2787
  );


  and
  g2970
  (
    n3001,
    n2845,
    n2820,
    n1912,
    n2752
  );


  or
  g2971
  (
    n2966,
    n2761,
    n2739,
    n2936,
    n2735
  );


  or
  g2972
  (
    n2956,
    n2862,
    n2837,
    n2760,
    n2903
  );


  nor
  g2973
  (
    n2987,
    n2946,
    n2718,
    n2825,
    n2723
  );


  nor
  g2974
  (
    n3000,
    n2923,
    n2912,
    n2781,
    n2758
  );


  xor
  g2975
  (
    n3008,
    n2883,
    n2745,
    n2780,
    n2766
  );


  xor
  g2976
  (
    n2974,
    n2926,
    n2884,
    n2731,
    n2919
  );


  xnor
  g2977
  (
    n2986,
    n2804,
    n2713,
    n2882,
    n2754
  );


  and
  g2978
  (
    n3013,
    n2747,
    n2831,
    n2894,
    n2872
  );


  nand
  g2979
  (
    n2985,
    n2910,
    n2892,
    n2801,
    n2717
  );


  xor
  g2980
  (
    n2996,
    n2813,
    n2942,
    n2846,
    n2847
  );


  and
  g2981
  (
    n2962,
    n2815,
    n2878,
    n2791,
    n2728
  );


  nand
  g2982
  (
    n2973,
    n2917,
    n2708,
    n2764,
    n2950
  );


  and
  g2983
  (
    n2990,
    n2748,
    n2868,
    n2726,
    n2779
  );


  and
  g2984
  (
    n3024,
    n2973,
    n2980,
    n2998,
    n2989
  );


  xor
  g2985
  (
    n3022,
    n2993,
    n2970,
    n3013,
    n2964
  );


  or
  g2986
  (
    n3027,
    n2982,
    n2977,
    n3009,
    n3012
  );


  nor
  g2987
  (
    n3026,
    n3014,
    n2971,
    n3016,
    n3002
  );


  nor
  g2988
  (
    n3031,
    n3005,
    n2965,
    n2992,
    n3008
  );


  and
  g2989
  (
    n3025,
    n2955,
    n2954,
    n2969,
    n3000
  );


  nand
  g2990
  (
    n3018,
    n2975,
    n2990,
    n3010,
    n2986
  );


  and
  g2991
  (
    n3017,
    n2966,
    n2974,
    n2997,
    n2999
  );


  xnor
  g2992
  (
    n3021,
    n2984,
    n2983,
    n2979,
    n2953
  );


  xor
  g2993
  (
    n3023,
    n2981,
    n2978,
    n2958,
    n2959
  );


  nand
  g2994
  (
    n3030,
    n3003,
    n2994,
    n2961,
    n2996
  );


  nand
  g2995
  (
    n3029,
    n2960,
    n3001,
    n2995,
    n2985
  );


  and
  g2996
  (
    n3019,
    n2988,
    n2972,
    n2957,
    n2987
  );


  nand
  g2997
  (
    n3020,
    n2976,
    n2991,
    n2963,
    n3006
  );


  or
  g2998
  (
    n3032,
    n2962,
    n2967,
    n3004,
    n3015
  );


  nor
  g2999
  (
    n3028,
    n2956,
    n3011,
    n3007,
    n2968
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n2857,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n2972,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n1155,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n2138,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n691,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n2467,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n475,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n693,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n709,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n2004,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n865,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1009,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n2763,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1107,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n954,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n2106,
    KeyNOTWire_0_15
  );


endmodule

