// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_976_2713 written by SynthGen on 2021/05/24 19:48:32
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_976_2713 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27,
 n968, n970, n975, n972, n986, n967, n980, n978,
 n966, n984, n985, n981, n974, n983, n976, n979,
 n969, n989, n971, n982, n988, n977, n991, n1001,
 n999, n1000, n1002, n998, n1003);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27;

output n968, n970, n975, n972, n986, n967, n980, n978,
 n966, n984, n985, n981, n974, n983, n976, n979,
 n969, n989, n971, n982, n988, n977, n991, n1001,
 n999, n1000, n1002, n998, n1003;

wire n28, n29, n30, n31, n32, n33, n34, n35,
 n36, n37, n38, n39, n40, n41, n42, n43,
 n44, n45, n46, n47, n48, n49, n50, n51,
 n52, n53, n54, n55, n56, n57, n58, n59,
 n60, n61, n62, n63, n64, n65, n66, n67,
 n68, n69, n70, n71, n72, n73, n74, n75,
 n76, n77, n78, n79, n80, n81, n82, n83,
 n84, n85, n86, n87, n88, n89, n90, n91,
 n92, n93, n94, n95, n96, n97, n98, n99,
 n100, n101, n102, n103, n104, n105, n106, n107,
 n108, n109, n110, n111, n112, n113, n114, n115,
 n116, n117, n118, n119, n120, n121, n122, n123,
 n124, n125, n126, n127, n128, n129, n130, n131,
 n132, n133, n134, n135, n136, n137, n138, n139,
 n140, n141, n142, n143, n144, n145, n146, n147,
 n148, n149, n150, n151, n152, n153, n154, n155,
 n156, n157, n158, n159, n160, n161, n162, n163,
 n164, n165, n166, n167, n168, n169, n170, n171,
 n172, n173, n174, n175, n176, n177, n178, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n189, n190, n191, n192, n193, n194, n195,
 n196, n197, n198, n199, n200, n201, n202, n203,
 n204, n205, n206, n207, n208, n209, n210, n211,
 n212, n213, n214, n215, n216, n217, n218, n219,
 n220, n221, n222, n223, n224, n225, n226, n227,
 n228, n229, n230, n231, n232, n233, n234, n235,
 n236, n237, n238, n239, n240, n241, n242, n243,
 n244, n245, n246, n247, n248, n249, n250, n251,
 n252, n253, n254, n255, n256, n257, n258, n259,
 n260, n261, n262, n263, n264, n265, n266, n267,
 n268, n269, n270, n271, n272, n273, n274, n275,
 n276, n277, n278, n279, n280, n281, n282, n283,
 n284, n285, n286, n287, n288, n289, n290, n291,
 n292, n293, n294, n295, n296, n297, n298, n299,
 n300, n301, n302, n303, n304, n305, n306, n307,
 n308, n309, n310, n311, n312, n313, n314, n315,
 n316, n317, n318, n319, n320, n321, n322, n323,
 n324, n325, n326, n327, n328, n329, n330, n331,
 n332, n333, n334, n335, n336, n337, n338, n339,
 n340, n341, n342, n343, n344, n345, n346, n347,
 n348, n349, n350, n351, n352, n353, n354, n355,
 n356, n357, n358, n359, n360, n361, n362, n363,
 n364, n365, n366, n367, n368, n369, n370, n371,
 n372, n373, n374, n375, n376, n377, n378, n379,
 n380, n381, n382, n383, n384, n385, n386, n387,
 n388, n389, n390, n391, n392, n393, n394, n395,
 n396, n397, n398, n399, n400, n401, n402, n403,
 n404, n405, n406, n407, n408, n409, n410, n411,
 n412, n413, n414, n415, n416, n417, n418, n419,
 n420, n421, n422, n423, n424, n425, n426, n427,
 n428, n429, n430, n431, n432, n433, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n634, n635,
 n636, n637, n638, n639, n640, n641, n642, n643,
 n644, n645, n646, n647, n648, n649, n650, n651,
 n652, n653, n654, n655, n656, n657, n658, n659,
 n660, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685, n686, n687, n688, n689, n690, n691,
 n692, n693, n694, n695, n696, n697, n698, n699,
 n700, n701, n702, n703, n704, n705, n706, n707,
 n708, n709, n710, n711, n712, n713, n714, n715,
 n716, n717, n718, n719, n720, n721, n722, n723,
 n724, n725, n726, n727, n728, n729, n730, n731,
 n732, n733, n734, n735, n736, n737, n738, n739,
 n740, n741, n742, n743, n744, n745, n746, n747,
 n748, n749, n750, n751, n752, n753, n754, n755,
 n756, n757, n758, n759, n760, n761, n762, n763,
 n764, n765, n766, n767, n768, n769, n770, n771,
 n772, n773, n774, n775, n776, n777, n778, n779,
 n780, n781, n782, n783, n784, n785, n786, n787,
 n788, n789, n790, n791, n792, n793, n794, n795,
 n796, n797, n798, n799, n800, n801, n802, n803,
 n804, n805, n806, n807, n808, n809, n810, n811,
 n812, n813, n814, n815, n816, n817, n818, n819,
 n820, n821, n822, n823, n824, n825, n826, n827,
 n828, n829, n830, n831, n832, n833, n834, n835,
 n836, n837, n838, n839, n840, n841, n842, n843,
 n844, n845, n846, n847, n848, n849, n850, n851,
 n852, n853, n854, n855, n856, n857, n858, n859,
 n860, n861, n862, n863, n864, n865, n866, n867,
 n868, n869, n870, n871, n872, n873, n874, n875,
 n876, n877, n878, n879, n880, n881, n882, n883,
 n884, n885, n886, n887, n888, n889, n890, n891,
 n892, n893, n894, n895, n896, n897, n898, n899,
 n900, n901, n902, n903, n904, n905, n906, n907,
 n908, n909, n910, n911, n912, n913, n914, n915,
 n916, n917, n918, n919, n920, n921, n922, n923,
 n924, n925, n926, n927, n928, n929, n930, n931,
 n932, n933, n934, n935, n936, n937, n938, n939,
 n940, n941, n942, n943, n944, n945, n946, n947,
 n948, n949, n950, n951, n952, n953, n954, n955,
 n956, n957, n958, n959, n960, n961, n962, n963,
 n964, n965, n973, n987, n990, n992, n993, n994,
 n995, n996, n997;

buf  g0 (n42, n17);
buf  g1 (n77, n13);
buf  g2 (n53, n5);
not  g3 (n37, n14);
buf  g4 (n78, n9);
not  g5 (n32, n13);
not  g6 (n36, n9);
buf  g7 (n55, n4);
not  g8 (n79, n14);
buf  g9 (n63, n7);
not  g10 (n28, n7);
not  g11 (n34, n17);
not  g12 (n40, n10);
buf  g13 (n31, n4);
buf  g14 (n64, n12);
not  g15 (n71, n12);
not  g16 (n82, n12);
not  g17 (n62, n11);
buf  g18 (n66, n8);
buf  g19 (n59, n18);
not  g20 (n72, n14);
not  g21 (n45, n3);
not  g22 (n81, n11);
not  g23 (n51, n12);
not  g24 (n30, n13);
buf  g25 (n33, n16);
not  g26 (n48, n10);
not  g27 (n56, n2);
not  g28 (n44, n19);
buf  g29 (n69, n13);
buf  g30 (n80, n18);
not  g31 (n43, n19);
buf  g32 (n41, n16);
buf  g33 (n60, n6);
buf  g34 (n67, n15);
not  g35 (n52, n3);
not  g36 (n73, n1);
not  g37 (n54, n8);
not  g38 (n39, n17);
not  g39 (n68, n5);
not  g40 (n35, n16);
buf  g41 (n29, n2);
buf  g42 (n47, n11);
not  g43 (n46, n10);
not  g44 (n75, n15);
buf  g45 (n65, n11);
buf  g46 (n76, n18);
buf  g47 (n70, n16);
buf  g48 (n38, n14);
not  g49 (n57, n18);
buf  g50 (n50, n1);
not  g51 (n61, n15);
not  g52 (n49, n6);
not  g53 (n74, n17);
not  g54 (n83, n10);
buf  g55 (n58, n15);
buf  g56 (n165, n54);
buf  g57 (n116, n48);
not  g58 (n146, n51);
buf  g59 (n163, n31);
buf  g60 (n90, n29);
buf  g61 (n153, n39);
buf  g62 (n157, n47);
buf  g63 (n161, n54);
not  g64 (n105, n30);
not  g65 (n143, n65);
not  g66 (n117, n49);
not  g67 (n131, n34);
not  g68 (n127, n62);
not  g69 (n132, n45);
not  g70 (n122, n28);
buf  g71 (n98, n28);
buf  g72 (n108, n37);
buf  g73 (n151, n61);
buf  g74 (n104, n68);
buf  g75 (n130, n46);
buf  g76 (n112, n40);
not  g77 (n140, n50);
buf  g78 (n110, n39);
not  g79 (n92, n32);
buf  g80 (n152, n43);
buf  g81 (n135, n41);
buf  g82 (n111, n33);
buf  g83 (n102, n36);
not  g84 (n134, n48);
not  g85 (n148, n49);
not  g86 (n149, n37);
not  g87 (n89, n56);
buf  g88 (n100, n61);
not  g89 (n106, n44);
not  g90 (n164, n56);
not  g91 (n147, n67);
buf  g92 (n138, n58);
buf  g93 (n109, n57);
buf  g94 (n126, n57);
buf  g95 (n97, n32);
not  g96 (n136, n46);
not  g97 (n154, n30);
buf  g98 (n124, n58);
not  g99 (n119, n50);
buf  g100 (n128, n38);
not  g101 (n120, n45);
not  g102 (n145, n52);
not  g103 (n107, n38);
buf  g104 (n166, n62);
not  g105 (n142, n51);
not  g106 (n144, n42);
not  g107 (n88, n47);
buf  g108 (n101, n53);
not  g109 (n113, n33);
not  g110 (n133, n67);
buf  g111 (n159, n66);
buf  g112 (n94, n53);
buf  g113 (n118, n60);
buf  g114 (n91, n63);
not  g115 (n125, n63);
buf  g116 (n150, n55);
buf  g117 (n129, n64);
buf  g118 (n86, n41);
not  g119 (n121, n65);
buf  g120 (n160, n60);
buf  g121 (n84, n44);
not  g122 (n96, n42);
not  g123 (n85, n35);
buf  g124 (n162, n34);
buf  g125 (n115, n59);
buf  g126 (n99, n31);
not  g127 (n95, n64);
buf  g128 (n103, n36);
buf  g129 (n156, n35);
buf  g130 (n93, n68);
buf  g131 (n139, n55);
not  g132 (n155, n43);
not  g133 (n123, n52);
not  g134 (n158, n29);
buf  g135 (n137, n66);
not  g136 (n114, n40);
buf  g137 (n141, n69);
not  g138 (n87, n59);
not  g139 (n226, n98);
not  g140 (n237, n138);
buf  g141 (n173, n161);
not  g142 (n280, n127);
buf  g143 (n246, n150);
buf  g144 (n261, n144);
buf  g145 (n214, n87);
buf  g146 (n180, n120);
not  g147 (n232, n155);
not  g148 (n221, n140);
not  g149 (n259, n114);
not  g150 (n279, n99);
not  g151 (n270, n143);
not  g152 (n168, n90);
buf  g153 (n216, n111);
not  g154 (n217, n155);
not  g155 (n222, n147);
not  g156 (n231, n138);
buf  g157 (n182, n106);
not  g158 (n169, n117);
buf  g159 (n178, n151);
not  g160 (n273, n131);
buf  g161 (n204, n104);
buf  g162 (n252, n133);
buf  g163 (n256, n156);
not  g164 (n170, n136);
buf  g165 (n268, n153);
buf  g166 (n251, n159);
not  g167 (n236, n140);
not  g168 (n206, n154);
buf  g169 (n271, n148);
buf  g170 (n265, n159);
not  g171 (n275, n108);
not  g172 (n201, n84);
not  g173 (n192, n137);
buf  g174 (n185, n88);
not  g175 (n183, n96);
not  g176 (n200, n93);
not  g177 (n278, n103);
not  g178 (n228, n110);
not  g179 (n195, n142);
not  g180 (n172, n148);
not  g181 (n171, n163);
buf  g182 (n235, n121);
not  g183 (n197, n145);
not  g184 (n238, n131);
buf  g185 (n230, n154);
buf  g186 (n225, n136);
buf  g187 (n167, n134);
not  g188 (n220, n129);
buf  g189 (n277, n153);
not  g190 (n208, n132);
not  g191 (n244, n124);
not  g192 (n202, n123);
buf  g193 (n209, n145);
not  g194 (n219, n139);
buf  g195 (n207, n146);
buf  g196 (n218, n113);
not  g197 (n260, n132);
buf  g198 (n198, n150);
not  g199 (n240, n101);
not  g200 (n239, n107);
buf  g201 (n247, n149);
buf  g202 (n186, n160);
buf  g203 (n262, n133);
not  g204 (n263, n102);
buf  g205 (n176, n141);
not  g206 (n223, n152);
not  g207 (n210, n92);
not  g208 (n233, n128);
buf  g209 (n184, n105);
buf  g210 (n264, n85);
not  g211 (n224, n157);
buf  g212 (n242, n86);
buf  g213 (n199, n162);
buf  g214 (n211, n112);
not  g215 (n253, n95);
buf  g216 (n248, n158);
buf  g217 (n258, n118);
buf  g218 (n193, n100);
not  g219 (n241, n139);
buf  g220 (n205, n89);
not  g221 (n177, n97);
not  g222 (n203, n147);
buf  g223 (n255, n160);
not  g224 (n257, n134);
buf  g225 (n249, n149);
buf  g226 (n250, n161);
buf  g227 (n196, n130);
buf  g228 (n269, n157);
not  g229 (n266, n162);
not  g230 (n272, n91);
buf  g231 (n245, n125);
not  g232 (n175, n156);
not  g233 (n229, n116);
buf  g234 (n274, n122);
not  g235 (n189, n152);
buf  g236 (n190, n135);
buf  g237 (n234, n144);
not  g238 (n267, n126);
buf  g239 (n194, n130);
buf  g240 (n243, n151);
buf  g241 (n227, n115);
buf  g242 (n254, n119);
buf  g243 (n213, n109);
buf  g244 (n187, n135);
buf  g245 (n215, n141);
buf  g246 (n181, n143);
not  g247 (n276, n129);
not  g248 (n212, n142);
buf  g249 (n179, n146);
not  g250 (n174, n94);
not  g251 (n191, n158);
buf  g252 (n188, n137);
buf  g253 (n300, n168);
not  g254 (n289, n171);
buf  g255 (n292, n177);
not  g256 (n296, n176);
not  g257 (n291, n174);
not  g258 (n293, n169);
not  g259 (n282, n176);
not  g260 (n301, n175);
buf  g261 (n283, n170);
buf  g262 (n299, n171);
buf  g263 (n288, n169);
not  g264 (n298, n172);
buf  g265 (n297, n174);
not  g266 (n290, n168);
buf  g267 (n287, n175);
buf  g268 (n302, n167);
not  g269 (n285, n170);
buf  g270 (n294, n172);
buf  g271 (n295, n173);
buf  g272 (n286, n167);
not  g273 (n284, n173);
not  g274 (n281, n177);
not  g275 (n309, n292);
not  g276 (n315, n286);
not  g277 (n307, n285);
not  g278 (n311, n293);
buf  g279 (n305, n287);
not  g280 (n317, n291);
buf  g281 (n312, n281);
buf  g282 (n306, n296);
not  g283 (n308, n178);
buf  g284 (n304, n179);
nor  g285 (n310, n180, n294);
or   g286 (n314, n295, n282);
xnor g287 (n313, n288, n180);
xor  g288 (n316, n178, n179);
and  g289 (n303, n284, n283);
xnor g290 (n318, n290, n289);
not  g291 (n357, n307);
buf  g292 (n371, n318);
buf  g293 (n346, n306);
not  g294 (n339, n308);
buf  g295 (n323, n311);
buf  g296 (n364, n303);
buf  g297 (n335, n310);
buf  g298 (n324, n306);
not  g299 (n347, n312);
not  g300 (n329, n304);
buf  g301 (n328, n311);
buf  g302 (n320, n310);
buf  g303 (n340, n305);
not  g304 (n363, n314);
not  g305 (n350, n312);
buf  g306 (n369, n315);
not  g307 (n336, n307);
not  g308 (n334, n318);
buf  g309 (n337, n308);
buf  g310 (n360, n315);
buf  g311 (n368, n303);
not  g312 (n319, n314);
buf  g313 (n372, n303);
not  g314 (n355, n317);
buf  g315 (n365, n313);
not  g316 (n381, n304);
buf  g317 (n341, n313);
not  g318 (n327, n304);
buf  g319 (n378, n316);
buf  g320 (n366, n307);
buf  g321 (n353, n311);
not  g322 (n348, n305);
buf  g323 (n351, n314);
buf  g324 (n321, n313);
not  g325 (n343, n305);
buf  g326 (n332, n303);
not  g327 (n370, n317);
buf  g328 (n377, n316);
not  g329 (n326, n305);
buf  g330 (n349, n317);
not  g331 (n376, n306);
not  g332 (n345, n315);
buf  g333 (n359, n315);
not  g334 (n361, n312);
buf  g335 (n338, n308);
buf  g336 (n379, n314);
not  g337 (n367, n313);
not  g338 (n333, n308);
not  g339 (n322, n309);
not  g340 (n358, n317);
not  g341 (n352, n309);
buf  g342 (n342, n304);
not  g343 (n344, n307);
not  g344 (n375, n311);
not  g345 (n354, n312);
not  g346 (n374, n318);
buf  g347 (n380, n310);
not  g348 (n331, n309);
buf  g349 (n330, n310);
not  g350 (n373, n316);
buf  g351 (n325, n309);
not  g352 (n356, n306);
buf  g353 (n362, n316);
not  g354 (n393, n187);
buf  g355 (n415, n339);
not  g356 (n403, n344);
not  g357 (n390, n337);
buf  g358 (n417, n325);
buf  g359 (n407, n346);
buf  g360 (n401, n333);
not  g361 (n397, n331);
not  g362 (n414, n182);
not  g363 (n400, n193);
not  g364 (n394, n181);
buf  g365 (n416, n341);
buf  g366 (n404, n322);
buf  g367 (n385, n192);
buf  g368 (n413, n334);
not  g369 (n409, n335);
buf  g370 (n388, n186);
buf  g371 (n418, n352);
buf  g372 (n402, n330);
buf  g373 (n384, n345);
buf  g374 (n411, n338);
buf  g375 (n391, n323);
not  g376 (n386, n183);
not  g377 (n412, n343);
not  g378 (n383, n332);
buf  g379 (n382, n328);
buf  g380 (n408, n342);
not  g381 (n406, n192);
and  g382 (n395, n185, n326, n336);
nor  g383 (n398, n190, n340, n188, n182);
xnor g384 (n399, n354, n181, n187, n347);
xnor g385 (n410, n324, n190, n321, n185);
nor  g386 (n392, n355, n320, n191, n353);
xnor g387 (n389, n183, n184, n348, n188);
or   g388 (n405, n350, n319, n184, n329);
or   g389 (n387, n189, n191, n186, n327);
nand g390 (n396, n351, n189, n349, n193);
nand g391 (n429, n393, n24, n395, n394);
and  g392 (n452, n383, n297, n20, n399);
or   g393 (n444, n359, n378, n393, n398);
and  g394 (n435, n394, n22, n383);
nor  g395 (n433, n298, n367, n383, n392);
xnor g396 (n460, n383, n24, n358, n22);
xnor g397 (n441, n370, n26, n378, n364);
xor  g398 (n451, n26, n386, n362, n374);
nor  g399 (n456, n20, n21, n375, n376);
nor  g400 (n427, n363, n362, n396, n357);
and  g401 (n436, n25, n400, n377, n356);
or   g402 (n426, n392, n24, n373, n397);
nand g403 (n442, n21, n19, n360, n385);
and  g404 (n453, n389, n365, n397, n381);
xnor g405 (n458, n373, n23, n361, n385);
or   g406 (n421, n23, n398, n395, n25);
nor  g407 (n446, n24, n374, n392, n388);
and  g408 (n434, n388, n359, n20, n360);
nand g409 (n457, n391, n372, n198, n377);
nor  g410 (n430, n21, n384, n386, n26);
nor  g411 (n432, n387, n300, n381, n197);
xnor g412 (n455, n392, n197, n380, n379);
xnor g413 (n459, n387, n382, n21, n388);
xor  g414 (n439, n371, n389, n366, n368);
xor  g415 (n425, n194, n386, n363, n391);
xnor g416 (n419, n380, n26, n395, n25);
and  g417 (n447, n398, n399, n369, n384);
xnor g418 (n420, n23, n299, n391, n393);
xnor g419 (n454, n390, n364, n361, n393);
xor  g420 (n448, n382, n385, n375, n379);
and  g421 (n437, n23, n368, n196, n387);
nor  g422 (n428, n398, n195, n382, n390);
xor  g423 (n438, n365, n399, n386, n384);
xor  g424 (n449, n372, n397, n396);
nor  g425 (n440, n389, n196, n382, n390);
or   g426 (n450, n25, n376, n396, n399);
xor  g427 (n431, n389, n194, n367, n385);
or   g428 (n424, n19, n371, n384, n20);
xor  g429 (n423, n387, n400, n395, n394);
or   g430 (n422, n388, n369, n397, n22);
nand g431 (n445, n391, n366, n394, n370);
or   g432 (n443, n301, n390, n302, n195);
xnor g433 (n474, n412, n411, n437);
and  g434 (n469, n404, n405, n428, n400);
xnor g435 (n478, n408, n425, n405, n414);
nor  g436 (n483, n422, n405, n424, n403);
xor  g437 (n462, n414, n433, n420, n409);
nor  g438 (n475, n432, n411, n405, n409);
nor  g439 (n476, n401, n406, n418, n408);
nand g440 (n481, n409, n401, n418, n443);
nand g441 (n473, n415, n414, n416, n413);
nor  g442 (n463, n418, n415, n426, n404);
xor  g443 (n479, n403, n414, n415, n412);
or   g444 (n471, n417, n408, n402);
xor  g445 (n485, n407, n406, n401, n417);
nand g446 (n464, n439, n407, n431, n413);
or   g447 (n465, n412, n430, n409, n436);
nand g448 (n468, n403, n406, n412, n416);
xnor g449 (n484, n413, n417, n402, n408);
or   g450 (n470, n438, n442, n417, n418);
and  g451 (n466, n401, n429, n406, n404);
or   g452 (n480, n407, n403, n416, n421);
and  g453 (n467, n435, n400, n427, n419);
nor  g454 (n472, n434, n411, n407, n404);
xor  g455 (n461, n415, n410, n441, n423);
xnor g456 (n477, n410, n413, n440, n402);
or   g457 (n482, n410, n410, n416, n318);
buf  g458 (n507, n466);
buf  g459 (n508, n470);
not  g460 (n509, n468);
buf  g461 (n511, n463);
buf  g462 (n499, n470);
not  g463 (n501, n465);
buf  g464 (n498, n469);
buf  g465 (n503, n467);
not  g466 (n504, n466);
not  g467 (n487, n462);
buf  g468 (n506, n469);
not  g469 (n497, n461);
buf  g470 (n494, n462);
not  g471 (n505, n469);
not  g472 (n502, n469);
buf  g473 (n486, n464);
buf  g474 (n492, n468);
not  g475 (n496, n467);
not  g476 (n491, n464);
buf  g477 (n493, n463);
not  g478 (n510, n470);
not  g479 (n513, n468);
buf  g480 (n489, n471);
not  g481 (n495, n468);
buf  g482 (n514, n461);
buf  g483 (n490, n465);
not  g484 (n512, n471);
buf  g485 (n500, n470);
not  g486 (n488, n467);
not  g487 (n515, n486);
not  g488 (n522, n487);
buf  g489 (n518, n472);
buf  g490 (n520, n472);
buf  g491 (n526, n472);
buf  g492 (n525, n488);
buf  g493 (n516, n488);
not  g494 (n524, n471);
xor  g495 (n521, n487, n472, n473, n471);
xor  g496 (n523, n488, n487, n474);
xnor g497 (n519, n473, n486, n474);
nor  g498 (n517, n486, n473, n488);
not  g499 (n530, n496);
not  g500 (n549, n453);
not  g501 (n561, n496);
buf  g502 (n543, n449);
buf  g503 (n538, n448);
buf  g504 (n551, n454);
buf  g505 (n554, n494);
buf  g506 (n533, n444);
buf  g507 (n529, n200);
not  g508 (n536, n519);
buf  g509 (n558, n494);
xnor g510 (n539, n494, n520, n491);
xnor g511 (n531, n525, n451, n490, n515);
and  g512 (n528, n497, n498, n446, n526);
xor  g513 (n559, n202, n523, n492, n445);
nand g514 (n552, n201, n521, n497, n493);
or   g515 (n560, n492, n456, n491, n495);
xor  g516 (n556, n457, n526, n497, n490);
xnor g517 (n557, n517, n489, n518, n495);
or   g518 (n546, n497, n498, n525, n526);
nand g519 (n553, n522, n494, n499, n492);
nor  g520 (n555, n493, n496, n199, n489);
nand g521 (n542, n447, n490, n521, n523);
xor  g522 (n532, n199, n499, n524);
and  g523 (n540, n499, n459, n460, n455);
and  g524 (n535, n516, n452, n517, n492);
xnor g525 (n534, n493, n450, n521, n518);
nand g526 (n527, n496, n522, n198, n489);
or   g527 (n547, n163, n525, n515, n200);
xnor g528 (n548, n519, n491, n495, n516);
xnor g529 (n550, n522, n526, n491, n490);
and  g530 (n545, n498, n458, n164, n489);
xor  g531 (n541, n493, n524, n201, n498);
xor  g532 (n537, n495, n522, n523, n524);
nand g533 (n544, n523, n525, n520, n524);
not  g534 (n616, n551);
not  g535 (n585, n550);
not  g536 (n659, n530);
not  g537 (n603, n548);
not  g538 (n581, n531);
buf  g539 (n656, n550);
buf  g540 (n649, n534);
buf  g541 (n576, n529);
not  g542 (n650, n540);
not  g543 (n583, n531);
buf  g544 (n622, n547);
not  g545 (n634, n538);
buf  g546 (n580, n536);
buf  g547 (n567, n545);
buf  g548 (n600, n546);
not  g549 (n602, n551);
not  g550 (n609, n538);
not  g551 (n648, n547);
buf  g552 (n658, n538);
not  g553 (n593, n533);
not  g554 (n618, n543);
not  g555 (n575, n551);
buf  g556 (n662, n532);
not  g557 (n654, n534);
not  g558 (n570, n529);
buf  g559 (n626, n536);
buf  g560 (n646, n538);
buf  g561 (n571, n541);
not  g562 (n615, n528);
buf  g563 (n655, n550);
buf  g564 (n577, n547);
not  g565 (n630, n548);
buf  g566 (n610, n534);
buf  g567 (n617, n549);
not  g568 (n613, n527);
not  g569 (n606, n536);
not  g570 (n599, n544);
buf  g571 (n657, n530);
not  g572 (n574, n545);
buf  g573 (n564, n536);
buf  g574 (n627, n543);
buf  g575 (n637, n550);
buf  g576 (n601, n545);
buf  g577 (n647, n532);
not  g578 (n653, n544);
buf  g579 (n623, n546);
not  g580 (n628, n541);
not  g581 (n621, n546);
not  g582 (n652, n548);
buf  g583 (n586, n529);
buf  g584 (n639, n549);
buf  g585 (n596, n540);
not  g586 (n614, n537);
not  g587 (n632, n531);
buf  g588 (n578, n535);
buf  g589 (n619, n541);
buf  g590 (n631, n532);
buf  g591 (n604, n535);
not  g592 (n608, n530);
not  g593 (n591, n551);
buf  g594 (n629, n533);
buf  g595 (n565, n544);
buf  g596 (n611, n552);
buf  g597 (n612, n552);
buf  g598 (n638, n552);
not  g599 (n589, n535);
buf  g600 (n605, n549);
buf  g601 (n572, n537);
buf  g602 (n640, n534);
not  g603 (n663, n532);
not  g604 (n620, n528);
not  g605 (n592, n527);
buf  g606 (n562, n535);
buf  g607 (n598, n530);
buf  g608 (n666, n527);
not  g609 (n590, n533);
not  g610 (n587, n549);
not  g611 (n633, n541);
not  g612 (n642, n531);
not  g613 (n563, n540);
not  g614 (n569, n539);
not  g615 (n643, n547);
buf  g616 (n661, n542);
not  g617 (n597, n544);
not  g618 (n641, n528);
buf  g619 (n644, n529);
buf  g620 (n645, n540);
buf  g621 (n595, n537);
not  g622 (n636, n543);
not  g623 (n660, n539);
not  g624 (n566, n533);
buf  g625 (n573, n553);
buf  g626 (n624, n543);
not  g627 (n664, n537);
buf  g628 (n651, n553);
not  g629 (n568, n539);
not  g630 (n582, n528);
not  g631 (n625, n552);
buf  g632 (n667, n548);
buf  g633 (n607, n539);
not  g634 (n665, n545);
not  g635 (n588, n546);
buf  g636 (n635, n542);
buf  g637 (n579, n542);
buf  g638 (n594, n542);
buf  g639 (n584, n527);
xor  g640 (n683, n506, n503, n567, n589);
and  g641 (n677, n574, n507, n555, n483);
xor  g642 (n713, n561, n590, n508, n481);
or   g643 (n680, n556, n503, n513, n479);
xnor g644 (n711, n502, n511, n509, n481);
nand g645 (n679, n580, n594, n505, n586);
xor  g646 (n706, n553, n555, n481, n587);
nor  g647 (n712, n502, n582, n575, n506);
or   g648 (n696, n476, n561, n514, n502);
xor  g649 (n700, n563, n559, n478, n477);
xor  g650 (n707, n560, n484, n508, n581);
or   g651 (n715, n500, n582, n506, n556);
xnor g652 (n695, n558, n594, n482, n500);
xor  g653 (n716, n593, n511, n514, n508);
and  g654 (n694, n568, n588, n579, n505);
xor  g655 (n678, n554, n507, n592, n566);
or   g656 (n681, n564, n554, n583, n476);
and  g657 (n671, n480, n572, n514);
xnor g658 (n684, n513, n500, n571, n564);
and  g659 (n718, n596, n503, n482, n559);
and  g660 (n669, n595, n568, n475, n512);
nand g661 (n686, n569, n573, n559, n476);
xnor g662 (n688, n475, n567, n500, n509);
nand g663 (n697, n587, n584, n554, n575);
nand g664 (n672, n586, n477, n596, n505);
nor  g665 (n708, n565, n562, n555, n502);
nand g666 (n685, n565, n585, n501);
nor  g667 (n674, n510, n511, n479, n579);
xor  g668 (n670, n480, n510, n591, n474);
xor  g669 (n673, n513, n558, n504, n501);
nand g670 (n692, n503, n557, n569, n511);
nor  g671 (n668, n556, n580, n509, n584);
nand g672 (n710, n509, n475, n557, n478);
nand g673 (n717, n483, n560, n482, n504);
or   g674 (n702, n576, n570, n571, n513);
xnor g675 (n704, n572, n560, n581, n561);
nand g676 (n705, n480, n476, n478, n477);
xnor g677 (n693, n570, n501, n588, n477);
xor  g678 (n689, n597, n583, n557, n593);
nand g679 (n714, n504, n510, n589, n559);
or   g680 (n699, n563, n595, n482, n558);
nand g681 (n675, n590, n573, n562, n592);
and  g682 (n709, n507, n555, n557, n591);
xor  g683 (n703, n553, n556, n576, n479);
xnor g684 (n682, n566, n501, n483, n505);
xor  g685 (n687, n507, n474, n561, n578);
xnor g686 (n691, n574, n483, n554, n512);
xor  g687 (n701, n560, n475, n504, n480);
nor  g688 (n676, n479, n512, n577);
or   g689 (n690, n478, n506, n481, n510);
nor  g690 (n698, n578, n512, n508, n558);
buf  g691 (n732, n614);
buf  g692 (n722, n629);
buf  g693 (n745, n603);
buf  g694 (n749, n670);
not  g695 (n739, n676);
not  g696 (n734, n608);
nor  g697 (n741, n612, n679);
nor  g698 (n742, n626, n673);
xor  g699 (n748, n613, n598, n601, n612);
or   g700 (n747, n627, n610, n607, n680);
or   g701 (n736, n626, n621, n630, n676);
xor  g702 (n743, n674, n608, n675, n680);
or   g703 (n733, n633, n631, n617);
nand g704 (n738, n603, n670, n629, n617);
or   g705 (n724, n610, n619, n607, n621);
nor  g706 (n750, n683, n674, n679, n682);
nand g707 (n746, n598, n630, n616, n597);
xor  g708 (n740, n609, n611, n619, n615);
or   g709 (n731, n682, n620, n675, n611);
and  g710 (n726, n614, n622, n618, n623);
and  g711 (n728, n625, n681, n632, n620);
nor  g712 (n720, n605, n600, n623, n602);
xor  g713 (n729, n628, n599, n615, n678);
xor  g714 (n735, n668, n605, n613, n600);
or   g715 (n719, n632, n627, n672, n677);
nor  g716 (n730, n618, n606, n677, n683);
nand g717 (n744, n668, n624, n633, n681);
and  g718 (n727, n609, n602, n604);
xor  g719 (n725, n606, n625, n628, n624);
xnor g720 (n723, n634, n669, n601);
xor  g721 (n721, n672, n673, n671, n678);
nand g722 (n737, n622, n671, n616, n599);
or   g723 (n761, n686, n166, n690, n689);
nand g724 (n770, n717, n69, n699, n165);
xor  g725 (n778, n705, n734, n724, n728);
or   g726 (n756, n700, n73, n699, n712);
xnor g727 (n765, n705, n701, n725, n702);
and  g728 (n763, n695, n74, n720, n688);
or   g729 (n773, n72, n697, n691, n706);
and  g730 (n780, n716, n710, n687, n715);
xnor g731 (n753, n731, n693, n165, n716);
or   g732 (n766, n702, n733, n730, n732);
or   g733 (n759, n698, n719, n714, n703);
and  g734 (n768, n697, n701, n709, n691);
nand g735 (n775, n717, n685, n716, n729);
nand g736 (n769, n728, n717, n709, n712);
and  g737 (n777, n727, n726, n715, n692);
xnor g738 (n767, n733, n721, n723, n695);
nand g739 (n758, n70, n72, n696, n71);
nand g740 (n774, n75, n700, n694, n704);
xor  g741 (n757, n708, n715, n726, n75);
nor  g742 (n776, n729, n76, n720, n164);
nor  g743 (n755, n730, n71, n732, n684);
xnor g744 (n760, n722, n686, n711, n713);
and  g745 (n764, n689, n707, n714);
xnor g746 (n754, n74, n708, n713, n727);
nand g747 (n779, n723, n703, n719, n73);
xor  g748 (n771, n731, n684, n715, n724);
and  g749 (n772, n706, n711, n693, n70);
xnor g750 (n781, n704, n690, n77, n721);
and  g751 (n752, n687, n725, n698, n710);
xnor g752 (n751, n688, n76, n694, n716);
and  g753 (n762, n722, n685, n692, n696);
or   g754 (n786, n652, n646, n657, n662);
and  g755 (n791, n758, n637, n767, n660);
xor  g756 (n790, n635, n665, n765, n657);
xor  g757 (n796, n640, n766, n639, n666);
nand g758 (n802, n761, n650, n753, n653);
nand g759 (n800, n667, n648, n637, n764);
xnor g760 (n804, n649, n659, n634, n772);
xnor g761 (n782, n762, n754, n643, n647);
xnor g762 (n799, n771, n770, n642, n769);
nand g763 (n784, n773, n651, n645);
nand g764 (n789, n640, n203, n760, n755);
xnor g765 (n794, n661, n658, n756, n638);
xor  g766 (n787, n648, n636, n644, n752);
or   g767 (n801, n642, n653, n664, n655);
or   g768 (n785, n646, n661, n649, n757);
xnor g769 (n793, n656, n641, n659, n663);
nand g770 (n788, n638, n768, n654, n663);
xor  g771 (n783, n644, n660, n667, n647);
nand g772 (n795, n651, n639, n666, n662);
nand g773 (n792, n641, n202, n759, n665);
xnor g774 (n798, n664, n650, n751, n643);
nand g775 (n797, n636, n654, n656, n655);
and  g776 (n803, n635, n652, n763, n658);
not  g777 (n806, n790);
not  g778 (n811, n799);
buf  g779 (n832, n206);
buf  g780 (n825, n796);
buf  g781 (n808, n217);
not  g782 (n830, n206);
xor  g783 (n827, n782, n222, n212);
xnor g784 (n819, n799, n205, n220);
nor  g785 (n820, n803, n718, n222);
xor  g786 (n815, n792, n783, n785);
nand g787 (n833, n205, n804, n218);
and  g788 (n824, n804, n203, n798);
or   g789 (n821, n214, n204, n801);
or   g790 (n805, n214, n717, n786);
xor  g791 (n810, n212, n789, n718);
xnor g792 (n828, n224, n217, n207);
nor  g793 (n826, n221, n802, n223);
and  g794 (n813, n784, n213, n221);
xor  g795 (n823, n788, n223, n216);
xor  g796 (n829, n794, n215);
xor  g797 (n809, n787, n219, n216);
xnor g798 (n818, n718, n207, n209);
xor  g799 (n812, n213, n718, n219);
nand g800 (n817, n208, n802, n800);
or   g801 (n814, n791, n224, n220);
and  g802 (n807, n795, n793, n210);
or   g803 (n822, n204, n208, n218);
nand g804 (n834, n209, n800, n803);
nor  g805 (n816, n798, n797, n211);
nor  g806 (n831, n211, n210, n801);
xor  g807 (n837, n741, n747, n750, n746);
nor  g808 (n842, n739, n485, n814);
nor  g809 (n847, n747, n807, n739, n736);
xor  g810 (n839, n737, n748, n741);
xor  g811 (n835, n744, n740, n748, n742);
nand g812 (n852, n225, n806, n743, n739);
and  g813 (n843, n750, n741, n813, n738);
or   g814 (n849, n749, n735, n736);
nand g815 (n845, n735, n816, n815, n806);
nor  g816 (n841, n811, n748, n746);
nand g817 (n846, n737, n745, n750, n749);
nor  g818 (n857, n747, n742, n810, n485);
and  g819 (n856, n809, n742, n807, n808);
xnor g820 (n853, n745, n745, n735, n741);
nor  g821 (n844, n484, n809, n744, n746);
nor  g822 (n850, n739, n750, n747, n812);
or   g823 (n854, n738, n743, n484);
nand g824 (n840, n812, n735, n749, n745);
nor  g825 (n848, n808, n740, n737, n805);
or   g826 (n836, n811, n805, n749, n740);
nand g827 (n858, n814, n737, n484, n738);
xnor g828 (n855, n743, n742, n740, n736);
nand g829 (n838, n813, n744, n810);
xnor g830 (n851, n734, n815, n816, n738);
and  g831 (n927, n238, n826, n80, n835);
nor  g832 (n867, n250, n27, n274, n857);
or   g833 (n932, n270, n27, n278, n263);
and  g834 (n887, n230, n829, n855, n841);
nand g835 (n897, n854, n849, n842, n853);
or   g836 (n914, n853, n846, n280, n830);
nand g837 (n920, n832, n259, n827, n853);
or   g838 (n921, n79, n269, n240);
nand g839 (n869, n774, n265, n273, n827);
or   g840 (n915, n828, n852, n256, n260);
or   g841 (n879, n246, n276, n239, n258);
xor  g842 (n865, n819, n228, n241, n858);
nand g843 (n868, n849, n262, n858, n259);
xor  g844 (n931, n244, n279, n272, n858);
or   g845 (n859, n279, n850, n280);
nor  g846 (n878, n250, n280, n258, n271);
nor  g847 (n898, n839, n828, n779, n276);
and  g848 (n902, n232, n837, n236, n265);
nand g849 (n892, n261, n823, n852, n271);
xor  g850 (n910, n778, n81, n226, n266);
nor  g851 (n894, n855, n848, n825, n79);
xnor g852 (n895, n838, n242, n274, n260);
or   g853 (n901, n279, n264, n275, n278);
nor  g854 (n886, n822, n851, n857, n846);
nor  g855 (n900, n843, n237, n829, n239);
nor  g856 (n907, n848, n256, n244, n260);
xor  g857 (n871, n234, n272, n260, n840);
or   g858 (n875, n837, n280, n233, n817);
and  g859 (n924, n781, n836, n858, n818);
xnor g860 (n863, n266, n272, n234, n851);
xnor g861 (n872, n241, n845, n228, n245);
or   g862 (n870, n854, n255, n842, n833);
or   g863 (n899, n847, n819, n841, n817);
nand g864 (n905, n81, n830, n855, n836);
nor  g865 (n911, n261, n823, n263, n246);
nor  g866 (n874, n834, n275, n831);
or   g867 (n926, n826, n857, n251, n847);
xor  g868 (n888, n818, n277, n267, n851);
xor  g869 (n884, n267, n78, n856, n831);
or   g870 (n929, n236, n846, n258, n833);
xnor g871 (n873, n850, n852, n856, n263);
nor  g872 (n860, n845, n226, n248, n259);
and  g873 (n925, n242, n232, n265, n829);
or   g874 (n861, n843, n857, n279, n827);
xor  g875 (n866, n820, n251, n822, n845);
nand g876 (n885, n833, n776, n821, n249);
xor  g877 (n916, n267, n831, n834, n252);
nand g878 (n882, n854, n775, n832, n830);
nand g879 (n880, n276, n272, n267, n265);
xnor g880 (n919, n82, n273, n277, n485);
xor  g881 (n904, n270, n840, n238, n849);
xnor g882 (n889, n269, n273, n276, n253);
xor  g883 (n935, n832, n227, n835, n847);
or   g884 (n922, n247, n247, n263, n243);
and  g885 (n877, n231, n839, n824, n254);
nand g886 (n933, n821, n229, n853, n262);
nand g887 (n876, n845, n834, n233, n277);
xor  g888 (n923, n847, n848, n254);
xor  g889 (n893, n271, n257, n844, n824);
nor  g890 (n862, n838, n249, n849, n830);
and  g891 (n890, n844, n828, n237, n833);
or   g892 (n896, n227, n78, n266, n856);
nor  g893 (n903, n261, n245, n832, n225);
or   g894 (n930, n275, n780, n278, n268);
and  g895 (n909, n850, n264, n856, n844);
and  g896 (n934, n274, n80, n278, n820);
nand g897 (n928, n231, n229, n27, n855);
and  g898 (n891, n268, n262, n266, n827);
or   g899 (n883, n270, n230, n243, n852);
and  g900 (n881, n851, n264, n277, n252);
or   g901 (n908, n77, n235, n248, n271);
xnor g902 (n864, n269, n834, n828, n273);
and  g903 (n913, n846, n253, n264, n261);
xnor g904 (n918, n854, n262, n235, n829);
nor  g905 (n917, n274, n777, n831, n268);
or   g906 (n912, n825, n82, n268, n270);
and  g907 (n906, n255, n240, n257, n259);
not  g908 (n950, n869);
not  g909 (n936, n870);
buf  g910 (n961, n881);
buf  g911 (n938, n882);
buf  g912 (n946, n867);
buf  g913 (n941, n859);
not  g914 (n955, n880);
buf  g915 (n963, n885);
not  g916 (n965, n876);
buf  g917 (n943, n887);
not  g918 (n953, n872);
buf  g919 (n964, n886);
buf  g920 (n959, n862);
not  g921 (n962, n888);
not  g922 (n954, n863);
not  g923 (n958, n873);
not  g924 (n940, n884);
not  g925 (n945, n879);
buf  g926 (n957, n878);
buf  g927 (n949, n877);
not  g928 (n937, n860);
not  g929 (n942, n875);
buf  g930 (n951, n871);
buf  g931 (n947, n864);
buf  g932 (n960, n866);
buf  g933 (n944, n883);
buf  g934 (n948, n868);
buf  g935 (n952, n874);
buf  g936 (n956, n861);
not  g937 (n939, n865);
xnor g938 (n975, n936, n922, n895, n959);
xnor g939 (n987, n946, n907, n913, n957);
nor  g940 (n979, n960, n941, n942, n954);
xnor g941 (n973, n904, n936, n940, n950);
nor  g942 (n971, n940, n945, n960, n890);
or   g943 (n969, n910, n897, n937, n956);
and  g944 (n984, n908, n915, n921, n898);
nand g945 (n980, n949, n943, n942, n952);
and  g946 (n989, n953, n949, n914, n939);
xnor g947 (n966, n950, n961, n891, n901);
nand g948 (n974, n948, n954, n937, n945);
xor  g949 (n983, n951, n944, n946, n952);
and  g950 (n972, n959, n951, n903, n902);
and  g951 (n985, n938, n899, n959, n900);
xor  g952 (n970, n906, n919, n912, n961);
and  g953 (n967, n956, n959, n894, n917);
xnor g954 (n976, n916, n943, n960, n958);
or   g955 (n981, n958, n947, n905, n961);
and  g956 (n977, n939, n911, n918, n955);
nor  g957 (n968, n893, n892, n961, n944);
nand g958 (n982, n957, n889, n953, n941);
or   g959 (n978, n962, n920, n938, n947);
xnor g960 (n986, n948, n962, n958, n960);
and  g961 (n988, n955, n896, n958, n909);
or   g962 (n990, n988, n962, n963);
buf  g963 (n991, n990);
not  g964 (n992, n990);
xor  g965 (n993, n963, n992);
xnor g966 (n996, n964, n965, n963);
xnor g967 (n994, n965, n964);
nor  g968 (n995, n965, n993);
and  g969 (n997, n965, n964, n963, n993);
and  g970 (n1001, n934, n926, n931, n924);
nand g971 (n1000, n933, n83, n994);
or   g972 (n1003, n927, n995, n935, n27);
xnor g973 (n998, n923, n930, n997);
xor  g974 (n1002, n932, n929, n928, n996);
or   g975 (n999, n166, n996, n989, n925);
endmodule
