

module Stat_850_1638
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n545,
  n665,
  n664,
  n681,
  n689,
  n657,
  n666,
  n674,
  n672,
  n663,
  n662,
  n669,
  n694,
  n684,
  n690,
  n678,
  n685,
  n844,
  n841,
  n879,
  n878,
  n877
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n545;output n665;output n664;output n681;output n689;output n657;output n666;output n674;output n672;output n663;output n662;output n669;output n694;output n684;output n690;output n678;output n685;output n844;output n841;output n879;output n878;output n877;
  wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n658;wire n659;wire n660;wire n661;wire n667;wire n668;wire n670;wire n671;wire n673;wire n675;wire n676;wire n677;wire n679;wire n680;wire n682;wire n683;wire n686;wire n687;wire n688;wire n691;wire n692;wire n693;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n842;wire n843;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyNOTWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    n122,
    n28
  );


  buf
  g1
  (
    n42,
    n17
  );


  buf
  g2
  (
    n51,
    n12
  );


  buf
  g3
  (
    n114,
    n9
  );


  buf
  g4
  (
    n120,
    n16
  );


  not
  g5
  (
    n92,
    n1
  );


  not
  g6
  (
    n104,
    n28
  );


  buf
  g7
  (
    n128,
    n29
  );


  not
  g8
  (
    n80,
    n18
  );


  not
  g9
  (
    n60,
    n19
  );


  buf
  g10
  (
    n68,
    n22
  );


  not
  g11
  (
    n65,
    n29
  );


  not
  g12
  (
    n31,
    n12
  );


  buf
  g13
  (
    n102,
    n22
  );


  buf
  g14
  (
    n126,
    n26
  );


  not
  g15
  (
    n39,
    n11
  );


  buf
  g16
  (
    n100,
    n16
  );


  buf
  g17
  (
    n58,
    n10
  );


  not
  g18
  (
    n91,
    n13
  );


  buf
  g19
  (
    n124,
    n22
  );


  not
  g20
  (
    n106,
    n26
  );


  buf
  g21
  (
    n83,
    n25
  );


  buf
  g22
  (
    n136,
    n14
  );


  not
  g23
  (
    n73,
    n24
  );


  not
  g24
  (
    n86,
    n4
  );


  not
  g25
  (
    n57,
    n21
  );


  not
  g26
  (
    n129,
    n4
  );


  buf
  g27
  (
    n118,
    n19
  );


  buf
  g28
  (
    n112,
    n2
  );


  not
  g29
  (
    n137,
    n21
  );


  not
  g30
  (
    n109,
    n11
  );


  not
  g31
  (
    n99,
    n24
  );


  not
  g32
  (
    n139,
    n15
  );


  not
  g33
  (
    n33,
    n27
  );


  not
  g34
  (
    n79,
    n7
  );


  not
  g35
  (
    n37,
    n22
  );


  buf
  g36
  (
    n145,
    n4
  );


  not
  g37
  (
    n141,
    n1
  );


  buf
  g38
  (
    n101,
    n14
  );


  not
  g39
  (
    n96,
    n18
  );


  buf
  g40
  (
    n95,
    n17
  );


  not
  g41
  (
    n108,
    n4
  );


  buf
  g42
  (
    n135,
    n23
  );


  not
  g43
  (
    n64,
    n27
  );


  not
  g44
  (
    n40,
    n10
  );


  not
  g45
  (
    n63,
    n1
  );


  buf
  g46
  (
    n69,
    n16
  );


  buf
  g47
  (
    n82,
    n11
  );


  buf
  g48
  (
    KeyWire_0_13,
    n1
  );


  not
  g49
  (
    n75,
    n8
  );


  not
  g50
  (
    n130,
    n3
  );


  buf
  g51
  (
    n47,
    n8
  );


  buf
  g52
  (
    n94,
    n20
  );


  not
  g53
  (
    n132,
    n13
  );


  not
  g54
  (
    n105,
    n3
  );


  not
  g55
  (
    n133,
    n15
  );


  not
  g56
  (
    n35,
    n12
  );


  not
  g57
  (
    n54,
    n20
  );


  not
  g58
  (
    n61,
    n23
  );


  not
  g59
  (
    n134,
    n17
  );


  not
  g60
  (
    n76,
    n19
  );


  buf
  g61
  (
    n62,
    n29
  );


  not
  g62
  (
    n74,
    n12
  );


  buf
  g63
  (
    n113,
    n2
  );


  not
  g64
  (
    n87,
    n20
  );


  not
  g65
  (
    n119,
    n18
  );


  not
  g66
  (
    n89,
    n10
  );


  buf
  g67
  (
    n111,
    n3
  );


  not
  g68
  (
    n59,
    n24
  );


  buf
  g69
  (
    n78,
    n21
  );


  not
  g70
  (
    n121,
    n17
  );


  buf
  g71
  (
    n41,
    n7
  );


  buf
  g72
  (
    n45,
    n20
  );


  not
  g73
  (
    n127,
    n6
  );


  buf
  g74
  (
    n77,
    n23
  );


  buf
  g75
  (
    KeyWire_0_21,
    n28
  );


  buf
  g76
  (
    n53,
    n9
  );


  not
  g77
  (
    n34,
    n13
  );


  buf
  g78
  (
    n56,
    n18
  );


  buf
  g79
  (
    n71,
    n29
  );


  buf
  g80
  (
    n46,
    n7
  );


  buf
  g81
  (
    n98,
    n28
  );


  buf
  g82
  (
    n67,
    n9
  );


  buf
  g83
  (
    n103,
    n9
  );


  not
  g84
  (
    n97,
    n8
  );


  buf
  g85
  (
    n55,
    n15
  );


  not
  g86
  (
    n90,
    n6
  );


  not
  g87
  (
    n142,
    n21
  );


  buf
  g88
  (
    n123,
    n15
  );


  not
  g89
  (
    KeyWire_0_50,
    n6
  );


  buf
  g90
  (
    n52,
    n16
  );


  buf
  g91
  (
    n38,
    n23
  );


  buf
  g92
  (
    n70,
    n13
  );


  not
  g93
  (
    n36,
    n7
  );


  buf
  g94
  (
    n110,
    n25
  );


  not
  g95
  (
    n88,
    n14
  );


  buf
  g96
  (
    KeyWire_0_55,
    n25
  );


  not
  g97
  (
    n43,
    n10
  );


  not
  g98
  (
    n50,
    n2
  );


  not
  g99
  (
    n84,
    n6
  );


  not
  g100
  (
    n30,
    n26
  );


  buf
  g101
  (
    n48,
    n5
  );


  buf
  g102
  (
    KeyWire_0_26,
    n19
  );


  buf
  g103
  (
    n138,
    n24
  );


  not
  g104
  (
    n66,
    n25
  );


  buf
  g105
  (
    n44,
    n11
  );


  not
  g106
  (
    n81,
    n5
  );


  not
  g107
  (
    n107,
    n27
  );


  not
  g108
  (
    n85,
    n2
  );


  not
  g109
  (
    n72,
    n3
  );


  buf
  g110
  (
    n125,
    n27
  );


  buf
  g111
  (
    n115,
    n26
  );


  buf
  g112
  (
    n140,
    n14
  );


  not
  g113
  (
    n93,
    n5
  );


  not
  g114
  (
    n117,
    n5
  );


  not
  g115
  (
    n116,
    n8
  );


  buf
  g116
  (
    n264,
    n85
  );


  not
  g117
  (
    n504,
    n46
  );


  not
  g118
  (
    n290,
    n65
  );


  buf
  g119
  (
    n278,
    n136
  );


  not
  g120
  (
    n425,
    n126
  );


  buf
  g121
  (
    KeyWire_0_1,
    n63
  );


  not
  g122
  (
    n353,
    n48
  );


  buf
  g123
  (
    n246,
    n120
  );


  not
  g124
  (
    n429,
    n55
  );


  buf
  g125
  (
    n177,
    n70
  );


  not
  g126
  (
    n398,
    n94
  );


  buf
  g127
  (
    n159,
    n71
  );


  not
  g128
  (
    n415,
    n34
  );


  buf
  g129
  (
    KeyWire_0_33,
    n118
  );


  buf
  g130
  (
    n265,
    n31
  );


  buf
  g131
  (
    n389,
    n90
  );


  buf
  g132
  (
    n288,
    n42
  );


  buf
  g133
  (
    n251,
    n132
  );


  buf
  g134
  (
    n487,
    n54
  );


  buf
  g135
  (
    n303,
    n92
  );


  buf
  g136
  (
    n319,
    n107
  );


  not
  g137
  (
    n191,
    n106
  );


  buf
  g138
  (
    n181,
    n64
  );


  not
  g139
  (
    n481,
    n114
  );


  buf
  g140
  (
    n395,
    n52
  );


  not
  g141
  (
    n227,
    n71
  );


  buf
  g142
  (
    n205,
    n89
  );


  not
  g143
  (
    n493,
    n120
  );


  buf
  g144
  (
    n506,
    n76
  );


  not
  g145
  (
    n318,
    n44
  );


  buf
  g146
  (
    n469,
    n82
  );


  buf
  g147
  (
    n369,
    n42
  );


  not
  g148
  (
    n382,
    n131
  );


  buf
  g149
  (
    n234,
    n115
  );


  not
  g150
  (
    n189,
    n47
  );


  buf
  g151
  (
    n454,
    n126
  );


  buf
  g152
  (
    KeyWire_0_54,
    n108
  );


  buf
  g153
  (
    n414,
    n36
  );


  not
  g154
  (
    n341,
    n83
  );


  buf
  g155
  (
    n249,
    n120
  );


  buf
  g156
  (
    n151,
    n79
  );


  buf
  g157
  (
    n476,
    n96
  );


  buf
  g158
  (
    KeyWire_0_22,
    n108
  );


  buf
  g159
  (
    n295,
    n85
  );


  buf
  g160
  (
    n328,
    n115
  );


  buf
  g161
  (
    n445,
    n65
  );


  not
  g162
  (
    n148,
    n45
  );


  not
  g163
  (
    n453,
    n69
  );


  not
  g164
  (
    n326,
    n135
  );


  buf
  g165
  (
    n195,
    n133
  );


  buf
  g166
  (
    n464,
    n56
  );


  buf
  g167
  (
    n339,
    n31
  );


  buf
  g168
  (
    n233,
    n97
  );


  not
  g169
  (
    n491,
    n40
  );


  not
  g170
  (
    n173,
    n113
  );


  buf
  g171
  (
    n505,
    n109
  );


  not
  g172
  (
    n309,
    n123
  );


  not
  g173
  (
    n291,
    n70
  );


  buf
  g174
  (
    n252,
    n101
  );


  buf
  g175
  (
    n190,
    n134
  );


  buf
  g176
  (
    n242,
    n88
  );


  not
  g177
  (
    n200,
    n129
  );


  buf
  g178
  (
    n374,
    n110
  );


  buf
  g179
  (
    n272,
    n61
  );


  buf
  g180
  (
    n457,
    n98
  );


  buf
  g181
  (
    KeyWire_0_39,
    n131
  );


  buf
  g182
  (
    n243,
    n49
  );


  buf
  g183
  (
    n416,
    n123
  );


  buf
  g184
  (
    n178,
    n136
  );


  buf
  g185
  (
    n510,
    n122
  );


  not
  g186
  (
    n312,
    n58
  );


  buf
  g187
  (
    n381,
    n122
  );


  not
  g188
  (
    n509,
    n33
  );


  buf
  g189
  (
    n495,
    n30
  );


  not
  g190
  (
    n376,
    n38
  );


  buf
  g191
  (
    n314,
    n95
  );


  buf
  g192
  (
    n410,
    n130
  );


  buf
  g193
  (
    KeyWire_0_60,
    n69
  );


  buf
  g194
  (
    n462,
    n117
  );


  buf
  g195
  (
    n490,
    n125
  );


  buf
  g196
  (
    n322,
    n131
  );


  buf
  g197
  (
    n473,
    n38
  );


  not
  g198
  (
    n474,
    n88
  );


  buf
  g199
  (
    n332,
    n121
  );


  not
  g200
  (
    n176,
    n67
  );


  buf
  g201
  (
    n180,
    n80
  );


  not
  g202
  (
    KeyWire_0_51,
    n73
  );


  not
  g203
  (
    n185,
    n45
  );


  buf
  g204
  (
    n241,
    n68
  );


  not
  g205
  (
    n197,
    n109
  );


  buf
  g206
  (
    n406,
    n75
  );


  buf
  g207
  (
    n432,
    n136
  );


  buf
  g208
  (
    n373,
    n53
  );


  buf
  g209
  (
    n263,
    n57
  );


  buf
  g210
  (
    n239,
    n69
  );


  not
  g211
  (
    n289,
    n118
  );


  buf
  g212
  (
    n400,
    n74
  );


  buf
  g213
  (
    n350,
    n114
  );


  not
  g214
  (
    n223,
    n142
  );


  not
  g215
  (
    KeyWire_0_5,
    n102
  );


  not
  g216
  (
    n359,
    n82
  );


  not
  g217
  (
    n270,
    n59
  );


  buf
  g218
  (
    n431,
    n104
  );


  not
  g219
  (
    n346,
    n44
  );


  buf
  g220
  (
    n340,
    n75
  );


  buf
  g221
  (
    n379,
    n76
  );


  buf
  g222
  (
    n163,
    n124
  );


  not
  g223
  (
    n330,
    n122
  );


  not
  g224
  (
    n167,
    n135
  );


  buf
  g225
  (
    n160,
    n81
  );


  buf
  g226
  (
    KeyWire_0_34,
    n102
  );


  not
  g227
  (
    n372,
    n45
  );


  buf
  g228
  (
    n394,
    n131
  );


  buf
  g229
  (
    n286,
    n83
  );


  buf
  g230
  (
    KeyWire_0_31,
    n108
  );


  buf
  g231
  (
    n370,
    n35
  );


  buf
  g232
  (
    n184,
    n97
  );


  not
  g233
  (
    n323,
    n91
  );


  buf
  g234
  (
    n337,
    n77
  );


  buf
  g235
  (
    n217,
    n63
  );


  not
  g236
  (
    n214,
    n70
  );


  buf
  g237
  (
    n298,
    n95
  );


  not
  g238
  (
    n203,
    n55
  );


  buf
  g239
  (
    n480,
    n30
  );


  not
  g240
  (
    n364,
    n135
  );


  buf
  g241
  (
    KeyWire_0_45,
    n44
  );


  buf
  g242
  (
    n206,
    n60
  );


  buf
  g243
  (
    n231,
    n112
  );


  buf
  g244
  (
    n164,
    n99
  );


  buf
  g245
  (
    n449,
    n80
  );


  not
  g246
  (
    n393,
    n119
  );


  not
  g247
  (
    n236,
    n110
  );


  not
  g248
  (
    n418,
    n31
  );


  buf
  g249
  (
    n315,
    n130
  );


  buf
  g250
  (
    n402,
    n40
  );


  buf
  g251
  (
    n198,
    n55
  );


  buf
  g252
  (
    n501,
    n72
  );


  buf
  g253
  (
    n477,
    n49
  );


  not
  g254
  (
    n237,
    n138
  );


  buf
  g255
  (
    n489,
    n32
  );


  buf
  g256
  (
    n363,
    n139
  );


  buf
  g257
  (
    n256,
    n112
  );


  not
  g258
  (
    n301,
    n95
  );


  buf
  g259
  (
    n387,
    n101
  );


  not
  g260
  (
    n209,
    n77
  );


  not
  g261
  (
    n368,
    n140
  );


  buf
  g262
  (
    n225,
    n117
  );


  not
  g263
  (
    n348,
    n137
  );


  not
  g264
  (
    n448,
    n116
  );


  buf
  g265
  (
    n169,
    n94
  );


  not
  g266
  (
    n497,
    n129
  );


  not
  g267
  (
    n150,
    n104
  );


  not
  g268
  (
    n193,
    n129
  );


  not
  g269
  (
    n441,
    n74
  );


  buf
  g270
  (
    n170,
    n138
  );


  buf
  g271
  (
    n187,
    n127
  );


  not
  g272
  (
    n384,
    n84
  );


  not
  g273
  (
    n212,
    n58
  );


  buf
  g274
  (
    n321,
    n57
  );


  buf
  g275
  (
    n333,
    n139
  );


  not
  g276
  (
    n267,
    n114
  );


  buf
  g277
  (
    KeyWire_0_56,
    n51
  );


  not
  g278
  (
    n467,
    n47
  );


  buf
  g279
  (
    n349,
    n59
  );


  buf
  g280
  (
    n335,
    n32
  );


  not
  g281
  (
    n463,
    n140
  );


  not
  g282
  (
    n262,
    n66
  );


  buf
  g283
  (
    n213,
    n90
  );


  not
  g284
  (
    n443,
    n124
  );


  buf
  g285
  (
    n275,
    n60
  );


  not
  g286
  (
    n354,
    n93
  );


  not
  g287
  (
    n345,
    n86
  );


  buf
  g288
  (
    n343,
    n54
  );


  buf
  g289
  (
    n451,
    n87
  );


  buf
  g290
  (
    n274,
    n118
  );


  not
  g291
  (
    n488,
    n110
  );


  buf
  g292
  (
    n404,
    n105
  );


  buf
  g293
  (
    n156,
    n141
  );


  not
  g294
  (
    n292,
    n39
  );


  buf
  g295
  (
    n498,
    n119
  );


  buf
  g296
  (
    n287,
    n135
  );


  buf
  g297
  (
    n468,
    n66
  );


  buf
  g298
  (
    n413,
    n93
  );


  buf
  g299
  (
    n500,
    n98
  );


  buf
  g300
  (
    n316,
    n88
  );


  buf
  g301
  (
    n279,
    n121
  );


  buf
  g302
  (
    n153,
    n50
  );


  buf
  g303
  (
    n260,
    n133
  );


  buf
  g304
  (
    n157,
    n121
  );


  buf
  g305
  (
    n507,
    n92
  );


  buf
  g306
  (
    n307,
    n128
  );


  not
  g307
  (
    n365,
    n79
  );


  not
  g308
  (
    n380,
    n125
  );


  buf
  g309
  (
    n434,
    n41
  );


  not
  g310
  (
    KeyWire_0_27,
    n46
  );


  buf
  g311
  (
    n494,
    n37
  );


  buf
  g312
  (
    n229,
    n113
  );


  not
  g313
  (
    n149,
    n125
  );


  not
  g314
  (
    n447,
    n106
  );


  not
  g315
  (
    n317,
    n123
  );


  not
  g316
  (
    n427,
    n129
  );


  not
  g317
  (
    n304,
    n81
  );


  not
  g318
  (
    n329,
    n43
  );


  buf
  g319
  (
    KeyWire_0_24,
    n91
  );


  not
  g320
  (
    n168,
    n89
  );


  not
  g321
  (
    n503,
    n72
  );


  not
  g322
  (
    n492,
    n97
  );


  not
  g323
  (
    KeyWire_0_36,
    n81
  );


  buf
  g324
  (
    n285,
    n62
  );


  not
  g325
  (
    n352,
    n122
  );


  not
  g326
  (
    n155,
    n102
  );


  not
  g327
  (
    n201,
    n52
  );


  not
  g328
  (
    n331,
    n37
  );


  not
  g329
  (
    n338,
    n126
  );


  buf
  g330
  (
    n367,
    n132
  );


  buf
  g331
  (
    KeyWire_0_29,
    n53
  );


  not
  g332
  (
    KeyWire_0_49,
    n92
  );


  buf
  g333
  (
    n261,
    n46
  );


  not
  g334
  (
    n228,
    n30
  );


  buf
  g335
  (
    n158,
    n127
  );


  buf
  g336
  (
    n479,
    n130
  );


  buf
  g337
  (
    n240,
    n141
  );


  buf
  g338
  (
    n302,
    n68
  );


  buf
  g339
  (
    n421,
    n104
  );


  buf
  g340
  (
    n409,
    n67
  );


  not
  g341
  (
    n356,
    n39
  );


  not
  g342
  (
    n280,
    n60
  );


  not
  g343
  (
    n255,
    n36
  );


  not
  g344
  (
    n433,
    n123
  );


  buf
  g345
  (
    n147,
    n93
  );


  buf
  g346
  (
    n483,
    n96
  );


  not
  g347
  (
    n269,
    n43
  );


  not
  g348
  (
    n336,
    n134
  );


  not
  g349
  (
    n375,
    n107
  );


  buf
  g350
  (
    n162,
    n119
  );


  buf
  g351
  (
    n388,
    n140
  );


  buf
  g352
  (
    n161,
    n53
  );


  buf
  g353
  (
    n440,
    n94
  );


  buf
  g354
  (
    n397,
    n67
  );


  not
  g355
  (
    n324,
    n106
  );


  not
  g356
  (
    n320,
    n115
  );


  not
  g357
  (
    n423,
    n51
  );


  buf
  g358
  (
    KeyWire_0_46,
    n49
  );


  buf
  g359
  (
    n276,
    n57
  );


  not
  g360
  (
    n230,
    n139
  );


  not
  g361
  (
    n299,
    n120
  );


  buf
  g362
  (
    n412,
    n117
  );


  not
  g363
  (
    n424,
    n62
  );


  buf
  g364
  (
    n253,
    n87
  );


  not
  g365
  (
    n199,
    n119
  );


  buf
  g366
  (
    n186,
    n124
  );


  buf
  g367
  (
    n419,
    n68
  );


  not
  g368
  (
    n254,
    n134
  );


  buf
  g369
  (
    n293,
    n76
  );


  buf
  g370
  (
    n436,
    n33
  );


  buf
  g371
  (
    n460,
    n133
  );


  buf
  g372
  (
    n407,
    n124
  );


  buf
  g373
  (
    n238,
    n113
  );


  buf
  g374
  (
    n439,
    n118
  );


  buf
  g375
  (
    n207,
    n87
  );


  not
  g376
  (
    KeyWire_0_41,
    n99
  );


  not
  g377
  (
    n386,
    n130
  );


  buf
  g378
  (
    n216,
    n58
  );


  buf
  g379
  (
    n311,
    n117
  );


  buf
  g380
  (
    n461,
    n34
  );


  buf
  g381
  (
    n366,
    n63
  );


  buf
  g382
  (
    n174,
    n100
  );


  buf
  g383
  (
    n371,
    n139
  );


  not
  g384
  (
    KeyWire_0_8,
    n62
  );


  buf
  g385
  (
    n358,
    n71
  );


  buf
  g386
  (
    n456,
    n132
  );


  buf
  g387
  (
    n484,
    n43
  );


  buf
  g388
  (
    n188,
    n54
  );


  not
  g389
  (
    KeyWire_0_11,
    n78
  );


  not
  g390
  (
    n172,
    n100
  );


  not
  g391
  (
    n259,
    n75
  );


  not
  g392
  (
    n417,
    n48
  );


  not
  g393
  (
    n245,
    n132
  );


  buf
  g394
  (
    n194,
    n73
  );


  not
  g395
  (
    n152,
    n116
  );


  buf
  g396
  (
    n486,
    n84
  );


  not
  g397
  (
    n266,
    n37
  );


  not
  g398
  (
    n478,
    n34
  );


  buf
  g399
  (
    n257,
    n86
  );


  not
  g400
  (
    n277,
    n61
  );


  not
  g401
  (
    n235,
    n128
  );


  buf
  g402
  (
    KeyWire_0_48,
    n61
  );


  buf
  g403
  (
    n232,
    n64
  );


  buf
  g404
  (
    n472,
    n133
  );


  buf
  g405
  (
    n396,
    n66
  );


  buf
  g406
  (
    n357,
    n138
  );


  not
  g407
  (
    KeyWire_0_57,
    n115
  );


  not
  g408
  (
    n175,
    n36
  );


  not
  g409
  (
    n401,
    n48
  );


  not
  g410
  (
    n281,
    n89
  );


  not
  g411
  (
    n306,
    n134
  );


  not
  g412
  (
    n248,
    n83
  );


  buf
  g413
  (
    n247,
    n73
  );


  not
  g414
  (
    n452,
    n111
  );


  buf
  g415
  (
    n378,
    n126
  );


  buf
  g416
  (
    n385,
    n82
  );


  not
  g417
  (
    n210,
    n41
  );


  buf
  g418
  (
    n344,
    n113
  );


  buf
  g419
  (
    KeyWire_0_18,
    n33
  );


  buf
  g420
  (
    n196,
    n127
  );


  buf
  g421
  (
    n165,
    n112
  );


  not
  g422
  (
    n446,
    n105
  );


  not
  g423
  (
    KeyWire_0_16,
    n136
  );


  buf
  g424
  (
    n296,
    n99
  );


  not
  g425
  (
    n218,
    n74
  );


  buf
  g426
  (
    n399,
    n77
  );


  buf
  g427
  (
    n300,
    n65
  );


  not
  g428
  (
    n171,
    n128
  );


  not
  g429
  (
    n244,
    n35
  );


  buf
  g430
  (
    n466,
    n56
  );


  not
  g431
  (
    n166,
    n42
  );


  buf
  g432
  (
    n405,
    n107
  );


  buf
  g433
  (
    n475,
    n103
  );


  buf
  g434
  (
    n283,
    n116
  );


  not
  g435
  (
    n146,
    n56
  );


  buf
  g436
  (
    n438,
    n100
  );


  buf
  g437
  (
    n362,
    n137
  );


  not
  g438
  (
    n297,
    n35
  );


  not
  g439
  (
    n511,
    n103
  );


  buf
  g440
  (
    n271,
    n137
  );


  buf
  g441
  (
    n284,
    n78
  );


  buf
  g442
  (
    n435,
    n32
  );


  not
  g443
  (
    n360,
    n86
  );


  not
  g444
  (
    KeyWire_0_44,
    n98
  );


  not
  g445
  (
    n208,
    n39
  );


  not
  g446
  (
    n294,
    n51
  );


  not
  g447
  (
    n221,
    n91
  );


  not
  g448
  (
    n377,
    n41
  );


  not
  g449
  (
    n430,
    n138
  );


  not
  g450
  (
    n222,
    n111
  );


  not
  g451
  (
    n282,
    n50
  );


  not
  g452
  (
    n444,
    n114
  );


  buf
  g453
  (
    n342,
    n101
  );


  buf
  g454
  (
    n459,
    n78
  );


  not
  g455
  (
    n420,
    n137
  );


  buf
  g456
  (
    n391,
    n127
  );


  buf
  g457
  (
    KeyWire_0_40,
    n38
  );


  buf
  g458
  (
    n471,
    n141
  );


  buf
  g459
  (
    n458,
    n40
  );


  not
  g460
  (
    KeyWire_0_6,
    n103
  );


  buf
  g461
  (
    n403,
    n96
  );


  buf
  g462
  (
    n183,
    n90
  );


  buf
  g463
  (
    n392,
    n141
  );


  buf
  g464
  (
    n224,
    n52
  );


  not
  g465
  (
    n465,
    n116
  );


  buf
  g466
  (
    n334,
    n47
  );


  not
  g467
  (
    n154,
    n85
  );


  buf
  g468
  (
    n211,
    n84
  );


  not
  g469
  (
    n499,
    n121
  );


  not
  g470
  (
    n426,
    n64
  );


  not
  g471
  (
    n250,
    n79
  );


  not
  g472
  (
    n202,
    n111
  );


  buf
  g473
  (
    KeyWire_0_58,
    n140
  );


  not
  g474
  (
    n182,
    n72
  );


  buf
  g475
  (
    n361,
    n109
  );


  buf
  g476
  (
    n437,
    n80
  );


  not
  g477
  (
    n485,
    n125
  );


  buf
  g478
  (
    n422,
    n50
  );


  not
  g479
  (
    n204,
    n59
  );


  buf
  g480
  (
    n220,
    n105
  );


  not
  g481
  (
    n390,
    n128
  );


  not
  g482
  (
    n545,
    n167
  );


  buf
  g483
  (
    n527,
    n196
  );


  buf
  g484
  (
    n513,
    n172
  );


  not
  g485
  (
    n546,
    n168
  );


  not
  g486
  (
    n535,
    n193
  );


  not
  g487
  (
    n559,
    n184
  );


  buf
  g488
  (
    n549,
    n199
  );


  not
  g489
  (
    n518,
    n175
  );


  buf
  g490
  (
    n548,
    n142
  );


  buf
  g491
  (
    n539,
    n169
  );


  buf
  g492
  (
    n567,
    n143
  );


  not
  g493
  (
    n525,
    n194
  );


  buf
  g494
  (
    n515,
    n173
  );


  buf
  g495
  (
    n514,
    n182
  );


  not
  g496
  (
    n555,
    n177
  );


  buf
  g497
  (
    n537,
    n180
  );


  not
  g498
  (
    n544,
    n202
  );


  buf
  g499
  (
    n516,
    n156
  );


  not
  g500
  (
    n566,
    n197
  );


  buf
  g501
  (
    n521,
    n149
  );


  buf
  g502
  (
    n531,
    n178
  );


  buf
  g503
  (
    n520,
    n148
  );


  buf
  g504
  (
    n526,
    n166
  );


  not
  g505
  (
    n551,
    n170
  );


  buf
  g506
  (
    n530,
    n174
  );


  not
  g507
  (
    n556,
    n151
  );


  not
  g508
  (
    n542,
    n162
  );


  buf
  g509
  (
    n558,
    n154
  );


  not
  g510
  (
    n568,
    n160
  );


  not
  g511
  (
    n543,
    n181
  );


  not
  g512
  (
    n565,
    n143
  );


  not
  g513
  (
    n561,
    n147
  );


  not
  g514
  (
    n560,
    n150
  );


  buf
  g515
  (
    n528,
    n155
  );


  buf
  g516
  (
    n557,
    n157
  );


  buf
  g517
  (
    n529,
    n189
  );


  not
  g518
  (
    n533,
    n195
  );


  not
  g519
  (
    n519,
    n158
  );


  buf
  g520
  (
    n540,
    n171
  );


  not
  g521
  (
    n512,
    n163
  );


  not
  g522
  (
    KeyWire_0_42,
    n142
  );


  not
  g523
  (
    n562,
    n143
  );


  buf
  g524
  (
    n547,
    n165
  );


  not
  g525
  (
    n536,
    n153
  );


  buf
  g526
  (
    n523,
    n191
  );


  buf
  g527
  (
    KeyWire_0_47,
    n190
  );


  not
  g528
  (
    n563,
    n187
  );


  buf
  g529
  (
    n524,
    n159
  );


  buf
  g530
  (
    n517,
    n146
  );


  not
  g531
  (
    n532,
    n176
  );


  not
  g532
  (
    n552,
    n200
  );


  not
  g533
  (
    n541,
    n185
  );


  not
  g534
  (
    n553,
    n201
  );


  not
  g535
  (
    n538,
    n186
  );


  buf
  g536
  (
    n534,
    n152
  );


  xor
  g537
  (
    n522,
    n198,
    n142,
    n183,
    n164
  );


  nor
  g538
  (
    n564,
    n192,
    n161,
    n179,
    n188
  );


  or
  g539
  (
    n584,
    n293,
    n266,
    n344,
    n352
  );


  nor
  g540
  (
    n605,
    n526,
    n279,
    n231,
    n304
  );


  and
  g541
  (
    n610,
    n283,
    n312,
    n285,
    n214
  );


  nand
  g542
  (
    n595,
    n558,
    n237,
    n289,
    n358
  );


  and
  g543
  (
    n620,
    n338,
    n353,
    n333,
    n342
  );


  xnor
  g544
  (
    n613,
    n223,
    n367,
    n291,
    n315
  );


  and
  g545
  (
    KeyWire_0_43,
    n259,
    n528,
    n356,
    n542
  );


  xnor
  g546
  (
    n573,
    n539,
    n536,
    n242,
    n300
  );


  xor
  g547
  (
    n621,
    n343,
    n271,
    n205,
    n560
  );


  xnor
  g548
  (
    KeyWire_0_53,
    n238,
    n253,
    n233,
    n221
  );


  nand
  g549
  (
    n600,
    n217,
    n545,
    n518,
    n227
  );


  or
  g550
  (
    KeyWire_0_0,
    n296,
    n257,
    n243,
    n314
  );


  xnor
  g551
  (
    n570,
    n555,
    n287,
    n282,
    n290
  );


  nand
  g552
  (
    n577,
    n360,
    n345,
    n224,
    n340
  );


  nor
  g553
  (
    n611,
    n322,
    n361,
    n218,
    n260
  );


  and
  g554
  (
    n585,
    n341,
    n335,
    n543,
    n363
  );


  xor
  g555
  (
    n624,
    n359,
    n349,
    n562,
    n228
  );


  nand
  g556
  (
    n598,
    n209,
    n294,
    n225,
    n522
  );


  nor
  g557
  (
    n616,
    n313,
    n521,
    n557,
    n255
  );


  nor
  g558
  (
    n578,
    n258,
    n531,
    n321,
    n339
  );


  nand
  g559
  (
    n575,
    n320,
    n541,
    n272,
    n229
  );


  xor
  g560
  (
    n581,
    n206,
    n203,
    n527,
    n309
  );


  nor
  g561
  (
    n576,
    n368,
    n537,
    n327,
    n216
  );


  xor
  g562
  (
    n604,
    n547,
    n311,
    n269,
    n292
  );


  nor
  g563
  (
    n612,
    n324,
    n204,
    n317,
    n332
  );


  nand
  g564
  (
    n582,
    n535,
    n240,
    n355,
    n236
  );


  nor
  g565
  (
    n607,
    n303,
    n346,
    n328,
    n370
  );


  xor
  g566
  (
    n571,
    n251,
    n334,
    n366,
    n515
  );


  and
  g567
  (
    n569,
    n273,
    n220,
    n230,
    n530
  );


  or
  g568
  (
    n579,
    n210,
    n533,
    n544,
    n365
  );


  nand
  g569
  (
    n617,
    n245,
    n263,
    n329,
    n532
  );


  nand
  g570
  (
    n590,
    n278,
    n280,
    n553,
    n241
  );


  nor
  g571
  (
    n586,
    n323,
    n554,
    n252,
    n523
  );


  nor
  g572
  (
    n588,
    n548,
    n564,
    n219,
    n288
  );


  nor
  g573
  (
    n574,
    n212,
    n546,
    n566,
    n270
  );


  or
  g574
  (
    n608,
    n350,
    n357,
    n549,
    n275
  );


  xnor
  g575
  (
    n597,
    n551,
    n516,
    n308,
    n276
  );


  and
  g576
  (
    n594,
    n232,
    n215,
    n354,
    n297
  );


  nor
  g577
  (
    n572,
    n568,
    n298,
    n550,
    n281
  );


  nor
  g578
  (
    n615,
    n525,
    n306,
    n336,
    n301
  );


  nand
  g579
  (
    n583,
    n519,
    n267,
    n325,
    n302
  );


  or
  g580
  (
    n592,
    n246,
    n567,
    n362,
    n305
  );


  nor
  g581
  (
    n622,
    n234,
    n286,
    n226,
    n211
  );


  xor
  g582
  (
    n614,
    n307,
    n277,
    n208,
    n316
  );


  nand
  g583
  (
    n601,
    n239,
    n351,
    n310,
    n319
  );


  or
  g584
  (
    n580,
    n249,
    n369,
    n563,
    n347
  );


  nand
  g585
  (
    KeyWire_0_12,
    n348,
    n540,
    n235,
    n364
  );


  xnor
  g586
  (
    n623,
    n268,
    n244,
    n331,
    n262
  );


  xor
  g587
  (
    n596,
    n330,
    n265,
    n256,
    n299
  );


  or
  g588
  (
    n599,
    n517,
    n213,
    n514,
    n524
  );


  nor
  g589
  (
    n593,
    n538,
    n284,
    n337,
    n254
  );


  nand
  g590
  (
    KeyWire_0_28,
    n261,
    n529,
    n556,
    n247
  );


  nor
  g591
  (
    n618,
    n326,
    n561,
    n250,
    n222
  );


  xor
  g592
  (
    n619,
    n264,
    n274,
    n295,
    n318
  );


  or
  g593
  (
    n591,
    n520,
    n559,
    n248,
    n534
  );


  and
  g594
  (
    n602,
    n513,
    n552,
    n207,
    n565
  );


  not
  g595
  (
    n634,
    n579
  );


  buf
  g596
  (
    n630,
    n577
  );


  not
  g597
  (
    n633,
    n582
  );


  not
  g598
  (
    n627,
    n575
  );


  not
  g599
  (
    n636,
    n574
  );


  not
  g600
  (
    n631,
    n569
  );


  buf
  g601
  (
    n628,
    n583
  );


  not
  g602
  (
    n625,
    n580
  );


  buf
  g603
  (
    n638,
    n572
  );


  not
  g604
  (
    n632,
    n571
  );


  not
  g605
  (
    n629,
    n578
  );


  buf
  g606
  (
    n626,
    n573
  );


  not
  g607
  (
    n635,
    n570
  );


  not
  g608
  (
    n639,
    n576
  );


  buf
  g609
  (
    n637,
    n581
  );


  xnor
  g610
  (
    n641,
    n608,
    n636,
    n627
  );


  nand
  g611
  (
    n651,
    n631,
    n605,
    n613,
    n598
  );


  and
  g612
  (
    n655,
    n629,
    n594,
    n604,
    n607
  );


  and
  g613
  (
    n647,
    n610,
    n601,
    n633,
    n596
  );


  nand
  g614
  (
    n650,
    n615,
    n590,
    n618,
    n595
  );


  and
  g615
  (
    n644,
    n617,
    n597,
    n612,
    n635
  );


  nand
  g616
  (
    n652,
    n634,
    n639,
    n586,
    n592
  );


  nand
  g617
  (
    n646,
    n637,
    n618,
    n609,
    n625
  );


  xor
  g618
  (
    n654,
    n613,
    n599,
    n611,
    n615
  );


  or
  g619
  (
    n640,
    n600,
    n612,
    n609,
    n614
  );


  xnor
  g620
  (
    n653,
    n611,
    n607,
    n606,
    n593
  );


  or
  g621
  (
    n642,
    n591,
    n639,
    n585,
    n614
  );


  or
  g622
  (
    n648,
    n628,
    n626,
    n616,
    n603
  );


  nor
  g623
  (
    n643,
    n610,
    n630,
    n588,
    n608
  );


  xnor
  g624
  (
    n649,
    n589,
    n616,
    n584,
    n587
  );


  nor
  g625
  (
    n645,
    n602,
    n632,
    n638,
    n617
  );


  or
  g626
  (
    n678,
    n422,
    n452,
    n650,
    n457
  );


  nand
  g627
  (
    n660,
    n400,
    n410,
    n652,
    n648
  );


  xnor
  g628
  (
    n671,
    n469,
    n448,
    n644,
    n412
  );


  nand
  g629
  (
    n685,
    n377,
    n381,
    n655,
    n483
  );


  nor
  g630
  (
    n681,
    n462,
    n374,
    n144,
    n641
  );


  xor
  g631
  (
    n690,
    n464,
    n456,
    n440,
    n406
  );


  and
  g632
  (
    n657,
    n425,
    n391,
    n450,
    n644
  );


  xor
  g633
  (
    n659,
    n646,
    n468,
    n396,
    n649
  );


  or
  g634
  (
    n684,
    n482,
    n471,
    n640,
    n475
  );


  xor
  g635
  (
    KeyWire_0_37,
    n461,
    n655,
    n435,
    n652
  );


  xor
  g636
  (
    n661,
    n472,
    n648,
    n418,
    n417
  );


  xnor
  g637
  (
    n692,
    n402,
    n654,
    n407,
    n423
  );


  nand
  g638
  (
    n694,
    n487,
    n653,
    n420,
    n654
  );


  xnor
  g639
  (
    n664,
    n426,
    n647,
    n389,
    n395
  );


  xor
  g640
  (
    KeyWire_0_61,
    n411,
    n458,
    n649,
    n652
  );


  nand
  g641
  (
    n687,
    n489,
    n492,
    n373,
    n442
  );


  nor
  g642
  (
    KeyWire_0_10,
    n653,
    n470,
    n421,
    n399
  );


  nor
  g643
  (
    n691,
    n651,
    n398,
    n642,
    n409
  );


  nor
  g644
  (
    n693,
    n380,
    n424,
    n378,
    n653
  );


  nand
  g645
  (
    n668,
    n651,
    n466,
    n428,
    n642
  );


  xor
  g646
  (
    n695,
    n655,
    n416,
    n397,
    n437
  );


  xor
  g647
  (
    n665,
    n478,
    n491,
    n390,
    n405
  );


  xor
  g648
  (
    KeyWire_0_38,
    n379,
    n485,
    n413,
    n376
  );


  xnor
  g649
  (
    n662,
    n443,
    n473,
    n388,
    n414
  );


  xnor
  g650
  (
    n679,
    n449,
    n652,
    n654,
    n467
  );


  xnor
  g651
  (
    n682,
    n476,
    n143,
    n641,
    n393
  );


  or
  g652
  (
    n667,
    n460,
    n415,
    n372,
    n385
  );


  nor
  g653
  (
    n680,
    n384,
    n144,
    n484,
    n651
  );


  nor
  g654
  (
    n686,
    n646,
    n650,
    n432,
    n651
  );


  and
  g655
  (
    n666,
    n446,
    n490,
    n488,
    n383
  );


  xor
  g656
  (
    n676,
    n654,
    n441,
    n419,
    n645
  );


  nand
  g657
  (
    KeyWire_0_2,
    n144,
    n444,
    n451,
    n647
  );


  xnor
  g658
  (
    KeyWire_0_30,
    n479,
    n427,
    n392,
    n655
  );


  or
  g659
  (
    n673,
    n431,
    n486,
    n408,
    n447
  );


  and
  g660
  (
    n697,
    n455,
    n429,
    n387,
    n401
  );


  nand
  g661
  (
    n683,
    n453,
    n465,
    n480,
    n394
  );


  xor
  g662
  (
    n688,
    n371,
    n645,
    n436,
    n653
  );


  and
  g663
  (
    n663,
    n454,
    n474,
    n439,
    n404
  );


  nor
  g664
  (
    n689,
    n459,
    n375,
    n640,
    n386
  );


  or
  g665
  (
    n672,
    n438,
    n477,
    n382,
    n643
  );


  xnor
  g666
  (
    n658,
    n433,
    n643,
    n445,
    n463
  );


  and
  g667
  (
    n669,
    n430,
    n481,
    n403,
    n434
  );


  buf
  g668
  (
    n706,
    n678
  );


  not
  g669
  (
    n698,
    n620
  );


  buf
  g670
  (
    n700,
    n144
  );


  not
  g671
  (
    n701,
    n676
  );


  not
  g672
  (
    n705,
    n619
  );


  buf
  g673
  (
    n699,
    n620
  );


  not
  g674
  (
    n703,
    n621
  );


  not
  g675
  (
    n704,
    n672
  );


  xnor
  g676
  (
    n702,
    n679,
    n677
  );


  xor
  g677
  (
    n708,
    n145,
    n675,
    n619,
    n682
  );


  nor
  g678
  (
    n707,
    n674,
    n681,
    n680,
    n673
  );


  buf
  g679
  (
    n712,
    n707
  );


  not
  g680
  (
    n710,
    n708
  );


  buf
  g681
  (
    n717,
    n706
  );


  buf
  g682
  (
    n713,
    n701
  );


  buf
  g683
  (
    n723,
    n145
  );


  buf
  g684
  (
    n724,
    n705
  );


  buf
  g685
  (
    n719,
    n145
  );


  not
  g686
  (
    n709,
    n702
  );


  buf
  g687
  (
    n711,
    n705
  );


  not
  g688
  (
    n718,
    n145
  );


  not
  g689
  (
    n714,
    n688
  );


  buf
  g690
  (
    n722,
    n698
  );


  buf
  g691
  (
    n720,
    n685
  );


  or
  g692
  (
    n716,
    n684,
    n686,
    n704
  );


  xnor
  g693
  (
    n721,
    n706,
    n708,
    n707,
    n687
  );


  or
  g694
  (
    n715,
    n700,
    n699,
    n703,
    n683
  );


  buf
  g695
  (
    n725,
    n709
  );


  buf
  g696
  (
    KeyWire_0_25,
    n717
  );


  buf
  g697
  (
    n770,
    n710
  );


  buf
  g698
  (
    n738,
    n720
  );


  buf
  g699
  (
    n751,
    n493
  );


  not
  g700
  (
    n731,
    n718
  );


  buf
  g701
  (
    n756,
    n720
  );


  buf
  g702
  (
    KeyWire_0_17,
    n506
  );


  buf
  g703
  (
    n752,
    n509
  );


  not
  g704
  (
    n753,
    n716
  );


  buf
  g705
  (
    n769,
    n499
  );


  not
  g706
  (
    n754,
    n720
  );


  not
  g707
  (
    n748,
    n502
  );


  not
  g708
  (
    KeyWire_0_15,
    n710
  );


  not
  g709
  (
    n768,
    n717
  );


  not
  g710
  (
    n739,
    n498
  );


  buf
  g711
  (
    n755,
    n503
  );


  not
  g712
  (
    n732,
    n497
  );


  not
  g713
  (
    n760,
    n712
  );


  not
  g714
  (
    n774,
    n721
  );


  buf
  g715
  (
    n730,
    n716
  );


  buf
  g716
  (
    n728,
    n714
  );


  buf
  g717
  (
    n737,
    n494
  );


  buf
  g718
  (
    n765,
    n712
  );


  buf
  g719
  (
    n776,
    n511
  );


  buf
  g720
  (
    n763,
    n495
  );


  buf
  g721
  (
    n736,
    n715
  );


  buf
  g722
  (
    n758,
    n711
  );


  nor
  g723
  (
    KeyWire_0_35,
    n709,
    n496
  );


  xor
  g724
  (
    n746,
    n510,
    n721
  );


  xor
  g725
  (
    KeyWire_0_52,
    n715,
    n713
  );


  nor
  g726
  (
    n745,
    n711,
    n508
  );


  or
  g727
  (
    n775,
    n714,
    n715
  );


  xnor
  g728
  (
    n741,
    n718,
    n711
  );


  xor
  g729
  (
    n767,
    n714,
    n717
  );


  or
  g730
  (
    n735,
    n718,
    n710
  );


  nor
  g731
  (
    n734,
    n713,
    n709
  );


  xnor
  g732
  (
    n747,
    n711,
    n718
  );


  xnor
  g733
  (
    n771,
    n510,
    n716
  );


  nor
  g734
  (
    n761,
    n721,
    n508
  );


  nand
  g735
  (
    n759,
    n719,
    n507
  );


  xor
  g736
  (
    n727,
    n714,
    n717
  );


  or
  g737
  (
    KeyWire_0_63,
    n504,
    n712
  );


  xor
  g738
  (
    n726,
    n715,
    n500
  );


  nor
  g739
  (
    n762,
    n511,
    n709
  );


  xnor
  g740
  (
    n743,
    n509,
    n720
  );


  and
  g741
  (
    n729,
    n712,
    n501
  );


  or
  g742
  (
    n766,
    n713,
    n721
  );


  and
  g743
  (
    n740,
    n716,
    n505
  );


  not
  g744
  (
    n773,
    n719
  );


  and
  g745
  (
    n733,
    n719,
    n507
  );


  and
  g746
  (
    n757,
    n713,
    n710
  );


  not
  g747
  (
    n780,
    n740
  );


  not
  g748
  (
    n787,
    n729
  );


  buf
  g749
  (
    n786,
    n747
  );


  buf
  g750
  (
    n800,
    n736
  );


  buf
  g751
  (
    n779,
    n725
  );


  not
  g752
  (
    n790,
    n755
  );


  buf
  g753
  (
    KeyWire_0_32,
    n743
  );


  not
  g754
  (
    n804,
    n745
  );


  not
  g755
  (
    n792,
    n739
  );


  not
  g756
  (
    KeyWire_0_4,
    n622
  );


  buf
  g757
  (
    n803,
    n752
  );


  not
  g758
  (
    n795,
    n733
  );


  nand
  g759
  (
    n801,
    n738,
    n622,
    n623,
    n757
  );


  nor
  g760
  (
    n783,
    n725,
    n735,
    n732,
    n737
  );


  and
  g761
  (
    n798,
    n750,
    n734,
    n737
  );


  and
  g762
  (
    n789,
    n624,
    n756,
    n727,
    n726
  );


  and
  g763
  (
    n802,
    n753,
    n756,
    n728,
    n748
  );


  xnor
  g764
  (
    n793,
    n753,
    n730,
    n735,
    n743
  );


  nand
  g765
  (
    n781,
    n741,
    n726,
    n751,
    n742
  );


  xnor
  g766
  (
    n784,
    n750,
    n623,
    n746,
    n624
  );


  and
  g767
  (
    n788,
    n741,
    n749,
    n728
  );


  xnor
  g768
  (
    n785,
    n736,
    n738,
    n746,
    n727
  );


  nand
  g769
  (
    n797,
    n729,
    n755,
    n733,
    n754
  );


  nor
  g770
  (
    n777,
    n739,
    n759,
    n731,
    n744
  );


  nand
  g771
  (
    n782,
    n731,
    n751,
    n757,
    n740
  );


  or
  g772
  (
    n796,
    n742,
    n758,
    n745,
    n747
  );


  nand
  g773
  (
    KeyWire_0_23,
    n730,
    n752,
    n758,
    n754
  );


  or
  g774
  (
    n791,
    n744,
    n732,
    n621,
    n748
  );


  not
  g775
  (
    n823,
    n786
  );


  not
  g776
  (
    n827,
    n760
  );


  buf
  g777
  (
    n826,
    n787
  );


  not
  g778
  (
    n825,
    n800
  );


  not
  g779
  (
    n816,
    n782
  );


  not
  g780
  (
    n808,
    n789
  );


  buf
  g781
  (
    n813,
    n764
  );


  not
  g782
  (
    n824,
    n761
  );


  not
  g783
  (
    n811,
    n784
  );


  buf
  g784
  (
    n817,
    n762
  );


  buf
  g785
  (
    KeyWire_0_59,
    n780
  );


  buf
  g786
  (
    KeyWire_0_62,
    n762
  );


  not
  g787
  (
    n815,
    n790
  );


  buf
  g788
  (
    n812,
    n785
  );


  not
  g789
  (
    n810,
    n763
  );


  not
  g790
  (
    n809,
    n759
  );


  buf
  g791
  (
    n818,
    n779
  );


  not
  g792
  (
    n807,
    n760
  );


  not
  g793
  (
    n806,
    n796
  );


  not
  g794
  (
    n814,
    n795
  );


  nor
  g795
  (
    n828,
    n792,
    n788
  );


  and
  g796
  (
    n819,
    n777,
    n781,
    n761,
    n793
  );


  nand
  g797
  (
    n821,
    n783,
    n799,
    n794,
    n778
  );


  or
  g798
  (
    n822,
    n763,
    n798,
    n791,
    n797
  );


  xnor
  g799
  (
    n843,
    n804,
    n808,
    n809,
    n815
  );


  xor
  g800
  (
    n830,
    n805,
    n818,
    n811,
    n691
  );


  nor
  g801
  (
    n842,
    n814,
    n724,
    n809,
    n813
  );


  nand
  g802
  (
    n829,
    n817,
    n816,
    n724,
    n812
  );


  xor
  g803
  (
    n846,
    n811,
    n816
  );


  nand
  g804
  (
    n847,
    n724,
    n722,
    n814
  );


  and
  g805
  (
    n833,
    n816,
    n805,
    n723,
    n807
  );


  or
  g806
  (
    n844,
    n810,
    n805,
    n817
  );


  xor
  g807
  (
    KeyWire_0_19,
    n815,
    n723,
    n817
  );


  or
  g808
  (
    n838,
    n689,
    n803,
    n807,
    n694
  );


  or
  g809
  (
    KeyWire_0_14,
    n801,
    n812,
    n807,
    n802
  );


  xor
  g810
  (
    n837,
    n812,
    n724,
    n723,
    n806
  );


  xor
  g811
  (
    n841,
    n722,
    n810,
    n814
  );


  xor
  g812
  (
    n831,
    n813,
    n808,
    n815,
    n814
  );


  xnor
  g813
  (
    n834,
    n818,
    n813,
    n806
  );


  nand
  g814
  (
    n840,
    n809,
    n693,
    n806,
    n690
  );


  nor
  g815
  (
    n832,
    n808,
    n809,
    n812,
    n806
  );


  and
  g816
  (
    n845,
    n722,
    n807,
    n723,
    n811
  );


  xnor
  g817
  (
    n835,
    n810,
    n815,
    n808,
    n692
  );


  xnor
  g818
  (
    n859,
    n824,
    n837,
    n835,
    n820
  );


  nor
  g819
  (
    n864,
    n767,
    n819,
    n768
  );


  or
  g820
  (
    n852,
    n821,
    n826,
    n831
  );


  nand
  g821
  (
    n855,
    n768,
    n823,
    n822,
    n825
  );


  nand
  g822
  (
    n857,
    n820,
    n846,
    n827,
    n839
  );


  xor
  g823
  (
    n848,
    n764,
    n828,
    n840,
    n827
  );


  nor
  g824
  (
    n858,
    n827,
    n823,
    n828,
    n844
  );


  nor
  g825
  (
    n853,
    n824,
    n828,
    n836,
    n821
  );


  and
  g826
  (
    n854,
    n767,
    n822,
    n818,
    n766
  );


  or
  g827
  (
    KeyWire_0_7,
    n825,
    n826,
    n841,
    n820
  );


  xor
  g828
  (
    n860,
    n825,
    n826,
    n821,
    n842
  );


  nor
  g829
  (
    n861,
    n823,
    n819,
    n822,
    n838
  );


  xnor
  g830
  (
    n863,
    n828,
    n833,
    n834,
    n847
  );


  xnor
  g831
  (
    n856,
    n818,
    n765,
    n822,
    n827
  );


  nand
  g832
  (
    n862,
    n824,
    n821,
    n843,
    n820
  );


  nor
  g833
  (
    KeyWire_0_3,
    n765,
    n766,
    n824,
    n832
  );


  and
  g834
  (
    n849,
    n823,
    n819,
    n845,
    n825
  );


  nand
  g835
  (
    n865,
    n773,
    n862,
    n855,
    n863
  );


  nand
  g836
  (
    n870,
    n775,
    n775,
    n772,
    n774
  );


  nor
  g837
  (
    n866,
    n776,
    n774,
    n771,
    n773
  );


  xor
  g838
  (
    n869,
    n772,
    n861,
    n774,
    n771
  );


  or
  g839
  (
    n867,
    n775,
    n852,
    n854,
    n848
  );


  nand
  g840
  (
    n871,
    n860,
    n857,
    n776,
    n859
  );


  nor
  g841
  (
    KeyWire_0_20,
    n858,
    n769,
    n851
  );


  xnor
  g842
  (
    n876,
    n696,
    n776,
    n853,
    n769
  );


  nand
  g843
  (
    n873,
    n849,
    n774,
    n770
  );


  and
  g844
  (
    n872,
    n771,
    n864,
    n776,
    n770
  );


  nor
  g845
  (
    n874,
    n850,
    n772,
    n695,
    n773
  );


  xor
  g846
  (
    n868,
    n773,
    n856,
    n697,
    n775
  );


  or
  g847
  (
    n878,
    n870,
    n874,
    n873,
    n871
  );


  and
  g848
  (
    n879,
    n865,
    n875,
    n876,
    n867
  );


  and
  g849
  (
    KeyWire_0_9,
    n868,
    n872,
    n866,
    n869
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n587,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n179,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n674,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n851,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n794,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n325,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n268,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n850,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n310,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n877,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n696,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n215,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n606,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n32,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n839,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n749,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n355,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n772,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n508,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n836,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n875,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n131,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n450,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n778,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n482,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n742,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n143,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n470,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n589,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n219,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n656,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n408,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n799,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n305,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n455,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n744,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n428,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n677,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n675,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n496,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n308,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n313,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n550,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n609,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n442,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n258,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n411,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n554,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n502,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n351,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n49,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n327,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n764,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n603,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n192,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n144,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n273,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n347,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n383,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n820,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n226,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n670,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n805,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n750,
    KeyNOTWire_0_63
  );


endmodule


