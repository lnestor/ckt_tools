// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_56 written by SynthGen on 2021/04/05 11:22:31
module MyModule( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n10, n105, n120, n101, n102, n104, n117, n122,
 n116, n123, n108, n99, n97, n121, n115, n95,
 n93, n107, n118, n98, n113, n106, n96, n109,
 n112, n114, n100, n128, n129, n130, n132, n131);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output nCHANGED, n105, n120, n101, n102, n104, n117, n122,
 n116, n123, n108, n99, n97, n121, n115, n95,
 n93, n107, n118, n98, n113, n106, n96, n109,
 n112, n114, n100, n128, n129, n130, n132, n131;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n94, n103, n110, n111,
 n119, n124, n125, n126, n127;

not  g0 (n52, n20);
not  g1 (n76, n28);
not  g2 (n36, n19);
not  g3 (n60, n19);
not  g4 (n64, n12);
not  g5 (n42, n18);
buf  g6 (n44, n25);
not  g7 (n71, n28);
not  g8 (n68, n25);
not  g9 (n34, n17);
buf  g10 (n47, n6);
buf  g11 (n35, n22);
not  g12 (n54, n23);
not  g13 (n81, n22);
not  g14 (n69, n16);
not  g15 (n58, n20);
not  g16 (n80, n23);
buf  g17 (n51, n3);
buf  g18 (n59, n25);
not  g19 (n33, n27);
buf  g20 (n46, n7);
buf  g21 (n67, n2);
not  g22 (n63, n26);
buf  g23 (n56, n24);
not  g24 (n78, n13);
not  g25 (n40, n15);
buf  g26 (n66, n11);
buf  g27 (n70, n22);
buf  g28 (n48, n24);
not  g29 (n37, n26);
buf  g30 (n72, n27);
buf  g31 (n65, n24);
buf  g32 (n57, n18);
buf  g33 (n41, n21);
buf  g34 (n82, n21);
buf  g35 (n61, n4);
buf  g36 (n49, n9);
not  g37 (n83, n20);
buf  g38 (n74, n27);
buf  g39 (n75, n21);
not  g40 (n38, n19);
buf  g41 (n43, n14);
buf  g42 (n84, n29);
buf  g43 (n77, n10);
buf  g44 (n79, n29);
buf  g45 (n62, n28);
not  g46 (n53, n23);
not  g47 (n73, n1);
not  g48 (n45, n5);
buf  g49 (n39, n8);
not  g50 (n55, n26);
not  g51 (n50, n18);
buf  g52 (n85, n35);
buf  g53 (n88, n34);
not  g54 (n86, n36);
buf  g55 (n87, n37);
not  g56 (n90, n33);
buf  g57 (n89, n38);
not  g58 (n92, n39);
buf  g59 (n91, n40);
xor  g60 (n121, n68, n82, n74, n85);
nor  g61 (n104, n57, n84, n75, n59);
nor  g62 (n117, n75, n88, n83, n42);
and  g63 (n99, n86, n56, n46, n71);
xor  g64 (n98, n63, n86, n91, n62);
nor  g65 (n107, n73, n79, n67);
xnor g66 (n110, n82, n83, n89, n81);
nand g67 (n111, n90, n85, n92, n78);
nand g68 (n113, n67, n70, n87, n78);
xnor g69 (n108, n74, n84, n77, n91);
or   g70 (n122, n76, n61, n73, n79);
xor  g71 (n112, n53, n92, n65, n89);
nand g72 (n105, n80, n72, n63);
nand g73 (n123, n77, n69);
nand g74 (n109, n75, n91, n86, n48);
and  g75 (n116, n89, n71, n77, n52);
and  g76 (n124, n91, n85, n54, n60);
nand g77 (n94, n62, n61, n87);
xnor g78 (n101, n71, n59, n50, n58);
nor  g79 (n96, n72, n79, n51, n88);
nor  g80 (n103, n65, n70, n76, n49);
xnor g81 (n97, n84, n90, n62, n80);
or   g82 (n118, n45, n66, n64, n90);
nor  g83 (n95, n66, n41, n47, n78);
nor  g84 (n102, n60, n43, n87, n89);
and  g85 (n100, n90, n61, n64, n83);
or   g86 (n114, n68, n55, n81, n72);
or   g87 (n119, n92, n73, n74, n85);
xor  g88 (n115, n76, n82, n60, n59);
or   g89 (n93, n64, n70, n68, n80);
xor  g90 (n106, n44, n92, n86, n88);
xnor g91 (n120, n81, n66, n65, n88);
not  g92 (n127, n121);
not  g93 (n126, n120);
not  g94 (n125, n119);
xnor g95 (n128, n123, n122, n127, n30);
and  g96 (n131, n126, n29, n31);
nor  g97 (n130, n125, n126, n30);
nand g98 (n129, n124, n32);
and  g99 (n132, n31, n127, n126);
buf g100 (nCHANGED, n10);
endmodule
