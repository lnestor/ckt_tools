

module Stat_100_51
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n129,
  n105,
  n102,
  n114,
  n120,
  n106,
  n119,
  n117,
  n108,
  n109,
  n124,
  n132,
  n103,
  n131,
  n116,
  n123,
  n104,
  n121,
  n111,
  n113,
  n125,
  n127,
  n122,
  n110,
  n130,
  n115,
  n118,
  n126,
  n112,
  n101,
  n128,
  n107
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n129;output n105;output n102;output n114;output n120;output n106;output n119;output n117;output n108;output n109;output n124;output n132;output n103;output n131;output n116;output n123;output n104;output n121;output n111;output n113;output n125;output n127;output n122;output n110;output n130;output n115;output n118;output n126;output n112;output n101;output n128;output n107;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n41,
    n22
  );


  and
  g1
  (
    n36,
    n24,
    n31,
    n5,
    n19
  );


  xnor
  g2
  (
    n39,
    n26,
    n20,
    n16,
    n1
  );


  and
  g3
  (
    KeyWire_0_25,
    n4,
    n2,
    n17,
    n21
  );


  xor
  g4
  (
    n35,
    n29,
    n9,
    n15,
    n8
  );


  xor
  g5
  (
    n40,
    n11,
    n6,
    n3,
    n30
  );


  and
  g6
  (
    KeyWire_0_28,
    n28,
    n27,
    n18,
    n31
  );


  xor
  g7
  (
    n38,
    n14,
    n10,
    n7,
    n23
  );


  or
  g8
  (
    KeyWire_0_26,
    n13,
    n12,
    n31,
    n25
  );


  not
  g9
  (
    n43,
    n35
  );


  not
  g10
  (
    n46,
    n36
  );


  not
  g11
  (
    n49,
    n37
  );


  buf
  g12
  (
    KeyWire_0_31,
    n40
  );


  not
  g13
  (
    KeyWire_0_8,
    n39
  );


  buf
  g14
  (
    n42,
    n33
  );


  buf
  g15
  (
    n47,
    n34
  );


  buf
  g16
  (
    KeyWire_0_29,
    n38
  );


  not
  g17
  (
    n65,
    n46
  );


  buf
  g18
  (
    n68,
    n44
  );


  buf
  g19
  (
    n76,
    n42
  );


  buf
  g20
  (
    KeyWire_0_0,
    n43
  );


  buf
  g21
  (
    n75,
    n45
  );


  not
  g22
  (
    KeyWire_0_2,
    n47
  );


  buf
  g23
  (
    n67,
    n43
  );


  buf
  g24
  (
    n77,
    n46
  );


  buf
  g25
  (
    n56,
    n41
  );


  not
  g26
  (
    n52,
    n44
  );


  buf
  g27
  (
    n66,
    n44
  );


  buf
  g28
  (
    n62,
    n47
  );


  buf
  g29
  (
    n55,
    n46
  );


  not
  g30
  (
    n54,
    n46
  );


  buf
  g31
  (
    KeyWire_0_4,
    n45
  );


  buf
  g32
  (
    n53,
    n49
  );


  buf
  g33
  (
    n78,
    n49
  );


  not
  g34
  (
    n73,
    n42
  );


  buf
  g35
  (
    n50,
    n47
  );


  not
  g36
  (
    n61,
    n43
  );


  not
  g37
  (
    n70,
    n42
  );


  buf
  g38
  (
    n59,
    n48
  );


  buf
  g39
  (
    KeyWire_0_18,
    n45
  );


  buf
  g40
  (
    KeyWire_0_19,
    n42
  );


  not
  g41
  (
    n74,
    n44
  );


  not
  g42
  (
    n58,
    n48
  );


  not
  g43
  (
    n71,
    n48
  );


  buf
  g44
  (
    n72,
    n45
  );


  not
  g45
  (
    n69,
    n32
  );


  nand
  g46
  (
    KeyWire_0_9,
    n32,
    n48,
    n43,
    n47
  );


  not
  g47
  (
    KeyWire_0_6,
    n54
  );


  not
  g48
  (
    n89,
    n51
  );


  buf
  g49
  (
    KeyWire_0_17,
    n32
  );


  buf
  g50
  (
    KeyWire_0_5,
    n55
  );


  buf
  g51
  (
    n82,
    n49
  );


  buf
  g52
  (
    n92,
    n50
  );


  not
  g53
  (
    n96,
    n52
  );


  buf
  g54
  (
    KeyWire_0_12,
    n54
  );


  buf
  g55
  (
    n81,
    n54
  );


  buf
  g56
  (
    n83,
    n52
  );


  not
  g57
  (
    n87,
    n53
  );


  not
  g58
  (
    n85,
    n55
  );


  buf
  g59
  (
    KeyWire_0_23,
    n50
  );


  buf
  g60
  (
    n80,
    n49
  );


  buf
  g61
  (
    KeyWire_0_20,
    n53
  );


  not
  g62
  (
    n94,
    n51
  );


  not
  g63
  (
    KeyWire_0_27,
    n55
  );


  buf
  g64
  (
    KeyWire_0_15,
    n52
  );


  not
  g65
  (
    n84,
    n53
  );


  buf
  g66
  (
    n99,
    n51
  );


  xor
  g67
  (
    KeyWire_0_7,
    n55,
    n50,
    n53,
    n54
  );


  and
  g68
  (
    n109,
    n93,
    n70,
    n99,
    n79
  );


  nor
  g69
  (
    KeyWire_0_22,
    n60,
    n77,
    n64,
    n73
  );


  nand
  g70
  (
    KeyWire_0_1,
    n63,
    n68,
    n56,
    n82
  );


  or
  g71
  (
    n107,
    n60,
    n67,
    n78,
    n62
  );


  xor
  g72
  (
    n122,
    n65,
    n56,
    n99,
    n76
  );


  or
  g73
  (
    n132,
    n74,
    n96,
    n67,
    n57
  );


  xor
  g74
  (
    n111,
    n69,
    n62,
    n74,
    n98
  );


  xor
  g75
  (
    KeyWire_0_13,
    n71,
    n58,
    n99,
    n62
  );


  xor
  g76
  (
    n102,
    n61,
    n71,
    n75,
    n64
  );


  or
  g77
  (
    KeyWire_0_10,
    n67,
    n75,
    n87,
    n79
  );


  xnor
  g78
  (
    n123,
    n59,
    n77,
    n96,
    n71
  );


  xor
  g79
  (
    n110,
    n97,
    n76,
    n57,
    n78
  );


  nor
  g80
  (
    n117,
    n63,
    n66,
    n62,
    n98
  );


  and
  g81
  (
    n127,
    n76,
    n65,
    n75,
    n66
  );


  and
  g82
  (
    n106,
    n64,
    n97,
    n70,
    n84
  );


  and
  g83
  (
    n130,
    n89,
    n59,
    n58,
    n69
  );


  or
  g84
  (
    KeyWire_0_11,
    n85,
    n100,
    n61,
    n57
  );


  nor
  g85
  (
    KeyWire_0_14,
    n98,
    n61,
    n88,
    n97
  );


  nand
  g86
  (
    n131,
    n91,
    n90,
    n58,
    n56
  );


  nor
  g87
  (
    KeyWire_0_21,
    n94,
    n68,
    n67,
    n78
  );


  nor
  g88
  (
    KeyWire_0_24,
    n70,
    n81,
    n68,
    n71
  );


  and
  g89
  (
    KeyWire_0_30,
    n78,
    n72,
    n77,
    n92
  );


  nand
  g90
  (
    n113,
    n66,
    n69,
    n73,
    n79
  );


  xnor
  g91
  (
    n101,
    n69,
    n59,
    n58,
    n68
  );


  xor
  g92
  (
    n103,
    n100,
    n60,
    n63
  );


  xor
  g93
  (
    n129,
    n95,
    n57,
    n66,
    n74
  );


  and
  g94
  (
    n118,
    n70,
    n61,
    n86,
    n73
  );


  nand
  g95
  (
    n115,
    n65,
    n83,
    n79,
    n100
  );


  xor
  g96
  (
    KeyWire_0_3,
    n64,
    n72,
    n77,
    n73
  );


  xor
  g97
  (
    n126,
    n63,
    n56,
    n75,
    n59
  );


  xor
  g98
  (
    n125,
    n80,
    n95,
    n72,
    n74
  );


  xor
  g99
  (
    KeyWire_0_16,
    n76,
    n72,
    n96,
    n65
  );


  xnor
  KeyGate_0_0
  (
    n64,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n124,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n57,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n112,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n51,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n90,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n93,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n88,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n48,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n79,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n114,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n116,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n100,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n108,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n128,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n91,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n120,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n86,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n63,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n60,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n97,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n121,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n119,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n95,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n105,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n37,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n34,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n98,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n33,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n44,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n104,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n45,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


