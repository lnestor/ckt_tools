

module Stat_100_43
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n108,
  n118,
  n127,
  n131,
  n124,
  n115,
  n125,
  n116,
  n101,
  n126,
  n129,
  n111,
  n112,
  n110,
  n120,
  n123,
  n104,
  n130,
  n113,
  n132,
  n128,
  n102,
  n114,
  n119,
  n109,
  n121,
  n122,
  n105,
  n106,
  n107,
  n117,
  n103
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n108;output n118;output n127;output n131;output n124;output n115;output n125;output n116;output n101;output n126;output n129;output n111;output n112;output n110;output n120;output n123;output n104;output n130;output n113;output n132;output n128;output n102;output n114;output n119;output n109;output n121;output n122;output n105;output n106;output n107;output n117;output n103;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  not
  g0
  (
    KeyWire_0_10,
    n3
  );


  not
  g1
  (
    n46,
    n4
  );


  not
  g2
  (
    n33,
    n2
  );


  buf
  g3
  (
    n39,
    n2
  );


  not
  g4
  (
    KeyWire_0_9,
    n2
  );


  not
  g5
  (
    n47,
    n1
  );


  not
  g6
  (
    KeyWire_0_7,
    n1
  );


  not
  g7
  (
    n35,
    n3
  );


  not
  g8
  (
    n36,
    n3
  );


  not
  g9
  (
    n37,
    n3
  );


  not
  g10
  (
    n40,
    n4
  );


  not
  g11
  (
    KeyWire_0_11,
    n1
  );


  buf
  g12
  (
    KeyWire_0_13,
    n4
  );


  not
  g13
  (
    n41,
    n1
  );


  buf
  g14
  (
    n42,
    n2
  );


  buf
  g15
  (
    KeyWire_0_15,
    n7
  );


  not
  g16
  (
    n76,
    n44
  );


  not
  g17
  (
    n49,
    n24
  );


  not
  g18
  (
    n57,
    n27
  );


  not
  g19
  (
    n63,
    n38
  );


  buf
  g20
  (
    n73,
    n35
  );


  or
  g21
  (
    n79,
    n12,
    n9,
    n13
  );


  xnor
  g22
  (
    n89,
    n34,
    n24,
    n8,
    n7
  );


  nand
  g23
  (
    n88,
    n38,
    n5,
    n22,
    n21
  );


  xor
  g24
  (
    KeyWire_0_5,
    n29,
    n11,
    n31,
    n39
  );


  xor
  g25
  (
    n51,
    n37,
    n30,
    n20,
    n43
  );


  and
  g26
  (
    n92,
    n23,
    n20,
    n14,
    n44
  );


  xnor
  g27
  (
    n48,
    n27,
    n10,
    n34,
    n15
  );


  nand
  g28
  (
    n71,
    n39,
    n19,
    n17,
    n37
  );


  nand
  g29
  (
    n72,
    n34,
    n15,
    n29,
    n31
  );


  xnor
  g30
  (
    n64,
    n41,
    n37,
    n6,
    n26
  );


  nor
  g31
  (
    n75,
    n22,
    n22,
    n30,
    n35
  );


  nand
  g32
  (
    n77,
    n29,
    n44,
    n18,
    n17
  );


  nand
  g33
  (
    KeyWire_0_4,
    n33,
    n29,
    n10,
    n17
  );


  xor
  g34
  (
    n53,
    n43,
    n28,
    n41,
    n14
  );


  or
  g35
  (
    n81,
    n32,
    n21,
    n42,
    n26
  );


  or
  g36
  (
    KeyWire_0_6,
    n17,
    n12,
    n30,
    n26
  );


  nand
  g37
  (
    n61,
    n16,
    n9,
    n26,
    n43
  );


  xor
  g38
  (
    n52,
    n31,
    n42,
    n20,
    n30
  );


  xnor
  g39
  (
    n82,
    n21,
    n19,
    n6,
    n5
  );


  and
  g40
  (
    KeyWire_0_12,
    n45,
    n16,
    n9,
    n23
  );


  xor
  g41
  (
    n86,
    n18,
    n18,
    n24,
    n36
  );


  xor
  g42
  (
    n80,
    n44,
    n11,
    n5,
    n25
  );


  nor
  g43
  (
    n67,
    n45,
    n40,
    n19,
    n42
  );


  and
  g44
  (
    n62,
    n25,
    n12,
    n38,
    n22
  );


  xor
  g45
  (
    n87,
    n32,
    n42,
    n8,
    n35
  );


  nor
  g46
  (
    n83,
    n40,
    n14,
    n15,
    n7
  );


  and
  g47
  (
    n66,
    n23,
    n15,
    n37,
    n32
  );


  and
  g48
  (
    n90,
    n28,
    n5,
    n25,
    n41
  );


  nand
  g49
  (
    n68,
    n16,
    n23,
    n31,
    n34
  );


  and
  g50
  (
    n50,
    n16,
    n45,
    n6,
    n10
  );


  or
  g51
  (
    n59,
    n39,
    n9,
    n25,
    n7
  );


  nor
  g52
  (
    n60,
    n36,
    n40,
    n35,
    n38
  );


  xor
  g53
  (
    n54,
    n14,
    n28,
    n36
  );


  nor
  g54
  (
    n58,
    n21,
    n40,
    n27,
    n43
  );


  nand
  g55
  (
    n69,
    n41,
    n8,
    n28
  );


  nand
  g56
  (
    n70,
    n18,
    n27,
    n11
  );


  xnor
  g57
  (
    n65,
    n12,
    n13,
    n24
  );


  nand
  g58
  (
    n85,
    n39,
    n4,
    n10,
    n6
  );


  and
  g59
  (
    n74,
    n20,
    n45,
    n19,
    n32
  );


  buf
  g60
  (
    n97,
    n51
  );


  not
  g61
  (
    n100,
    n47
  );


  not
  g62
  (
    n95,
    n48
  );


  not
  g63
  (
    n99,
    n50
  );


  xor
  g64
  (
    n96,
    n47,
    n58,
    n46
  );


  nand
  g65
  (
    n93,
    n47,
    n49,
    n57,
    n53
  );


  xnor
  g66
  (
    n94,
    n56,
    n46,
    n52
  );


  nor
  g67
  (
    n98,
    n47,
    n59,
    n54,
    n55
  );


  or
  g68
  (
    n102,
    n90,
    n75,
    n87,
    n83
  );


  xor
  g69
  (
    n104,
    n96,
    n90,
    n79,
    n89
  );


  xnor
  g70
  (
    n106,
    n67,
    n72,
    n60,
    n90
  );


  nand
  g71
  (
    KeyWire_0_2,
    n81,
    n61,
    n84,
    n93
  );


  nor
  g72
  (
    n113,
    n85,
    n73,
    n77,
    n93
  );


  xnor
  g73
  (
    n122,
    n97,
    n80,
    n83,
    n89
  );


  xor
  g74
  (
    n109,
    n85,
    n95,
    n99,
    n90
  );


  xor
  g75
  (
    n118,
    n99,
    n89,
    n77,
    n68
  );


  or
  g76
  (
    n117,
    n75,
    n74,
    n78,
    n92
  );


  xnor
  g77
  (
    n125,
    n81,
    n76,
    n72,
    n85
  );


  nor
  g78
  (
    n123,
    n85,
    n77,
    n82,
    n92
  );


  nor
  g79
  (
    KeyWire_0_3,
    n89,
    n76,
    n70,
    n64
  );


  nand
  g80
  (
    n128,
    n100,
    n74,
    n96,
    n95
  );


  xnor
  g81
  (
    n129,
    n83,
    n75,
    n93,
    n73
  );


  xnor
  g82
  (
    n107,
    n96,
    n88,
    n95,
    n79
  );


  xnor
  g83
  (
    KeyWire_0_14,
    n80,
    n65,
    n81,
    n73
  );


  xor
  g84
  (
    n112,
    n86,
    n87,
    n91,
    n97
  );


  or
  g85
  (
    n111,
    n100,
    n82,
    n66,
    n72
  );


  nor
  g86
  (
    n126,
    n100,
    n96,
    n93,
    n92
  );


  xnor
  g87
  (
    n116,
    n94,
    n95,
    n62,
    n86
  );


  or
  g88
  (
    n131,
    n79,
    n78,
    n98,
    n81
  );


  nand
  g89
  (
    KeyWire_0_8,
    n84,
    n94,
    n72,
    n88
  );


  xor
  g90
  (
    n105,
    n91,
    n77,
    n97,
    n71
  );


  xnor
  g91
  (
    n110,
    n98,
    n86,
    n99,
    n97
  );


  xor
  g92
  (
    n124,
    n91,
    n82,
    n74,
    n76
  );


  or
  g93
  (
    KeyWire_0_0,
    n94,
    n94,
    n87,
    n76
  );


  xnor
  g94
  (
    n115,
    n86,
    n88,
    n78,
    n82
  );


  nand
  g95
  (
    n108,
    n63,
    n73,
    n99,
    n80
  );


  and
  g96
  (
    n103,
    n74,
    n79,
    n84,
    n91
  );


  nand
  g97
  (
    n119,
    n92,
    n88,
    n80,
    n98
  );


  and
  g98
  (
    KeyWire_0_1,
    n87,
    n75,
    n100,
    n69
  );


  or
  g99
  (
    n120,
    n83,
    n84,
    n98,
    n78
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n132,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n121,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n130,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n114,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n56,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n78,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n91,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n38,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n101,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n44,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n43,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n45,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n84,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n34,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n127,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n55,
    KeyNOTWire_0_15
  );


endmodule


