

module Stat_100_41
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n131,
  n117,
  n108,
  n125,
  n121,
  n130,
  n118,
  n102,
  n116,
  n110,
  n124,
  n128,
  n122,
  n114,
  n104,
  n109,
  n113,
  n123,
  n101,
  n127,
  n105,
  n119,
  n103,
  n120,
  n106,
  n132,
  n129,
  n107,
  n126,
  n111,
  n115
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n112;output n131;output n117;output n108;output n125;output n121;output n130;output n118;output n102;output n116;output n110;output n124;output n128;output n122;output n114;output n104;output n109;output n113;output n123;output n101;output n127;output n105;output n119;output n103;output n120;output n106;output n132;output n129;output n107;output n126;output n111;output n115;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;

  not
  g0
  (
    KeyWire_0_12,
    n4
  );


  not
  g1
  (
    n39,
    n2
  );


  not
  g2
  (
    n34,
    n3
  );


  buf
  g3
  (
    n42,
    n3
  );


  buf
  g4
  (
    n35,
    n2
  );


  not
  g5
  (
    n41,
    n1
  );


  buf
  g6
  (
    KeyWire_0_11,
    n3
  );


  not
  g7
  (
    n38,
    n4
  );


  buf
  g8
  (
    n36,
    n1
  );


  not
  g9
  (
    n43,
    n1
  );


  buf
  g10
  (
    n33,
    n2
  );


  not
  g11
  (
    n44,
    n4
  );


  not
  g12
  (
    KeyWire_0_8,
    n13
  );


  buf
  g13
  (
    n66,
    n15
  );


  buf
  g14
  (
    n76,
    n27
  );


  not
  g15
  (
    n72,
    n8
  );


  not
  g16
  (
    n51,
    n31
  );


  not
  g17
  (
    n73,
    n33
  );


  buf
  g18
  (
    n71,
    n31
  );


  not
  g19
  (
    n75,
    n19
  );


  or
  g20
  (
    n61,
    n11,
    n21,
    n18,
    n42
  );


  nor
  g21
  (
    n64,
    n22,
    n41,
    n36,
    n18
  );


  nand
  g22
  (
    KeyWire_0_4,
    n35,
    n17,
    n25,
    n20
  );


  nand
  g23
  (
    n45,
    n37,
    n39,
    n42,
    n43
  );


  nor
  g24
  (
    n80,
    n22,
    n19,
    n35,
    n44
  );


  or
  g25
  (
    n74,
    n18,
    n13,
    n7,
    n28
  );


  xor
  g26
  (
    KeyWire_0_5,
    n43,
    n30,
    n39,
    n38
  );


  xor
  g27
  (
    n49,
    n29,
    n24,
    n6,
    n26
  );


  nor
  g28
  (
    n65,
    n40,
    n14,
    n9,
    n11
  );


  and
  g29
  (
    n50,
    n7,
    n16,
    n10,
    n19
  );


  or
  g30
  (
    n58,
    n9,
    n35,
    n16,
    n42
  );


  and
  g31
  (
    n69,
    n29,
    n41,
    n37,
    n20
  );


  and
  g32
  (
    n53,
    n37,
    n44,
    n23,
    n27
  );


  nand
  g33
  (
    n63,
    n32,
    n25,
    n34,
    n5
  );


  and
  g34
  (
    n52,
    n14,
    n38,
    n44,
    n8
  );


  xor
  g35
  (
    n55,
    n9,
    n23,
    n22,
    n15
  );


  and
  g36
  (
    n70,
    n17,
    n6,
    n33,
    n43
  );


  nand
  g37
  (
    n47,
    n12,
    n24,
    n5,
    n26
  );


  or
  g38
  (
    n79,
    n24,
    n16,
    n32,
    n13
  );


  and
  g39
  (
    n48,
    n29,
    n11,
    n7,
    n26
  );


  nand
  g40
  (
    n46,
    n30,
    n36,
    n40,
    n6
  );


  nor
  g41
  (
    n56,
    n30,
    n39,
    n21,
    n10
  );


  nand
  g42
  (
    KeyWire_0_13,
    n25,
    n10,
    n41,
    n31
  );


  nand
  g43
  (
    n67,
    n14,
    n15,
    n5,
    n8
  );


  nor
  g44
  (
    KeyWire_0_1,
    n38,
    n27,
    n36,
    n32
  );


  and
  g45
  (
    n68,
    n17,
    n34,
    n33,
    n20
  );


  xor
  g46
  (
    n77,
    n28,
    n23,
    n12,
    n40
  );


  xor
  g47
  (
    n62,
    n34,
    n21,
    n12,
    n28
  );


  buf
  g48
  (
    KeyWire_0_6,
    n45
  );


  not
  g49
  (
    n84,
    n49
  );


  buf
  g50
  (
    KeyWire_0_7,
    n48
  );


  buf
  g51
  (
    n92,
    n45
  );


  buf
  g52
  (
    n83,
    n46
  );


  buf
  g53
  (
    n91,
    n48
  );


  buf
  g54
  (
    n85,
    n46
  );


  not
  g55
  (
    n90,
    n50
  );


  buf
  g56
  (
    n82,
    n50
  );


  buf
  g57
  (
    n89,
    n49
  );


  buf
  g58
  (
    n94,
    n51
  );


  not
  g59
  (
    KeyWire_0_15,
    n51
  );


  buf
  g60
  (
    n86,
    n48
  );


  buf
  g61
  (
    n100,
    n50
  );


  not
  g62
  (
    n98,
    n46
  );


  buf
  g63
  (
    KeyWire_0_0,
    n45
  );


  buf
  g64
  (
    n87,
    n47
  );


  not
  g65
  (
    n97,
    n47
  );


  not
  g66
  (
    n99,
    n47
  );


  not
  g67
  (
    KeyWire_0_14,
    n49
  );


  or
  g68
  (
    KeyWire_0_9,
    n97,
    n64,
    n98,
    n70
  );


  xnor
  g69
  (
    n102,
    n60,
    n80,
    n95
  );


  or
  g70
  (
    n125,
    n78,
    n74,
    n71,
    n77
  );


  or
  g71
  (
    n130,
    n57,
    n63,
    n69,
    n99
  );


  xnor
  g72
  (
    n121,
    n88,
    n56,
    n72,
    n58
  );


  or
  g73
  (
    n128,
    n70,
    n91,
    n94,
    n60
  );


  or
  g74
  (
    n113,
    n71,
    n54,
    n51,
    n59
  );


  nand
  g75
  (
    n115,
    n86,
    n94,
    n62
  );


  nand
  g76
  (
    n129,
    n82,
    n75,
    n52,
    n61
  );


  and
  g77
  (
    n112,
    n62,
    n85,
    n54,
    n75
  );


  xor
  g78
  (
    n108,
    n59,
    n79,
    n68,
    n91
  );


  xor
  g79
  (
    n114,
    n69,
    n92,
    n53,
    n65
  );


  xor
  g80
  (
    KeyWire_0_2,
    n83,
    n91,
    n60,
    n68
  );


  nand
  g81
  (
    n104,
    n74,
    n72,
    n89,
    n65
  );


  xor
  g82
  (
    n105,
    n68,
    n64,
    n81,
    n92
  );


  xnor
  g83
  (
    n110,
    n53,
    n92,
    n99,
    n98
  );


  or
  g84
  (
    n101,
    n56,
    n56,
    n61,
    n66
  );


  nand
  g85
  (
    n106,
    n65,
    n99,
    n93,
    n74
  );


  nand
  g86
  (
    n118,
    n73,
    n55,
    n78,
    n76
  );


  xnor
  g87
  (
    n123,
    n95,
    n87,
    n71,
    n55
  );


  nor
  g88
  (
    n107,
    n97,
    n70,
    n84,
    n79
  );


  nor
  g89
  (
    n103,
    n58,
    n77,
    n66,
    n52
  );


  nand
  g90
  (
    n122,
    n63,
    n80,
    n59,
    n93
  );


  nand
  g91
  (
    n109,
    n64,
    n72,
    n100,
    n57
  );


  nor
  g92
  (
    n126,
    n58,
    n67,
    n73,
    n66
  );


  xor
  g93
  (
    KeyWire_0_10,
    n100,
    n73,
    n80,
    n96
  );


  and
  g94
  (
    n124,
    n54,
    n67,
    n90,
    n61
  );


  xnor
  g95
  (
    n111,
    n76,
    n75,
    n52,
    n53
  );


  or
  g96
  (
    n132,
    n67,
    n93,
    n96,
    n78
  );


  or
  g97
  (
    n131,
    n98,
    n96,
    n94,
    n79
  );


  nor
  g98
  (
    n116,
    n69,
    n97,
    n57,
    n100
  );


  or
  g99
  (
    KeyWire_0_3,
    n55,
    n76,
    n63,
    n77
  );


  xnor
  KeyGate_0_0
  (
    n93,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n57,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n119,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n127,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n78,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n60,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n96,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n81,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n59,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n120,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n117,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n37,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n40,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n54,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n95,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n88,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


