

module Stat_393_1615
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n153,
  n158,
  n151,
  n140,
  n155,
  n354,
  n381,
  n386,
  n383,
  n391,
  n395,
  n399,
  n390,
  n389,
  n408,
  n406,
  n405,
  n402,
  n404,
  n407,
  n410,
  n401,
  n411,
  n400,
  n409,
  n403
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n153;output n158;output n151;output n140;output n155;output n354;output n381;output n386;output n383;output n391;output n395;output n399;output n390;output n389;output n408;output n406;output n405;output n402;output n404;output n407;output n410;output n401;output n411;output n400;output n409;output n403;
  wire n19;wire n20;wire n21;wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n152;wire n154;wire n156;wire n157;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n382;wire n384;wire n385;wire n387;wire n388;wire n392;wire n393;wire n394;wire n396;wire n397;wire n398;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    KeyWire_0_47,
    n3
  );


  buf
  g1
  (
    n33,
    n6
  );


  not
  g2
  (
    n49,
    n2
  );


  buf
  g3
  (
    n44,
    n2
  );


  buf
  g4
  (
    KeyWire_0_50,
    n4
  );


  not
  g5
  (
    n21,
    n4
  );


  not
  g6
  (
    n23,
    n6
  );


  buf
  g7
  (
    n27,
    n5
  );


  buf
  g8
  (
    n25,
    n6
  );


  not
  g9
  (
    n42,
    n5
  );


  not
  g10
  (
    n46,
    n8
  );


  buf
  g11
  (
    n48,
    n8
  );


  buf
  g12
  (
    n22,
    n7
  );


  not
  g13
  (
    KeyWire_0_35,
    n2
  );


  not
  g14
  (
    n47,
    n3
  );


  buf
  g15
  (
    n34,
    n7
  );


  not
  g16
  (
    n28,
    n4
  );


  buf
  g17
  (
    n36,
    n7
  );


  not
  g18
  (
    n26,
    n5
  );


  buf
  g19
  (
    KeyWire_0_60,
    n5
  );


  not
  g20
  (
    n19,
    n3
  );


  not
  g21
  (
    n35,
    n1
  );


  buf
  g22
  (
    n24,
    n4
  );


  not
  g23
  (
    n43,
    n3
  );


  buf
  g24
  (
    n41,
    n1
  );


  buf
  g25
  (
    n20,
    n6
  );


  buf
  g26
  (
    KeyWire_0_49,
    n2
  );


  not
  g27
  (
    n40,
    n1
  );


  not
  g28
  (
    KeyWire_0_25,
    n1
  );


  buf
  g29
  (
    n32,
    n8
  );


  buf
  g30
  (
    n39,
    n7
  );


  buf
  g31
  (
    n75,
    n26
  );


  buf
  g32
  (
    n62,
    n24
  );


  not
  g33
  (
    n53,
    n24
  );


  buf
  g34
  (
    n69,
    n23
  );


  buf
  g35
  (
    n72,
    n20
  );


  buf
  g36
  (
    n71,
    n22
  );


  not
  g37
  (
    n79,
    n19
  );


  not
  g38
  (
    KeyWire_0_4,
    n22
  );


  buf
  g39
  (
    n60,
    n21
  );


  not
  g40
  (
    n56,
    n20
  );


  buf
  g41
  (
    KeyWire_0_7,
    n23
  );


  not
  g42
  (
    KeyWire_0_0,
    n20
  );


  not
  g43
  (
    n58,
    n23
  );


  not
  g44
  (
    n65,
    n21
  );


  buf
  g45
  (
    n67,
    n25
  );


  not
  g46
  (
    n52,
    n24
  );


  buf
  g47
  (
    n66,
    n19
  );


  buf
  g48
  (
    n76,
    n25
  );


  buf
  g49
  (
    n63,
    n21
  );


  not
  g50
  (
    n59,
    n21
  );


  not
  g51
  (
    KeyWire_0_13,
    n23
  );


  not
  g52
  (
    n68,
    n22
  );


  buf
  g53
  (
    n73,
    n20
  );


  not
  g54
  (
    n57,
    n22
  );


  not
  g55
  (
    n54,
    n24
  );


  buf
  g56
  (
    n51,
    n19
  );


  not
  g57
  (
    n77,
    n26
  );


  not
  g58
  (
    n61,
    n25
  );


  not
  g59
  (
    n64,
    n19
  );


  buf
  g60
  (
    n74,
    n25
  );


  buf
  g61
  (
    n86,
    n60
  );


  not
  g62
  (
    n99,
    n54
  );


  not
  g63
  (
    n97,
    n61
  );


  not
  g64
  (
    KeyWire_0_3,
    n62
  );


  buf
  g65
  (
    n106,
    n52
  );


  buf
  g66
  (
    n107,
    n53
  );


  not
  g67
  (
    n83,
    n58
  );


  buf
  g68
  (
    n131,
    n58
  );


  not
  g69
  (
    n111,
    n51
  );


  buf
  g70
  (
    n113,
    n57
  );


  not
  g71
  (
    n88,
    n55
  );


  not
  g72
  (
    n121,
    n57
  );


  not
  g73
  (
    n82,
    n57
  );


  not
  g74
  (
    n119,
    n53
  );


  not
  g75
  (
    n114,
    n50
  );


  buf
  g76
  (
    n98,
    n50
  );


  not
  g77
  (
    KeyWire_0_6,
    n52
  );


  not
  g78
  (
    n103,
    n51
  );


  buf
  g79
  (
    n128,
    n53
  );


  buf
  g80
  (
    n129,
    n54
  );


  not
  g81
  (
    KeyWire_0_40,
    n51
  );


  not
  g82
  (
    n90,
    n52
  );


  buf
  g83
  (
    n104,
    n53
  );


  not
  g84
  (
    n123,
    n56
  );


  buf
  g85
  (
    n117,
    n62
  );


  buf
  g86
  (
    n80,
    n61
  );


  buf
  g87
  (
    KeyWire_0_1,
    n54
  );


  buf
  g88
  (
    n120,
    n59
  );


  buf
  g89
  (
    KeyWire_0_16,
    n52
  );


  not
  g90
  (
    n93,
    n60
  );


  buf
  g91
  (
    n125,
    n56
  );


  buf
  g92
  (
    n109,
    n58
  );


  not
  g93
  (
    n94,
    n60
  );


  buf
  g94
  (
    n100,
    n50
  );


  not
  g95
  (
    n126,
    n59
  );


  not
  g96
  (
    n81,
    n59
  );


  buf
  g97
  (
    n127,
    n62
  );


  not
  g98
  (
    n130,
    n57
  );


  buf
  g99
  (
    n91,
    n58
  );


  not
  g100
  (
    n118,
    n59
  );


  not
  g101
  (
    n116,
    n61
  );


  buf
  g102
  (
    n101,
    n51
  );


  buf
  g103
  (
    n84,
    n62
  );


  not
  g104
  (
    n102,
    n56
  );


  not
  g105
  (
    n124,
    n56
  );


  buf
  g106
  (
    n85,
    n50
  );


  buf
  g107
  (
    n96,
    n60
  );


  not
  g108
  (
    n87,
    n55
  );


  buf
  g109
  (
    n89,
    n55
  );


  buf
  g110
  (
    n112,
    n61
  );


  not
  g111
  (
    n122,
    n55
  );


  not
  g112
  (
    n95,
    n54
  );


  not
  g113
  (
    n146,
    n99
  );


  not
  g114
  (
    n133,
    n81
  );


  not
  g115
  (
    n132,
    n101
  );


  buf
  g116
  (
    KeyWire_0_14,
    n94
  );


  not
  g117
  (
    n147,
    n88
  );


  not
  g118
  (
    KeyWire_0_48,
    n81
  );


  and
  g119
  (
    n158,
    n86,
    n92
  );


  nor
  g120
  (
    n153,
    n97,
    n88,
    n98,
    n92
  );


  xor
  g121
  (
    n148,
    n87,
    n84,
    n82,
    n93
  );


  xnor
  g122
  (
    n137,
    n96,
    n101,
    n85,
    n93
  );


  and
  g123
  (
    n145,
    n84,
    n88,
    n100,
    n80
  );


  nor
  g124
  (
    KeyWire_0_44,
    n98,
    n86,
    n94,
    n91
  );


  or
  g125
  (
    KeyWire_0_42,
    n84,
    n90,
    n97,
    n95
  );


  nor
  g126
  (
    n151,
    n88,
    n87,
    n89,
    n83
  );


  and
  g127
  (
    n152,
    n97,
    n95,
    n90
  );


  xnor
  g128
  (
    n134,
    n94,
    n81,
    n97,
    n80
  );


  or
  g129
  (
    n138,
    n86,
    n89,
    n96,
    n90
  );


  xor
  g130
  (
    n143,
    n98,
    n80,
    n86,
    n87
  );


  nand
  g131
  (
    KeyWire_0_5,
    n83,
    n96,
    n98,
    n99
  );


  or
  g132
  (
    n156,
    n91,
    n99,
    n90,
    n87
  );


  nor
  g133
  (
    n155,
    n100,
    n82,
    n91,
    n94
  );


  or
  g134
  (
    n135,
    n85,
    n92,
    n83,
    n82
  );


  or
  g135
  (
    KeyWire_0_21,
    n91,
    n96,
    n92,
    n84
  );


  nand
  g136
  (
    n154,
    n89,
    n85,
    n100,
    n83
  );


  or
  g137
  (
    n142,
    n82,
    n100,
    n89,
    n93
  );


  xnor
  g138
  (
    n136,
    n95,
    n93,
    n85,
    n101
  );


  nor
  g139
  (
    n149,
    n101,
    n81,
    n99,
    n80
  );


  not
  g140
  (
    n165,
    n146
  );


  not
  g141
  (
    n167,
    n144
  );


  buf
  g142
  (
    n163,
    n137
  );


  buf
  g143
  (
    KeyWire_0_58,
    n138
  );


  buf
  g144
  (
    KeyWire_0_24,
    n142
  );


  not
  g145
  (
    n159,
    n145
  );


  not
  g146
  (
    n168,
    n143
  );


  buf
  g147
  (
    n166,
    n139
  );


  not
  g148
  (
    n161,
    n140
  );


  buf
  g149
  (
    n164,
    n141
  );


  buf
  g150
  (
    n185,
    n167
  );


  buf
  g151
  (
    n202,
    n9
  );


  not
  g152
  (
    n190,
    n8
  );


  not
  g153
  (
    n173,
    n14
  );


  buf
  g154
  (
    n204,
    n11
  );


  buf
  g155
  (
    n199,
    n163
  );


  buf
  g156
  (
    n180,
    n10
  );


  not
  g157
  (
    n186,
    n15
  );


  not
  g158
  (
    n206,
    n160
  );


  buf
  g159
  (
    n169,
    n165
  );


  not
  g160
  (
    n183,
    n13
  );


  not
  g161
  (
    n175,
    n12
  );


  buf
  g162
  (
    KeyWire_0_10,
    n166
  );


  buf
  g163
  (
    n181,
    n166
  );


  not
  g164
  (
    n192,
    n168
  );


  buf
  g165
  (
    n176,
    n164
  );


  buf
  g166
  (
    n198,
    n167
  );


  not
  g167
  (
    n205,
    n167
  );


  buf
  g168
  (
    n172,
    n166
  );


  not
  g169
  (
    KeyWire_0_29,
    n161
  );


  not
  g170
  (
    n182,
    n168
  );


  not
  g171
  (
    KeyWire_0_23,
    n9
  );


  buf
  g172
  (
    n178,
    n159
  );


  not
  g173
  (
    KeyWire_0_41,
    n166
  );


  buf
  g174
  (
    n197,
    n10
  );


  not
  g175
  (
    n188,
    n168
  );


  buf
  g176
  (
    n196,
    n161
  );


  buf
  g177
  (
    n203,
    n167
  );


  and
  g178
  (
    n189,
    n164,
    n161,
    n162,
    n11
  );


  and
  g179
  (
    n187,
    n163,
    n9,
    n160,
    n161
  );


  nand
  g180
  (
    n193,
    n162,
    n13,
    n10
  );


  and
  g181
  (
    n171,
    n160,
    n165,
    n16
  );


  nor
  g182
  (
    KeyWire_0_43,
    n14,
    n15,
    n12,
    n162
  );


  xnor
  g183
  (
    n174,
    n14,
    n11,
    n160,
    n9
  );


  nor
  g184
  (
    n177,
    n163,
    n164,
    n15
  );


  xnor
  g185
  (
    n195,
    n13,
    n10,
    n12,
    n164
  );


  xnor
  g186
  (
    KeyWire_0_34,
    n168,
    n159,
    n12,
    n11
  );


  nor
  g187
  (
    KeyWire_0_62,
    n163,
    n165,
    n162,
    n14
  );


  not
  g188
  (
    n209,
    n170
  );


  not
  g189
  (
    n214,
    n177
  );


  buf
  g190
  (
    n215,
    n177
  );


  buf
  g191
  (
    n213,
    n174
  );


  not
  g192
  (
    n208,
    n171
  );


  not
  g193
  (
    n211,
    n176
  );


  not
  g194
  (
    n212,
    n169
  );


  buf
  g195
  (
    KeyWire_0_46,
    n175
  );


  buf
  g196
  (
    n210,
    n173
  );


  not
  g197
  (
    n216,
    n172
  );


  buf
  g198
  (
    n244,
    n207
  );


  not
  g199
  (
    n235,
    n67
  );


  buf
  g200
  (
    KeyWire_0_11,
    n73
  );


  buf
  g201
  (
    n237,
    n68
  );


  not
  g202
  (
    n250,
    n69
  );


  not
  g203
  (
    n255,
    n66
  );


  not
  g204
  (
    n240,
    n215
  );


  buf
  g205
  (
    n219,
    n16
  );


  not
  g206
  (
    n226,
    n213
  );


  buf
  g207
  (
    n223,
    n64
  );


  buf
  g208
  (
    n227,
    n71
  );


  not
  g209
  (
    n221,
    n71
  );


  xor
  g210
  (
    n247,
    n65,
    n216,
    n209
  );


  or
  g211
  (
    n218,
    n65,
    n64,
    n73
  );


  nor
  g212
  (
    n234,
    n70,
    n16,
    n213
  );


  nor
  g213
  (
    n231,
    n209,
    n208,
    n68
  );


  or
  g214
  (
    n241,
    n215,
    n70,
    n73
  );


  or
  g215
  (
    n224,
    n75,
    n207,
    n76
  );


  xor
  g216
  (
    n251,
    n75,
    n215,
    n16
  );


  or
  g217
  (
    n245,
    n63,
    n69,
    n75
  );


  xor
  g218
  (
    KeyWire_0_9,
    n207,
    n66,
    n70
  );


  nand
  g219
  (
    n236,
    n73,
    n211,
    n213
  );


  nor
  g220
  (
    n253,
    n63,
    n216,
    n74
  );


  or
  g221
  (
    n239,
    n211,
    n210,
    n214
  );


  nor
  g222
  (
    n222,
    n64,
    n67,
    n207
  );


  xor
  g223
  (
    n249,
    n69,
    n67,
    n212
  );


  xnor
  g224
  (
    n256,
    n214,
    n72,
    n211
  );


  nor
  g225
  (
    KeyWire_0_28,
    n70,
    n212,
    n65
  );


  and
  g226
  (
    n230,
    n68,
    n210,
    n208
  );


  nor
  g227
  (
    n254,
    n209,
    n212,
    n75
  );


  and
  g228
  (
    n217,
    n72,
    n63,
    n68
  );


  xnor
  g229
  (
    KeyWire_0_31,
    n71,
    n76,
    n212
  );


  xor
  g230
  (
    KeyWire_0_17,
    n211,
    n213,
    n64
  );


  nor
  g231
  (
    n232,
    n67,
    n74,
    n208
  );


  xor
  g232
  (
    n220,
    n208,
    n69,
    n210
  );


  or
  g233
  (
    n248,
    n63,
    n65,
    n74
  );


  xor
  g234
  (
    KeyWire_0_53,
    n74,
    n72,
    n210
  );


  or
  g235
  (
    n252,
    n71,
    n72,
    n66
  );


  or
  g236
  (
    n242,
    n216,
    n209,
    n214
  );


  nand
  g237
  (
    n225,
    n214,
    n215,
    n66,
    n216
  );


  or
  g238
  (
    KeyWire_0_26,
    n121,
    n106,
    n39,
    n47
  );


  nor
  g239
  (
    n285,
    n102,
    n104,
    n43,
    n38
  );


  nor
  g240
  (
    n280,
    n48,
    n231,
    n105
  );


  xor
  g241
  (
    n311,
    n44,
    n111,
    n120,
    n42
  );


  nor
  g242
  (
    n281,
    n114,
    n28,
    n232,
    n37
  );


  nand
  g243
  (
    n315,
    n127,
    n117,
    n243,
    n42
  );


  nand
  g244
  (
    n291,
    n34,
    n109,
    n107,
    n238
  );


  and
  g245
  (
    n265,
    n42,
    n239,
    n242,
    n45
  );


  xor
  g246
  (
    n275,
    n109,
    n104,
    n110,
    n31
  );


  xnor
  g247
  (
    n278,
    n243,
    n30,
    n125
  );


  xnor
  g248
  (
    n313,
    n127,
    n39,
    n106,
    n26
  );


  and
  g249
  (
    n304,
    n34,
    n104,
    n123,
    n40
  );


  nand
  g250
  (
    KeyWire_0_56,
    n242,
    n27,
    n249,
    n102
  );


  and
  g251
  (
    n268,
    n233,
    n248,
    n41,
    n226
  );


  xnor
  g252
  (
    n296,
    n49,
    n36,
    n33,
    n112
  );


  and
  g253
  (
    n297,
    n124,
    n113,
    n128,
    n245
  );


  and
  g254
  (
    n321,
    n124,
    n118,
    n43,
    n225
  );


  or
  g255
  (
    n324,
    n229,
    n111,
    n248,
    n116
  );


  nand
  g256
  (
    n274,
    n120,
    n49,
    n226,
    n123
  );


  or
  g257
  (
    n272,
    n35,
    n105,
    n220,
    n225
  );


  nand
  g258
  (
    n258,
    n238,
    n217,
    n37,
    n41
  );


  nor
  g259
  (
    KeyWire_0_57,
    n30,
    n42,
    n113,
    n114
  );


  nor
  g260
  (
    n312,
    n106,
    n118,
    n109,
    n112
  );


  and
  g261
  (
    n314,
    n122,
    n103,
    n33,
    n107
  );


  xnor
  g262
  (
    n320,
    n221,
    n44,
    n35,
    n227
  );


  nor
  g263
  (
    n307,
    n46,
    n232,
    n121,
    n250
  );


  xor
  g264
  (
    n282,
    n28,
    n28,
    n249,
    n107
  );


  nand
  g265
  (
    n295,
    n237,
    n219,
    n28,
    n39
  );


  nor
  g266
  (
    n273,
    n244,
    n118,
    n46,
    n116
  );


  xor
  g267
  (
    n305,
    n120,
    n102,
    n112,
    n223
  );


  nand
  g268
  (
    n289,
    n246,
    n218,
    n108,
    n41
  );


  or
  g269
  (
    n283,
    n250,
    n111,
    n105,
    n121
  );


  or
  g270
  (
    KeyWire_0_27,
    n34,
    n247,
    n43,
    n112
  );


  xnor
  g271
  (
    n292,
    n32,
    n106,
    n122,
    n37
  );


  or
  g272
  (
    n316,
    n125,
    n29,
    n43,
    n240
  );


  and
  g273
  (
    n290,
    n111,
    n128,
    n32,
    n224
  );


  xnor
  g274
  (
    n294,
    n115,
    n115,
    n37,
    n117
  );


  nand
  g275
  (
    n260,
    n127,
    n116,
    n45,
    n40
  );


  nor
  g276
  (
    n276,
    n230,
    n48,
    n115,
    n39
  );


  or
  g277
  (
    KeyWire_0_54,
    n102,
    n117,
    n27,
    n122
  );


  nor
  g278
  (
    n302,
    n114,
    n126,
    n241,
    n245
  );


  nor
  g279
  (
    n303,
    n239,
    n103,
    n44
  );


  xnor
  g280
  (
    n257,
    n33,
    n45,
    n47,
    n123
  );


  xor
  g281
  (
    n308,
    n48,
    n129,
    n40,
    n38
  );


  and
  g282
  (
    n277,
    n109,
    n48,
    n27,
    n44
  );


  nand
  g283
  (
    n301,
    n46,
    n47,
    n27,
    n129
  );


  xor
  g284
  (
    KeyWire_0_61,
    n105,
    n32,
    n228,
    n119
  );


  xnor
  g285
  (
    n306,
    n224,
    n113,
    n116,
    n108
  );


  or
  g286
  (
    n261,
    n30,
    n31,
    n228,
    n123
  );


  xor
  g287
  (
    n318,
    n241,
    n222,
    n121,
    n46
  );


  or
  g288
  (
    n287,
    n247,
    n36,
    n113,
    n35
  );


  xor
  g289
  (
    KeyWire_0_8,
    n119,
    n108,
    n47,
    n115
  );


  nor
  g290
  (
    n298,
    n110,
    n244,
    n120,
    n36
  );


  or
  g291
  (
    n323,
    n235,
    n219,
    n110,
    n128
  );


  nand
  g292
  (
    n269,
    n119,
    n104,
    n40,
    n32
  );


  xor
  g293
  (
    n300,
    n246,
    n218,
    n33,
    n29
  );


  xnor
  g294
  (
    KeyWire_0_15,
    n236,
    n45,
    n125,
    n35
  );


  and
  g295
  (
    n271,
    n223,
    n38,
    n126,
    n110
  );


  or
  g296
  (
    n322,
    n36,
    n229,
    n30,
    n26
  );


  and
  g297
  (
    n310,
    n29,
    n122,
    n103,
    n31
  );


  nor
  g298
  (
    n270,
    n127,
    n41,
    n34,
    n118
  );


  nor
  g299
  (
    n267,
    n108,
    n29,
    n117,
    n217
  );


  nand
  g300
  (
    n259,
    n220,
    n126,
    n234,
    n222
  );


  xnor
  g301
  (
    n286,
    n38,
    n114,
    n234,
    n49
  );


  xnor
  g302
  (
    n279,
    n236,
    n49,
    n233,
    n128
  );


  and
  g303
  (
    n288,
    n227,
    n124,
    n235,
    n221
  );


  nand
  g304
  (
    KeyWire_0_12,
    n119,
    n126,
    n107,
    n31
  );


  and
  g305
  (
    n317,
    n124,
    n240,
    n237,
    n230
  );


  not
  g306
  (
    n334,
    n268
  );


  not
  g307
  (
    n327,
    n265
  );


  buf
  g308
  (
    n326,
    n262
  );


  buf
  g309
  (
    n330,
    n259
  );


  not
  g310
  (
    n328,
    n257
  );


  not
  g311
  (
    n329,
    n261
  );


  not
  g312
  (
    n331,
    n266
  );


  not
  g313
  (
    n332,
    n267
  );


  buf
  g314
  (
    n336,
    n258
  );


  buf
  g315
  (
    n333,
    n260
  );


  buf
  g316
  (
    KeyWire_0_32,
    n263
  );


  not
  g317
  (
    n325,
    n264
  );


  nand
  g318
  (
    n345,
    n79,
    n329,
    n326,
    n131
  );


  nand
  g319
  (
    n338,
    n328,
    n77,
    n330
  );


  or
  g320
  (
    n346,
    n129,
    n79,
    n76,
    n325
  );


  and
  g321
  (
    n344,
    n78,
    n129,
    n77,
    n149
  );


  xor
  g322
  (
    n343,
    n334,
    n78,
    n131
  );


  nor
  g323
  (
    n341,
    n152,
    n150,
    n130
  );


  and
  g324
  (
    n337,
    n130,
    n131,
    n331,
    n76
  );


  and
  g325
  (
    KeyWire_0_22,
    n130,
    n151,
    n79,
    n332
  );


  nand
  g326
  (
    KeyWire_0_55,
    n327,
    n79,
    n147,
    n77
  );


  xor
  g327
  (
    KeyWire_0_36,
    n333,
    n78,
    n148,
    n131
  );


  or
  g328
  (
    n353,
    n194,
    n186,
    n340,
    n188
  );


  nand
  g329
  (
    n354,
    n179,
    n343,
    n341,
    n188
  );


  nand
  g330
  (
    KeyWire_0_20,
    n344,
    n346,
    n180,
    n338
  );


  or
  g331
  (
    n351,
    n180,
    n189,
    n183,
    n182
  );


  xnor
  g332
  (
    n355,
    n192,
    n190,
    n181,
    n185
  );


  xnor
  g333
  (
    n350,
    n191,
    n339,
    n342,
    n193
  );


  xor
  g334
  (
    n356,
    n345,
    n192,
    n193,
    n191
  );


  xor
  g335
  (
    n357,
    n179,
    n337,
    n183,
    n187
  );


  xnor
  g336
  (
    n352,
    n346,
    n184,
    n182,
    n178
  );


  nand
  g337
  (
    n347,
    n184,
    n185,
    n186,
    n181
  );


  and
  g338
  (
    n348,
    n190,
    n178,
    n189,
    n187
  );


  not
  g339
  (
    n361,
    n158
  );


  buf
  g340
  (
    KeyWire_0_37,
    n153
  );


  buf
  g341
  (
    n365,
    n155
  );


  buf
  g342
  (
    n360,
    n352
  );


  not
  g343
  (
    n363,
    n195
  );


  or
  g344
  (
    KeyWire_0_19,
    n196,
    n194
  );


  nand
  g345
  (
    n358,
    n156,
    n357,
    n356,
    n195
  );


  and
  g346
  (
    KeyWire_0_52,
    n157,
    n354,
    n349,
    n351
  );


  xnor
  g347
  (
    n362,
    n353,
    n197,
    n355,
    n348
  );


  xnor
  g348
  (
    n364,
    n350,
    n154,
    n197,
    n196
  );


  and
  g349
  (
    KeyWire_0_51,
    n364,
    n253,
    n17,
    n204
  );


  or
  g350
  (
    n379,
    n17,
    n200,
    n18,
    n204
  );


  and
  g351
  (
    n375,
    n367,
    n251,
    n199,
    n361
  );


  and
  g352
  (
    n371,
    n256,
    n17,
    n202,
    n206
  );


  and
  g353
  (
    KeyWire_0_33,
    n17,
    n362,
    n18,
    n255
  );


  and
  g354
  (
    n372,
    n205,
    n365,
    n199,
    n252
  );


  xnor
  g355
  (
    n369,
    n203,
    n255,
    n201
  );


  or
  g356
  (
    n374,
    n256,
    n363,
    n203,
    n252
  );


  and
  g357
  (
    KeyWire_0_2,
    n359,
    n360,
    n200,
    n198
  );


  xor
  g358
  (
    KeyWire_0_45,
    n358,
    n366,
    n367,
    n253
  );


  or
  g359
  (
    n376,
    n202,
    n254,
    n366
  );


  xnor
  g360
  (
    KeyWire_0_39,
    n251,
    n198,
    n205,
    n206
  );


  xor
  g361
  (
    n383,
    n378,
    n379,
    n282,
    n289
  );


  nand
  g362
  (
    n392,
    n318,
    n299,
    n371,
    n283
  );


  nor
  g363
  (
    n384,
    n287,
    n271,
    n314,
    n376
  );


  xnor
  g364
  (
    n398,
    n305,
    n372,
    n374,
    n324
  );


  xnor
  g365
  (
    n391,
    n290,
    n296,
    n378,
    n306
  );


  nor
  g366
  (
    n389,
    n284,
    n288,
    n373,
    n320
  );


  nor
  g367
  (
    n396,
    n301,
    n291,
    n274,
    n18
  );


  nor
  g368
  (
    n394,
    n377,
    n293,
    n275,
    n298
  );


  xnor
  g369
  (
    n399,
    n373,
    n369,
    n368,
    n319
  );


  xnor
  g370
  (
    n382,
    n276,
    n308,
    n323,
    n280
  );


  nand
  g371
  (
    KeyWire_0_30,
    n269,
    n311,
    n321,
    n375
  );


  or
  g372
  (
    n380,
    n323,
    n313,
    n310,
    n377
  );


  and
  g373
  (
    n388,
    n316,
    n278,
    n315,
    n273
  );


  and
  g374
  (
    n397,
    n302,
    n312,
    n304,
    n295
  );


  nand
  g375
  (
    n385,
    n375,
    n285,
    n303,
    n307
  );


  xnor
  g376
  (
    n387,
    n270,
    n272,
    n297,
    n376
  );


  xor
  g377
  (
    n381,
    n281,
    n370,
    n18,
    n292
  );


  xor
  g378
  (
    n386,
    n374,
    n309,
    n317,
    n322
  );


  or
  g379
  (
    KeyWire_0_63,
    n372,
    n294,
    n300,
    n277
  );


  xnor
  g380
  (
    n393,
    n324,
    n286,
    n279,
    n379
  );


  buf
  g381
  (
    n403,
    n398
  );


  buf
  g382
  (
    KeyWire_0_38,
    n395
  );


  buf
  g383
  (
    n409,
    n336
  );


  not
  g384
  (
    n405,
    n396
  );


  not
  g385
  (
    n408,
    n397
  );


  not
  g386
  (
    KeyWire_0_18,
    n394
  );


  not
  g387
  (
    n407,
    n389
  );


  buf
  g388
  (
    n411,
    n388
  );


  buf
  g389
  (
    n404,
    n335
  );


  buf
  g390
  (
    n410,
    n390
  );


  not
  g391
  (
    n401,
    n392
  );


  xor
  g392
  (
    KeyWire_0_59,
    n391,
    n393,
    n399
  );


  xor
  KeyGate_0_0
  (
    n70,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n110,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n378,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n92,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n55,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n150,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n115,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n50,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n293,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n233,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n170,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n246,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n309,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n78,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n144,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n299,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n108,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n228,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n402,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n366,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n349,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n141,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n339,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n194,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n160,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n37,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n264,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n263,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n243,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n201,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n390,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n229,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n335,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n370,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n184,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n31,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n342,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n359,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n406,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n377,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n105,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n200,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n139,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n191,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n140,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n368,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n207,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n38,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n157,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n30,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n29,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n373,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n367,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n238,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n319,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n340,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n266,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n262,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n162,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n400,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n45,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n284,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n179,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n395,
    KeyNOTWire_0_63
  );


endmodule


