

module Stat_1928_79_6
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n1028,
  n1009,
  n1003,
  n1006,
  n1032,
  n1008,
  n1005,
  n1015,
  n1011,
  n1026,
  n1022,
  n1010,
  n1030,
  n1014,
  n1012,
  n1020,
  n1025,
  n1017,
  n1019,
  n1021,
  n1027,
  n1029,
  n1013,
  n1004,
  n1024,
  n1031,
  n1632,
  n1630,
  n1629,
  n1634,
  n1628,
  n1637,
  n1639,
  n1643,
  n1640,
  n1641,
  n1638,
  n1735,
  n1733,
  n1732,
  n1737,
  n1938,
  n1940,
  n1945,
  n1949,
  n1957,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1028;
  output n1009;
  output n1003;
  output n1006;
  output n1032;
  output n1008;
  output n1005;
  output n1015;
  output n1011;
  output n1026;
  output n1022;
  output n1010;
  output n1030;
  output n1014;
  output n1012;
  output n1020;
  output n1025;
  output n1017;
  output n1019;
  output n1021;
  output n1027;
  output n1029;
  output n1013;
  output n1004;
  output n1024;
  output n1031;
  output n1632;
  output n1630;
  output n1629;
  output n1634;
  output n1628;
  output n1637;
  output n1639;
  output n1643;
  output n1640;
  output n1641;
  output n1638;
  output n1735;
  output n1733;
  output n1732;
  output n1737;
  output n1938;
  output n1940;
  output n1945;
  output n1949;
  output n1957;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1007;
  wire n1016;
  wire n1018;
  wire n1023;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1631;
  wire n1633;
  wire n1635;
  wire n1636;
  wire n1642;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1734;
  wire n1736;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1939;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;

  buf
  g0
  (
    n44,
    n11
  );


  buf
  g1
  (
    n121,
    n1
  );


  not
  g2
  (
    n60,
    n29
  );


  not
  g3
  (
    n133,
    n20
  );


  not
  g4
  (
    n74,
    n12
  );


  not
  g5
  (
    n76,
    n22
  );


  not
  g6
  (
    n99,
    n23
  );


  buf
  g7
  (
    n53,
    n6
  );


  not
  g8
  (
    n91,
    n21
  );


  not
  g9
  (
    n96,
    n21
  );


  not
  g10
  (
    n142,
    n18
  );


  buf
  g11
  (
    n83,
    n28
  );


  not
  g12
  (
    n135,
    n27
  );


  not
  g13
  (
    n86,
    n9
  );


  not
  g14
  (
    n84,
    n18
  );


  not
  g15
  (
    n89,
    n4
  );


  buf
  g16
  (
    n72,
    n1
  );


  buf
  g17
  (
    n143,
    n23
  );


  not
  g18
  (
    n110,
    n20
  );


  not
  g19
  (
    n128,
    n24
  );


  buf
  g20
  (
    n69,
    n6
  );


  buf
  g21
  (
    n126,
    n5
  );


  not
  g22
  (
    n112,
    n13
  );


  buf
  g23
  (
    n129,
    n16
  );


  buf
  g24
  (
    n55,
    n16
  );


  buf
  g25
  (
    n108,
    n2
  );


  not
  g26
  (
    n88,
    n12
  );


  buf
  g27
  (
    n87,
    n19
  );


  not
  g28
  (
    n113,
    n14
  );


  not
  g29
  (
    n90,
    n3
  );


  buf
  g30
  (
    KeyWire_0_3,
    n28
  );


  buf
  g31
  (
    n35,
    n27
  );


  buf
  g32
  (
    n82,
    n11
  );


  not
  g33
  (
    n145,
    n24
  );


  not
  g34
  (
    n52,
    n27
  );


  not
  g35
  (
    n34,
    n12
  );


  not
  g36
  (
    n41,
    n2
  );


  buf
  g37
  (
    n98,
    n24
  );


  not
  g38
  (
    n124,
    n29
  );


  buf
  g39
  (
    n104,
    n28
  );


  buf
  g40
  (
    n36,
    n26
  );


  not
  g41
  (
    n63,
    n4
  );


  not
  g42
  (
    n95,
    n7
  );


  buf
  g43
  (
    n94,
    n8
  );


  not
  g44
  (
    n138,
    n9
  );


  buf
  g45
  (
    n127,
    n15
  );


  not
  g46
  (
    n73,
    n24
  );


  buf
  g47
  (
    n77,
    n20
  );


  buf
  g48
  (
    n132,
    n14
  );


  not
  g49
  (
    n58,
    n25
  );


  not
  g50
  (
    n119,
    n14
  );


  not
  g51
  (
    n40,
    n8
  );


  buf
  g52
  (
    n51,
    n21
  );


  not
  g53
  (
    n118,
    n22
  );


  buf
  g54
  (
    n62,
    n25
  );


  buf
  g55
  (
    n131,
    n1
  );


  not
  g56
  (
    n106,
    n2
  );


  not
  g57
  (
    n144,
    n12
  );


  buf
  g58
  (
    n67,
    n17
  );


  buf
  g59
  (
    n61,
    n29
  );


  not
  g60
  (
    n120,
    n26
  );


  not
  g61
  (
    n46,
    n19
  );


  not
  g62
  (
    n66,
    n10
  );


  not
  g63
  (
    n48,
    n26
  );


  not
  g64
  (
    n30,
    n5
  );


  buf
  g65
  (
    n80,
    n3
  );


  not
  g66
  (
    n123,
    n17
  );


  buf
  g67
  (
    n54,
    n10
  );


  buf
  g68
  (
    n140,
    n10
  );


  not
  g69
  (
    n117,
    n6
  );


  buf
  g70
  (
    n101,
    n13
  );


  not
  g71
  (
    n43,
    n16
  );


  buf
  g72
  (
    n65,
    n5
  );


  not
  g73
  (
    n111,
    n13
  );


  buf
  g74
  (
    n141,
    n7
  );


  not
  g75
  (
    n81,
    n22
  );


  not
  g76
  (
    n47,
    n22
  );


  not
  g77
  (
    n103,
    n18
  );


  buf
  g78
  (
    n136,
    n6
  );


  buf
  g79
  (
    n59,
    n4
  );


  not
  g80
  (
    n64,
    n19
  );


  buf
  g81
  (
    n85,
    n9
  );


  buf
  g82
  (
    n137,
    n18
  );


  not
  g83
  (
    n134,
    n8
  );


  buf
  g84
  (
    n49,
    n8
  );


  not
  g85
  (
    KeyWire_0_5,
    n11
  );


  not
  g86
  (
    n114,
    n5
  );


  buf
  g87
  (
    n32,
    n2
  );


  buf
  g88
  (
    n107,
    n20
  );


  buf
  g89
  (
    n93,
    n15
  );


  not
  g90
  (
    n125,
    n11
  );


  buf
  g91
  (
    n37,
    n17
  );


  buf
  g92
  (
    n78,
    n13
  );


  buf
  g93
  (
    n116,
    n7
  );


  not
  g94
  (
    n105,
    n9
  );


  not
  g95
  (
    n31,
    n15
  );


  buf
  g96
  (
    n122,
    n17
  );


  not
  g97
  (
    n50,
    n21
  );


  buf
  g98
  (
    n68,
    n23
  );


  not
  g99
  (
    n70,
    n14
  );


  buf
  g100
  (
    n42,
    n25
  );


  not
  g101
  (
    n97,
    n1
  );


  not
  g102
  (
    n109,
    n29
  );


  not
  g103
  (
    n71,
    n3
  );


  buf
  g104
  (
    n45,
    n19
  );


  not
  g105
  (
    n56,
    n27
  );


  not
  g106
  (
    n39,
    n10
  );


  not
  g107
  (
    n100,
    n16
  );


  buf
  g108
  (
    n57,
    n23
  );


  buf
  g109
  (
    n75,
    n3
  );


  buf
  g110
  (
    n139,
    n7
  );


  buf
  g111
  (
    n33,
    n15
  );


  not
  g112
  (
    n115,
    n28
  );


  not
  g113
  (
    n38,
    n26
  );


  not
  g114
  (
    n92,
    n4
  );


  buf
  g115
  (
    n79,
    n25
  );


  buf
  g116
  (
    n236,
    n50
  );


  not
  g117
  (
    n484,
    n59
  );


  not
  g118
  (
    n393,
    n40
  );


  not
  g119
  (
    n304,
    n121
  );


  not
  g120
  (
    n274,
    n66
  );


  not
  g121
  (
    n388,
    n128
  );


  buf
  g122
  (
    n255,
    n113
  );


  not
  g123
  (
    KeyWire_0_10,
    n51
  );


  not
  g124
  (
    n413,
    n96
  );


  buf
  g125
  (
    n381,
    n131
  );


  buf
  g126
  (
    n222,
    n40
  );


  buf
  g127
  (
    n161,
    n74
  );


  buf
  g128
  (
    n359,
    n48
  );


  buf
  g129
  (
    n476,
    n62
  );


  buf
  g130
  (
    n415,
    n87
  );


  not
  g131
  (
    n455,
    n46
  );


  not
  g132
  (
    n224,
    n130
  );


  buf
  g133
  (
    n208,
    n95
  );


  buf
  g134
  (
    n325,
    n124
  );


  buf
  g135
  (
    n344,
    n95
  );


  not
  g136
  (
    n181,
    n96
  );


  not
  g137
  (
    n347,
    n111
  );


  not
  g138
  (
    n187,
    n76
  );


  not
  g139
  (
    n363,
    n90
  );


  buf
  g140
  (
    n361,
    n92
  );


  not
  g141
  (
    n147,
    n137
  );


  not
  g142
  (
    n301,
    n30
  );


  not
  g143
  (
    n308,
    n65
  );


  not
  g144
  (
    n399,
    n86
  );


  buf
  g145
  (
    n220,
    n101
  );


  buf
  g146
  (
    n350,
    n53
  );


  not
  g147
  (
    n316,
    n138
  );


  buf
  g148
  (
    n414,
    n45
  );


  not
  g149
  (
    n151,
    n140
  );


  buf
  g150
  (
    n149,
    n82
  );


  not
  g151
  (
    n309,
    n52
  );


  not
  g152
  (
    n279,
    n137
  );


  not
  g153
  (
    n375,
    n120
  );


  not
  g154
  (
    n370,
    n97
  );


  not
  g155
  (
    n230,
    n56
  );


  buf
  g156
  (
    n449,
    n126
  );


  buf
  g157
  (
    n186,
    n98
  );


  buf
  g158
  (
    n379,
    n136
  );


  not
  g159
  (
    n157,
    n88
  );


  buf
  g160
  (
    n268,
    n37
  );


  not
  g161
  (
    n214,
    n97
  );


  not
  g162
  (
    n232,
    n64
  );


  not
  g163
  (
    n465,
    n57
  );


  not
  g164
  (
    n299,
    n127
  );


  not
  g165
  (
    n217,
    n141
  );


  not
  g166
  (
    n258,
    n64
  );


  buf
  g167
  (
    n302,
    n68
  );


  buf
  g168
  (
    n273,
    n41
  );


  not
  g169
  (
    n262,
    n31
  );


  not
  g170
  (
    n456,
    n134
  );


  not
  g171
  (
    n153,
    n60
  );


  not
  g172
  (
    n470,
    n116
  );


  buf
  g173
  (
    n430,
    n100
  );


  buf
  g174
  (
    n196,
    n30
  );


  buf
  g175
  (
    n202,
    n61
  );


  not
  g176
  (
    n227,
    n135
  );


  not
  g177
  (
    n332,
    n45
  );


  not
  g178
  (
    n211,
    n73
  );


  buf
  g179
  (
    n297,
    n139
  );


  buf
  g180
  (
    n405,
    n131
  );


  buf
  g181
  (
    n247,
    n122
  );


  not
  g182
  (
    n374,
    n83
  );


  buf
  g183
  (
    n246,
    n46
  );


  buf
  g184
  (
    n263,
    n58
  );


  buf
  g185
  (
    n152,
    n32
  );


  buf
  g186
  (
    n183,
    n126
  );


  buf
  g187
  (
    n432,
    n103
  );


  buf
  g188
  (
    n180,
    n123
  );


  buf
  g189
  (
    n174,
    n104
  );


  buf
  g190
  (
    n369,
    n33
  );


  not
  g191
  (
    n280,
    n38
  );


  not
  g192
  (
    n435,
    n98
  );


  not
  g193
  (
    n283,
    n108
  );


  buf
  g194
  (
    n445,
    n56
  );


  not
  g195
  (
    n321,
    n128
  );


  not
  g196
  (
    n178,
    n42
  );


  buf
  g197
  (
    n295,
    n141
  );


  not
  g198
  (
    n160,
    n92
  );


  buf
  g199
  (
    n451,
    n54
  );


  not
  g200
  (
    n253,
    n72
  );


  not
  g201
  (
    n356,
    n86
  );


  buf
  g202
  (
    n320,
    n79
  );


  buf
  g203
  (
    n158,
    n65
  );


  not
  g204
  (
    n225,
    n78
  );


  buf
  g205
  (
    n286,
    n112
  );


  not
  g206
  (
    n221,
    n53
  );


  not
  g207
  (
    n310,
    n37
  );


  buf
  g208
  (
    n318,
    n125
  );


  buf
  g209
  (
    n446,
    n141
  );


  buf
  g210
  (
    n327,
    n56
  );


  not
  g211
  (
    n210,
    n116
  );


  not
  g212
  (
    n342,
    n129
  );


  not
  g213
  (
    n226,
    n133
  );


  not
  g214
  (
    n471,
    n72
  );


  not
  g215
  (
    n441,
    n81
  );


  not
  g216
  (
    n172,
    n52
  );


  not
  g217
  (
    n329,
    n111
  );


  not
  g218
  (
    n336,
    n113
  );


  not
  g219
  (
    n385,
    n113
  );


  buf
  g220
  (
    n163,
    n74
  );


  not
  g221
  (
    n339,
    n44
  );


  buf
  g222
  (
    n287,
    n64
  );


  not
  g223
  (
    n315,
    n73
  );


  buf
  g224
  (
    n194,
    n72
  );


  not
  g225
  (
    n452,
    n94
  );


  buf
  g226
  (
    n311,
    n77
  );


  buf
  g227
  (
    n398,
    n69
  );


  buf
  g228
  (
    n387,
    n50
  );


  not
  g229
  (
    n249,
    n61
  );


  buf
  g230
  (
    n397,
    n60
  );


  not
  g231
  (
    n298,
    n134
  );


  not
  g232
  (
    n337,
    n66
  );


  buf
  g233
  (
    n468,
    n41
  );


  buf
  g234
  (
    n235,
    n67
  );


  buf
  g235
  (
    n303,
    n38
  );


  not
  g236
  (
    n475,
    n52
  );


  buf
  g237
  (
    n464,
    n68
  );


  buf
  g238
  (
    n453,
    n51
  );


  not
  g239
  (
    n219,
    n141
  );


  buf
  g240
  (
    n358,
    n86
  );


  buf
  g241
  (
    n477,
    n97
  );


  buf
  g242
  (
    n155,
    n138
  );


  not
  g243
  (
    n390,
    n120
  );


  not
  g244
  (
    n469,
    n93
  );


  not
  g245
  (
    n335,
    n107
  );


  not
  g246
  (
    n392,
    n131
  );


  buf
  g247
  (
    n443,
    n107
  );


  buf
  g248
  (
    n270,
    n116
  );


  not
  g249
  (
    n307,
    n118
  );


  not
  g250
  (
    n467,
    n49
  );


  buf
  g251
  (
    n371,
    n76
  );


  not
  g252
  (
    n402,
    n62
  );


  buf
  g253
  (
    n164,
    n69
  );


  buf
  g254
  (
    n238,
    n128
  );


  not
  g255
  (
    n457,
    n86
  );


  not
  g256
  (
    n326,
    n108
  );


  not
  g257
  (
    n150,
    n77
  );


  not
  g258
  (
    n296,
    n47
  );


  not
  g259
  (
    n460,
    n137
  );


  buf
  g260
  (
    n400,
    n96
  );


  buf
  g261
  (
    n423,
    n43
  );


  not
  g262
  (
    n418,
    n41
  );


  not
  g263
  (
    n345,
    n54
  );


  buf
  g264
  (
    n179,
    n47
  );


  buf
  g265
  (
    n166,
    n69
  );


  not
  g266
  (
    n482,
    n98
  );


  not
  g267
  (
    n473,
    n130
  );


  not
  g268
  (
    n319,
    n112
  );


  buf
  g269
  (
    n188,
    n122
  );


  not
  g270
  (
    n324,
    n70
  );


  buf
  g271
  (
    n368,
    n49
  );


  buf
  g272
  (
    n323,
    n75
  );


  not
  g273
  (
    n406,
    n59
  );


  buf
  g274
  (
    n293,
    n78
  );


  not
  g275
  (
    n412,
    n115
  );


  not
  g276
  (
    n284,
    n94
  );


  buf
  g277
  (
    n447,
    n57
  );


  buf
  g278
  (
    n256,
    n76
  );


  not
  g279
  (
    n190,
    n129
  );


  buf
  g280
  (
    n189,
    n99
  );


  not
  g281
  (
    n349,
    n35
  );


  buf
  g282
  (
    n448,
    n89
  );


  buf
  g283
  (
    n191,
    n102
  );


  not
  g284
  (
    n313,
    n32
  );


  not
  g285
  (
    n250,
    n138
  );


  buf
  g286
  (
    n428,
    n106
  );


  buf
  g287
  (
    n213,
    n70
  );


  not
  g288
  (
    n360,
    n74
  );


  buf
  g289
  (
    n401,
    n44
  );


  buf
  g290
  (
    n410,
    n118
  );


  not
  g291
  (
    n276,
    n93
  );


  not
  g292
  (
    n472,
    n125
  );


  buf
  g293
  (
    n156,
    n126
  );


  not
  g294
  (
    n197,
    n39
  );


  buf
  g295
  (
    n317,
    n108
  );


  buf
  g296
  (
    n277,
    n127
  );


  buf
  g297
  (
    n409,
    n100
  );


  not
  g298
  (
    n239,
    n60
  );


  not
  g299
  (
    n193,
    n84
  );


  not
  g300
  (
    n200,
    n105
  );


  buf
  g301
  (
    n395,
    n44
  );


  not
  g302
  (
    n427,
    n79
  );


  buf
  g303
  (
    n290,
    n135
  );


  buf
  g304
  (
    n328,
    n121
  );


  not
  g305
  (
    n248,
    n53
  );


  buf
  g306
  (
    n272,
    n53
  );


  buf
  g307
  (
    n289,
    n55
  );


  buf
  g308
  (
    n377,
    n37
  );


  buf
  g309
  (
    n278,
    n136
  );


  buf
  g310
  (
    n404,
    n127
  );


  not
  g311
  (
    n266,
    n64
  );


  not
  g312
  (
    n165,
    n37
  );


  buf
  g313
  (
    n267,
    n72
  );


  buf
  g314
  (
    n426,
    n132
  );


  buf
  g315
  (
    n234,
    n89
  );


  not
  g316
  (
    n338,
    n123
  );


  buf
  g317
  (
    n177,
    n58
  );


  buf
  g318
  (
    n378,
    n48
  );


  buf
  g319
  (
    n162,
    n85
  );


  not
  g320
  (
    n480,
    n91
  );


  buf
  g321
  (
    n173,
    n48
  );


  not
  g322
  (
    n416,
    n92
  );


  not
  g323
  (
    n271,
    n105
  );


  buf
  g324
  (
    n474,
    n32
  );


  not
  g325
  (
    n312,
    n41
  );


  buf
  g326
  (
    n260,
    n122
  );


  not
  g327
  (
    n192,
    n83
  );


  not
  g328
  (
    n433,
    n140
  );


  buf
  g329
  (
    n171,
    n36
  );


  buf
  g330
  (
    n244,
    n117
  );


  buf
  g331
  (
    n228,
    n73
  );


  not
  g332
  (
    n285,
    n132
  );


  not
  g333
  (
    n252,
    n103
  );


  not
  g334
  (
    n351,
    n106
  );


  buf
  g335
  (
    n366,
    n125
  );


  buf
  g336
  (
    n251,
    n42
  );


  not
  g337
  (
    n365,
    n81
  );


  buf
  g338
  (
    n241,
    n93
  );


  buf
  g339
  (
    n485,
    n83
  );


  buf
  g340
  (
    n463,
    n66
  );


  not
  g341
  (
    n431,
    n40
  );


  buf
  g342
  (
    n176,
    n33
  );


  buf
  g343
  (
    n450,
    n109
  );


  not
  g344
  (
    n434,
    n103
  );


  buf
  g345
  (
    n386,
    n38
  );


  buf
  g346
  (
    n408,
    n107
  );


  buf
  g347
  (
    n354,
    n82
  );


  not
  g348
  (
    n364,
    n138
  );


  not
  g349
  (
    n148,
    n133
  );


  not
  g350
  (
    n185,
    n36
  );


  not
  g351
  (
    n259,
    n48
  );


  buf
  g352
  (
    n292,
    n60
  );


  not
  g353
  (
    n206,
    n140
  );


  not
  g354
  (
    n146,
    n59
  );


  not
  g355
  (
    n478,
    n51
  );


  buf
  g356
  (
    n380,
    n105
  );


  not
  g357
  (
    n243,
    n43
  );


  buf
  g358
  (
    n201,
    n83
  );


  buf
  g359
  (
    n240,
    n115
  );


  not
  g360
  (
    n422,
    n61
  );


  not
  g361
  (
    n175,
    n125
  );


  buf
  g362
  (
    n454,
    n78
  );


  not
  g363
  (
    n403,
    n47
  );


  not
  g364
  (
    n184,
    n30
  );


  not
  g365
  (
    n352,
    n102
  );


  not
  g366
  (
    n341,
    n45
  );


  not
  g367
  (
    n411,
    n38
  );


  buf
  g368
  (
    n466,
    n117
  );


  buf
  g369
  (
    n182,
    n132
  );


  buf
  g370
  (
    n438,
    n129
  );


  not
  g371
  (
    n362,
    n123
  );


  buf
  g372
  (
    n444,
    n109
  );


  buf
  g373
  (
    n417,
    n80
  );


  not
  g374
  (
    n215,
    n34
  );


  buf
  g375
  (
    n216,
    n104
  );


  buf
  g376
  (
    n442,
    n50
  );


  not
  g377
  (
    n481,
    n35
  );


  not
  g378
  (
    n384,
    n78
  );


  not
  g379
  (
    n209,
    n94
  );


  buf
  g380
  (
    n396,
    n142
  );


  not
  g381
  (
    n340,
    n87
  );


  not
  g382
  (
    n372,
    n121
  );


  buf
  g383
  (
    n343,
    n112
  );


  buf
  g384
  (
    n195,
    n80
  );


  not
  g385
  (
    n257,
    n119
  );


  not
  g386
  (
    n233,
    n55
  );


  buf
  g387
  (
    n169,
    n33
  );


  buf
  g388
  (
    n373,
    n137
  );


  buf
  g389
  (
    n218,
    n34
  );


  buf
  g390
  (
    n306,
    n93
  );


  buf
  g391
  (
    n294,
    n119
  );


  not
  g392
  (
    n281,
    n58
  );


  not
  g393
  (
    n275,
    n34
  );


  not
  g394
  (
    n154,
    n55
  );


  buf
  g395
  (
    n419,
    n117
  );


  not
  g396
  (
    n461,
    n36
  );


  not
  g397
  (
    n159,
    n59
  );


  not
  g398
  (
    n367,
    n103
  );


  buf
  g399
  (
    n330,
    n120
  );


  buf
  g400
  (
    n254,
    n52
  );


  not
  g401
  (
    n203,
    n47
  );


  not
  g402
  (
    n261,
    n54
  );


  not
  g403
  (
    n291,
    n98
  );


  not
  g404
  (
    n420,
    n139
  );


  not
  g405
  (
    n264,
    n81
  );


  not
  g406
  (
    n439,
    n122
  );


  not
  g407
  (
    n483,
    n85
  );


  not
  g408
  (
    n167,
    n140
  );


  not
  g409
  (
    n348,
    n102
  );


  buf
  g410
  (
    n357,
    n111
  );


  not
  g411
  (
    n391,
    n90
  );


  buf
  g412
  (
    n245,
    n100
  );


  not
  g413
  (
    n459,
    n65
  );


  buf
  g414
  (
    n331,
    n99
  );


  buf
  g415
  (
    n440,
    n63
  );


  buf
  g416
  (
    n436,
    n77
  );


  not
  g417
  (
    n346,
    n121
  );


  and
  g418
  (
    n389,
    n30,
    n70
  );


  or
  g419
  (
    n314,
    n84,
    n85
  );


  nand
  g420
  (
    n223,
    n87,
    n70,
    n111,
    n81
  );


  or
  g421
  (
    n424,
    n35,
    n71,
    n57,
    n87
  );


  nor
  g422
  (
    n212,
    n43,
    n91,
    n119,
    n34
  );


  and
  g423
  (
    n198,
    n57,
    n95,
    n124,
    n69
  );


  xor
  g424
  (
    n168,
    n114,
    n136,
    n39,
    n90
  );


  and
  g425
  (
    n353,
    n63,
    n56,
    n91,
    n82
  );


  or
  g426
  (
    n407,
    n90,
    n77,
    n49,
    n99
  );


  nor
  g427
  (
    n265,
    n108,
    n104,
    n75,
    n128
  );


  and
  g428
  (
    n231,
    n131,
    n45,
    n118,
    n136
  );


  xor
  g429
  (
    n376,
    n58,
    n42,
    n91,
    n68
  );


  nand
  g430
  (
    n458,
    n43,
    n74,
    n133,
    n124
  );


  xor
  g431
  (
    n242,
    n32,
    n46,
    n75,
    n88
  );


  nand
  g432
  (
    n355,
    n84,
    n89,
    n85,
    n88
  );


  xnor
  g433
  (
    n334,
    n80,
    n99,
    n76,
    n112
  );


  and
  g434
  (
    n237,
    n67,
    n110,
    n126,
    n124
  );


  xnor
  g435
  (
    n300,
    n106,
    n71,
    n82,
    n109
  );


  xor
  g436
  (
    n205,
    n46,
    n71,
    n142,
    n61
  );


  xnor
  g437
  (
    n269,
    n75,
    n54,
    n67,
    n134
  );


  or
  g438
  (
    n462,
    n110,
    n39,
    n113,
    n65
  );


  nand
  g439
  (
    n421,
    n84,
    n139,
    n79,
    n73
  );


  nor
  g440
  (
    n305,
    n100,
    n44,
    n114,
    n95
  );


  and
  g441
  (
    n288,
    n110,
    n104,
    n133,
    n80
  );


  nor
  g442
  (
    n394,
    n117,
    n139,
    n66,
    n35
  );


  or
  g443
  (
    n383,
    n62,
    n107,
    n105,
    n116
  );


  nor
  g444
  (
    n170,
    n120,
    n92,
    n130,
    n79
  );


  or
  g445
  (
    n479,
    n33,
    n40,
    n36,
    n94
  );


  nand
  g446
  (
    n333,
    n88,
    n63,
    n50,
    n132
  );


  nor
  g447
  (
    n322,
    n135,
    n123,
    n106,
    n118
  );


  or
  g448
  (
    n382,
    n96,
    n101,
    n31
  );


  nand
  g449
  (
    n429,
    n102,
    n109,
    n134,
    n49
  );


  xor
  g450
  (
    n199,
    n115,
    n71,
    n55,
    n62
  );


  and
  g451
  (
    n282,
    n129,
    n115,
    n97,
    n67
  );


  xnor
  g452
  (
    n437,
    n101,
    n119,
    n114
  );


  nand
  g453
  (
    n207,
    n89,
    n110,
    n63,
    n135
  );


  xor
  g454
  (
    n425,
    n101,
    n127,
    n31,
    n51
  );


  xnor
  g455
  (
    n204,
    n42,
    n68,
    n39,
    n130
  );


  buf
  g456
  (
    n694,
    n404
  );


  buf
  g457
  (
    n744,
    n398
  );


  buf
  g458
  (
    n778,
    n404
  );


  not
  g459
  (
    n734,
    n423
  );


  buf
  g460
  (
    n768,
    n401
  );


  buf
  g461
  (
    n736,
    n384
  );


  not
  g462
  (
    n611,
    n427
  );


  not
  g463
  (
    n870,
    n167
  );


  not
  g464
  (
    n587,
    n265
  );


  not
  g465
  (
    KeyWire_0_1,
    n207
  );


  buf
  g466
  (
    n505,
    n279
  );


  buf
  g467
  (
    n780,
    n193
  );


  not
  g468
  (
    n843,
    n386
  );


  buf
  g469
  (
    n729,
    n316
  );


  not
  g470
  (
    n650,
    n413
  );


  not
  g471
  (
    n579,
    n394
  );


  not
  g472
  (
    n837,
    n250
  );


  buf
  g473
  (
    n871,
    n396
  );


  not
  g474
  (
    n687,
    n390
  );


  not
  g475
  (
    n743,
    n253
  );


  not
  g476
  (
    n765,
    n262
  );


  buf
  g477
  (
    n798,
    n405
  );


  buf
  g478
  (
    n707,
    n175
  );


  not
  g479
  (
    n868,
    n194
  );


  buf
  g480
  (
    n544,
    n376
  );


  buf
  g481
  (
    n790,
    n391
  );


  buf
  g482
  (
    n561,
    n156
  );


  not
  g483
  (
    n677,
    n417
  );


  not
  g484
  (
    n488,
    n293
  );


  buf
  g485
  (
    n819,
    n407
  );


  buf
  g486
  (
    n844,
    n411
  );


  not
  g487
  (
    n704,
    n273
  );


  not
  g488
  (
    n738,
    n405
  );


  not
  g489
  (
    n892,
    n386
  );


  not
  g490
  (
    n716,
    n351
  );


  buf
  g491
  (
    n532,
    n161
  );


  not
  g492
  (
    n583,
    n359
  );


  not
  g493
  (
    n821,
    n274
  );


  not
  g494
  (
    n801,
    n423
  );


  not
  g495
  (
    n570,
    n393
  );


  not
  g496
  (
    n697,
    n245
  );


  not
  g497
  (
    n847,
    n246
  );


  buf
  g498
  (
    n572,
    n260
  );


  not
  g499
  (
    n889,
    n395
  );


  not
  g500
  (
    n664,
    n409
  );


  not
  g501
  (
    n711,
    n223
  );


  buf
  g502
  (
    n826,
    n409
  );


  not
  g503
  (
    n761,
    n390
  );


  buf
  g504
  (
    n618,
    n339
  );


  buf
  g505
  (
    n688,
    n251
  );


  not
  g506
  (
    n635,
    n237
  );


  not
  g507
  (
    n856,
    n415
  );


  buf
  g508
  (
    n537,
    n181
  );


  buf
  g509
  (
    n574,
    n389
  );


  buf
  g510
  (
    KeyWire_0_0,
    n416
  );


  not
  g511
  (
    n540,
    n312
  );


  buf
  g512
  (
    n846,
    n195
  );


  not
  g513
  (
    n756,
    n426
  );


  buf
  g514
  (
    n838,
    n426
  );


  buf
  g515
  (
    n816,
    n399
  );


  buf
  g516
  (
    n810,
    n154
  );


  not
  g517
  (
    n634,
    n384
  );


  not
  g518
  (
    n735,
    n390
  );


  buf
  g519
  (
    n865,
    n390
  );


  buf
  g520
  (
    n722,
    n210
  );


  buf
  g521
  (
    n516,
    n290
  );


  buf
  g522
  (
    n667,
    n385
  );


  buf
  g523
  (
    n828,
    n428
  );


  buf
  g524
  (
    n695,
    n203
  );


  buf
  g525
  (
    n550,
    n352
  );


  buf
  g526
  (
    n669,
    n340
  );


  not
  g527
  (
    n513,
    n247
  );


  not
  g528
  (
    n775,
    n187
  );


  buf
  g529
  (
    n519,
    n220
  );


  not
  g530
  (
    n774,
    n403
  );


  not
  g531
  (
    n749,
    n304
  );


  not
  g532
  (
    n725,
    n377
  );


  buf
  g533
  (
    n526,
    n170
  );


  buf
  g534
  (
    n642,
    n147
  );


  buf
  g535
  (
    n811,
    n397
  );


  buf
  g536
  (
    n896,
    n424
  );


  buf
  g537
  (
    n829,
    n363
  );


  not
  g538
  (
    n872,
    n311
  );


  buf
  g539
  (
    n733,
    n149
  );


  not
  g540
  (
    n580,
    n177
  );


  buf
  g541
  (
    n739,
    n309
  );


  not
  g542
  (
    n556,
    n392
  );


  not
  g543
  (
    n804,
    n257
  );


  buf
  g544
  (
    n602,
    n426
  );


  buf
  g545
  (
    n782,
    n383
  );


  not
  g546
  (
    n612,
    n414
  );


  buf
  g547
  (
    n569,
    n180
  );


  not
  g548
  (
    n663,
    n414
  );


  buf
  g549
  (
    n900,
    n422
  );


  buf
  g550
  (
    n632,
    n345
  );


  buf
  g551
  (
    n575,
    n393
  );


  buf
  g552
  (
    n496,
    n353
  );


  buf
  g553
  (
    n533,
    n409
  );


  not
  g554
  (
    n806,
    n252
  );


  not
  g555
  (
    n636,
    n396
  );


  buf
  g556
  (
    n509,
    n385
  );


  not
  g557
  (
    n795,
    n416
  );


  buf
  g558
  (
    n495,
    n291
  );


  not
  g559
  (
    n709,
    n360
  );


  buf
  g560
  (
    n820,
    n423
  );


  not
  g561
  (
    n771,
    n163
  );


  not
  g562
  (
    n622,
    n402
  );


  not
  g563
  (
    n607,
    n385
  );


  buf
  g564
  (
    n620,
    n242
  );


  not
  g565
  (
    n873,
    n238
  );


  not
  g566
  (
    n777,
    n403
  );


  buf
  g567
  (
    n755,
    n389
  );


  not
  g568
  (
    n623,
    n387
  );


  buf
  g569
  (
    n718,
    n399
  );


  not
  g570
  (
    n888,
    n401
  );


  buf
  g571
  (
    n728,
    n427
  );


  buf
  g572
  (
    n874,
    n424
  );


  buf
  g573
  (
    n672,
    n400
  );


  buf
  g574
  (
    n747,
    n406
  );


  not
  g575
  (
    n813,
    n162
  );


  not
  g576
  (
    n676,
    n296
  );


  not
  g577
  (
    n603,
    n278
  );


  not
  g578
  (
    n880,
    n188
  );


  buf
  g579
  (
    n646,
    n399
  );


  not
  g580
  (
    n818,
    n189
  );


  buf
  g581
  (
    n593,
    n408
  );


  buf
  g582
  (
    n742,
    n281
  );


  not
  g583
  (
    n521,
    n349
  );


  not
  g584
  (
    n489,
    n157
  );


  buf
  g585
  (
    n643,
    n153
  );


  not
  g586
  (
    n770,
    n357
  );


  not
  g587
  (
    n604,
    n411
  );


  not
  g588
  (
    n702,
    n179
  );


  buf
  g589
  (
    n668,
    n419
  );


  not
  g590
  (
    n898,
    n323
  );


  not
  g591
  (
    n754,
    n343
  );


  not
  g592
  (
    n701,
    n307
  );


  buf
  g593
  (
    n654,
    n225
  );


  not
  g594
  (
    n705,
    n411
  );


  buf
  g595
  (
    n784,
    n425
  );


  buf
  g596
  (
    n762,
    n308
  );


  not
  g597
  (
    n527,
    n303
  );


  not
  g598
  (
    n767,
    n422
  );


  buf
  g599
  (
    n730,
    n319
  );


  not
  g600
  (
    n609,
    n356
  );


  buf
  g601
  (
    n662,
    n428
  );


  buf
  g602
  (
    n524,
    n218
  );


  not
  g603
  (
    n564,
    n403
  );


  buf
  g604
  (
    n599,
    n322
  );


  not
  g605
  (
    n605,
    n213
  );


  not
  g606
  (
    n682,
    n239
  );


  buf
  g607
  (
    n535,
    n405
  );


  buf
  g608
  (
    n842,
    n152
  );


  buf
  g609
  (
    n582,
    n346
  );


  buf
  g610
  (
    n512,
    n151
  );


  not
  g611
  (
    n753,
    n350
  );


  not
  g612
  (
    n504,
    n324
  );


  buf
  g613
  (
    n671,
    n327
  );


  buf
  g614
  (
    n867,
    n371
  );


  buf
  g615
  (
    n853,
    n400
  );


  buf
  g616
  (
    n502,
    n396
  );


  not
  g617
  (
    n789,
    n249
  );


  buf
  g618
  (
    n510,
    n336
  );


  buf
  g619
  (
    n503,
    n417
  );


  buf
  g620
  (
    n538,
    n227
  );


  buf
  g621
  (
    n759,
    n413
  );


  buf
  g622
  (
    n800,
    n155
  );


  not
  g623
  (
    n520,
    n320
  );


  not
  g624
  (
    n491,
    n298
  );


  not
  g625
  (
    n893,
    n334
  );


  not
  g626
  (
    n823,
    n384
  );


  buf
  g627
  (
    n490,
    n190
  );


  buf
  g628
  (
    n629,
    n420
  );


  buf
  g629
  (
    n792,
    n241
  );


  buf
  g630
  (
    n661,
    n410
  );


  not
  g631
  (
    n670,
    n372
  );


  not
  g632
  (
    n547,
    n263
  );


  not
  g633
  (
    n536,
    n410
  );


  buf
  g634
  (
    n831,
    n416
  );


  buf
  g635
  (
    n560,
    n386
  );


  buf
  g636
  (
    n827,
    n407
  );


  not
  g637
  (
    n608,
    n276
  );


  buf
  g638
  (
    n657,
    n184
  );


  buf
  g639
  (
    n684,
    n285
  );


  buf
  g640
  (
    n788,
    n292
  );


  buf
  g641
  (
    n568,
    n318
  );


  buf
  g642
  (
    n731,
    n268
  );


  not
  g643
  (
    n857,
    n295
  );


  buf
  g644
  (
    n653,
    n289
  );


  buf
  g645
  (
    n647,
    n418
  );


  not
  g646
  (
    n760,
    n196
  );


  buf
  g647
  (
    n786,
    n174
  );


  buf
  g648
  (
    n641,
    n400
  );


  not
  g649
  (
    n703,
    n169
  );


  not
  g650
  (
    n522,
    n172
  );


  not
  g651
  (
    n508,
    n412
  );


  not
  g652
  (
    n894,
    n389
  );


  not
  g653
  (
    n895,
    n407
  );


  buf
  g654
  (
    n617,
    n421
  );


  not
  g655
  (
    n854,
    n277
  );


  buf
  g656
  (
    n863,
    n406
  );


  buf
  g657
  (
    n499,
    n325
  );


  not
  g658
  (
    n876,
    n414
  );


  buf
  g659
  (
    n683,
    n214
  );


  buf
  g660
  (
    n713,
    n420
  );


  buf
  g661
  (
    n825,
    n321
  );


  not
  g662
  (
    n884,
    n397
  );


  not
  g663
  (
    n793,
    n226
  );


  buf
  g664
  (
    n883,
    n398
  );


  not
  g665
  (
    n652,
    n408
  );


  not
  g666
  (
    n737,
    n310
  );


  not
  g667
  (
    KeyWire_0_9,
    n148
  );


  not
  g668
  (
    n757,
    n422
  );


  buf
  g669
  (
    n645,
    n424
  );


  not
  g670
  (
    n591,
    n219
  );


  buf
  g671
  (
    n809,
    n393
  );


  buf
  g672
  (
    n781,
    n229
  );


  not
  g673
  (
    n808,
    n178
  );


  not
  g674
  (
    n553,
    n171
  );


  buf
  g675
  (
    n594,
    n305
  );


  buf
  g676
  (
    n691,
    n266
  );


  not
  g677
  (
    n835,
    n410
  );


  buf
  g678
  (
    n833,
    n301
  );


  not
  g679
  (
    n500,
    n287
  );


  not
  g680
  (
    n518,
    n370
  );


  not
  g681
  (
    n541,
    n333
  );


  not
  g682
  (
    n890,
    n387
  );


  buf
  g683
  (
    n710,
    n355
  );


  not
  g684
  (
    n858,
    n388
  );


  not
  g685
  (
    n861,
    n389
  );


  not
  g686
  (
    n534,
    n366
  );


  buf
  g687
  (
    n830,
    n420
  );


  buf
  g688
  (
    n769,
    n168
  );


  not
  g689
  (
    n673,
    n407
  );


  buf
  g690
  (
    n891,
    n381
  );


  buf
  g691
  (
    n552,
    n259
  );


  not
  g692
  (
    n610,
    n330
  );


  buf
  g693
  (
    n581,
    n215
  );


  buf
  g694
  (
    n764,
    n335
  );


  not
  g695
  (
    n839,
    n234
  );


  not
  g696
  (
    n794,
    n392
  );


  not
  g697
  (
    n746,
    n269
  );


  buf
  g698
  (
    n659,
    n337
  );


  buf
  g699
  (
    n555,
    n361
  );


  buf
  g700
  (
    n562,
    n342
  );


  buf
  g701
  (
    n866,
    n386
  );


  buf
  g702
  (
    n748,
    n198
  );


  not
  g703
  (
    n766,
    n314
  );


  buf
  g704
  (
    n752,
    n255
  );


  buf
  g705
  (
    n660,
    n385
  );


  not
  g706
  (
    n805,
    n424
  );


  buf
  g707
  (
    n625,
    n412
  );


  not
  g708
  (
    n577,
    n397
  );


  buf
  g709
  (
    n644,
    n419
  );


  not
  g710
  (
    n741,
    n329
  );


  not
  g711
  (
    n523,
    n186
  );


  not
  g712
  (
    n595,
    n421
  );


  not
  g713
  (
    n848,
    n422
  );


  buf
  g714
  (
    n542,
    n197
  );


  not
  g715
  (
    n675,
    n415
  );


  buf
  g716
  (
    n649,
    n425
  );


  not
  g717
  (
    n708,
    n400
  );


  not
  g718
  (
    n530,
    n406
  );


  buf
  g719
  (
    n726,
    n224
  );


  buf
  g720
  (
    n578,
    n373
  );


  not
  g721
  (
    n627,
    n300
  );


  buf
  g722
  (
    n517,
    n331
  );


  buf
  g723
  (
    n565,
    n399
  );


  buf
  g724
  (
    n686,
    n272
  );


  not
  g725
  (
    n814,
    n209
  );


  not
  g726
  (
    n601,
    n379
  );


  buf
  g727
  (
    n897,
    n280
  );


  not
  g728
  (
    n590,
    n254
  );


  buf
  g729
  (
    n834,
    n176
  );


  not
  g730
  (
    n548,
    n394
  );


  buf
  g731
  (
    n557,
    n212
  );


  not
  g732
  (
    n740,
    n317
  );


  not
  g733
  (
    n514,
    n425
  );


  not
  g734
  (
    n549,
    n391
  );


  buf
  g735
  (
    n850,
    n396
  );


  not
  g736
  (
    n717,
    n358
  );


  not
  g737
  (
    n855,
    n202
  );


  buf
  g738
  (
    n696,
    n294
  );


  not
  g739
  (
    n515,
    n408
  );


  not
  g740
  (
    n878,
    n418
  );


  buf
  g741
  (
    n706,
    n362
  );


  not
  g742
  (
    n885,
    n423
  );


  not
  g743
  (
    n674,
    n200
  );


  buf
  g744
  (
    n586,
    n221
  );


  buf
  g745
  (
    n724,
    n387
  );


  not
  g746
  (
    n638,
    n412
  );


  not
  g747
  (
    n531,
    n326
  );


  not
  g748
  (
    n751,
    n159
  );


  buf
  g749
  (
    n877,
    n313
  );


  not
  g750
  (
    n807,
    n404
  );


  not
  g751
  (
    n699,
    n282
  );


  buf
  g752
  (
    n773,
    n419
  );


  not
  g753
  (
    n822,
    n374
  );


  not
  g754
  (
    n614,
    n270
  );


  buf
  g755
  (
    n589,
    n231
  );


  not
  g756
  (
    n681,
    n344
  );


  not
  g757
  (
    n630,
    n387
  );


  buf
  g758
  (
    n529,
    n417
  );


  not
  g759
  (
    n640,
    n204
  );


  buf
  g760
  (
    n576,
    n388
  );


  not
  g761
  (
    n869,
    n182
  );


  not
  g762
  (
    n723,
    n401
  );


  buf
  g763
  (
    n597,
    n418
  );


  not
  g764
  (
    n815,
    n367
  );


  not
  g765
  (
    n656,
    n375
  );


  not
  g766
  (
    n639,
    n414
  );


  buf
  g767
  (
    n700,
    n427
  );


  not
  g768
  (
    n507,
    n185
  );


  buf
  g769
  (
    n501,
    n315
  );


  not
  g770
  (
    n616,
    n395
  );


  buf
  g771
  (
    n692,
    n397
  );


  buf
  g772
  (
    n679,
    n415
  );


  not
  g773
  (
    n860,
    n398
  );


  buf
  g774
  (
    n882,
    n164
  );


  not
  g775
  (
    n797,
    n267
  );


  buf
  g776
  (
    n841,
    n402
  );


  buf
  g777
  (
    n779,
    n165
  );


  not
  g778
  (
    n628,
    n283
  );


  buf
  g779
  (
    n685,
    n415
  );


  buf
  g780
  (
    n836,
    n425
  );


  not
  g781
  (
    n812,
    n417
  );


  buf
  g782
  (
    n799,
    n408
  );


  not
  g783
  (
    n758,
    n302
  );


  not
  g784
  (
    n732,
    n388
  );


  not
  g785
  (
    n763,
    n240
  );


  buf
  g786
  (
    n633,
    n392
  );


  buf
  g787
  (
    n545,
    n393
  );


  not
  g788
  (
    n680,
    n416
  );


  not
  g789
  (
    n487,
    n392
  );


  not
  g790
  (
    n651,
    n230
  );


  buf
  g791
  (
    n498,
    n286
  );


  not
  g792
  (
    n624,
    n232
  );


  not
  g793
  (
    n566,
    n158
  );


  buf
  g794
  (
    n772,
    n297
  );


  not
  g795
  (
    n497,
    n211
  );


  not
  g796
  (
    n621,
    n394
  );


  not
  g797
  (
    n783,
    n412
  );


  not
  g798
  (
    n719,
    n328
  );


  buf
  g799
  (
    n849,
    n192
  );


  buf
  g800
  (
    n539,
    n199
  );


  buf
  g801
  (
    n592,
    n348
  );


  not
  g802
  (
    n720,
    n338
  );


  not
  g803
  (
    n558,
    n403
  );


  not
  g804
  (
    n859,
    n391
  );


  not
  g805
  (
    n824,
    n365
  );


  buf
  g806
  (
    n666,
    n391
  );


  buf
  g807
  (
    n588,
    n368
  );


  not
  g808
  (
    n506,
    n428
  );


  buf
  g809
  (
    n875,
    n208
  );


  buf
  g810
  (
    n886,
    n413
  );


  not
  g811
  (
    n840,
    n306
  );


  not
  g812
  (
    n693,
    n288
  );


  buf
  g813
  (
    n546,
    n256
  );


  not
  g814
  (
    n492,
    n341
  );


  buf
  g815
  (
    n585,
    n216
  );


  not
  g816
  (
    n862,
    n236
  );


  buf
  g817
  (
    n787,
    n347
  );


  buf
  g818
  (
    n714,
    n402
  );


  not
  g819
  (
    n803,
    n404
  );


  not
  g820
  (
    n802,
    n418
  );


  not
  g821
  (
    n899,
    n406
  );


  buf
  g822
  (
    n600,
    n150
  );


  not
  g823
  (
    n690,
    n410
  );


  not
  g824
  (
    n637,
    n426
  );


  buf
  g825
  (
    n776,
    n244
  );


  not
  g826
  (
    n615,
    n419
  );


  buf
  g827
  (
    n887,
    n388
  );


  buf
  g828
  (
    n832,
    n201
  );


  buf
  g829
  (
    n712,
    n369
  );


  buf
  g830
  (
    n493,
    n146
  );


  not
  g831
  (
    n750,
    n183
  );


  buf
  g832
  (
    n573,
    n261
  );


  buf
  g833
  (
    n598,
    n284
  );


  not
  g834
  (
    n689,
    n166
  );


  buf
  g835
  (
    n881,
    n354
  );


  buf
  g836
  (
    n785,
    n395
  );


  buf
  g837
  (
    n626,
    n217
  );


  not
  g838
  (
    n791,
    n380
  );


  buf
  g839
  (
    n528,
    n409
  );


  buf
  g840
  (
    n551,
    n160
  );


  not
  g841
  (
    n554,
    n421
  );


  buf
  g842
  (
    n796,
    n411
  );


  not
  g843
  (
    n613,
    n243
  );


  not
  g844
  (
    n631,
    n248
  );


  not
  g845
  (
    n678,
    n275
  );


  buf
  g846
  (
    n715,
    n332
  );


  buf
  g847
  (
    n559,
    n394
  );


  not
  g848
  (
    n494,
    n206
  );


  buf
  g849
  (
    n619,
    n233
  );


  buf
  g850
  (
    n852,
    n382
  );


  buf
  g851
  (
    n745,
    n191
  );


  not
  g852
  (
    n606,
    n258
  );


  not
  g853
  (
    n567,
    n235
  );


  buf
  g854
  (
    n525,
    n421
  );


  not
  g855
  (
    n698,
    n395
  );


  buf
  g856
  (
    n584,
    n228
  );


  not
  g857
  (
    n817,
    n364
  );


  not
  g858
  (
    n879,
    n205
  );


  not
  g859
  (
    n655,
    n402
  );


  buf
  g860
  (
    n511,
    n413
  );


  not
  g861
  (
    n864,
    n405
  );


  buf
  g862
  (
    n596,
    n378
  );


  buf
  g863
  (
    n543,
    n401
  );


  not
  g864
  (
    n486,
    n222
  );


  buf
  g865
  (
    n721,
    n420
  );


  not
  g866
  (
    n851,
    n384
  );


  buf
  g867
  (
    n571,
    n271
  );


  buf
  g868
  (
    n845,
    n173
  );


  buf
  g869
  (
    n648,
    n299
  );


  nor
  g870
  (
    n665,
    n398,
    n264,
    n428,
    n427
  );


  not
  g871
  (
    n971,
    n507
  );


  not
  g872
  (
    n990,
    n580
  );


  buf
  g873
  (
    n978,
    n553
  );


  buf
  g874
  (
    n970,
    n546
  );


  buf
  g875
  (
    n911,
    n494
  );


  not
  g876
  (
    n965,
    n554
  );


  buf
  g877
  (
    n995,
    n490
  );


  not
  g878
  (
    n1002,
    n583
  );


  not
  g879
  (
    n916,
    n536
  );


  not
  g880
  (
    n950,
    n581
  );


  not
  g881
  (
    n951,
    n533
  );


  buf
  g882
  (
    n964,
    n585
  );


  not
  g883
  (
    n992,
    n543
  );


  not
  g884
  (
    n979,
    n556
  );


  buf
  g885
  (
    n943,
    n529
  );


  not
  g886
  (
    n901,
    n565
  );


  buf
  g887
  (
    n927,
    n551
  );


  buf
  g888
  (
    n920,
    n515
  );


  not
  g889
  (
    n981,
    n535
  );


  buf
  g890
  (
    n905,
    n509
  );


  buf
  g891
  (
    n994,
    n549
  );


  not
  g892
  (
    n993,
    n517
  );


  buf
  g893
  (
    n949,
    n538
  );


  buf
  g894
  (
    n945,
    n492
  );


  not
  g895
  (
    n963,
    n504
  );


  not
  g896
  (
    n968,
    n545
  );


  buf
  g897
  (
    n915,
    n486
  );


  not
  g898
  (
    n926,
    n510
  );


  not
  g899
  (
    n934,
    n491
  );


  buf
  g900
  (
    n919,
    n557
  );


  not
  g901
  (
    n947,
    n495
  );


  buf
  g902
  (
    n910,
    n587
  );


  buf
  g903
  (
    n912,
    n572
  );


  not
  g904
  (
    n976,
    n567
  );


  buf
  g905
  (
    n983,
    n539
  );


  not
  g906
  (
    n998,
    n571
  );


  not
  g907
  (
    n942,
    n552
  );


  not
  g908
  (
    n957,
    n576
  );


  buf
  g909
  (
    n972,
    n577
  );


  buf
  g910
  (
    n953,
    n511
  );


  buf
  g911
  (
    n958,
    n518
  );


  not
  g912
  (
    n975,
    n498
  );


  not
  g913
  (
    n997,
    n534
  );


  not
  g914
  (
    n967,
    n582
  );


  not
  g915
  (
    n1001,
    n531
  );


  not
  g916
  (
    n908,
    n569
  );


  buf
  g917
  (
    n961,
    n542
  );


  buf
  g918
  (
    n955,
    n516
  );


  not
  g919
  (
    n952,
    n520
  );


  not
  g920
  (
    n902,
    n521
  );


  not
  g921
  (
    n924,
    n586
  );


  buf
  g922
  (
    n914,
    n548
  );


  not
  g923
  (
    n966,
    n560
  );


  not
  g924
  (
    n969,
    n574
  );


  not
  g925
  (
    n921,
    n532
  );


  buf
  g926
  (
    n960,
    n506
  );


  buf
  g927
  (
    n1000,
    n530
  );


  buf
  g928
  (
    n913,
    n513
  );


  buf
  g929
  (
    n936,
    n555
  );


  not
  g930
  (
    n903,
    n489
  );


  not
  g931
  (
    n980,
    n575
  );


  buf
  g932
  (
    n918,
    n505
  );


  buf
  g933
  (
    n904,
    n525
  );


  not
  g934
  (
    n988,
    n514
  );


  not
  g935
  (
    n946,
    n566
  );


  not
  g936
  (
    n948,
    n558
  );


  not
  g937
  (
    n932,
    n564
  );


  not
  g938
  (
    n974,
    n537
  );


  not
  g939
  (
    n907,
    n528
  );


  buf
  g940
  (
    n933,
    n527
  );


  buf
  g941
  (
    n923,
    n561
  );


  not
  g942
  (
    n938,
    n487
  );


  not
  g943
  (
    n956,
    n496
  );


  not
  g944
  (
    n985,
    n540
  );


  buf
  g945
  (
    n929,
    n500
  );


  buf
  g946
  (
    n922,
    n544
  );


  buf
  g947
  (
    n996,
    n522
  );


  not
  g948
  (
    n930,
    n501
  );


  not
  g949
  (
    n940,
    n493
  );


  not
  g950
  (
    n928,
    n570
  );


  not
  g951
  (
    n986,
    n488
  );


  not
  g952
  (
    n987,
    n568
  );


  not
  g953
  (
    n925,
    n559
  );


  buf
  g954
  (
    n977,
    n541
  );


  buf
  g955
  (
    n959,
    n573
  );


  not
  g956
  (
    n935,
    n579
  );


  buf
  g957
  (
    n989,
    n524
  );


  buf
  g958
  (
    n991,
    n502
  );


  buf
  g959
  (
    KeyWire_0_6,
    n547
  );


  buf
  g960
  (
    n931,
    n508
  );


  buf
  g961
  (
    n937,
    n578
  );


  buf
  g962
  (
    n954,
    n497
  );


  buf
  g963
  (
    n909,
    n584
  );


  buf
  g964
  (
    n984,
    n512
  );


  not
  g965
  (
    n906,
    n526
  );


  buf
  g966
  (
    n973,
    n550
  );


  not
  g967
  (
    n939,
    n523
  );


  buf
  g968
  (
    n962,
    n562
  );


  not
  g969
  (
    n982,
    n519
  );


  not
  g970
  (
    n999,
    n503
  );


  buf
  g971
  (
    n941,
    n563
  );


  not
  g972
  (
    n917,
    n499
  );


  nor
  g973
  (
    n1024,
    n902,
    n908,
    n921
  );


  xor
  g974
  (
    n1010,
    n906,
    n919,
    n904,
    n914
  );


  or
  g975
  (
    n1031,
    n929,
    n923,
    n924,
    n915
  );


  or
  g976
  (
    n1026,
    n429,
    n912,
    n906,
    n929
  );


  nand
  g977
  (
    n1008,
    n929,
    n922,
    n909,
    n913
  );


  and
  g978
  (
    n1022,
    n921,
    n910,
    n906,
    n905
  );


  nand
  g979
  (
    n1015,
    n901,
    n916,
    n910,
    n907
  );


  nand
  g980
  (
    n1007,
    n916,
    n928,
    n918,
    n919
  );


  or
  g981
  (
    n1014,
    n429,
    n908,
    n906,
    n921
  );


  nor
  g982
  (
    n1013,
    n918,
    n915,
    n907,
    n925
  );


  xnor
  g983
  (
    n1021,
    n925,
    n910,
    n903,
    n928
  );


  nand
  g984
  (
    n1028,
    n918,
    n921,
    n902,
    n924
  );


  or
  g985
  (
    n1005,
    n909,
    n903,
    n914,
    n913
  );


  nor
  g986
  (
    n1003,
    n930,
    n919,
    n908,
    n903
  );


  xor
  g987
  (
    n1025,
    n905,
    n912,
    n926,
    n920
  );


  and
  g988
  (
    n1023,
    n904,
    n920,
    n902,
    n913
  );


  and
  g989
  (
    n1006,
    n901,
    n922,
    n917
  );


  or
  g990
  (
    n1020,
    n909,
    n912,
    n922,
    n911
  );


  and
  g991
  (
    n1012,
    n926,
    n917,
    n911
  );


  and
  g992
  (
    n1009,
    n928,
    n907,
    n927,
    n915
  );


  xor
  g993
  (
    n1019,
    n913,
    n927,
    n905,
    n911
  );


  xnor
  g994
  (
    n1016,
    n926,
    n925,
    n923,
    n903
  );


  xnor
  g995
  (
    n1032,
    n914,
    n928,
    n923,
    n912
  );


  or
  g996
  (
    n1017,
    n916,
    n905,
    n909,
    n926
  );


  and
  g997
  (
    n1004,
    n922,
    n901,
    n920,
    n923
  );


  xor
  g998
  (
    n1027,
    n929,
    n907,
    n915,
    n916
  );


  or
  g999
  (
    n1030,
    n910,
    n918,
    n904,
    n902
  );


  nand
  g1000
  (
    n1018,
    n914,
    n919,
    n920,
    n924
  );


  and
  g1001
  (
    n1029,
    n925,
    n927,
    n924
  );


  and
  g1002
  (
    n1011,
    n917,
    n901,
    n904,
    n930
  );


  buf
  g1003
  (
    n1035,
    n1030
  );


  buf
  g1004
  (
    n1034,
    n1032
  );


  not
  g1005
  (
    n1033,
    n1031
  );


  not
  g1006
  (
    n1036,
    n1029
  );


  nor
  g1007
  (
    n1044,
    n441,
    n429,
    n434,
    n432
  );


  nor
  g1008
  (
    n1045,
    n436,
    n431,
    n1033
  );


  xor
  g1009
  (
    n1041,
    n1036,
    n430,
    n439,
    n437
  );


  nand
  g1010
  (
    n1049,
    n438,
    n431,
    n1034,
    n435
  );


  xor
  g1011
  (
    n1051,
    n440,
    n1033,
    n433,
    n439
  );


  and
  g1012
  (
    n1037,
    n434,
    n432,
    n435
  );


  nand
  g1013
  (
    n1043,
    n441,
    n434,
    n1036,
    n438
  );


  or
  g1014
  (
    n1047,
    n437,
    n439,
    n1035,
    n1034
  );


  xnor
  g1015
  (
    n1048,
    n1035,
    n438,
    n433
  );


  nand
  g1016
  (
    n1042,
    n430,
    n440,
    n439
  );


  nor
  g1017
  (
    n1052,
    n436,
    n1033,
    n1036,
    n433
  );


  and
  g1018
  (
    n1038,
    n437,
    n436,
    n430
  );


  and
  g1019
  (
    n1046,
    n436,
    n435,
    n1035
  );


  xor
  g1020
  (
    n1040,
    n433,
    n429,
    n440,
    n1036
  );


  xnor
  g1021
  (
    n1039,
    n1034,
    n432,
    n431
  );


  xnor
  g1022
  (
    n1050,
    n432,
    n1034,
    n434,
    n437
  );


  xnor
  g1023
  (
    n1076,
    n718,
    n632,
    n1049,
    n593
  );


  xnor
  g1024
  (
    n1066,
    n1041,
    n736,
    n734,
    n694
  );


  nand
  g1025
  (
    n1073,
    n1045,
    n1045,
    n592,
    n678
  );


  and
  g1026
  (
    n1098,
    n696,
    n710,
    n743,
    n760
  );


  nand
  g1027
  (
    n1095,
    n607,
    n711,
    n1043,
    n724
  );


  nand
  g1028
  (
    n1086,
    n716,
    n1045,
    n1037,
    n657
  );


  xnor
  g1029
  (
    n1078,
    n722,
    n733,
    n762,
    n1038
  );


  xor
  g1030
  (
    n1088,
    n640,
    n641,
    n1047,
    n658
  );


  xnor
  g1031
  (
    n1058,
    n609,
    n625,
    n706,
    n1038
  );


  nand
  g1032
  (
    n1093,
    n613,
    n766,
    n590,
    n699
  );


  xor
  g1033
  (
    n1089,
    n631,
    n611,
    n708,
    n673
  );


  nor
  g1034
  (
    n1094,
    n660,
    n1049,
    n712,
    n633
  );


  xnor
  g1035
  (
    n1069,
    n667,
    n603,
    n1040,
    n753
  );


  or
  g1036
  (
    n1071,
    n707,
    n644,
    n1050,
    n1044
  );


  or
  g1037
  (
    n1092,
    n627,
    n680,
    n1051,
    n765
  );


  or
  g1038
  (
    n1075,
    n1041,
    n630,
    n747,
    n648
  );


  nand
  g1039
  (
    n1068,
    n705,
    n1042,
    n1040,
    n765
  );


  nand
  g1040
  (
    n1061,
    n721,
    n1041,
    n727,
    n758
  );


  nor
  g1041
  (
    n1084,
    n1052,
    n672,
    n684,
    n689
  );


  or
  g1042
  (
    n1072,
    n742,
    n709,
    n1038,
    n600
  );


  xnor
  g1043
  (
    n1107,
    n703,
    n701,
    n601,
    n763
  );


  xor
  g1044
  (
    n1083,
    n638,
    n754,
    n682,
    n697
  );


  or
  g1045
  (
    n1057,
    n739,
    n617,
    n723,
    n634
  );


  and
  g1046
  (
    n1087,
    n1040,
    n1049,
    n1039,
    n647
  );


  xor
  g1047
  (
    n1114,
    n741,
    n760,
    n650,
    n702
  );


  xor
  g1048
  (
    n1106,
    n1043,
    n676,
    n693,
    n1037
  );


  xor
  g1049
  (
    n1091,
    n1047,
    n665,
    n764,
    n738
  );


  nand
  g1050
  (
    n1105,
    n1039,
    n756,
    n1051,
    n1042
  );


  nand
  g1051
  (
    n1065,
    n626,
    n704,
    n1047,
    n728
  );


  nor
  g1052
  (
    n1113,
    n1045,
    n674,
    n614,
    n687
  );


  nand
  g1053
  (
    n1060,
    n616,
    n1043,
    n654,
    n602
  );


  and
  g1054
  (
    n1062,
    n620,
    n615,
    n1042,
    n1046
  );


  nor
  g1055
  (
    n1064,
    n763,
    n1039,
    n597,
    n594
  );


  and
  g1056
  (
    n1103,
    n717,
    n1048,
    n731,
    n757
  );


  nand
  g1057
  (
    n1101,
    n596,
    n621,
    n1046,
    n761
  );


  xor
  g1058
  (
    n1111,
    n675,
    n692,
    n649,
    n653
  );


  nor
  g1059
  (
    n1096,
    n1047,
    n691,
    n588,
    n599
  );


  xor
  g1060
  (
    KeyWire_0_7,
    n730,
    n1046,
    n748
  );


  or
  g1061
  (
    n1100,
    n666,
    n1044,
    n656,
    n695
  );


  or
  g1062
  (
    n1070,
    n668,
    n713,
    n1042,
    n762
  );


  or
  g1063
  (
    n1053,
    n604,
    n661,
    n619,
    n726
  );


  and
  g1064
  (
    n1110,
    n759,
    n686,
    n1037,
    n683
  );


  nand
  g1065
  (
    n1112,
    n670,
    n635,
    n1038,
    n690
  );


  nor
  g1066
  (
    n1108,
    n745,
    n681,
    n685,
    n643
  );


  xor
  g1067
  (
    n1055,
    n740,
    n598,
    n637,
    n749
  );


  nand
  g1068
  (
    n1079,
    n664,
    n729,
    n715,
    n1039
  );


  xnor
  g1069
  (
    n1102,
    n744,
    n606,
    n618,
    n1048
  );


  and
  g1070
  (
    n1109,
    n605,
    n759,
    n764,
    n1052
  );


  xor
  g1071
  (
    n1077,
    n623,
    n720,
    n761,
    n688
  );


  and
  g1072
  (
    n1063,
    n642,
    n639,
    n591,
    n610
  );


  xor
  g1073
  (
    n1080,
    n1040,
    n1048,
    n636
  );


  and
  g1074
  (
    n1059,
    n752,
    n1044,
    n629,
    n608
  );


  xor
  g1075
  (
    n1056,
    n1044,
    n700,
    n663,
    n612
  );


  nor
  g1076
  (
    n1074,
    n645,
    n659,
    n1050,
    n622
  );


  and
  g1077
  (
    n1081,
    n669,
    n655,
    n735,
    n746
  );


  and
  g1078
  (
    n1085,
    n589,
    n1043,
    n1050,
    n755
  );


  xnor
  g1079
  (
    n1054,
    n1041,
    n737,
    n671,
    n1051
  );


  xor
  g1080
  (
    n1099,
    n1037,
    n714,
    n732,
    n651
  );


  or
  g1081
  (
    n1104,
    n725,
    n662,
    n646,
    n750
  );


  and
  g1082
  (
    n1082,
    n624,
    n719,
    n679,
    n1050
  );


  xor
  g1083
  (
    n1067,
    n595,
    n751,
    n1051,
    n1049
  );


  xor
  g1084
  (
    n1090,
    n677,
    n698,
    n628,
    n652
  );


  not
  g1085
  (
    n1195,
    n940
  );


  not
  g1086
  (
    n1167,
    n1103
  );


  not
  g1087
  (
    n1158,
    n967
  );


  buf
  g1088
  (
    n1177,
    n932
  );


  not
  g1089
  (
    n1192,
    n967
  );


  not
  g1090
  (
    n1129,
    n1092
  );


  not
  g1091
  (
    n1131,
    n1112
  );


  buf
  g1092
  (
    n1193,
    n1083
  );


  not
  g1093
  (
    n1219,
    n968
  );


  not
  g1094
  (
    KeyWire_0_12,
    n985
  );


  not
  g1095
  (
    n1135,
    n1103
  );


  not
  g1096
  (
    n1202,
    n1096
  );


  nand
  g1097
  (
    n1152,
    n1085,
    n955,
    n964,
    n936
  );


  xor
  g1098
  (
    n1139,
    n1107,
    n954,
    n938,
    n145
  );


  xnor
  g1099
  (
    n1205,
    n145,
    n946,
    n977,
    n1106
  );


  xnor
  g1100
  (
    n1170,
    n999,
    n1109,
    n951
  );


  nand
  g1101
  (
    n1126,
    n947,
    n975,
    n949,
    n942
  );


  and
  g1102
  (
    n1175,
    n956,
    n1097,
    n976,
    n1056
  );


  and
  g1103
  (
    n1220,
    n941,
    n970,
    n984,
    n935
  );


  xnor
  g1104
  (
    n1117,
    n968,
    n962,
    n936,
    n966
  );


  nor
  g1105
  (
    n1200,
    n938,
    n1079,
    n960,
    n1104
  );


  and
  g1106
  (
    n1125,
    n992,
    n1090,
    n1111,
    n1100
  );


  nand
  g1107
  (
    n1197,
    n933,
    n983,
    n987,
    n999
  );


  or
  g1108
  (
    n1119,
    n970,
    n983,
    n988,
    n945
  );


  xor
  g1109
  (
    n1181,
    n950,
    n1106,
    n935,
    n939
  );


  nand
  g1110
  (
    n1130,
    n983,
    n984,
    n1100,
    n980
  );


  xor
  g1111
  (
    n1183,
    n975,
    n970,
    n932,
    n957
  );


  nor
  g1112
  (
    n1147,
    n951,
    n1102,
    n932,
    n1075
  );


  and
  g1113
  (
    n1180,
    n987,
    n953,
    n1089,
    n145
  );


  or
  g1114
  (
    n1186,
    n930,
    n948,
    n979,
    n1107
  );


  or
  g1115
  (
    n1168,
    n990,
    n980,
    n142,
    n1088
  );


  nand
  g1116
  (
    n1194,
    n1110,
    n986,
    n949
  );


  nand
  g1117
  (
    n1128,
    n994,
    n1091,
    n935,
    n1112
  );


  xor
  g1118
  (
    n1190,
    n978,
    n974,
    n933,
    n940
  );


  nand
  g1119
  (
    n1206,
    n956,
    n144,
    n963,
    n978
  );


  xnor
  g1120
  (
    n1123,
    n989,
    n949,
    n950,
    n948
  );


  or
  g1121
  (
    n1155,
    n953,
    n934,
    n1110,
    n1074
  );


  xor
  g1122
  (
    n1133,
    n960,
    n934,
    n1111,
    n931
  );


  xor
  g1123
  (
    n1188,
    n991,
    n1080,
    n1112,
    n941
  );


  xor
  g1124
  (
    n1145,
    n1093,
    n958,
    n961,
    n1061
  );


  or
  g1125
  (
    n1162,
    n972,
    n978,
    n1108,
    n964
  );


  nand
  g1126
  (
    n1146,
    n1000,
    n959,
    n1070,
    n1065
  );


  and
  g1127
  (
    n1127,
    n944,
    n1101,
    n966,
    n931
  );


  xnor
  g1128
  (
    n1151,
    n1100,
    n997,
    n1001,
    n989
  );


  and
  g1129
  (
    n1150,
    n976,
    n977,
    n943,
    n1084
  );


  nor
  g1130
  (
    n1134,
    n1066,
    n933,
    n947,
    n945
  );


  xnor
  g1131
  (
    n1138,
    n939,
    n1100,
    n1110,
    n988
  );


  nand
  g1132
  (
    n1185,
    n993,
    n974,
    n933,
    n1110
  );


  xor
  g1133
  (
    n1215,
    n937,
    n971,
    n1102,
    n948
  );


  and
  g1134
  (
    n1149,
    n938,
    n938,
    n985,
    n994
  );


  nor
  g1135
  (
    n1174,
    n937,
    n1057,
    n982,
    n942
  );


  nand
  g1136
  (
    n1169,
    n955,
    n1099,
    n946,
    n935
  );


  or
  g1137
  (
    n1121,
    n1113,
    n943,
    n954,
    n965
  );


  and
  g1138
  (
    n1212,
    n1104,
    n1106,
    n954,
    n943
  );


  nor
  g1139
  (
    n1120,
    n967,
    n1000,
    n930,
    n1112
  );


  or
  g1140
  (
    n1141,
    n973,
    n1076,
    n958,
    n1077
  );


  nor
  g1141
  (
    n1217,
    n950,
    n143,
    n1105,
    n963
  );


  xnor
  g1142
  (
    n1144,
    n997,
    n1114,
    n972,
    n1107
  );


  and
  g1143
  (
    n1140,
    n1107,
    n963,
    n975,
    n995
  );


  nor
  g1144
  (
    n1184,
    n959,
    n1068,
    n1072,
    n989
  );


  and
  g1145
  (
    n1223,
    n945,
    n971,
    n947,
    n975
  );


  or
  g1146
  (
    n1163,
    n1001,
    n1060,
    n952,
    n999
  );


  xnor
  g1147
  (
    n1225,
    n957,
    n945,
    n962,
    n1053
  );


  nor
  g1148
  (
    n1203,
    n953,
    n987,
    n972,
    n934
  );


  and
  g1149
  (
    n1142,
    n1114,
    n958,
    n992,
    n981
  );


  xor
  g1150
  (
    n1156,
    n950,
    n1108,
    n969,
    n993
  );


  nand
  g1151
  (
    n1178,
    n961,
    n1062,
    n959,
    n1105
  );


  and
  g1152
  (
    n1179,
    n145,
    n981,
    n979,
    n1109
  );


  nor
  g1153
  (
    n1154,
    n979,
    n965,
    n976,
    n984
  );


  xnor
  g1154
  (
    n1160,
    n1086,
    n1099,
    n993,
    n992
  );


  xor
  g1155
  (
    n1209,
    n1000,
    n1104,
    n1099,
    n957
  );


  and
  g1156
  (
    n1166,
    n983,
    n961,
    n1101
  );


  and
  g1157
  (
    n1208,
    n939,
    n998,
    n974,
    n1103
  );


  or
  g1158
  (
    n1124,
    n951,
    n992,
    n143,
    n995
  );


  nor
  g1159
  (
    n1199,
    n984,
    n941,
    n142,
    n990
  );


  xor
  g1160
  (
    n1218,
    n957,
    n991,
    n969,
    n1101
  );


  nand
  g1161
  (
    n1132,
    n1097,
    n144,
    n995,
    n965
  );


  xor
  g1162
  (
    n1171,
    n936,
    n963,
    n949,
    n934
  );


  and
  g1163
  (
    n1161,
    n977,
    n982,
    n974,
    n946
  );


  xnor
  g1164
  (
    n1187,
    n1064,
    n968,
    n1054,
    n961
  );


  xor
  g1165
  (
    n1191,
    n996,
    n998,
    n955,
    n973
  );


  nand
  g1166
  (
    n1157,
    n1001,
    n990,
    n993,
    n944
  );


  xor
  g1167
  (
    n1182,
    n1113,
    n1082,
    n1059,
    n954
  );


  nand
  g1168
  (
    n1115,
    n981,
    n985,
    n998,
    n971
  );


  or
  g1169
  (
    n1196,
    n1071,
    n987,
    n981,
    n996
  );


  nand
  g1170
  (
    n1148,
    n1099,
    n982,
    n947,
    n976
  );


  or
  g1171
  (
    n1118,
    n943,
    n937,
    n996,
    n952
  );


  or
  g1172
  (
    n1201,
    n942,
    n1105,
    n982,
    n986
  );


  and
  g1173
  (
    n1153,
    n144,
    n979,
    n1069,
    n964
  );


  nor
  g1174
  (
    n1213,
    n1113,
    n1094,
    n958,
    n940
  );


  nor
  g1175
  (
    n1137,
    n994,
    n931,
    n937,
    n1081
  );


  xor
  g1176
  (
    n1216,
    n1108,
    n1114,
    n931,
    n1073
  );


  and
  g1177
  (
    n1143,
    n997,
    n956,
    n967,
    n941
  );


  xnor
  g1178
  (
    n1224,
    n1105,
    n971,
    n953,
    n960
  );


  xnor
  g1179
  (
    n1164,
    n965,
    n143,
    n968,
    n1098
  );


  nand
  g1180
  (
    n1226,
    n948,
    n989,
    n944,
    n960
  );


  nand
  g1181
  (
    n1172,
    n1063,
    n1111,
    n991,
    n1113
  );


  and
  g1182
  (
    n1198,
    n973,
    n940,
    n144,
    n978
  );


  and
  g1183
  (
    n1222,
    n990,
    n994,
    n969
  );


  xor
  g1184
  (
    n1122,
    n951,
    n955,
    n946,
    n1078
  );


  xor
  g1185
  (
    n1173,
    n1104,
    n1095,
    n962,
    n988
  );


  nand
  g1186
  (
    n1176,
    n966,
    n1108,
    n972,
    n986
  );


  xnor
  g1187
  (
    n1189,
    n997,
    n995,
    n936,
    n1098
  );


  nor
  g1188
  (
    n1214,
    n991,
    n1000,
    n1102,
    n973
  );


  nor
  g1189
  (
    n1211,
    n956,
    n970,
    n962,
    n1087
  );


  nand
  g1190
  (
    n1136,
    n1114,
    n939,
    n1102,
    n143
  );


  or
  g1191
  (
    n1221,
    n966,
    n1109,
    n988,
    n952
  );


  or
  g1192
  (
    n1204,
    n952,
    n996,
    n999,
    n1103
  );


  nor
  g1193
  (
    n1165,
    n959,
    n985,
    n1055,
    n964
  );


  and
  g1194
  (
    n1159,
    n942,
    n1067,
    n980
  );


  or
  g1195
  (
    n1116,
    n977,
    n1058,
    n932,
    n1001
  );


  xnor
  g1196
  (
    n1207,
    n1111,
    n998,
    n944,
    n1106
  );


  not
  g1197
  (
    n1246,
    n1119
  );


  buf
  g1198
  (
    n1235,
    n1116
  );


  buf
  g1199
  (
    n1253,
    n1121
  );


  buf
  g1200
  (
    n1240,
    n1122
  );


  not
  g1201
  (
    n1236,
    n1116
  );


  not
  g1202
  (
    n1251,
    n1116
  );


  buf
  g1203
  (
    n1257,
    n1117
  );


  buf
  g1204
  (
    n1231,
    n1119
  );


  buf
  g1205
  (
    n1245,
    n1116
  );


  buf
  g1206
  (
    n1254,
    n1120
  );


  buf
  g1207
  (
    n1248,
    n1122
  );


  buf
  g1208
  (
    n1230,
    n1119
  );


  not
  g1209
  (
    n1229,
    n1118
  );


  not
  g1210
  (
    n1237,
    n1115
  );


  buf
  g1211
  (
    KeyWire_0_15,
    n1115
  );


  buf
  g1212
  (
    n1239,
    n1118
  );


  not
  g1213
  (
    n1250,
    n1121
  );


  not
  g1214
  (
    n1234,
    n1120
  );


  buf
  g1215
  (
    n1252,
    n1115
  );


  not
  g1216
  (
    n1232,
    n1118
  );


  not
  g1217
  (
    n1249,
    n1119
  );


  not
  g1218
  (
    n1227,
    n1121
  );


  buf
  g1219
  (
    n1243,
    n1122
  );


  buf
  g1220
  (
    n1233,
    n1121
  );


  buf
  g1221
  (
    n1238,
    n1115
  );


  buf
  g1222
  (
    n1228,
    n1120
  );


  not
  g1223
  (
    n1258,
    n1117
  );


  buf
  g1224
  (
    n1255,
    n1117
  );


  not
  g1225
  (
    n1244,
    n1120
  );


  buf
  g1226
  (
    n1242,
    n1117
  );


  not
  g1227
  (
    n1256,
    n1122
  );


  buf
  g1228
  (
    n1241,
    n1118
  );


  xor
  g1229
  (
    n1383,
    n864,
    n861,
    n783,
    n1235
  );


  nand
  g1230
  (
    n1342,
    n1227,
    n1258,
    n849,
    n797
  );


  and
  g1231
  (
    n1356,
    n859,
    n850,
    n1237,
    n823
  );


  xor
  g1232
  (
    n1327,
    n781,
    n1250,
    n837,
    n802
  );


  nand
  g1233
  (
    n1359,
    n851,
    n803,
    n1227,
    n1248
  );


  and
  g1234
  (
    n1345,
    n1245,
    n775,
    n842,
    n806
  );


  nand
  g1235
  (
    n1380,
    n779,
    n841,
    n817,
    n865
  );


  nand
  g1236
  (
    n1381,
    n1230,
    n780,
    n790,
    n1244
  );


  nor
  g1237
  (
    n1349,
    n811,
    n1234,
    n800,
    n776
  );


  or
  g1238
  (
    n1325,
    n766,
    n802,
    n840,
    n796
  );


  xnor
  g1239
  (
    n1353,
    n1256,
    n1227,
    n847,
    n835
  );


  xor
  g1240
  (
    n1310,
    n1256,
    n1257,
    n829,
    n786
  );


  or
  g1241
  (
    n1301,
    n805,
    n811,
    n833,
    n789
  );


  xnor
  g1242
  (
    n1360,
    n799,
    n803,
    n1242,
    n782
  );


  nor
  g1243
  (
    n1376,
    n804,
    n1243,
    n1240,
    n823
  );


  xnor
  g1244
  (
    n1296,
    n783,
    n1239,
    n781,
    n1255
  );


  or
  g1245
  (
    n1317,
    n845,
    n1251,
    n846,
    n1228
  );


  nand
  g1246
  (
    n1280,
    n770,
    n1245,
    n838,
    n811
  );


  xnor
  g1247
  (
    n1322,
    n774,
    n1249,
    n1256,
    n781
  );


  nor
  g1248
  (
    n1299,
    n842,
    n829,
    n857,
    n788
  );


  xor
  g1249
  (
    n1330,
    n824,
    n1241,
    n789,
    n863
  );


  nand
  g1250
  (
    n1328,
    n818,
    n1247,
    n768,
    n819
  );


  xnor
  g1251
  (
    n1265,
    n862,
    n804,
    n822,
    n797
  );


  nand
  g1252
  (
    n1331,
    n864,
    n847,
    n778,
    n818
  );


  nor
  g1253
  (
    n1282,
    n1245,
    n850,
    n1248,
    n774
  );


  nand
  g1254
  (
    n1373,
    n820,
    n1243,
    n832,
    n801
  );


  nor
  g1255
  (
    n1273,
    n799,
    n848,
    n1235,
    n861
  );


  xnor
  g1256
  (
    n1275,
    n799,
    n810,
    n785,
    n805
  );


  or
  g1257
  (
    n1308,
    n842,
    n849,
    n844,
    n855
  );


  or
  g1258
  (
    n1361,
    n811,
    n830,
    n855,
    n1232
  );


  nand
  g1259
  (
    n1290,
    n798,
    n778,
    n1229,
    n1253
  );


  or
  g1260
  (
    n1269,
    n846,
    n795,
    n842,
    n803
  );


  or
  g1261
  (
    n1287,
    n817,
    n861,
    n795,
    n1243
  );


  xor
  g1262
  (
    n1371,
    n1245,
    n1239,
    n826,
    n1256
  );


  nor
  g1263
  (
    n1319,
    n790,
    n814,
    n819,
    n860
  );


  nor
  g1264
  (
    n1365,
    n839,
    n1239,
    n1246,
    n1227
  );


  xnor
  g1265
  (
    n1315,
    n857,
    n853,
    n802,
    n837
  );


  or
  g1266
  (
    n1369,
    n826,
    n836,
    n801,
    n1253
  );


  xnor
  g1267
  (
    n1261,
    n824,
    n1255,
    n821,
    n786
  );


  nor
  g1268
  (
    n1320,
    n1246,
    n810,
    n827
  );


  or
  g1269
  (
    n1292,
    n816,
    n814,
    n828,
    n833
  );


  xor
  g1270
  (
    n1362,
    n1237,
    n779,
    n854,
    n783
  );


  and
  g1271
  (
    n1277,
    n836,
    n863,
    n1257,
    n851
  );


  or
  g1272
  (
    n1333,
    n820,
    n844,
    n798,
    n848
  );


  or
  g1273
  (
    n1309,
    n849,
    n865,
    n800,
    n807
  );


  xor
  g1274
  (
    n1337,
    n1251,
    n812,
    n857,
    n1236
  );


  nor
  g1275
  (
    n1270,
    n807,
    n1244,
    n1231,
    n1252
  );


  or
  g1276
  (
    n1289,
    n860,
    n835,
    n797,
    n840
  );


  nand
  g1277
  (
    n1374,
    n843,
    n776,
    n1229,
    n1231
  );


  and
  g1278
  (
    n1283,
    n832,
    n782,
    n837
  );


  nor
  g1279
  (
    n1363,
    n828,
    n793,
    n1258,
    n1241
  );


  and
  g1280
  (
    n1268,
    n775,
    n1248,
    n820,
    n792
  );


  xor
  g1281
  (
    n1368,
    n1247,
    n863,
    n809,
    n860
  );


  and
  g1282
  (
    n1302,
    n1238,
    n776,
    n834,
    n792
  );


  xnor
  g1283
  (
    n1298,
    n1237,
    n816,
    n803,
    n1250
  );


  nor
  g1284
  (
    n1281,
    n859,
    n841,
    n853,
    n770
  );


  or
  g1285
  (
    n1306,
    n796,
    n843,
    n794,
    n795
  );


  and
  g1286
  (
    n1355,
    n863,
    n833,
    n1251,
    n1257
  );


  xnor
  g1287
  (
    n1357,
    n822,
    n794,
    n820,
    n824
  );


  and
  g1288
  (
    n1329,
    n1252,
    n812,
    n840,
    n787
  );


  xnor
  g1289
  (
    n1284,
    n830,
    n856,
    n808,
    n777
  );


  nor
  g1290
  (
    n1263,
    n1243,
    n1233,
    n840,
    n780
  );


  or
  g1291
  (
    n1339,
    n1244,
    n1240,
    n848,
    n791
  );


  nor
  g1292
  (
    n1285,
    n771,
    n853,
    n864,
    n846
  );


  nand
  g1293
  (
    n1384,
    n784,
    n832,
    n1250,
    n800
  );


  nor
  g1294
  (
    n1267,
    n847,
    n819,
    n785,
    n834
  );


  xnor
  g1295
  (
    n1336,
    n829,
    n787,
    n844,
    n1238
  );


  xnor
  g1296
  (
    n1286,
    n828,
    n1246,
    n839,
    n1231
  );


  or
  g1297
  (
    n1266,
    n851,
    n796,
    n806,
    n823
  );


  and
  g1298
  (
    n1378,
    n836,
    n1253,
    n769,
    n779
  );


  nor
  g1299
  (
    n1338,
    n794,
    n809,
    n784,
    n834
  );


  nand
  g1300
  (
    n1291,
    n1254,
    n772,
    n1257,
    n1229
  );


  xnor
  g1301
  (
    n1259,
    n1241,
    n862,
    n806,
    n1251
  );


  and
  g1302
  (
    n1326,
    n1258,
    n847,
    n1232,
    n793
  );


  and
  g1303
  (
    n1335,
    n831,
    n857,
    n769,
    n866
  );


  nand
  g1304
  (
    n1385,
    n1242,
    n817,
    n1247,
    n1236
  );


  and
  g1305
  (
    n1344,
    n805,
    n865,
    n848,
    n822
  );


  nand
  g1306
  (
    n1311,
    n792,
    n854,
    n1248,
    n1249
  );


  or
  g1307
  (
    n1348,
    n818,
    n824,
    n853,
    n777
  );


  and
  g1308
  (
    n1278,
    n856,
    n816,
    n851,
    n800
  );


  xnor
  g1309
  (
    n1346,
    n862,
    n1242,
    n1247,
    n815
  );


  nand
  g1310
  (
    n1332,
    n828,
    n767,
    n787,
    n837
  );


  or
  g1311
  (
    n1323,
    n858,
    n780,
    n854,
    n1235
  );


  xor
  g1312
  (
    n1386,
    n781,
    n813,
    n852,
    n816
  );


  or
  g1313
  (
    n1288,
    n786,
    n821,
    n1258,
    n1237
  );


  xor
  g1314
  (
    n1297,
    n834,
    n831,
    n1238,
    n852
  );


  and
  g1315
  (
    n1343,
    n817,
    n1235,
    n778,
    n807
  );


  nor
  g1316
  (
    n1295,
    n1233,
    n779,
    n1249,
    n813
  );


  nor
  g1317
  (
    n1382,
    n846,
    n772,
    n798,
    n804
  );


  xor
  g1318
  (
    n1377,
    n1230,
    n774,
    n843,
    n1252
  );


  nor
  g1319
  (
    n1276,
    n810,
    n864,
    n792,
    n768
  );


  xnor
  g1320
  (
    n1262,
    n1236,
    n862,
    n1229,
    n861
  );


  or
  g1321
  (
    n1370,
    n795,
    n1246,
    n773,
    n813
  );


  or
  g1322
  (
    n1293,
    n776,
    n827,
    n821,
    n859
  );


  xnor
  g1323
  (
    n1264,
    n771,
    n774,
    n812,
    n1241
  );


  nor
  g1324
  (
    n1312,
    n812,
    n845,
    n805,
    n788
  );


  nand
  g1325
  (
    n1300,
    n841,
    n808,
    n793,
    n827
  );


  nor
  g1326
  (
    n1366,
    n858,
    n858,
    n850,
    n1255
  );


  nand
  g1327
  (
    n1321,
    n815,
    n1234,
    n1228,
    n823
  );


  and
  g1328
  (
    n1272,
    n808,
    n849,
    n1252,
    n844
  );


  or
  g1329
  (
    n1304,
    n791,
    n1254,
    n850,
    n797
  );


  and
  g1330
  (
    n1350,
    n1238,
    n1240,
    n777,
    n855
  );


  or
  g1331
  (
    n1314,
    n860,
    n1253,
    n787,
    n777
  );


  xnor
  g1332
  (
    n1279,
    n839,
    n804,
    n801,
    n835
  );


  or
  g1333
  (
    n1318,
    n790,
    n845,
    n865,
    n858
  );


  nand
  g1334
  (
    n1334,
    n852,
    n821,
    n833,
    n836
  );


  nand
  g1335
  (
    n1367,
    n1230,
    n784,
    n831,
    n796
  );


  nor
  g1336
  (
    n1358,
    n775,
    n838,
    n1240,
    n783
  );


  nand
  g1337
  (
    n1352,
    n832,
    n1242,
    n789,
    n1254
  );


  xnor
  g1338
  (
    n1379,
    n775,
    n809,
    n808,
    n818
  );


  nand
  g1339
  (
    n1372,
    n793,
    n815,
    n838,
    n782
  );


  nor
  g1340
  (
    n1307,
    n780,
    n1233,
    n841,
    n1232
  );


  nor
  g1341
  (
    n1347,
    n843,
    n814,
    n852,
    n1234
  );


  or
  g1342
  (
    n1375,
    n1249,
    n802,
    n1234,
    n1254
  );


  xor
  g1343
  (
    n1305,
    n825,
    n829,
    n819,
    n1232
  );


  nor
  g1344
  (
    n1271,
    n830,
    n807,
    n1228,
    n825
  );


  xnor
  g1345
  (
    n1313,
    n856,
    n838,
    n815,
    n790
  );


  xor
  g1346
  (
    n1324,
    n813,
    n799,
    n785,
    n773
  );


  and
  g1347
  (
    n1260,
    n809,
    n845,
    n767,
    n826
  );


  or
  g1348
  (
    n1351,
    n778,
    n801,
    n791,
    n822
  );


  xor
  g1349
  (
    n1274,
    n839,
    n814,
    n831,
    n825
  );


  nor
  g1350
  (
    n1316,
    n786,
    n856,
    n827,
    n784
  );


  or
  g1351
  (
    n1294,
    n791,
    n1255,
    n794,
    n1236
  );


  xnor
  g1352
  (
    n1341,
    n1231,
    n1239,
    n835,
    n1244
  );


  nor
  g1353
  (
    n1364,
    n789,
    n788,
    n830,
    n826
  );


  xor
  g1354
  (
    n1340,
    n798,
    n1250,
    n806,
    n825
  );


  xnor
  g1355
  (
    n1354,
    n859,
    n785,
    n855,
    n854
  );


  xor
  g1356
  (
    n1303,
    n1228,
    n1233,
    n1230,
    n788
  );


  not
  g1357
  (
    n1388,
    n1260
  );


  buf
  g1358
  (
    n1389,
    n1270
  );


  not
  g1359
  (
    n1393,
    n1002
  );


  not
  g1360
  (
    n1390,
    n1272
  );


  not
  g1361
  (
    KeyWire_0_2,
    n1264
  );


  buf
  g1362
  (
    n1395,
    n1271
  );


  nor
  g1363
  (
    n1387,
    n1259,
    n1266,
    n1261,
    n1269
  );


  xnor
  g1364
  (
    n1394,
    n1267,
    n1268,
    n1002,
    n1263
  );


  or
  g1365
  (
    n1391,
    n1262,
    n1002,
    n1265
  );


  buf
  g1366
  (
    n1396,
    n1387
  );


  and
  g1367
  (
    n1399,
    n1125,
    n1123,
    n1124
  );


  xnor
  g1368
  (
    n1397,
    n1123,
    n1396,
    n1124
  );


  nand
  g1369
  (
    n1398,
    n1124,
    n1396,
    n1123
  );


  or
  g1370
  (
    n1408,
    n1126,
    n1127,
    n442,
    n1125
  );


  nor
  g1371
  (
    n1411,
    n1399,
    n446,
    n1398,
    n1125
  );


  or
  g1372
  (
    n1409,
    n443,
    n1128,
    n1127,
    n1126
  );


  xor
  g1373
  (
    n1407,
    n445,
    n443,
    n442,
    n1126
  );


  or
  g1374
  (
    n1402,
    n445,
    n441,
    n1128,
    n1052
  );


  nand
  g1375
  (
    n1410,
    n1125,
    n445,
    n1399,
    n1052
  );


  nand
  g1376
  (
    n1405,
    n443,
    n441,
    n444,
    n1398
  );


  nand
  g1377
  (
    n1403,
    n1126,
    n1128,
    n445,
    n444
  );


  nand
  g1378
  (
    n1401,
    n1398,
    n443,
    n1397
  );


  or
  g1379
  (
    n1400,
    n1397,
    n444,
    n442,
    n1127
  );


  xor
  g1380
  (
    n1404,
    n1398,
    n1127,
    n444,
    n442
  );


  nor
  g1381
  (
    n1406,
    n1397,
    n1399,
    n1128
  );


  or
  g1382
  (
    n1428,
    n1404,
    n1304
  );


  xnor
  g1383
  (
    n1413,
    n1403,
    n1285
  );


  xor
  g1384
  (
    n1412,
    n1282,
    n1402
  );


  nand
  g1385
  (
    n1425,
    n1274,
    n1402
  );


  xnor
  g1386
  (
    n1431,
    n1302,
    n1283
  );


  nor
  g1387
  (
    n1415,
    n1288,
    n1303
  );


  xnor
  g1388
  (
    n1427,
    n1284,
    n1400
  );


  xnor
  g1389
  (
    n1426,
    n1400,
    n1299
  );


  and
  g1390
  (
    n1424,
    n1403,
    n1402
  );


  nor
  g1391
  (
    n1418,
    n1273,
    n1297
  );


  nor
  g1392
  (
    n1422,
    n1298,
    n1403
  );


  xor
  g1393
  (
    n1421,
    n1405,
    n1291
  );


  or
  g1394
  (
    n1432,
    n1289,
    n1278
  );


  xor
  g1395
  (
    n1430,
    n1401,
    n1277,
    n1402,
    n1405
  );


  xnor
  g1396
  (
    n1429,
    n1294,
    n1307,
    n1401,
    n1276
  );


  nand
  g1397
  (
    n1419,
    n1300,
    n1404,
    n1295
  );


  nand
  g1398
  (
    n1417,
    n1129,
    n1400,
    n1405,
    n1306
  );


  xor
  g1399
  (
    n1414,
    n1290,
    n1404,
    n1296,
    n1281
  );


  or
  g1400
  (
    n1423,
    n1401,
    n1293,
    n1279,
    n1129
  );


  nand
  g1401
  (
    n1416,
    n1275,
    n1280,
    n1286,
    n1292
  );


  and
  g1402
  (
    n1420,
    n1287,
    n1301,
    n1403,
    n1305
  );


  buf
  g1403
  (
    n1433,
    n1412
  );


  not
  g1404
  (
    n1436,
    n1433
  );


  buf
  g1405
  (
    n1437,
    n1433
  );


  buf
  g1406
  (
    n1435,
    n1433
  );


  buf
  g1407
  (
    n1434,
    n1433
  );


  buf
  g1408
  (
    n1446,
    n1315
  );


  not
  g1409
  (
    n1452,
    n1437
  );


  not
  g1410
  (
    n1447,
    n1435
  );


  buf
  g1411
  (
    n1443,
    n1434
  );


  not
  g1412
  (
    n1439,
    n1434
  );


  not
  g1413
  (
    n1448,
    n1434
  );


  buf
  g1414
  (
    n1441,
    n1310
  );


  buf
  g1415
  (
    n1449,
    n1313
  );


  not
  g1416
  (
    n1453,
    n1436
  );


  buf
  g1417
  (
    KeyWire_0_13,
    n1437
  );


  buf
  g1418
  (
    n1438,
    n1435
  );


  buf
  g1419
  (
    n1444,
    n1436
  );


  not
  g1420
  (
    n1445,
    n1312
  );


  and
  g1421
  (
    n1450,
    n1436,
    n1435,
    n1309,
    n1437
  );


  nand
  g1422
  (
    n1451,
    n1314,
    n1308,
    n1437,
    n1311
  );


  nor
  g1423
  (
    n1440,
    n1316,
    n1434,
    n1435,
    n1436
  );


  xor
  g1424
  (
    n1492,
    n463,
    n1442,
    n476,
    n1449
  );


  or
  g1425
  (
    n1480,
    n462,
    n1440,
    n484,
    n1134
  );


  or
  g1426
  (
    n1472,
    n467,
    n1130,
    n461,
    n480
  );


  nor
  g1427
  (
    n1508,
    n448,
    n1389,
    n465,
    n468
  );


  xnor
  g1428
  (
    n1499,
    n456,
    n474,
    n1451,
    n1444
  );


  or
  g1429
  (
    n1515,
    n458,
    n1133,
    n1453,
    n1440
  );


  and
  g1430
  (
    n1454,
    n1441,
    n455,
    n482,
    n478
  );


  xnor
  g1431
  (
    n1488,
    n1388,
    n1394,
    n459,
    n447
  );


  or
  g1432
  (
    n1501,
    n468,
    n453,
    n467,
    n1447
  );


  or
  g1433
  (
    n1455,
    n482,
    n474,
    n457,
    n1442
  );


  and
  g1434
  (
    n1514,
    n1448,
    n1448,
    n470,
    n471
  );


  or
  g1435
  (
    n1513,
    n1390,
    n1453,
    n1406,
    n1135
  );


  xor
  g1436
  (
    n1466,
    n1129,
    n462,
    n1450,
    n480
  );


  nor
  g1437
  (
    n1487,
    n447,
    n1406,
    n468,
    n449
  );


  nand
  g1438
  (
    n1475,
    n469,
    n1449,
    n481,
    n473
  );


  and
  g1439
  (
    n1507,
    n450,
    n468,
    n1441,
    n466
  );


  xnor
  g1440
  (
    n1503,
    n477,
    n475,
    n1447,
    n446
  );


  or
  g1441
  (
    n1457,
    n446,
    n1438,
    n463,
    n1441
  );


  nand
  g1442
  (
    n1459,
    n448,
    n465,
    n1446,
    n477
  );


  nor
  g1443
  (
    n1473,
    n453,
    n1132,
    n479
  );


  nor
  g1444
  (
    n1512,
    n1445,
    n1132,
    n452,
    n1438
  );


  nand
  g1445
  (
    n1500,
    n484,
    n448,
    n1440,
    n1449
  );


  and
  g1446
  (
    n1462,
    n452,
    n1132,
    n1439,
    n1133
  );


  nand
  g1447
  (
    n1511,
    n475,
    n476,
    n1442,
    n480
  );


  nand
  g1448
  (
    n1495,
    n456,
    n1446,
    n478
  );


  nand
  g1449
  (
    n1509,
    n1444,
    n475,
    n1443,
    n485
  );


  nand
  g1450
  (
    n1496,
    n1133,
    n1443,
    n451,
    n1392
  );


  and
  g1451
  (
    n1463,
    n454,
    n451,
    n1450
  );


  and
  g1452
  (
    n1458,
    n1450,
    n466,
    n1448
  );


  and
  g1453
  (
    n1504,
    n1448,
    n471,
    n460,
    n1452
  );


  xor
  g1454
  (
    n1517,
    n485,
    n464,
    n483,
    n473
  );


  xor
  g1455
  (
    n1498,
    n456,
    n1451,
    n455,
    n477
  );


  xnor
  g1456
  (
    n1468,
    n448,
    n452,
    n479,
    n1438
  );


  or
  g1457
  (
    n1479,
    n469,
    n1446,
    n1444,
    n484
  );


  xor
  g1458
  (
    n1491,
    n472,
    n446,
    n481,
    n1130
  );


  nor
  g1459
  (
    n1489,
    n465,
    n1445,
    n458,
    n454
  );


  xnor
  g1460
  (
    n1483,
    n481,
    n472,
    n483,
    n1452
  );


  or
  g1461
  (
    n1502,
    n450,
    n1449,
    n1442,
    n479
  );


  or
  g1462
  (
    n1474,
    n1450,
    n451,
    n482,
    n1134
  );


  nor
  g1463
  (
    n1490,
    n464,
    n449,
    n456,
    n470
  );


  nor
  g1464
  (
    n1510,
    n475,
    n1443,
    n1134
  );


  or
  g1465
  (
    n1486,
    n1406,
    n460,
    n454,
    n449
  );


  or
  g1466
  (
    n1460,
    n1131,
    n471,
    n469,
    n470
  );


  xor
  g1467
  (
    n1478,
    n1447,
    n1131,
    n459,
    n1453
  );


  or
  g1468
  (
    n1506,
    n458,
    n474,
    n478,
    n453
  );


  xor
  g1469
  (
    n1464,
    n450,
    n480,
    n1444,
    n463
  );


  or
  g1470
  (
    KeyWire_0_14,
    n470,
    n1453,
    n1441,
    n1133
  );


  xor
  g1471
  (
    n1493,
    n455,
    n472,
    n464,
    n1130
  );


  xnor
  g1472
  (
    n1471,
    n1447,
    n479,
    n461,
    n476
  );


  nor
  g1473
  (
    n1456,
    n484,
    n1130,
    n1439,
    n447
  );


  nor
  g1474
  (
    n1470,
    n482,
    n461,
    n1452,
    n472
  );


  xor
  g1475
  (
    n1505,
    n476,
    n465,
    n447,
    n471
  );


  or
  g1476
  (
    n1497,
    n473,
    n450,
    n454,
    n1129
  );


  or
  g1477
  (
    n1484,
    n459,
    n452,
    n1451,
    n474
  );


  xor
  g1478
  (
    n1467,
    n478,
    n483,
    n467,
    n453
  );


  nor
  g1479
  (
    n1485,
    n1391,
    n1451,
    n463,
    n1445
  );


  xnor
  g1480
  (
    n1461,
    n1393,
    n483,
    n449,
    n467
  );


  nand
  g1481
  (
    n1482,
    n1131,
    n1439,
    n464,
    n455
  );


  nor
  g1482
  (
    n1469,
    n1452,
    n469,
    n461,
    n457
  );


  xnor
  g1483
  (
    n1494,
    n457,
    n460,
    n1134,
    n1405
  );


  or
  g1484
  (
    n1481,
    n1440,
    n460,
    n473,
    n1131
  );


  nor
  g1485
  (
    n1516,
    n481,
    n1438,
    n462,
    n459
  );


  or
  g1486
  (
    n1465,
    n457,
    n1406,
    n1445,
    n1439
  );


  nand
  g1487
  (
    n1476,
    n458,
    n477,
    n466,
    n462
  );


  nand
  g1488
  (
    n1523,
    n880,
    n880,
    n867,
    n869
  );


  xnor
  g1489
  (
    n1527,
    n867,
    n871,
    n1455,
    n868
  );


  xnor
  g1490
  (
    n1533,
    n879,
    n866,
    n880,
    n867
  );


  or
  g1491
  (
    n1532,
    n869,
    n1469,
    n878,
    n879
  );


  nand
  g1492
  (
    n1531,
    n877,
    n870,
    n876,
    n1473
  );


  nand
  g1493
  (
    n1521,
    n880,
    n1460,
    n873,
    n1465
  );


  xnor
  g1494
  (
    n1520,
    n1459,
    n872,
    n866,
    n1464
  );


  xnor
  g1495
  (
    n1522,
    n873,
    n875,
    n872
  );


  nand
  g1496
  (
    n1536,
    n1471,
    n874,
    n870
  );


  nor
  g1497
  (
    n1518,
    n869,
    n878,
    n876,
    n875
  );


  xor
  g1498
  (
    n1519,
    n876,
    n1458,
    n866,
    n1466
  );


  nand
  g1499
  (
    n1535,
    n1470,
    n877,
    n1462,
    n870
  );


  nand
  g1500
  (
    n1534,
    n868,
    n870,
    n1463,
    n879
  );


  xor
  g1501
  (
    n1525,
    n872,
    n878,
    n1468,
    n1454
  );


  xor
  g1502
  (
    n1526,
    n872,
    n871,
    n875,
    n1472
  );


  xnor
  g1503
  (
    n1530,
    n873,
    n873,
    n1461,
    n1456
  );


  and
  g1504
  (
    n1537,
    n874,
    n485,
    n868,
    n871
  );


  nor
  g1505
  (
    n1529,
    n878,
    n869,
    n871,
    n1467
  );


  nand
  g1506
  (
    n1524,
    n1457,
    n868,
    n876,
    n877
  );


  xnor
  g1507
  (
    n1528,
    n879,
    n867,
    n877,
    n874
  );


  buf
  g1508
  (
    n1539,
    n1518
  );


  buf
  g1509
  (
    n1538,
    n1519
  );


  buf
  g1510
  (
    n1540,
    n1520
  );


  xor
  g1511
  (
    n1550,
    n1408,
    n1539,
    n1540
  );


  nand
  g1512
  (
    n1552,
    n1409,
    n1137,
    n1136
  );


  nand
  g1513
  (
    n1551,
    n1139,
    n1409,
    n1411
  );


  and
  g1514
  (
    n1543,
    n1410,
    n1138,
    n1411
  );


  nor
  g1515
  (
    n1548,
    n1136,
    n1540,
    n1135,
    n1538
  );


  nor
  g1516
  (
    n1541,
    n1410,
    n1135,
    n1538,
    n1408
  );


  xnor
  g1517
  (
    n1549,
    n1409,
    n1138,
    n1407
  );


  or
  g1518
  (
    n1545,
    n1407,
    n1137,
    n1538,
    n1410
  );


  or
  g1519
  (
    n1546,
    n1407,
    n1411,
    n1540
  );


  nor
  g1520
  (
    n1542,
    n1538,
    n1136,
    n1539
  );


  nor
  g1521
  (
    n1547,
    n1135,
    n1408,
    n1407,
    n1136
  );


  nand
  g1522
  (
    n1544,
    n1408,
    n1410,
    n1137,
    n1539
  );


  or
  g1523
  (
    n1557,
    n1330,
    n1351,
    n1418,
    n1545
  );


  or
  g1524
  (
    n1576,
    n1321,
    n1331,
    n1424,
    n1543
  );


  nand
  g1525
  (
    n1571,
    n1547,
    n1426,
    n1546,
    n1332
  );


  or
  g1526
  (
    n1564,
    n1550,
    n1421,
    n1428,
    n1319
  );


  nor
  g1527
  (
    n1560,
    n1552,
    n1422,
    n1551,
    n1423
  );


  and
  g1528
  (
    n1586,
    n1417,
    n1548,
    n1339,
    n1355
  );


  nor
  g1529
  (
    n1566,
    n1355,
    n1343,
    n1333,
    n1350
  );


  xor
  g1530
  (
    n1555,
    n1354,
    n1430,
    n1324
  );


  xnor
  g1531
  (
    n1583,
    n1357,
    n1423,
    n1338,
    n1542
  );


  and
  g1532
  (
    n1565,
    n1429,
    n1423,
    n1426,
    n1355
  );


  or
  g1533
  (
    n1573,
    n1323,
    n1348,
    n1431,
    n1428
  );


  and
  g1534
  (
    n1569,
    n1552,
    n1550,
    n1422,
    n1342
  );


  and
  g1535
  (
    n1554,
    n1547,
    n1549,
    n1548,
    n1432
  );


  and
  g1536
  (
    n1582,
    n1426,
    n1419,
    n1322,
    n1320
  );


  xnor
  g1537
  (
    n1585,
    n1354,
    n1424,
    n1344,
    n1317
  );


  or
  g1538
  (
    n1575,
    n1334,
    n1329,
    n1414,
    n1423
  );


  xor
  g1539
  (
    n1577,
    n1549,
    n1544,
    n1354,
    n1429
  );


  xor
  g1540
  (
    n1587,
    n1352,
    n1549,
    n1551,
    n1430
  );


  xnor
  g1541
  (
    n1579,
    n1426,
    n1552,
    n1413,
    n1356
  );


  nand
  g1542
  (
    n1581,
    n1428,
    n1427,
    n1541,
    n1346
  );


  and
  g1543
  (
    n1556,
    n1354,
    n1335,
    n1327,
    n1547
  );


  xor
  g1544
  (
    n1553,
    n1550,
    n1337,
    n1353,
    n1357
  );


  or
  g1545
  (
    n1572,
    n1318,
    n1431,
    n1356,
    n1548
  );


  xor
  g1546
  (
    n1562,
    n1340,
    n1541,
    n1430,
    n1427
  );


  nor
  g1547
  (
    n1561,
    n1427,
    n1345,
    n1356,
    n1420
  );


  xnor
  g1548
  (
    n1563,
    n1355,
    n1542,
    n1429,
    n1543
  );


  xor
  g1549
  (
    n1570,
    n1428,
    n1356,
    n1416,
    n1552
  );


  or
  g1550
  (
    n1584,
    n1548,
    n1549,
    n1328,
    n1422
  );


  xor
  g1551
  (
    n1578,
    n1429,
    n1431,
    n1544,
    n1425
  );


  nor
  g1552
  (
    n1574,
    n1336,
    n1550,
    n1432
  );


  and
  g1553
  (
    n1568,
    n1422,
    n1139,
    n1427,
    n1325
  );


  nor
  g1554
  (
    n1567,
    n1432,
    n1425,
    n1424,
    n1551
  );


  or
  g1555
  (
    n1558,
    n1431,
    n1349,
    n1546,
    n1545
  );


  or
  g1556
  (
    n1580,
    n1551,
    n1326,
    n1425,
    n1424
  );


  and
  g1557
  (
    n1559,
    n1341,
    n1415,
    n1425,
    n1347
  );


  buf
  g1558
  (
    n1592,
    n1557
  );


  buf
  g1559
  (
    n1591,
    n1562
  );


  buf
  g1560
  (
    n1588,
    n1565
  );


  not
  g1561
  (
    n1597,
    n1560
  );


  buf
  g1562
  (
    n1593,
    n1566
  );


  not
  g1563
  (
    n1590,
    n1559
  );


  and
  g1564
  (
    n1595,
    n1554,
    n1558
  );


  xor
  g1565
  (
    n1589,
    n1564,
    n1563
  );


  and
  g1566
  (
    n1594,
    n1553,
    n1555
  );


  or
  g1567
  (
    n1596,
    n1561,
    n1556
  );


  nor
  g1568
  (
    n1615,
    n896,
    n883,
    n1522,
    n892
  );


  and
  g1569
  (
    n1600,
    n894,
    n1594,
    n1139,
    n1595
  );


  xnor
  g1570
  (
    n1598,
    n884,
    n887,
    n891,
    n1589
  );


  xor
  g1571
  (
    n1606,
    n1524,
    n894,
    n890,
    n882
  );


  nand
  g1572
  (
    n1605,
    n888,
    n1590,
    n1591,
    n1594
  );


  and
  g1573
  (
    n1617,
    n881,
    n896,
    n890,
    n885
  );


  nor
  g1574
  (
    n1610,
    n894,
    n1592,
    n896,
    n887
  );


  or
  g1575
  (
    n1619,
    n1141,
    n884,
    n1594,
    n881
  );


  nand
  g1576
  (
    n1599,
    n893,
    n892,
    n898,
    n899
  );


  xor
  g1577
  (
    n1609,
    n1521,
    n898,
    n888
  );


  nor
  g1578
  (
    n1624,
    n884,
    n1592,
    n1591,
    n889
  );


  xnor
  g1579
  (
    n1608,
    n889,
    n1593,
    n893,
    n890
  );


  and
  g1580
  (
    n1601,
    n1140,
    n1588,
    n1592,
    n1595
  );


  xor
  g1581
  (
    n1611,
    n882,
    n885,
    n1140,
    n890
  );


  or
  g1582
  (
    n1625,
    n881,
    n895,
    n885
  );


  or
  g1583
  (
    n1612,
    n883,
    n897,
    n895,
    n881
  );


  or
  g1584
  (
    n1607,
    n885,
    n886,
    n883,
    n1594
  );


  xor
  g1585
  (
    n1620,
    n897,
    n898,
    n892,
    n1593
  );


  xnor
  g1586
  (
    n1603,
    n888,
    n891,
    n889,
    n1589
  );


  nor
  g1587
  (
    n1614,
    n1595,
    n1590,
    n895,
    n897
  );


  xnor
  g1588
  (
    n1602,
    n891,
    n1590,
    n1592,
    n893
  );


  and
  g1589
  (
    n1604,
    n887,
    n886,
    n896
  );


  and
  g1590
  (
    n1613,
    n888,
    n1590,
    n894,
    n1140
  );


  xnor
  g1591
  (
    n1618,
    n897,
    n891,
    n882,
    n889
  );


  or
  g1592
  (
    n1616,
    n1593,
    n1589,
    n882,
    n1140
  );


  and
  g1593
  (
    n1621,
    n883,
    n1589,
    n893,
    n884
  );


  xor
  g1594
  (
    n1623,
    n887,
    n886,
    n1139,
    n1523
  );


  and
  g1595
  (
    n1622,
    n1593,
    n1591,
    n892
  );


  buf
  g1596
  (
    n1626,
    n1599
  );


  buf
  g1597
  (
    n1627,
    n1598
  );


  xnor
  g1598
  (
    n1628,
    n1627,
    n1491,
    n1626
  );


  nand
  g1599
  (
    n1634,
    n1481,
    n1486,
    n1141,
    n1476
  );


  nor
  g1600
  (
    n1632,
    n1484,
    n1492,
    n1627,
    n1480
  );


  xor
  g1601
  (
    n1630,
    n1141,
    n1477,
    n1490,
    n1478
  );


  xnor
  g1602
  (
    n1631,
    n1626,
    n1488,
    n1482,
    n1627
  );


  nor
  g1603
  (
    n1633,
    n1479,
    n1474,
    n1487,
    n1475
  );


  and
  g1604
  (
    n1629,
    n1627,
    n1489,
    n1485,
    n1483
  );


  xor
  g1605
  (
    n1635,
    n1526,
    n1634,
    n1633,
    n1358
  );


  xnor
  g1606
  (
    n1636,
    n1358,
    n1357,
    n1525
  );


  xor
  g1607
  (
    n1638,
    n1635,
    n1145,
    n1636
  );


  xnor
  g1608
  (
    n1642,
    n1144,
    n1143,
    n1146
  );


  and
  g1609
  (
    n1643,
    n1636,
    n1358,
    n1635,
    n1146
  );


  nand
  g1610
  (
    n1641,
    n1143,
    n1142,
    n1635,
    n1146
  );


  xor
  g1611
  (
    n1637,
    n1141,
    n1145,
    n1142
  );


  xnor
  g1612
  (
    n1639,
    n1144,
    n1142,
    n1636
  );


  or
  g1613
  (
    n1640,
    n1144,
    n1144,
    n1143,
    n1145
  );


  buf
  g1614
  (
    n1644,
    n1643
  );


  nand
  g1615
  (
    n1646,
    n1644,
    n1147
  );


  nor
  g1616
  (
    n1645,
    n1146,
    n1148,
    n1147,
    n1644
  );


  xor
  g1617
  (
    n1647,
    n1645,
    n1595
  );


  nor
  g1618
  (
    n1650,
    n1151,
    n1149,
    n1148,
    n1150
  );


  nor
  g1619
  (
    n1648,
    n1150,
    n1647,
    n1149
  );


  nor
  g1620
  (
    n1651,
    n1148,
    n1150,
    n1647
  );


  xor
  g1621
  (
    n1649,
    n1150,
    n1149,
    n1148
  );


  and
  g1622
  (
    n1658,
    n1651,
    n1160,
    n1158,
    n1153
  );


  and
  g1623
  (
    n1656,
    n1155,
    n1157,
    n1159
  );


  nor
  g1624
  (
    n1664,
    n1160,
    n1152,
    n1161,
    n1649
  );


  xor
  g1625
  (
    n1659,
    n1160,
    n1151,
    n1161,
    n1648
  );


  xor
  g1626
  (
    n1655,
    n1152,
    n1159,
    n1154,
    n1153
  );


  nor
  g1627
  (
    n1666,
    n1161,
    n1153,
    n1152,
    n1160
  );


  or
  g1628
  (
    n1654,
    n1156,
    n1650,
    n485,
    n1649
  );


  nand
  g1629
  (
    n1667,
    n1162,
    n1151,
    n1650
  );


  nand
  g1630
  (
    n1657,
    n1651,
    n1650,
    n1156
  );


  xnor
  g1631
  (
    n1652,
    n1161,
    n1649,
    n1162,
    n1154
  );


  and
  g1632
  (
    n1653,
    n1648,
    n1158,
    n1156,
    n1157
  );


  nor
  g1633
  (
    n1661,
    n1159,
    n1155,
    n1152
  );


  or
  g1634
  (
    n1660,
    n1650,
    n1648,
    n1158,
    n1155
  );


  xor
  g1635
  (
    n1662,
    n1154,
    n1157,
    n1649,
    n1162
  );


  xnor
  g1636
  (
    n1663,
    n1158,
    n1651,
    n1153
  );


  or
  g1637
  (
    n1665,
    n1162,
    n1157,
    n1648,
    n1154
  );


  not
  g1638
  (
    n1669,
    n1655
  );


  and
  g1639
  (
    n1668,
    n1654,
    n1652
  );


  and
  g1640
  (
    n1671,
    n1657,
    n1659
  );


  or
  g1641
  (
    n1670,
    n1653,
    n1660,
    n1656,
    n1658
  );


  xnor
  g1642
  (
    n1675,
    n1668,
    n1669,
    n1671,
    n1363
  );


  nor
  g1643
  (
    n1678,
    n1670,
    n1670,
    n1361,
    n1363
  );


  xnor
  g1644
  (
    n1676,
    n1363,
    n1359
  );


  nand
  g1645
  (
    n1679,
    n1362,
    n1362,
    n1358,
    n1361
  );


  or
  g1646
  (
    n1673,
    n1360,
    n1362,
    n1361
  );


  or
  g1647
  (
    n1677,
    n1363,
    n1359,
    n1360,
    n1670
  );


  and
  g1648
  (
    n1674,
    n1671,
    n1362,
    n1360,
    n1364
  );


  nand
  g1649
  (
    n1672,
    n1364,
    n1670,
    n1646,
    n1360
  );


  xor
  g1650
  (
    n1680,
    n1672,
    n1596,
    n1597
  );


  nor
  g1651
  (
    n1681,
    n1596,
    n1597,
    n1674,
    n1673
  );


  nor
  g1652
  (
    n1682,
    n1597,
    n1675,
    n1596
  );


  xnor
  g1653
  (
    n1686,
    n1532,
    n1528,
    n1531,
    n1680
  );


  xor
  g1654
  (
    n1688,
    n1530,
    n1605,
    n1611,
    n1681
  );


  nor
  g1655
  (
    n1685,
    n1612,
    n1527,
    n1602,
    n1609
  );


  and
  g1656
  (
    n1689,
    n1603,
    n1606,
    n1533,
    n1682
  );


  nand
  g1657
  (
    n1690,
    n1534,
    n1537,
    n1536,
    n1682
  );


  or
  g1658
  (
    n1691,
    n1608,
    n1607,
    n1610,
    n1681
  );


  and
  g1659
  (
    n1684,
    n1681,
    n1682,
    n1613,
    n1535
  );


  nand
  g1660
  (
    n1687,
    n1614,
    n1604,
    n1529,
    n1615
  );


  nand
  g1661
  (
    n1683,
    n1600,
    n1681,
    n1682,
    n1601
  );


  nand
  g1662
  (
    n1692,
    n1684,
    n1683
  );


  nand
  g1663
  (
    n1693,
    n1671,
    n1692
  );


  xnor
  g1664
  (
    n1694,
    n1671,
    n899,
    n1692
  );


  or
  g1665
  (
    n1702,
    n1167,
    n1167,
    n1166,
    n1694
  );


  xor
  g1666
  (
    n1700,
    n1163,
    n1693,
    n1165,
    n1164
  );


  nand
  g1667
  (
    n1698,
    n1693,
    n1165,
    n1163
  );


  xnor
  g1668
  (
    n1696,
    n1166,
    n1694,
    n1168
  );


  and
  g1669
  (
    n1695,
    n1164,
    n1164,
    n1163,
    n1166
  );


  xor
  g1670
  (
    n1697,
    n1165,
    n1693,
    n1167
  );


  nor
  g1671
  (
    n1699,
    n1168,
    n1694,
    n1164,
    n1165
  );


  or
  g1672
  (
    n1701,
    n1693,
    n1694,
    n1166,
    n1168
  );


  nand
  g1673
  (
    n1713,
    n1698,
    n1500,
    n1504,
    n1511
  );


  and
  g1674
  (
    n1709,
    n1514,
    n1702,
    n1501,
    n1515
  );


  nand
  g1675
  (
    n1712,
    n1701,
    n1170,
    n1662,
    n1503
  );


  xnor
  g1676
  (
    n1703,
    n1699,
    n1702,
    n1169,
    n1701
  );


  xnor
  g1677
  (
    n1708,
    n1502,
    n1663,
    n1509,
    n1700
  );


  or
  g1678
  (
    n1707,
    n1661,
    n1169,
    n1170,
    n1515
  );


  xor
  g1679
  (
    n1717,
    n1697,
    n1497,
    n1517,
    n1513
  );


  or
  g1680
  (
    n1706,
    n1517,
    n1510,
    n1498,
    n1170
  );


  xor
  g1681
  (
    n1714,
    n1662,
    n1700,
    n1702,
    n1506
  );


  nor
  g1682
  (
    n1704,
    n1170,
    n1662,
    n1696,
    n1695
  );


  nor
  g1683
  (
    n1711,
    n1516,
    n1505,
    n1702,
    n1701
  );


  xnor
  g1684
  (
    n1710,
    n1169,
    n1662,
    n1517,
    n1507
  );


  xor
  g1685
  (
    n1716,
    n1169,
    n1661,
    n1499,
    n1508
  );


  nand
  g1686
  (
    n1715,
    n1512,
    n1494,
    n1701,
    n1661
  );


  nand
  g1687
  (
    n1705,
    n1495,
    n1493,
    n1516,
    n1496
  );


  xnor
  g1688
  (
    n1718,
    n1703,
    n1171
  );


  nor
  g1689
  (
    n1719,
    n1618,
    n1718,
    n1567
  );


  nand
  g1690
  (
    n1720,
    n1568,
    n1616,
    n1718,
    n1617
  );


  and
  g1691
  (
    n1721,
    n1719,
    n1364
  );


  not
  g1692
  (
    n1723,
    n1721
  );


  not
  g1693
  (
    n1722,
    n1721
  );


  and
  g1694
  (
    n1731,
    n1717,
    n1707,
    n1704,
    n1722
  );


  xor
  g1695
  (
    n1724,
    n1710,
    n1715,
    n1723
  );


  xor
  g1696
  (
    n1729,
    n1722,
    n1716,
    n1714,
    n1708
  );


  and
  g1697
  (
    n1726,
    n1715,
    n1723,
    n1722,
    n1709
  );


  or
  g1698
  (
    n1730,
    n1716,
    n1706,
    n1712,
    n1717
  );


  xor
  g1699
  (
    n1727,
    n1723,
    n1722,
    n1711,
    n1717
  );


  nor
  g1700
  (
    n1728,
    n1705,
    n1715,
    n1716,
    n1717
  );


  or
  g1701
  (
    n1725,
    n1716,
    n1715,
    n1714,
    n1713
  );


  nor
  g1702
  (
    n1734,
    n1727,
    n900,
    n1725,
    n1625
  );


  xnor
  g1703
  (
    n1733,
    n1726,
    n1623,
    n1620,
    n1622
  );


  nand
  g1704
  (
    n1732,
    n1724,
    n900,
    n899
  );


  or
  g1705
  (
    n1735,
    n900,
    n1621,
    n1624,
    n1619
  );


  xnor
  g1706
  (
    n1736,
    n1735,
    n1720
  );


  buf
  g1707
  (
    n1738,
    n1736
  );


  nand
  g1708
  (
    n1737,
    n1736,
    n1517,
    n1395
  );


  and
  g1709
  (
    n1739,
    n1738,
    n1364,
    n1171
  );


  nand
  g1710
  (
    n1740,
    n1739,
    n1663
  );


  xnor
  g1711
  (
    n1741,
    n1664,
    n1664,
    n1663,
    n1739
  );


  and
  g1712
  (
    n1747,
    n1176,
    n1740,
    n1173,
    n1172
  );


  nor
  g1713
  (
    n1743,
    n1740,
    n1172,
    n1176
  );


  nor
  g1714
  (
    n1742,
    n1740,
    n1175,
    n1177,
    n1174
  );


  or
  g1715
  (
    n1749,
    n1177,
    n1741,
    n1173,
    n1740
  );


  nand
  g1716
  (
    n1746,
    n1175,
    n1173,
    n1177,
    n1174
  );


  or
  g1717
  (
    n1748,
    n1171,
    n1175,
    n1174,
    n1741
  );


  and
  g1718
  (
    n1744,
    n1176,
    n1173,
    n1172,
    n1741
  );


  xnor
  g1719
  (
    n1745,
    n1175,
    n1741,
    n1174,
    n1172
  );


  nand
  g1720
  (
    n1750,
    n1179,
    n1180,
    n1178
  );


  and
  g1721
  (
    n1753,
    n1177,
    n1178,
    n1742
  );


  nand
  g1722
  (
    n1752,
    n1178,
    n1745,
    n1180,
    n1179
  );


  nand
  g1723
  (
    n1751,
    n1743,
    n1179,
    n1744
  );


  xor
  g1724
  (
    n1754,
    n1729,
    n1664,
    n1665
  );


  xor
  g1725
  (
    n1756,
    n1750,
    n1728,
    n1751
  );


  or
  g1726
  (
    n1755,
    n1730,
    n1729,
    n1752,
    n1666
  );


  and
  g1727
  (
    n1757,
    n1753,
    n1665
  );


  nand
  g1728
  (
    n1762,
    n1365,
    n1757,
    n1368,
    n1369
  );


  nand
  g1729
  (
    n1761,
    n1366,
    n1755,
    n1756,
    n1370
  );


  xor
  g1730
  (
    n1758,
    n1757,
    n1755,
    n1687,
    n1366
  );


  nand
  g1731
  (
    n1764,
    n1368,
    n1366,
    n1686,
    n1365
  );


  or
  g1732
  (
    n1760,
    n1365,
    n1369,
    n1367,
    n1757
  );


  nand
  g1733
  (
    n1759,
    n1368,
    n1370,
    n1754
  );


  or
  g1734
  (
    n1766,
    n1367,
    n1369,
    n1685,
    n1757
  );


  nor
  g1735
  (
    n1763,
    n1369,
    n1367,
    n1366,
    n1370
  );


  xnor
  g1736
  (
    n1765,
    n1368,
    n1367,
    n1756,
    n1365
  );


  buf
  g1737
  (
    n1767,
    n1759
  );


  not
  g1738
  (
    n1769,
    n1761
  );


  xor
  g1739
  (
    n1770,
    n1760,
    n1689
  );


  nor
  g1740
  (
    n1768,
    n1758,
    n1688,
    n1690,
    n1691
  );


  buf
  g1741
  (
    n1773,
    n1767
  );


  buf
  g1742
  (
    n1771,
    n1768
  );


  not
  g1743
  (
    n1772,
    n1767
  );


  not
  g1744
  (
    n1774,
    n1768
  );


  not
  g1745
  (
    n1775,
    n1767
  );


  not
  g1746
  (
    n1779,
    n1772
  );


  not
  g1747
  (
    n1777,
    n1181
  );


  not
  g1748
  (
    n1788,
    n1184
  );


  buf
  g1749
  (
    n1785,
    n1771
  );


  not
  g1750
  (
    n1784,
    n1569
  );


  not
  g1751
  (
    n1792,
    n1183
  );


  not
  g1752
  (
    n1790,
    n1775
  );


  buf
  g1753
  (
    n1780,
    n1182
  );


  or
  g1754
  (
    n1781,
    n1183,
    n1775,
    n1772,
    n1184
  );


  xor
  g1755
  (
    n1782,
    n1185,
    n1186,
    n1775
  );


  nor
  g1756
  (
    n1786,
    n1774,
    n1678,
    n1182,
    n1183
  );


  nand
  g1757
  (
    n1776,
    n1183,
    n1774
  );


  xnor
  g1758
  (
    n1793,
    n1186,
    n1773,
    n1679
  );


  and
  g1759
  (
    n1783,
    n1185,
    n1181,
    n1773
  );


  nand
  g1760
  (
    n1778,
    n1677,
    n1182,
    n1773,
    n1181
  );


  xnor
  g1761
  (
    n1787,
    n1184,
    n1184,
    n1676,
    n1182
  );


  nand
  g1762
  (
    n1791,
    n1186,
    n1772,
    n1180,
    n1185
  );


  or
  g1763
  (
    n1789,
    n1772,
    n1185,
    n1775,
    n1771
  );


  nor
  g1764
  (
    n1795,
    n1193,
    n1193,
    n1187,
    n1197
  );


  nand
  g1765
  (
    n1794,
    n1785,
    n1790,
    n1189,
    n1194
  );


  nor
  g1766
  (
    n1807,
    n1195,
    n1195,
    n1191,
    n1788
  );


  nor
  g1767
  (
    n1797,
    n1190,
    n1779,
    n1191,
    n1197
  );


  xnor
  g1768
  (
    n1808,
    n1191,
    n1787,
    n1783,
    n1792
  );


  nand
  g1769
  (
    n1810,
    n1190,
    n1188,
    n1782,
    n1198
  );


  or
  g1770
  (
    n1803,
    n1786,
    n1188,
    n1198
  );


  nand
  g1771
  (
    n1798,
    n1197,
    n1195,
    n1199,
    n1191
  );


  xnor
  g1772
  (
    n1805,
    n1190,
    n1198,
    n1777,
    n1784
  );


  nor
  g1773
  (
    n1809,
    n1187,
    n1776,
    n1189
  );


  xnor
  g1774
  (
    KeyWire_0_11,
    n1199,
    n1196,
    n1189,
    n1194
  );


  and
  g1775
  (
    n1802,
    n1791,
    n1193,
    n1781,
    n1192
  );


  nand
  g1776
  (
    n1801,
    n1193,
    n1194,
    n1187
  );


  or
  g1777
  (
    n1796,
    n1192,
    n1195,
    n1188,
    n1197
  );


  xor
  g1778
  (
    n1806,
    n1192,
    n1196,
    n1778
  );


  and
  g1779
  (
    n1800,
    n1196,
    n1199,
    n1780,
    n1190
  );


  or
  g1780
  (
    n1804,
    n1192,
    n1188,
    n1187,
    n1789
  );


  nor
  g1781
  (
    n1814,
    n1200,
    n1201,
    n1746,
    n1797
  );


  or
  g1782
  (
    n1813,
    n1794,
    n1748,
    n1795,
    n1749
  );


  nand
  g1783
  (
    n1812,
    n1200,
    n1201,
    n1199
  );


  xor
  g1784
  (
    n1811,
    n1200,
    n1200,
    n1796,
    n1747
  );


  not
  g1785
  (
    n1817,
    n1812
  );


  not
  g1786
  (
    n1816,
    n1813
  );


  buf
  g1787
  (
    n1815,
    n1811
  );


  buf
  g1788
  (
    n1818,
    n1814
  );


  buf
  g1789
  (
    n1819,
    n1814
  );


  not
  g1790
  (
    n1835,
    n1202
  );


  not
  g1791
  (
    n1826,
    n1212
  );


  buf
  g1792
  (
    n1822,
    n1816
  );


  not
  g1793
  (
    n1831,
    n1816
  );


  and
  g1794
  (
    n1838,
    n1211,
    n1212,
    n1819,
    n1818
  );


  nand
  g1795
  (
    n1827,
    n1204,
    n1207,
    n1211,
    n1818
  );


  nor
  g1796
  (
    n1824,
    n1204,
    n1208,
    n1211,
    n1201
  );


  nand
  g1797
  (
    n1836,
    n1210,
    n1203,
    n1202,
    n1206
  );


  nand
  g1798
  (
    n1832,
    n1210,
    n1202,
    n1205,
    n1208
  );


  nand
  g1799
  (
    n1833,
    n1210,
    n1209,
    n1818,
    n1211
  );


  or
  g1800
  (
    n1829,
    n1206,
    n1817,
    n1210,
    n1212
  );


  or
  g1801
  (
    n1821,
    n1209,
    n1208,
    n1815
  );


  xor
  g1802
  (
    n1825,
    n1209,
    n1212,
    n1207,
    n1819
  );


  and
  g1803
  (
    n1828,
    n1209,
    n1818,
    n1205,
    n1207
  );


  nand
  g1804
  (
    n1830,
    n1202,
    n1815,
    n1205
  );


  or
  g1805
  (
    n1823,
    n1204,
    n1207,
    n1817
  );


  xnor
  g1806
  (
    n1837,
    n1815,
    n1203,
    n1206
  );


  or
  g1807
  (
    n1820,
    n1203,
    n1206,
    n1819
  );


  or
  g1808
  (
    n1834,
    n1204,
    n1816,
    n1817
  );


  not
  g1809
  (
    n1845,
    n1821
  );


  not
  g1810
  (
    n1841,
    n1827
  );


  buf
  g1811
  (
    n1843,
    n1824
  );


  not
  g1812
  (
    n1839,
    n1820
  );


  not
  g1813
  (
    n1844,
    n1826
  );


  buf
  g1814
  (
    n1846,
    n1823
  );


  not
  g1815
  (
    n1840,
    n1822
  );


  buf
  g1816
  (
    n1842,
    n1825
  );


  nand
  g1817
  (
    n1859,
    n1802,
    n1384,
    n1381
  );


  xnor
  g1818
  (
    n1875,
    n1769,
    n1383,
    n1380,
    n1381
  );


  nor
  g1819
  (
    n1870,
    n1379,
    n1842,
    n1844,
    n1377
  );


  xnor
  g1820
  (
    KeyWire_0_4,
    n1666,
    n1844,
    n1371,
    n1379
  );


  or
  g1821
  (
    n1856,
    n1379,
    n1840,
    n1846,
    n1372
  );


  xor
  g1822
  (
    n1877,
    n1807,
    n1809,
    n1799,
    n1377
  );


  xnor
  g1823
  (
    n1848,
    n1842,
    n1730,
    n1376,
    n1381
  );


  and
  g1824
  (
    n1874,
    n1770,
    n1845,
    n1385,
    n1375
  );


  or
  g1825
  (
    n1850,
    n1731,
    n1839,
    n1378,
    n1842
  );


  xnor
  g1826
  (
    n1876,
    n1841,
    n1804,
    n1840,
    n1844
  );


  nor
  g1827
  (
    n1869,
    n1770,
    n1374,
    n1840,
    n1372
  );


  xor
  g1828
  (
    n1853,
    n1386,
    n1798,
    n1803,
    n1801
  );


  or
  g1829
  (
    n1857,
    n1386,
    n1843,
    n1845
  );


  nor
  g1830
  (
    n1863,
    n1846,
    n1378,
    n1371,
    n1372
  );


  nor
  g1831
  (
    n1852,
    n1841,
    n1846,
    n1769
  );


  or
  g1832
  (
    n1878,
    n1839,
    n1840,
    n1374,
    n1810
  );


  nand
  g1833
  (
    n1854,
    n1377,
    n1730,
    n1384,
    n1666
  );


  nand
  g1834
  (
    n1862,
    n1842,
    n1380,
    n1376,
    n1381
  );


  xor
  g1835
  (
    n1860,
    n1382,
    n1770,
    n1374,
    n1805
  );


  xnor
  g1836
  (
    n1872,
    n1373,
    n1845,
    n1382,
    n1839
  );


  or
  g1837
  (
    n1868,
    n1770,
    n1383,
    n1371,
    n1385
  );


  nor
  g1838
  (
    n1866,
    n1768,
    n1376,
    n1375,
    n1385
  );


  xor
  g1839
  (
    n1849,
    n1382,
    n1376,
    n1731,
    n1843
  );


  or
  g1840
  (
    n1867,
    n1375,
    n1374,
    n1373,
    n1769
  );


  xnor
  g1841
  (
    n1873,
    n1380,
    n1380,
    n1373,
    n1382
  );


  xor
  g1842
  (
    n1847,
    n1379,
    n1731,
    n1385,
    n1375
  );


  nand
  g1843
  (
    n1864,
    n1371,
    n1377,
    n1383,
    n1384
  );


  xor
  g1844
  (
    n1861,
    n1844,
    n1808,
    n1806,
    n1386
  );


  and
  g1845
  (
    n1851,
    n1800,
    n1378,
    n1843
  );


  nand
  g1846
  (
    n1858,
    n1730,
    n1386,
    n1843,
    n1839
  );


  xor
  g1847
  (
    n1865,
    n1768,
    n1769,
    n1841,
    n1373
  );


  or
  g1848
  (
    n1855,
    n1383,
    n1841,
    n1731,
    n1372
  );


  nand
  g1849
  (
    n1880,
    n1857,
    n1848,
    n1858,
    n1854
  );


  or
  g1850
  (
    n1879,
    n1858,
    n1855,
    n1853,
    n1857
  );


  or
  g1851
  (
    n1881,
    n1851,
    n1853,
    n1857
  );


  nor
  g1852
  (
    n1882,
    n1854,
    n1858,
    n1855,
    n1852
  );


  nand
  g1853
  (
    n1883,
    n1849,
    n1856,
    n1847
  );


  xnor
  g1854
  (
    n1884,
    n1858,
    n1851,
    n1850,
    n1852
  );


  buf
  g1855
  (
    n1890,
    n1883
  );


  buf
  g1856
  (
    n1885,
    n1884
  );


  not
  g1857
  (
    n1889,
    n1793
  );


  buf
  g1858
  (
    n1886,
    n1882
  );


  buf
  g1859
  (
    n1888,
    n1881
  );


  and
  g1860
  (
    n1887,
    n1859,
    n1880,
    n1879
  );


  xnor
  g1861
  (
    n1892,
    n1890,
    n1218,
    n1224,
    n1221
  );


  nand
  g1862
  (
    n1891,
    n1888,
    n1887,
    n1885,
    n1830
  );


  xor
  g1863
  (
    n1909,
    n1215,
    n1889,
    n1667,
    n1221
  );


  xor
  g1864
  (
    n1902,
    n1215,
    n1890,
    n1222,
    n1223
  );


  or
  g1865
  (
    n1894,
    n1833,
    n1226,
    n1217,
    n1835
  );


  xor
  g1866
  (
    n1895,
    n1889,
    n1888,
    n1220,
    n1887
  );


  nor
  g1867
  (
    n1893,
    n1225,
    n1217,
    n1219,
    n1886
  );


  nand
  g1868
  (
    n1911,
    n1222,
    n1832,
    n1219,
    n1213
  );


  xor
  g1869
  (
    n1905,
    n1885,
    n1888,
    n1222,
    n1215
  );


  or
  g1870
  (
    n1910,
    n1829,
    n1219,
    n1221,
    n1886
  );


  nand
  g1871
  (
    n1904,
    n1226,
    n1886,
    n1218,
    n1887
  );


  or
  g1872
  (
    n1907,
    n1220,
    n1834,
    n1219,
    n1216
  );


  and
  g1873
  (
    n1898,
    n1889,
    n1828,
    n1890,
    n1831
  );


  and
  g1874
  (
    n1896,
    n1216,
    n1223,
    n1213,
    n1217
  );


  and
  g1875
  (
    n1901,
    n1217,
    n1215,
    n1224,
    n1223
  );


  xnor
  g1876
  (
    n1912,
    n1220,
    n1667,
    n1886,
    n1888
  );


  nor
  g1877
  (
    KeyWire_0_8,
    n1889,
    n1837,
    n1213,
    n1887
  );


  nand
  g1878
  (
    n1906,
    n1218,
    n1226,
    n1885,
    n1667
  );


  xnor
  g1879
  (
    n1900,
    n1221,
    n1220,
    n1223,
    n1225
  );


  and
  g1880
  (
    n1897,
    n1218,
    n1216,
    n1890,
    n1225
  );


  xnor
  g1881
  (
    n1913,
    n1666,
    n1838,
    n1226,
    n1885
  );


  nor
  g1882
  (
    n1903,
    n1224,
    n1214
  );


  xnor
  g1883
  (
    n1914,
    n1225,
    n1667,
    n1836,
    n1224
  );


  nor
  g1884
  (
    n1908,
    n1213,
    n1216,
    n1222,
    n1214
  );


  xor
  g1885
  (
    n1921,
    n1859,
    n1864,
    n1580,
    n1765
  );


  xor
  g1886
  (
    n1922,
    n1906,
    n1908,
    n1901,
    n1864
  );


  or
  g1887
  (
    n1920,
    n1866,
    n1867,
    n1905,
    n1869
  );


  xor
  g1888
  (
    n1933,
    n1866,
    n1862,
    n1863,
    n1904
  );


  nand
  g1889
  (
    n1915,
    n1576,
    n1575,
    n1587,
    n1762
  );


  nand
  g1890
  (
    n1931,
    n1868,
    n1891,
    n1579,
    n1870
  );


  xor
  g1891
  (
    n1932,
    n1907,
    n1894,
    n1585,
    n1860
  );


  and
  g1892
  (
    n1937,
    n1583,
    n1860,
    n1865
  );


  or
  g1893
  (
    n1924,
    n1584,
    n1764,
    n1868,
    n1766
  );


  and
  g1894
  (
    n1917,
    n1863,
    n1863,
    n1903,
    n1895
  );


  or
  g1895
  (
    n1916,
    n1896,
    n1570,
    n1862,
    n1864
  );


  xnor
  g1896
  (
    n1927,
    n1862,
    n1869,
    n1893,
    n1571
  );


  xor
  g1897
  (
    n1926,
    n1897,
    n1909,
    n1911,
    n1900
  );


  and
  g1898
  (
    n1936,
    n1859,
    n1581,
    n1861,
    n1870
  );


  xnor
  g1899
  (
    n1928,
    n1910,
    n1869,
    n1899,
    n1586
  );


  and
  g1900
  (
    n1930,
    n1869,
    n1868,
    n1860,
    n1582
  );


  xnor
  g1901
  (
    n1925,
    n1861,
    n1574,
    n1867,
    n1865
  );


  or
  g1902
  (
    n1935,
    n1577,
    n1867,
    n1892,
    n1573
  );


  xnor
  g1903
  (
    n1918,
    n1862,
    n1867,
    n1861,
    n1763
  );


  nand
  g1904
  (
    n1919,
    n1866,
    n1865,
    n1870,
    n1912
  );


  and
  g1905
  (
    n1934,
    n1866,
    n1913,
    n1859,
    n1863
  );


  xnor
  g1906
  (
    n1929,
    n1868,
    n1578,
    n1865,
    n1861
  );


  nand
  g1907
  (
    n1923,
    n1902,
    n1864,
    n1898,
    n1572
  );


  nor
  g1908
  (
    n1938,
    n1872,
    n1871,
    n1873
  );


  xor
  g1909
  (
    n1940,
    n1870,
    n1917,
    n1872,
    n1918
  );


  xnor
  g1910
  (
    n1939,
    n1871,
    n1872,
    n1915
  );


  nor
  g1911
  (
    n1941,
    n1873,
    n1916,
    n1871
  );


  xnor
  g1912
  (
    n1943,
    n1873,
    n1874
  );


  nor
  g1913
  (
    n1942,
    n1941,
    n1874,
    n1940,
    n1875
  );


  nor
  g1914
  (
    n1944,
    n1875,
    n1942
  );


  xor
  g1915
  (
    n1945,
    n1875,
    n1944,
    n1876,
    n1877
  );


  xnor
  g1916
  (
    n1946,
    n1944,
    n1876,
    n1877
  );


  xor
  g1917
  (
    n1947,
    n1875,
    n1944,
    n1876
  );


  xnor
  g1918
  (
    n1948,
    n1921,
    n1923,
    n1924,
    n1920
  );


  or
  g1919
  (
    n1949,
    n1946,
    n1947,
    n1919,
    n1922
  );


  and
  g1920
  (
    n1950,
    n1878,
    n1878,
    n1877,
    n1949
  );


  and
  g1921
  (
    n1952,
    n1914,
    n1925,
    n1878,
    n1943
  );


  xnor
  g1922
  (
    n1951,
    n1950,
    n1950,
    n1943,
    n1878
  );


  xnor
  g1923
  (
    n1954,
    n1928,
    n1927,
    n1934,
    n1930
  );


  and
  g1924
  (
    n1955,
    n1952,
    n1931,
    n1926,
    n1951
  );


  nor
  g1925
  (
    n1953,
    n1952,
    n1936,
    n1937,
    n1932
  );


  xnor
  g1926
  (
    n1956,
    n1951,
    n1935,
    n1929,
    n1933
  );


  nand
  g1927
  (
    n1957,
    n1954,
    n1956,
    n1955,
    n1953
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n727,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n563,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1392,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n130,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1871,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n102,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n944,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1097,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n1899,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n658,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n229,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1799,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n1210,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1442,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1477,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1247,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule

