// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_2173_26_6 written by SynthGen on 2021/06/15 15:05:36
module Stat_2173_26_6( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45,
 n1805, n1807, n1798, n1810, n1804, n1806, n1802, n1801,
 n1808, n1811, n1800, n1809, n1803, n1823, n1819, n1830,
 n1828, n2195, n2217, n2210, n2212, n2215, n2206, n2199,
 n2200, n2198, n2213, n2211, n2207, n2194, n2196, n2218,
 n2214, n2202, n2204, n2193, n2201, n2192, n2203, n2208,
 n2197, n2209, n2205, n2216);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45;

output n1805, n1807, n1798, n1810, n1804, n1806, n1802, n1801,
 n1808, n1811, n1800, n1809, n1803, n1823, n1819, n1830,
 n1828, n2195, n2217, n2210, n2212, n2215, n2206, n2199,
 n2200, n2198, n2213, n2211, n2207, n2194, n2196, n2218,
 n2214, n2202, n2204, n2193, n2201, n2192, n2203, n2208,
 n2197, n2209, n2205, n2216;

wire n46, n47, n48, n49, n50, n51, n52, n53,
 n54, n55, n56, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n67, n68, n69,
 n70, n71, n72, n73, n74, n75, n76, n77,
 n78, n79, n80, n81, n82, n83, n84, n85,
 n86, n87, n88, n89, n90, n91, n92, n93,
 n94, n95, n96, n97, n98, n99, n100, n101,
 n102, n103, n104, n105, n106, n107, n108, n109,
 n110, n111, n112, n113, n114, n115, n116, n117,
 n118, n119, n120, n121, n122, n123, n124, n125,
 n126, n127, n128, n129, n130, n131, n132, n133,
 n134, n135, n136, n137, n138, n139, n140, n141,
 n142, n143, n144, n145, n146, n147, n148, n149,
 n150, n151, n152, n153, n154, n155, n156, n157,
 n158, n159, n160, n161, n162, n163, n164, n165,
 n166, n167, n168, n169, n170, n171, n172, n173,
 n174, n175, n176, n177, n178, n179, n180, n181,
 n182, n183, n184, n185, n186, n187, n188, n189,
 n190, n191, n192, n193, n194, n195, n196, n197,
 n198, n199, n200, n201, n202, n203, n204, n205,
 n206, n207, n208, n209, n210, n211, n212, n213,
 n214, n215, n216, n217, n218, n219, n220, n221,
 n222, n223, n224, n225, n226, n227, n228, n229,
 n230, n231, n232, n233, n234, n235, n236, n237,
 n238, n239, n240, n241, n242, n243, n244, n245,
 n246, n247, n248, n249, n250, n251, n252, n253,
 n254, n255, n256, n257, n258, n259, n260, n261,
 n262, n263, n264, n265, n266, n267, n268, n269,
 n270, n271, n272, n273, n274, n275, n276, n277,
 n278, n279, n280, n281, n282, n283, n284, n285,
 n286, n287, n288, n289, n290, n291, n292, n293,
 n294, n295, n296, n297, n298, n299, n300, n301,
 n302, n303, n304, n305, n306, n307, n308, n309,
 n310, n311, n312, n313, n314, n315, n316, n317,
 n318, n319, n320, n321, n322, n323, n324, n325,
 n326, n327, n328, n329, n330, n331, n332, n333,
 n334, n335, n336, n337, n338, n339, n340, n341,
 n342, n343, n344, n345, n346, n347, n348, n349,
 n350, n351, n352, n353, n354, n355, n356, n357,
 n358, n359, n360, n361, n362, n363, n364, n365,
 n366, n367, n368, n369, n370, n371, n372, n373,
 n374, n375, n376, n377, n378, n379, n380, n381,
 n382, n383, n384, n385, n386, n387, n388, n389,
 n390, n391, n392, n393, n394, n395, n396, n397,
 n398, n399, n400, n401, n402, n403, n404, n405,
 n406, n407, n408, n409, n410, n411, n412, n413,
 n414, n415, n416, n417, n418, n419, n420, n421,
 n422, n423, n424, n425, n426, n427, n428, n429,
 n430, n431, n432, n433, n434, n435, n436, n437,
 n438, n439, n440, n441, n442, n443, n444, n445,
 n446, n447, n448, n449, n450, n451, n452, n453,
 n454, n455, n456, n457, n458, n459, n460, n461,
 n462, n463, n464, n465, n466, n467, n468, n469,
 n470, n471, n472, n473, n474, n475, n476, n477,
 n478, n479, n480, n481, n482, n483, n484, n485,
 n486, n487, n488, n489, n490, n491, n492, n493,
 n494, n495, n496, n497, n498, n499, n500, n501,
 n502, n503, n504, n505, n506, n507, n508, n509,
 n510, n511, n512, n513, n514, n515, n516, n517,
 n518, n519, n520, n521, n522, n523, n524, n525,
 n526, n527, n528, n529, n530, n531, n532, n533,
 n534, n535, n536, n537, n538, n539, n540, n541,
 n542, n543, n544, n545, n546, n547, n548, n549,
 n550, n551, n552, n553, n554, n555, n556, n557,
 n558, n559, n560, n561, n562, n563, n564, n565,
 n566, n567, n568, n569, n570, n571, n572, n573,
 n574, n575, n576, n577, n578, n579, n580, n581,
 n582, n583, n584, n585, n586, n587, n588, n589,
 n590, n591, n592, n593, n594, n595, n596, n597,
 n598, n599, n600, n601, n602, n603, n604, n605,
 n606, n607, n608, n609, n610, n611, n612, n613,
 n614, n615, n616, n617, n618, n619, n620, n621,
 n622, n623, n624, n625, n626, n627, n628, n629,
 n630, n631, n632, n633, n634, n635, n636, n637,
 n638, n639, n640, n641, n642, n643, n644, n645,
 n646, n647, n648, n649, n650, n651, n652, n653,
 n654, n655, n656, n657, n658, n659, n660, n661,
 n662, n663, n664, n665, n666, n667, n668, n669,
 n670, n671, n672, n673, n674, n675, n676, n677,
 n678, n679, n680, n681, n682, n683, n684, n685,
 n686, n687, n688, n689, n690, n691, n692, n693,
 n694, n695, n696, n697, n698, n699, n700, n701,
 n702, n703, n704, n705, n706, n707, n708, n709,
 n710, n711, n712, n713, n714, n715, n716, n717,
 n718, n719, n720, n721, n722, n723, n724, n725,
 n726, n727, n728, n729, n730, n731, n732, n733,
 n734, n735, n736, n737, n738, n739, n740, n741,
 n742, n743, n744, n745, n746, n747, n748, n749,
 n750, n751, n752, n753, n754, n755, n756, n757,
 n758, n759, n760, n761, n762, n763, n764, n765,
 n766, n767, n768, n769, n770, n771, n772, n773,
 n774, n775, n776, n777, n778, n779, n780, n781,
 n782, n783, n784, n785, n786, n787, n788, n789,
 n790, n791, n792, n793, n794, n795, n796, n797,
 n798, n799, n800, n801, n802, n803, n804, n805,
 n806, n807, n808, n809, n810, n811, n812, n813,
 n814, n815, n816, n817, n818, n819, n820, n821,
 n822, n823, n824, n825, n826, n827, n828, n829,
 n830, n831, n832, n833, n834, n835, n836, n837,
 n838, n839, n840, n841, n842, n843, n844, n845,
 n846, n847, n848, n849, n850, n851, n852, n853,
 n854, n855, n856, n857, n858, n859, n860, n861,
 n862, n863, n864, n865, n866, n867, n868, n869,
 n870, n871, n872, n873, n874, n875, n876, n877,
 n878, n879, n880, n881, n882, n883, n884, n885,
 n886, n887, n888, n889, n890, n891, n892, n893,
 n894, n895, n896, n897, n898, n899, n900, n901,
 n902, n903, n904, n905, n906, n907, n908, n909,
 n910, n911, n912, n913, n914, n915, n916, n917,
 n918, n919, n920, n921, n922, n923, n924, n925,
 n926, n927, n928, n929, n930, n931, n932, n933,
 n934, n935, n936, n937, n938, n939, n940, n941,
 n942, n943, n944, n945, n946, n947, n948, n949,
 n950, n951, n952, n953, n954, n955, n956, n957,
 n958, n959, n960, n961, n962, n963, n964, n965,
 n966, n967, n968, n969, n970, n971, n972, n973,
 n974, n975, n976, n977, n978, n979, n980, n981,
 n982, n983, n984, n985, n986, n987, n988, n989,
 n990, n991, n992, n993, n994, n995, n996, n997,
 n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
 n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
 n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
 n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
 n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
 n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
 n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
 n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
 n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
 n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
 n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
 n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
 n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
 n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
 n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
 n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
 n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
 n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
 n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
 n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
 n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
 n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
 n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
 n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
 n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
 n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
 n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
 n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
 n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
 n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
 n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
 n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
 n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
 n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
 n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
 n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
 n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
 n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
 n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
 n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
 n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
 n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
 n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
 n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
 n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
 n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
 n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
 n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
 n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
 n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
 n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
 n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
 n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
 n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
 n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
 n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
 n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
 n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
 n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
 n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
 n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
 n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
 n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
 n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
 n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
 n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
 n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
 n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
 n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
 n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
 n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
 n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
 n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
 n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
 n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
 n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
 n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
 n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
 n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
 n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
 n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
 n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
 n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
 n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
 n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
 n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
 n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
 n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
 n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
 n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
 n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
 n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
 n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
 n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
 n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
 n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
 n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
 n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
 n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
 n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
 n1799, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1820, n1821, n1822, n1824, n1825, n1826, n1827, n1829,
 n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
 n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
 n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
 n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
 n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
 n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
 n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
 n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
 n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
 n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
 n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
 n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
 n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
 n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
 n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
 n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
 n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
 n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
 n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
 n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
 n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
 n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
 n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
 n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
 n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
 n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
 n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
 n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
 n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
 n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
 n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
 n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
 n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
 n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
 n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
 n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
 n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
 n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
 n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
 n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
 n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
 n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
 n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
 n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
 n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
 n2191;

buf  g0 (n55, n34);
buf  g1 (n219, n5);
buf  g2 (n179, n35);
not  g3 (n102, n26);
buf  g4 (n213, n36);
not  g5 (n95, n6);
buf  g6 (n157, n22);
not  g7 (n49, n3);
not  g8 (n181, n34);
not  g9 (n206, n45);
buf  g10 (n84, n35);
buf  g11 (n187, n4);
not  g12 (n138, n38);
buf  g13 (n106, n2);
buf  g14 (n225, n16);
not  g15 (n107, n1);
not  g16 (n130, n19);
not  g17 (n197, n28);
not  g18 (n113, n20);
not  g19 (n87, n43);
buf  g20 (n203, n8);
not  g21 (n153, n37);
buf  g22 (n224, n33);
not  g23 (n63, n16);
buf  g24 (n75, n43);
not  g25 (n204, n20);
not  g26 (n146, n27);
not  g27 (n103, n25);
not  g28 (n51, n45);
not  g29 (n46, n43);
buf  g30 (n62, n45);
not  g31 (n142, n36);
not  g32 (n116, n1);
buf  g33 (n221, n40);
buf  g34 (n156, n10);
buf  g35 (n111, n39);
buf  g36 (n91, n7);
buf  g37 (n140, n42);
not  g38 (n152, n32);
buf  g39 (n126, n9);
buf  g40 (n124, n39);
not  g41 (n210, n13);
not  g42 (n121, n13);
not  g43 (n99, n33);
buf  g44 (n76, n17);
not  g45 (n77, n21);
buf  g46 (n155, n31);
not  g47 (n200, n21);
buf  g48 (n85, n11);
not  g49 (n81, n11);
not  g50 (n175, n9);
not  g51 (n169, n6);
not  g52 (n158, n23);
buf  g53 (n207, n36);
not  g54 (n164, n10);
not  g55 (n141, n29);
buf  g56 (n56, n25);
buf  g57 (n89, n20);
not  g58 (n60, n24);
buf  g59 (n74, n33);
buf  g60 (n47, n35);
not  g61 (n59, n19);
buf  g62 (n122, n41);
not  g63 (n123, n31);
not  g64 (n61, n25);
buf  g65 (n185, n18);
buf  g66 (n165, n33);
not  g67 (n195, n27);
buf  g68 (n192, n36);
not  g69 (n150, n30);
not  g70 (n216, n42);
not  g71 (n57, n40);
buf  g72 (n105, n18);
buf  g73 (n131, n8);
not  g74 (n220, n2);
buf  g75 (n73, n7);
buf  g76 (n208, n44);
not  g77 (n163, n12);
buf  g78 (n199, n8);
buf  g79 (n64, n30);
not  g80 (n151, n21);
buf  g81 (n96, n32);
buf  g82 (n170, n4);
buf  g83 (n92, n24);
not  g84 (n129, n18);
buf  g85 (n180, n27);
not  g86 (n120, n30);
buf  g87 (n79, n4);
not  g88 (n88, n6);
not  g89 (n72, n26);
buf  g90 (n173, n17);
not  g91 (n83, n2);
buf  g92 (n135, n18);
not  g93 (n148, n22);
not  g94 (n94, n44);
not  g95 (n69, n4);
not  g96 (n159, n2);
buf  g97 (n191, n5);
not  g98 (n209, n17);
buf  g99 (n145, n29);
not  g100 (n65, n15);
buf  g101 (n127, n38);
not  g102 (n125, n41);
not  g103 (n167, n3);
buf  g104 (n110, n10);
not  g105 (n48, n28);
not  g106 (n147, n30);
buf  g107 (n100, n44);
not  g108 (n90, n38);
buf  g109 (n149, n34);
not  g110 (n54, n19);
buf  g111 (n201, n12);
not  g112 (n176, n12);
not  g113 (n186, n37);
buf  g114 (n136, n19);
buf  g115 (n172, n37);
buf  g116 (n214, n42);
buf  g117 (n82, n23);
buf  g118 (n196, n9);
buf  g119 (n108, n1);
not  g120 (n217, n6);
not  g121 (n194, n10);
buf  g122 (n162, n20);
not  g123 (n86, n22);
not  g124 (n154, n35);
not  g125 (n52, n23);
not  g126 (n109, n38);
buf  g127 (n222, n7);
not  g128 (n97, n17);
not  g129 (n177, n28);
not  g130 (n188, n21);
not  g131 (n118, n5);
buf  g132 (n114, n41);
not  g133 (n171, n39);
not  g134 (n161, n26);
buf  g135 (n66, n14);
buf  g136 (n132, n3);
buf  g137 (n137, n32);
not  g138 (n198, n15);
buf  g139 (n139, n45);
buf  g140 (n183, n22);
not  g141 (n184, n39);
not  g142 (n115, n5);
buf  g143 (n58, n27);
buf  g144 (n223, n11);
not  g145 (n101, n11);
buf  g146 (n215, n25);
buf  g147 (n168, n41);
not  g148 (n67, n23);
not  g149 (n70, n40);
not  g150 (n166, n14);
buf  g151 (n143, n31);
not  g152 (n174, n13);
buf  g153 (n190, n42);
buf  g154 (n133, n14);
buf  g155 (n98, n32);
not  g156 (n202, n8);
not  g157 (n211, n29);
not  g158 (n128, n24);
not  g159 (n193, n15);
buf  g160 (n117, n40);
not  g161 (n80, n14);
not  g162 (n144, n31);
buf  g163 (n112, n16);
not  g164 (n205, n9);
not  g165 (n189, n24);
buf  g166 (n182, n1);
buf  g167 (n218, n16);
not  g168 (n104, n13);
buf  g169 (n53, n15);
buf  g170 (n71, n7);
buf  g171 (n212, n37);
buf  g172 (n78, n3);
not  g173 (n178, n28);
not  g174 (n68, n12);
not  g175 (n160, n44);
buf  g176 (n50, n26);
not  g177 (n93, n34);
not  g178 (n134, n29);
not  g179 (n119, n43);
buf  g180 (n840, n137);
buf  g181 (n472, n68);
not  g182 (n349, n204);
not  g183 (n606, n50);
buf  g184 (n592, n203);
buf  g185 (n789, n148);
not  g186 (n231, n104);
buf  g187 (n395, n197);
not  g188 (n608, n211);
buf  g189 (n504, n168);
buf  g190 (n794, n112);
not  g191 (n392, n187);
not  g192 (n492, n152);
buf  g193 (n800, n201);
buf  g194 (n843, n219);
not  g195 (n748, n149);
buf  g196 (n279, n200);
not  g197 (n583, n153);
buf  g198 (n227, n121);
buf  g199 (n847, n177);
buf  g200 (n473, n143);
not  g201 (n904, n141);
not  g202 (n807, n136);
buf  g203 (n348, n156);
not  g204 (n620, n154);
buf  g205 (n300, n177);
buf  g206 (n921, n46);
buf  g207 (n574, n188);
buf  g208 (n350, n114);
not  g209 (n468, n143);
not  g210 (n282, n71);
not  g211 (n604, n92);
not  g212 (n917, n188);
not  g213 (n378, n194);
buf  g214 (n865, n189);
buf  g215 (n314, n112);
not  g216 (n514, n148);
not  g217 (n871, n133);
not  g218 (n321, n125);
buf  g219 (n796, n170);
buf  g220 (n544, n63);
buf  g221 (n648, n47);
buf  g222 (n833, n71);
not  g223 (n286, n91);
buf  g224 (n740, n215);
buf  g225 (n403, n78);
buf  g226 (n377, n120);
not  g227 (n554, n135);
buf  g228 (n393, n170);
buf  g229 (n541, n49);
not  g230 (n512, n79);
buf  g231 (n614, n89);
not  g232 (n438, n155);
not  g233 (n238, n100);
buf  g234 (n434, n190);
not  g235 (n640, n73);
buf  g236 (n889, n80);
not  g237 (n535, n166);
buf  g238 (n284, n203);
buf  g239 (n386, n144);
buf  g240 (n230, n82);
not  g241 (n382, n206);
buf  g242 (n240, n159);
not  g243 (n804, n86);
buf  g244 (n405, n149);
buf  g245 (n511, n48);
buf  g246 (n346, n210);
buf  g247 (n490, n146);
buf  g248 (n657, n81);
buf  g249 (n570, n184);
buf  g250 (n723, n163);
buf  g251 (n823, n153);
buf  g252 (n628, n106);
not  g253 (n337, n102);
not  g254 (n884, n158);
not  g255 (n241, n173);
not  g256 (n599, n195);
not  g257 (n582, n110);
not  g258 (n435, n121);
buf  g259 (n869, n161);
not  g260 (n295, n174);
buf  g261 (n462, n56);
not  g262 (n718, n121);
buf  g263 (n777, n49);
not  g264 (n715, n160);
not  g265 (n688, n151);
buf  g266 (n543, n216);
not  g267 (n782, n144);
buf  g268 (n754, n89);
buf  g269 (n360, n50);
buf  g270 (n338, n128);
buf  g271 (n335, n115);
buf  g272 (n870, n55);
not  g273 (n885, n218);
buf  g274 (n256, n117);
not  g275 (n485, n209);
buf  g276 (n562, n212);
buf  g277 (n533, n73);
not  g278 (n581, n76);
buf  g279 (n824, n202);
buf  g280 (n265, n192);
not  g281 (n703, n182);
buf  g282 (n345, n162);
not  g283 (n422, n59);
buf  g284 (n249, n76);
not  g285 (n817, n48);
buf  g286 (n302, n62);
not  g287 (n263, n74);
buf  g288 (n897, n217);
buf  g289 (n426, n46);
not  g290 (n766, n180);
not  g291 (n711, n83);
not  g292 (n523, n78);
buf  g293 (n311, n88);
buf  g294 (n589, n134);
not  g295 (n373, n184);
buf  g296 (n527, n208);
buf  g297 (n397, n193);
buf  g298 (n503, n167);
not  g299 (n465, n179);
not  g300 (n636, n105);
buf  g301 (n459, n134);
buf  g302 (n320, n123);
not  g303 (n344, n72);
not  g304 (n253, n95);
buf  g305 (n494, n213);
buf  g306 (n659, n120);
buf  g307 (n500, n99);
buf  g308 (n361, n47);
buf  g309 (n704, n102);
buf  g310 (n660, n113);
not  g311 (n600, n144);
buf  g312 (n742, n169);
buf  g313 (n552, n56);
not  g314 (n440, n63);
not  g315 (n773, n96);
buf  g316 (n625, n68);
not  g317 (n829, n199);
buf  g318 (n370, n146);
not  g319 (n647, n73);
buf  g320 (n291, n65);
buf  g321 (n612, n124);
buf  g322 (n880, n131);
not  g323 (n588, n161);
buf  g324 (n501, n107);
buf  g325 (n451, n130);
buf  g326 (n668, n108);
not  g327 (n329, n123);
not  g328 (n287, n109);
not  g329 (n285, n124);
not  g330 (n367, n205);
buf  g331 (n911, n201);
not  g332 (n530, n84);
not  g333 (n616, n187);
buf  g334 (n696, n216);
buf  g335 (n683, n69);
not  g336 (n551, n97);
not  g337 (n771, n131);
buf  g338 (n716, n142);
not  g339 (n774, n82);
buf  g340 (n858, n66);
buf  g341 (n483, n115);
not  g342 (n401, n127);
not  g343 (n493, n174);
not  g344 (n601, n199);
not  g345 (n733, n86);
buf  g346 (n729, n191);
buf  g347 (n784, n117);
buf  g348 (n330, n75);
buf  g349 (n860, n147);
buf  g350 (n839, n87);
buf  g351 (n863, n206);
not  g352 (n486, n123);
not  g353 (n596, n137);
buf  g354 (n467, n114);
buf  g355 (n228, n163);
not  g356 (n873, n101);
not  g357 (n255, n71);
buf  g358 (n707, n203);
buf  g359 (n567, n139);
not  g360 (n406, n142);
buf  g361 (n379, n198);
not  g362 (n728, n218);
buf  g363 (n236, n126);
not  g364 (n431, n209);
buf  g365 (n611, n213);
not  g366 (n566, n59);
buf  g367 (n399, n51);
not  g368 (n825, n134);
not  g369 (n832, n122);
buf  g370 (n470, n206);
buf  g371 (n506, n213);
buf  g372 (n540, n110);
buf  g373 (n734, n124);
not  g374 (n271, n57);
buf  g375 (n699, n201);
not  g376 (n430, n70);
not  g377 (n531, n211);
not  g378 (n791, n164);
buf  g379 (n864, n89);
buf  g380 (n257, n94);
not  g381 (n568, n207);
not  g382 (n388, n73);
buf  g383 (n821, n198);
not  g384 (n428, n118);
not  g385 (n595, n99);
not  g386 (n615, n168);
not  g387 (n635, n104);
not  g388 (n779, n55);
not  g389 (n900, n193);
buf  g390 (n914, n91);
not  g391 (n805, n133);
buf  g392 (n327, n214);
buf  g393 (n232, n219);
not  g394 (n664, n132);
buf  g395 (n651, n169);
buf  g396 (n902, n72);
not  g397 (n355, n212);
buf  g398 (n682, n167);
not  g399 (n621, n116);
buf  g400 (n436, n147);
not  g401 (n899, n158);
buf  g402 (n398, n84);
not  g403 (n505, n95);
not  g404 (n515, n101);
buf  g405 (n751, n110);
not  g406 (n895, n111);
buf  g407 (n624, n62);
not  g408 (n532, n70);
buf  g409 (n308, n129);
not  g410 (n809, n136);
buf  g411 (n549, n149);
not  g412 (n250, n76);
not  g413 (n632, n158);
buf  g414 (n433, n194);
buf  g415 (n247, n136);
not  g416 (n358, n105);
not  g417 (n915, n85);
buf  g418 (n266, n61);
buf  g419 (n708, n60);
not  g420 (n819, n129);
buf  g421 (n617, n93);
not  g422 (n852, n93);
buf  g423 (n571, n143);
buf  g424 (n908, n58);
buf  g425 (n686, n86);
buf  g426 (n627, n64);
not  g427 (n781, n135);
not  g428 (n747, n74);
buf  g429 (n815, n196);
not  g430 (n323, n202);
not  g431 (n484, n97);
not  g432 (n861, n203);
not  g433 (n396, n105);
not  g434 (n916, n159);
not  g435 (n736, n58);
not  g436 (n301, n89);
buf  g437 (n797, n207);
not  g438 (n480, n138);
buf  g439 (n679, n91);
buf  g440 (n464, n165);
buf  g441 (n260, n212);
buf  g442 (n529, n46);
buf  g443 (n721, n58);
not  g444 (n315, n188);
not  g445 (n439, n171);
buf  g446 (n363, n167);
buf  g447 (n811, n138);
not  g448 (n559, n156);
buf  g449 (n802, n61);
not  g450 (n394, n126);
buf  g451 (n425, n185);
not  g452 (n639, n128);
buf  g453 (n412, n93);
buf  g454 (n644, n209);
not  g455 (n709, n55);
buf  g456 (n387, n160);
not  g457 (n516, n80);
buf  g458 (n874, n76);
not  g459 (n385, n75);
buf  g460 (n297, n82);
not  g461 (n739, n156);
buf  g462 (n762, n51);
buf  g463 (n761, n206);
not  g464 (n489, n192);
buf  g465 (n691, n134);
not  g466 (n767, n74);
not  g467 (n769, n131);
not  g468 (n591, n162);
buf  g469 (n539, n113);
buf  g470 (n325, n186);
buf  g471 (n429, n186);
buf  g472 (n607, n98);
buf  g473 (n538, n77);
buf  g474 (n558, n150);
not  g475 (n354, n200);
not  g476 (n828, n65);
buf  g477 (n259, n175);
buf  g478 (n481, n111);
buf  g479 (n787, n132);
not  g480 (n509, n166);
not  g481 (n536, n147);
not  g482 (n866, n66);
not  g483 (n375, n84);
not  g484 (n643, n132);
not  g485 (n673, n50);
buf  g486 (n306, n68);
buf  g487 (n463, n122);
not  g488 (n909, n107);
not  g489 (n763, n112);
buf  g490 (n795, n60);
buf  g491 (n482, n130);
buf  g492 (n258, n116);
buf  g493 (n638, n129);
not  g494 (n339, n191);
buf  g495 (n730, n117);
not  g496 (n725, n177);
not  g497 (n898, n182);
not  g498 (n442, n155);
not  g499 (n706, n212);
not  g500 (n546, n141);
buf  g501 (n233, n179);
buf  g502 (n366, n137);
not  g503 (n652, n185);
buf  g504 (n893, n145);
buf  g505 (n423, n88);
not  g506 (n577, n55);
not  g507 (n573, n160);
not  g508 (n333, n172);
not  g509 (n813, n183);
buf  g510 (n666, n127);
not  g511 (n658, n103);
buf  g512 (n328, n217);
not  g513 (n288, n180);
buf  g514 (n522, n59);
buf  g515 (n758, n205);
buf  g516 (n471, n135);
not  g517 (n310, n52);
not  g518 (n383, n124);
not  g519 (n765, n195);
not  g520 (n835, n54);
buf  g521 (n694, n145);
not  g522 (n294, n163);
buf  g523 (n910, n211);
buf  g524 (n854, n145);
not  g525 (n879, n139);
not  g526 (n882, n90);
buf  g527 (n684, n200);
not  g528 (n896, n79);
buf  g529 (n603, n63);
not  g530 (n305, n57);
not  g531 (n623, n154);
buf  g532 (n553, n153);
buf  g533 (n520, n181);
buf  g534 (n332, n140);
buf  g535 (n410, n195);
buf  g536 (n365, n220);
not  g537 (n550, n165);
not  g538 (n645, n152);
not  g539 (n322, n133);
buf  g540 (n449, n149);
not  g541 (n919, n80);
not  g542 (n687, n195);
buf  g543 (n510, n157);
buf  g544 (n724, n132);
buf  g545 (n677, n189);
buf  g546 (n418, n140);
not  g547 (n752, n207);
buf  g548 (n799, n164);
not  g549 (n818, n193);
not  g550 (n400, n53);
not  g551 (n356, n155);
not  g552 (n743, n179);
buf  g553 (n404, n150);
buf  g554 (n312, n126);
buf  g555 (n547, n97);
not  g556 (n690, n168);
buf  g557 (n248, n175);
buf  g558 (n786, n199);
buf  g559 (n775, n161);
not  g560 (n534, n72);
buf  g561 (n602, n173);
not  g562 (n669, n127);
not  g563 (n229, n119);
buf  g564 (n409, n66);
not  g565 (n252, n150);
buf  g566 (n697, n192);
not  g567 (n458, n214);
buf  g568 (n918, n48);
not  g569 (n576, n54);
buf  g570 (n411, n50);
buf  g571 (n609, n77);
not  g572 (n655, n77);
not  g573 (n226, n166);
buf  g574 (n572, n62);
buf  g575 (n755, n94);
not  g576 (n319, n87);
buf  g577 (n672, n118);
not  g578 (n556, n104);
buf  g579 (n605, n178);
buf  g580 (n507, n151);
buf  g581 (n816, n96);
buf  g582 (n298, n98);
buf  g583 (n856, n86);
buf  g584 (n764, n144);
not  g585 (n836, n108);
not  g586 (n477, n160);
buf  g587 (n353, n70);
not  g588 (n334, n117);
not  g589 (n318, n130);
not  g590 (n678, n114);
not  g591 (n922, n174);
buf  g592 (n750, n178);
buf  g593 (n590, n183);
not  g594 (n780, n163);
not  g595 (n281, n184);
not  g596 (n712, n182);
buf  g597 (n267, n152);
buf  g598 (n663, n90);
buf  g599 (n331, n204);
buf  g600 (n476, n217);
not  g601 (n519, n53);
buf  g602 (n646, n152);
buf  g603 (n727, n180);
not  g604 (n391, n109);
buf  g605 (n857, n67);
buf  g606 (n675, n93);
not  g607 (n746, n95);
buf  g608 (n569, n99);
buf  g609 (n901, n168);
buf  g610 (n368, n201);
not  g611 (n637, n169);
buf  g612 (n380, n138);
not  g613 (n801, n61);
not  g614 (n749, n126);
not  g615 (n268, n54);
buf  g616 (n710, n159);
not  g617 (n670, n77);
buf  g618 (n649, n92);
not  g619 (n513, n87);
buf  g620 (n737, n135);
buf  g621 (n415, n92);
buf  g622 (n408, n46);
buf  g623 (n487, n141);
not  g624 (n785, n57);
not  g625 (n720, n106);
buf  g626 (n292, n91);
not  g627 (n390, n175);
not  g628 (n845, n62);
buf  g629 (n299, n193);
not  g630 (n537, n170);
buf  g631 (n525, n198);
not  g632 (n565, n164);
not  g633 (n316, n143);
buf  g634 (n894, n176);
buf  g635 (n347, n79);
buf  g636 (n244, n100);
not  g637 (n831, n166);
buf  g638 (n461, n98);
not  g639 (n447, n125);
not  g640 (n705, n64);
buf  g641 (n521, n177);
not  g642 (n665, n157);
not  g643 (n618, n56);
not  g644 (n594, n80);
not  g645 (n875, n85);
not  g646 (n806, n139);
not  g647 (n759, n94);
buf  g648 (n814, n190);
not  g649 (n726, n186);
not  g650 (n579, n176);
not  g651 (n474, n81);
not  g652 (n498, n119);
not  g653 (n876, n122);
buf  g654 (n270, n69);
not  g655 (n352, n184);
buf  g656 (n341, n161);
buf  g657 (n701, n51);
not  g658 (n309, n210);
not  g659 (n905, n142);
not  g660 (n757, n98);
not  g661 (n613, n121);
buf  g662 (n907, n95);
not  g663 (n584, n69);
not  g664 (n437, n150);
not  g665 (n671, n81);
not  g666 (n667, n100);
not  g667 (n783, n64);
not  g668 (n261, n151);
buf  g669 (n585, n140);
not  g670 (n676, n137);
buf  g671 (n488, n164);
buf  g672 (n455, n176);
buf  g673 (n661, n162);
not  g674 (n629, n96);
not  g675 (n402, n182);
buf  g676 (n906, n148);
not  g677 (n272, n172);
not  g678 (n820, n47);
not  g679 (n242, n70);
buf  g680 (n826, n174);
buf  g681 (n846, n88);
not  g682 (n851, n158);
not  g683 (n626, n178);
not  g684 (n741, n217);
buf  g685 (n853, n189);
buf  g686 (n810, n178);
buf  g687 (n364, n210);
not  g688 (n848, n66);
not  g689 (n307, n194);
buf  g690 (n444, n87);
not  g691 (n456, n82);
not  g692 (n280, n47);
buf  g693 (n838, n65);
not  g694 (n745, n111);
buf  g695 (n891, n109);
not  g696 (n384, n141);
not  g697 (n597, n208);
buf  g698 (n424, n53);
buf  g699 (n633, n94);
buf  g700 (n460, n202);
buf  g701 (n803, n92);
not  g702 (n689, n138);
not  g703 (n580, n190);
not  g704 (n417, n114);
buf  g705 (n867, n67);
buf  g706 (n413, n74);
not  g707 (n262, n171);
buf  g708 (n381, n53);
not  g709 (n475, n171);
buf  g710 (n738, n219);
not  g711 (n912, n204);
buf  g712 (n274, n68);
not  g713 (n296, n196);
buf  g714 (n685, n103);
not  g715 (n662, n147);
not  g716 (n888, n99);
not  g717 (n878, n156);
not  g718 (n371, n60);
not  g719 (n681, n102);
not  g720 (n732, n84);
not  g721 (n561, n197);
buf  g722 (n788, n90);
not  g723 (n598, n108);
buf  g724 (n479, n128);
buf  g725 (n326, n170);
not  g726 (n849, n145);
not  g727 (n692, n106);
not  g728 (n454, n120);
buf  g729 (n304, n172);
buf  g730 (n407, n49);
buf  g731 (n357, n185);
not  g732 (n822, n112);
not  g733 (n830, n96);
not  g734 (n842, n113);
not  g735 (n778, n208);
not  g736 (n441, n165);
not  g737 (n641, n162);
not  g738 (n837, n108);
buf  g739 (n693, n60);
not  g740 (n243, n122);
not  g741 (n448, n197);
buf  g742 (n526, n107);
buf  g743 (n563, n190);
not  g744 (n450, n214);
buf  g745 (n508, n209);
not  g746 (n290, n115);
not  g747 (n744, n67);
buf  g748 (n278, n169);
not  g749 (n827, n215);
buf  g750 (n275, n85);
buf  g751 (n887, n88);
not  g752 (n427, n180);
not  g753 (n445, n207);
buf  g754 (n443, n198);
buf  g755 (n735, n159);
not  g756 (n575, n52);
not  g757 (n234, n139);
not  g758 (n478, n188);
not  g759 (n560, n148);
buf  g760 (n698, n181);
not  g761 (n722, n194);
not  g762 (n517, n83);
not  g763 (n920, n183);
buf  g764 (n619, n140);
not  g765 (n756, n102);
not  g766 (n702, n127);
not  g767 (n622, n58);
not  g768 (n303, n179);
buf  g769 (n313, n118);
buf  g770 (n528, n101);
buf  g771 (n868, n51);
not  g772 (n245, n125);
buf  g773 (n420, n211);
not  g774 (n890, n113);
buf  g775 (n772, n205);
buf  g776 (n695, n205);
not  g777 (n656, n56);
not  g778 (n254, n204);
not  g779 (n336, n115);
buf  g780 (n872, n75);
buf  g781 (n239, n101);
not  g782 (n631, n106);
buf  g783 (n389, n157);
not  g784 (n768, n103);
buf  g785 (n419, n83);
buf  g786 (n630, n61);
buf  g787 (n235, n129);
buf  g788 (n793, n78);
buf  g789 (n653, n185);
not  g790 (n834, n200);
buf  g791 (n545, n119);
not  g792 (n883, n167);
not  g793 (n502, n192);
not  g794 (n555, n154);
not  g795 (n251, n107);
buf  g796 (n859, n154);
buf  g797 (n844, n49);
not  g798 (n277, n171);
buf  g799 (n416, n75);
not  g800 (n369, n146);
not  g801 (n753, n202);
not  g802 (n642, n213);
buf  g803 (n650, n48);
buf  g804 (n457, n172);
buf  g805 (n432, n146);
not  g806 (n542, n176);
not  g807 (n491, n119);
not  g808 (n414, n72);
buf  g809 (n564, n81);
not  g810 (n892, n215);
buf  g811 (n446, n175);
not  g812 (n452, n173);
buf  g813 (n237, n83);
not  g814 (n792, n109);
not  g815 (n674, n52);
not  g816 (n317, n183);
not  g817 (n841, n216);
not  g818 (n578, n64);
buf  g819 (n700, n215);
buf  g820 (n343, n52);
not  g821 (n770, n186);
not  g822 (n850, n218);
buf  g823 (n886, n125);
buf  g824 (n760, n128);
not  g825 (n790, n104);
buf  g826 (n812, n191);
not  g827 (n557, n67);
buf  g828 (n877, n208);
not  g829 (n264, n54);
buf  g830 (n374, n116);
buf  g831 (n283, n123);
not  g832 (n340, n90);
buf  g833 (n289, n63);
not  g834 (n469, n130);
not  g835 (n499, n151);
buf  g836 (n497, n71);
not  g837 (n610, n79);
buf  g838 (n776, n199);
not  g839 (n714, n187);
buf  g840 (n713, n116);
buf  g841 (n362, n181);
buf  g842 (n495, n216);
buf  g843 (n862, n85);
buf  g844 (n881, n133);
not  g845 (n808, n97);
buf  g846 (n453, n78);
buf  g847 (n246, n218);
not  g848 (n359, n197);
not  g849 (n276, n187);
not  g850 (n376, n105);
not  g851 (n903, n57);
buf  g852 (n587, n65);
not  g853 (n798, n100);
not  g854 (n548, n103);
not  g855 (n342, n111);
not  g856 (n731, n191);
buf  g857 (n351, n189);
buf  g858 (n855, n155);
buf  g859 (n324, n120);
not  g860 (n421, n181);
not  g861 (n913, n196);
not  g862 (n273, n59);
not  g863 (n466, n136);
not  g864 (n654, n214);
buf  g865 (n496, n157);
not  g866 (n269, n142);
not  g867 (n593, n210);
buf  g868 (n634, n118);
buf  g869 (n680, n69);
not  g870 (n719, n219);
buf  g871 (n293, n165);
not  g872 (n372, n173);
buf  g873 (n717, n131);
not  g874 (n524, n196);
buf  g875 (n518, n110);
not  g876 (n586, n153);
nor  g877 (n1133, n772, n403, n822, n422);
xnor g878 (n1206, n773, n390, n587, n868);
nor  g879 (n1225, n823, n584, n566, n871);
nand g880 (n1319, n373, n594, n262, n277);
nor  g881 (n925, n608, n639, n439, n579);
xor  g882 (n953, n723, n833, n706, n514);
xor  g883 (n1570, n369, n794, n635, n558);
xnor g884 (n1164, n809, n429, n765, n751);
nor  g885 (n941, n559, n441, n403, n440);
xnor g886 (n1350, n601, n878, n589, n403);
xnor g887 (n1349, n750, n577, n265, n664);
nand g888 (n1389, n639, n879, n847, n780);
nand g889 (n1260, n862, n640, n425, n716);
or   g890 (n1101, n452, n729, n445, n249);
or   g891 (n1420, n380, n448, n753, n557);
nor  g892 (n1191, n377, n549, n416, n840);
xnor g893 (n1279, n664, n454, n897, n529);
and  g894 (n1185, n578, n368, n855, n676);
nand g895 (n1076, n691, n853, n659, n643);
and  g896 (n1126, n449, n561, n345, n522);
xnor g897 (n1140, n264, n394, n429, n717);
nor  g898 (n1243, n600, n386, n435, n676);
or   g899 (n1504, n257, n853, n819, n792);
or   g900 (n1034, n792, n334, n921, n447);
xnor g901 (n1202, n235, n331, n680, n312);
nand g902 (n1304, n794, n369, n366, n799);
and  g903 (n960, n566, n311, n705, n899);
or   g904 (n1158, n648, n601, n329, n513);
xnor g905 (n1410, n817, n391, n908, n546);
xnor g906 (n1521, n641, n898, n873, n575);
nand g907 (n1314, n414, n413, n799, n457);
xnor g908 (n1439, n835, n825, n631, n327);
and  g909 (n1517, n816, n338, n748, n806);
nor  g910 (n1259, n838, n418, n872, n564);
xnor g911 (n1174, n576, n635, n708, n881);
nand g912 (n1338, n526, n813, n468, n804);
nor  g913 (n1151, n685, n536, n548, n280);
and  g914 (n1490, n358, n862, n661, n323);
or   g915 (n1532, n777, n422, n910, n314);
nand g916 (n974, n681, n256, n362, n903);
xnor g917 (n1115, n393, n385, n630, n833);
and  g918 (n1452, n889, n527, n496, n550);
xnor g919 (n1458, n834, n394, n343, n640);
xor  g920 (n1138, n252, n461, n381, n350);
nor  g921 (n1003, n918, n280, n754, n857);
and  g922 (n1057, n739, n488, n307, n399);
xnor g923 (n1274, n544, n388, n597, n759);
and  g924 (n954, n677, n593, n478, n344);
xnor g925 (n1406, n281, n747, n233, n330);
nor  g926 (n1568, n741, n574, n917, n748);
xnor g927 (n988, n299, n269, n666, n582);
xor  g928 (n1316, n410, n513, n229, n869);
nand g929 (n1413, n733, n746, n285, n699);
and  g930 (n1566, n740, n636, n668, n317);
xnor g931 (n1296, n392, n730, n329, n423);
or   g932 (n1007, n421, n374, n645, n408);
or   g933 (n977, n389, n650, n862, n849);
nor  g934 (n1105, n518, n818, n772, n492);
nand g935 (n1228, n468, n834, n432, n614);
xor  g936 (n1137, n637, n297, n600, n620);
and  g937 (n1496, n359, n539, n878, n412);
and  g938 (n1263, n774, n497, n516, n891);
xor  g939 (n1080, n846, n693, n831, n303);
or   g940 (n1553, n282, n397, n235, n548);
and  g941 (n950, n747, n845, n341, n752);
or   g942 (n1367, n518, n345, n811, n797);
or   g943 (n1069, n250, n605, n412, n228);
xor  g944 (n942, n526, n587, n240, n546);
and  g945 (n1294, n631, n841, n855, n884);
xor  g946 (n1336, n578, n731, n734, n883);
xnor g947 (n1574, n315, n827, n735, n854);
xnor g948 (n1363, n646, n871, n874, n906);
or   g949 (n1044, n487, n864, n506, n858);
xnor g950 (n1108, n854, n699, n876, n627);
xor  g951 (n1386, n688, n378, n613, n798);
and  g952 (n1214, n737, n474, n610, n467);
xnor g953 (n1258, n598, n479, n845, n914);
xor  g954 (n1128, n285, n776, n300, n485);
xor  g955 (n1447, n376, n560, n693, n333);
nor  g956 (n1313, n431, n734, n312, n362);
or   g957 (n982, n553, n491, n696, n236);
nor  g958 (n1280, n606, n790, n358, n289);
xor  g959 (n1453, n828, n272, n510, n551);
and  g960 (n1004, n642, n332, n520, n456);
and  g961 (n1329, n326, n802, n436, n899);
nand g962 (n975, n491, n426, n379, n628);
or   g963 (n952, n774, n718, n650, n712);
and  g964 (n1300, n827, n287, n666, n366);
xor  g965 (n1515, n860, n464, n655, n789);
xnor g966 (n1396, n646, n529, n244, n571);
xor  g967 (n1530, n298, n784, n455, n500);
and  g968 (n978, n306, n550, n821, n421);
nand g969 (n1110, n728, n787, n920, n591);
or   g970 (n1213, n416, n611, n702, n695);
nand g971 (n1184, n481, n591, n726, n868);
xnor g972 (n1006, n886, n451, n466, n759);
xnor g973 (n1579, n702, n411, n542, n798);
or   g974 (n1591, n392, n715, n796, n735);
xnor g975 (n973, n812, n358, n301, n526);
or   g976 (n1265, n556, n604, n850, n245);
xnor g977 (n1539, n351, n719, n315, n390);
xnor g978 (n1157, n414, n771, n691, n570);
and  g979 (n1286, n372, n604, n255, n712);
nand g980 (n1463, n897, n365, n427, n423);
or   g981 (n1502, n810, n393, n915, n396);
nor  g982 (n957, n801, n419, n494, n339);
or   g983 (n1564, n708, n739, n354, n897);
nor  g984 (n1156, n850, n378, n751, n704);
xnor g985 (n943, n670, n409, n347, n624);
nor  g986 (n1012, n431, n750, n639, n449);
xor  g987 (n1017, n438, n682, n589, n263);
xor  g988 (n985, n356, n626, n590, n404);
and  g989 (n1493, n838, n304, n802, n267);
and  g990 (n1498, n547, n708, n518, n306);
nand g991 (n1198, n418, n278, n562, n848);
nand g992 (n1374, n556, n756, n833, n460);
xor  g993 (n1008, n554, n485, n265, n748);
nand g994 (n1475, n655, n438, n844, n906);
xor  g995 (n1380, n243, n612, n355, n853);
nand g996 (n1289, n463, n584, n402, n568);
nand g997 (n939, n481, n814, n554, n673);
or   g998 (n1216, n657, n375, n868, n311);
xor  g999 (n999, n833, n866, n798, n600);
and  g1000 (n1510, n453, n243, n308, n547);
nor  g1001 (n1347, n555, n279, n913, n765);
or   g1002 (n1464, n309, n851, n686, n293);
xor  g1003 (n1045, n489, n262, n226, n296);
nor  g1004 (n1175, n880, n435, n611, n780);
nand g1005 (n962, n654, n556, n613, n860);
or   g1006 (n1064, n744, n764, n460, n911);
nor  g1007 (n1376, n846, n826, n675, n832);
and  g1008 (n1436, n584, n913, n308, n660);
xnor g1009 (n1288, n326, n784, n510, n720);
or   g1010 (n1520, n873, n807, n569, n539);
and  g1011 (n1311, n463, n576, n486, n643);
xor  g1012 (n1168, n396, n688, n500, n407);
nand g1013 (n1241, n621, n835, n365, n768);
xor  g1014 (n1283, n239, n896, n288, n326);
xnor g1015 (n1409, n760, n345, n344, n899);
nand g1016 (n1028, n482, n745, n643, n435);
nand g1017 (n1205, n631, n499, n400, n813);
nand g1018 (n1232, n438, n504, n580, n843);
nor  g1019 (n1527, n770, n774, n888, n726);
xnor g1020 (n1195, n476, n333, n648, n778);
nor  g1021 (n1589, n891, n314, n304, n581);
or   g1022 (n967, n419, n588, n331, n595);
and  g1023 (n955, n852, n773, n592, n263);
xnor g1024 (n1199, n479, n361, n364, n596);
xor  g1025 (n1122, n279, n783, n302, n448);
xnor g1026 (n1524, n783, n530, n477, n307);
xnor g1027 (n1285, n554, n375, n832, n527);
xor  g1028 (n986, n714, n468, n320, n623);
or   g1029 (n1472, n238, n352, n738, n690);
or   g1030 (n1114, n391, n482, n592, n862);
or   g1031 (n1573, n543, n557, n405, n631);
or   g1032 (n1340, n851, n856, n737, n363);
and  g1033 (n1266, n452, n430, n336, n528);
nor  g1034 (n1441, n739, n698, n567, n815);
nor  g1035 (n931, n350, n900, n773, n294);
xor  g1036 (n1016, n842, n743, n684, n817);
or   g1037 (n1405, n605, n809, n524, n751);
xnor g1038 (n1173, n782, n384, n894, n835);
xor  g1039 (n994, n586, n866, n673, n757);
nor  g1040 (n1081, n831, n791, n770, n237);
xnor g1041 (n1587, n515, n232, n384, n801);
or   g1042 (n1599, n473, n629, n907, n869);
or   g1043 (n1056, n550, n393, n654, n453);
xor  g1044 (n1430, n445, n657, n395, n642);
xnor g1045 (n1427, n277, n850, n540, n888);
xnor g1046 (n1455, n321, n480, n895, n815);
xnor g1047 (n1027, n779, n537, n798, n488);
xnor g1048 (n1144, n727, n266, n533, n763);
or   g1049 (n1495, n260, n359, n264, n680);
xor  g1050 (n1513, n323, n692, n735, n697);
nor  g1051 (n1569, n603, n887, n585, n779);
xor  g1052 (n1501, n786, n837, n629, n816);
xor  g1053 (n1014, n842, n560, n410, n454);
or   g1054 (n1362, n475, n744, n909, n711);
or   g1055 (n1567, n692, n654, n848, n894);
xor  g1056 (n1079, n271, n366, n432, n596);
and  g1057 (n928, n788, n337, n662, n493);
xor  g1058 (n1356, n907, n517, n651, n468);
xnor g1059 (n1369, n313, n834, n744, n317);
and  g1060 (n1167, n702, n585, n772, n275);
or   g1061 (n1196, n539, n825, n534, n253);
or   g1062 (n1107, n258, n332, n400, n714);
and  g1063 (n1431, n730, n409, n267, n680);
xor  g1064 (n1215, n430, n477, n408, n856);
xnor g1065 (n1402, n626, n385, n250, n696);
or   g1066 (n945, n503, n269, n578, n641);
xor  g1067 (n1200, n698, n858, n687, n857);
xor  g1068 (n1378, n765, n713, n480, n775);
and  g1069 (n1366, n749, n544, n335, n443);
xnor g1070 (n1090, n349, n303, n288, n310);
and  g1071 (n1013, n337, n521, n372);
xor  g1072 (n1118, n465, n837, n359, n786);
xnor g1073 (n1522, n390, n297, n767, n769);
xor  g1074 (n1476, n628, n607, n373, n562);
nand g1075 (n926, n731, n268, n424, n474);
nor  g1076 (n1075, n407, n460, n645, n609);
nor  g1077 (n1019, n656, n902, n671, n889);
nor  g1078 (n1234, n650, n405, n467, n599);
nor  g1079 (n1166, n261, n470, n723, n844);
nor  g1080 (n1204, n293, n677, n561, n778);
xor  g1081 (n1507, n390, n227, n695, n235);
nand g1082 (n1091, n265, n762, n572, n555);
xor  g1083 (n1368, n383, n305, n531, n890);
nand g1084 (n969, n523, n254, n377, n366);
xnor g1085 (n1211, n346, n731, n379, n625);
nand g1086 (n1361, n437, n459, n433, n484);
nand g1087 (n1559, n494, n427, n255, n460);
xor  g1088 (n1141, n447, n271, n693, n580);
nand g1089 (n1395, n382, n822, n871, n351);
xor  g1090 (n1163, n801, n634, n846, n880);
nor  g1091 (n1408, n884, n363, n802, n716);
nor  g1092 (n1322, n820, n916, n318, n391);
xor  g1093 (n1400, n542, n397, n768, n330);
and  g1094 (n1254, n675, n767, n290, n313);
nand g1095 (n1305, n609, n256, n667, n872);
xnor g1096 (n1565, n420, n774, n668, n401);
nand g1097 (n1015, n375, n722, n273, n692);
nand g1098 (n1301, n764, n890, n487, n605);
xor  g1099 (n1330, n493, n795, n713, n727);
nand g1100 (n1276, n417, n519, n507, n404);
xor  g1101 (n976, n337, n289, n686, n902);
nor  g1102 (n1433, n790, n720, n783, n658);
and  g1103 (n1106, n694, n753, n229, n661);
xnor g1104 (n1327, n610, n381, n704, n589);
nor  g1105 (n1482, n464, n565, n487, n302);
xnor g1106 (n1451, n462, n480, n768, n694);
xnor g1107 (n1207, n702, n353, n671, n803);
xor  g1108 (n1295, n618, n277, n399, n387);
xnor g1109 (n951, n551, n636, n633, n892);
and  g1110 (n1542, n339, n467, n720, n670);
xor  g1111 (n996, n426, n764, n258, n483);
xnor g1112 (n1360, n377, n657, n861, n571);
nand g1113 (n1180, n906, n674, n733, n339);
nor  g1114 (n1082, n551, n333, n867, n908);
xnor g1115 (n1201, n525, n888, n891, n315);
or   g1116 (n1217, n652, n517, n808, n788);
xnor g1117 (n1468, n427, n613, n737, n881);
xnor g1118 (n1548, n692, n770, n698, n450);
xnor g1119 (n1018, n544, n383, n749, n797);
xor  g1120 (n1197, n545, n409, n852, n709);
xnor g1121 (n1514, n852, n227, n482, n333);
xnor g1122 (n1268, n425, n635, n577, n325);
and  g1123 (n1237, n413, n776, n649, n698);
nor  g1124 (n1424, n767, n360, n247, n750);
xor  g1125 (n1519, n795, n591, n456, n746);
nand g1126 (n1139, n705, n893, n437, n821);
nand g1127 (n940, n457, n590, n898, n719);
nor  g1128 (n1323, n771, n296, n575, n856);
and  g1129 (n1040, n818, n863, n421, n533);
nor  g1130 (n972, n527, n790, n407, n272);
and  g1131 (n1425, n563, n760, n559, n327);
nor  g1132 (n938, n886, n839, n303, n498);
xor  g1133 (n948, n632, n568, n861, n890);
or   g1134 (n1357, n657, n679, n629, n733);
xor  g1135 (n944, n473, n588, n540, n452);
or   g1136 (n1443, n378, n714, n335, n857);
nand g1137 (n1052, n436, n682, n420, n367);
xor  g1138 (n1421, n914, n829, n421, n689);
or   g1139 (n1518, n532, n529, n309, n653);
or   g1140 (n1426, n824, n597, n662, n295);
or   g1141 (n1331, n496, n490, n890, n625);
nor  g1142 (n1562, n420, n253, n340, n370);
xnor g1143 (n1392, n393, n797, n419, n841);
nand g1144 (n1104, n885, n814, n248, n257);
xor  g1145 (n1030, n458, n429, n912, n623);
or   g1146 (n1147, n525, n474, n870, n775);
nand g1147 (n1454, n344, n820, n566, n661);
and  g1148 (n1024, n470, n573, n658, n731);
nand g1149 (n1146, n847, n741, n562, n616);
xnor g1150 (n1572, n595, n270, n552, n519);
xnor g1151 (n1481, n451, n381, n810, n717);
nand g1152 (n1236, n357, n603, n418, n596);
xor  g1153 (n1494, n767, n442, n761, n677);
xnor g1154 (n1470, n347, n764, n513, n601);
nand g1155 (n1066, n617, n349, n328, n307);
nand g1156 (n1130, n236, n598, n662, n573);
xnor g1157 (n1242, n858, n747, n824, n918);
xnor g1158 (n924, n800, n251, n380, n472);
xor  g1159 (n1328, n360, n541, n781, n533);
or   g1160 (n1538, n814, n344, n493, n370);
xor  g1161 (n1063, n340, n637, n529, n495);
xor  g1162 (n1089, n458, n832, n350, n638);
xor  g1163 (n1315, n432, n646, n401, n875);
xnor g1164 (n1172, n240, n825, n354, n282);
or   g1165 (n1483, n608, n683, n388, n700);
and  g1166 (n1193, n444, n536, n581, n465);
xnor g1167 (n1480, n289, n436, n507, n898);
xnor g1168 (n1125, n780, n242, n323, n428);
and  g1169 (n1512, n315, n470, n238, n622);
and  g1170 (n1046, n870, n609, n666, n907);
nor  g1171 (n1165, n442, n697, n392, n547);
or   g1172 (n1177, n361, n477, n651, n831);
and  g1173 (n1437, n573, n245, n644, n359);
xnor g1174 (n1403, n266, n905, n396, n664);
or   g1175 (n1473, n802, n497, n409, n595);
and  g1176 (n1229, n490, n917, n483, n555);
or   g1177 (n1337, n577, n226, n524, n254);
nor  g1178 (n1282, n669, n276, n244, n455);
xnor g1179 (n1062, n614, n382, n811, n894);
nand g1180 (n1287, n405, n589, n371, n512);
xnor g1181 (n1050, n247, n865, n867, n278);
xnor g1182 (n1404, n680, n541, n412, n535);
or   g1183 (n958, n775, n903, n911, n348);
nor  g1184 (n1256, n508, n763, n534, n426);
nand g1185 (n1529, n368, n336, n443, n459);
nor  g1186 (n1585, n919, n514, n415, n786);
or   g1187 (n1245, n813, n776, n395, n717);
nor  g1188 (n1597, n545, n518, n778, n406);
nand g1189 (n1541, n602, n848, n454, n632);
nand g1190 (n1278, n865, n627, n877, n678);
nor  g1191 (n934, n807, n757, n578, n387);
xor  g1192 (n964, n325, n548, n249, n679);
or   g1193 (n1466, n358, n346, n586, n822);
xor  g1194 (n1461, n353, n624, n832, n782);
xnor g1195 (n1555, n523, n864, n351, n647);
xnor g1196 (n1379, n771, n808, n515, n879);
nand g1197 (n1264, n252, n424, n311, n910);
nand g1198 (n1575, n712, n617, n439, n559);
or   g1199 (n1485, n836, n380, n484, n246);
or   g1200 (n1095, n898, n785, n525, n678);
and  g1201 (n1041, n441, n328, n914, n427);
xor  g1202 (n965, n464, n621, n757, n454);
or   g1203 (n992, n282, n456, n311, n706);
or   g1204 (n1230, n872, n404, n592, n511);
xnor g1205 (n1124, n755, n728, n295, n827);
or   g1206 (n1043, n442, n856, n528, n437);
nor  g1207 (n1239, n303, n543, n388, n618);
nand g1208 (n923, n234, n455, n640, n686);
xor  g1209 (n1194, n566, n343, n387, n896);
xor  g1210 (n1382, n714, n326, n398, n548);
nor  g1211 (n1536, n472, n583, n769, n753);
nor  g1212 (n1065, n625, n374, n233, n868);
nand g1213 (n1446, n309, n614, n322, n904);
nand g1214 (n1377, n557, n865, n352, n555);
and  g1215 (n1032, n716, n242, n503, n504);
and  g1216 (n1000, n875, n673, n641, n256);
and  g1217 (n1556, n261, n905, n451, n722);
xnor g1218 (n1142, n404, n506, n915, n707);
or   g1219 (n1332, n885, n406, n463, n553);
or   g1220 (n1321, n916, n732, n583, n649);
or   g1221 (n1250, n264, n318, n512, n516);
and  g1222 (n1253, n626, n251, n472, n398);
and  g1223 (n1035, n886, n645, n374, n859);
or   g1224 (n1031, n292, n807, n576, n894);
nand g1225 (n1523, n552, n588, n505, n659);
nand g1226 (n935, n493, n632, n634, n531);
xor  g1227 (n1364, n785, n509, n661, n319);
nand g1228 (n1341, n815, n686, n330, n825);
nor  g1229 (n1393, n301, n730, n701, n230);
nand g1230 (n1093, n820, n604, n462, n710);
nand g1231 (n1534, n844, n425, n652, n726);
xor  g1232 (n1134, n815, n527, n352, n287);
xor  g1233 (n1419, n349, n546, n234, n732);
xor  g1234 (n1129, n389, n819, n459, n792);
nand g1235 (n1171, n501, n738, n594, n579);
nor  g1236 (n1025, n643, n467, n800, n367);
xor  g1237 (n959, n494, n363, n550, n313);
xor  g1238 (n1552, n367, n490, n667, n564);
or   g1239 (n1576, n260, n809, n732, n874);
xnor g1240 (n1415, n376, n696, n305, n360);
xnor g1241 (n1486, n648, n787, n283, n415);
nand g1242 (n1203, n476, n386, n318, n777);
xor  g1243 (n1371, n884, n563, n912, n510);
xor  g1244 (n1235, n797, n469, n523, n722);
nor  g1245 (n1398, n919, n704, n855, n461);
nand g1246 (n1083, n339, n628, n299, n739);
nor  g1247 (n1391, n701, n455, n615, n374);
or   g1248 (n1223, n851, n549, n447, n479);
nand g1249 (n993, n706, n725, n766, n695);
xnor g1250 (n1212, n538, n877, n665, n519);
nor  g1251 (n1102, n663, n839, n249, n905);
or   g1252 (n981, n766, n274, n515, n288);
xnor g1253 (n1487, n783, n546, n620, n337);
nand g1254 (n1290, n666, n660, n231, n674);
nand g1255 (n1560, n495, n237, n875, n787);
nand g1256 (n1159, n500, n408, n639, n679);
xor  g1257 (n1150, n694, n689, n837, n655);
or   g1258 (n984, n490, n465, n813, n446);
and  g1259 (n1267, n414, n747, n400, n823);
xor  g1260 (n1477, n247, n754, n876, n544);
or   g1261 (n1072, n593, n864, n294, n439);
nor  g1262 (n1503, n402, n443, n902, n227);
nand g1263 (n1297, n568, n672, n828, n273);
xnor g1264 (n1500, n391, n512, n508, n304);
xor  g1265 (n1318, n859, n538, n394, n438);
nand g1266 (n1417, n317, n703, n538, n840);
or   g1267 (n1220, n452, n602, n532, n704);
xor  g1268 (n987, n793, n560, n703, n240);
nand g1269 (n1343, n457, n514, n866, n399);
xor  g1270 (n1038, n796, n556, n376, n519);
xor  g1271 (n946, n361, n448, n461, n823);
or   g1272 (n1578, n586, n745, n497, n756);
and  g1273 (n1160, n615, n761, n545, n824);
and  g1274 (n1149, n633, n443, n325, n693);
nand g1275 (n983, n520, n572, n892, n624);
and  g1276 (n1580, n371, n424, n638, n267);
nor  g1277 (n1275, n508, n710, n232, n649);
and  g1278 (n949, n794, n826, n780, n399);
nand g1279 (n1231, n801, n869, n811, n847);
xor  g1280 (n1308, n572, n756, n588, n501);
or   g1281 (n1143, n516, n242, n567, n701);
and  g1282 (n1255, n724, n688, n316, n507);
nor  g1283 (n1096, n920, n722, n611, n473);
and  g1284 (n1291, n649, n541, n330, n340);
or   g1285 (n1469, n370, n481, n346, n286);
xnor g1286 (n1059, n575, n335, n711, n919);
xnor g1287 (n1489, n632, n880, n322, n274);
xor  g1288 (n1186, n428, n834, n891, n279);
or   g1289 (n1387, n599, n745, n233, n671);
nand g1290 (n1348, n483, n317, n524, n830);
and  g1291 (n1136, n478, n430, n370, n342);
nand g1292 (n1112, n551, n343, n746, n481);
or   g1293 (n1592, n257, n499, n742, n314);
xnor g1294 (n1563, n842, n314, n284, n386);
nor  g1295 (n1246, n231, n362, n750, n610);
or   g1296 (n1414, n607, n373, n601, n759);
xnor g1297 (n1375, n626, n847, n530, n689);
or   g1298 (n1333, n464, n607, n587, n270);
nand g1299 (n1492, n717, n583, n501, n444);
or   g1300 (n1435, n660, n725, n604, n807);
nand g1301 (n1550, n281, n789, n724, n322);
xor  g1302 (n1384, n630, n752, n536, n697);
xnor g1303 (n991, n432, n498, n619, n700);
xnor g1304 (n1219, n849, n479, n319, n417);
xor  g1305 (n1586, n428, n565, n620, n699);
nor  g1306 (n1434, n684, n425, n896, n590);
or   g1307 (n1346, n355, n678, n280, n580);
nand g1308 (n1067, n695, n332, n408, n553);
and  g1309 (n1103, n721, n854, n496, n765);
or   g1310 (n1178, n412, n321, n484, n893);
nor  g1311 (n1528, n691, n900, n268, n392);
xnor g1312 (n1132, n561, n486, n338, n532);
nand g1313 (n1448, n685, n562, n694, n814);
or   g1314 (n1109, n610, n615, n471, n511);
and  g1315 (n1247, n323, n361, n806, n559);
and  g1316 (n990, n709, n474, n446, n595);
or   g1317 (n1462, n347, n720, n808, n842);
xnor g1318 (n1511, n348, n306, n896, n327);
and  g1319 (n1022, n473, n876, n715, n530);
xnor g1320 (n1182, n276, n741, n592, n640);
and  g1321 (n1508, n655, n729, n599, n517);
and  g1322 (n937, n642, n913, n745, n760);
nand g1323 (n929, n872, n910, n320, n465);
xnor g1324 (n1352, n402, n908, n709, n434);
or   g1325 (n1238, n670, n755, n441, n560);
or   g1326 (n1581, n449, n785, n737, n549);
and  g1327 (n1525, n851, n838, n569, n415);
xor  g1328 (n1001, n341, n434, n383, n489);
nand g1329 (n1183, n554, n499, n841, n902);
or   g1330 (n1261, n919, n684, n740, n696);
nand g1331 (n1385, n531, n328, n597, n724);
nor  g1332 (n1509, n348, n484, n685, n819);
xnor g1333 (n1119, n849, n607, n875, n381);
xnor g1334 (n1179, n522, n236, n585, n357);
xor  g1335 (n1499, n376, n517, n312, n573);
xor  g1336 (n1145, n677, n700, n676, n697);
xnor g1337 (n1516, n870, n647, n276, n510);
nor  g1338 (n1222, n884, n895, n488, n662);
or   g1339 (n1335, n582, n705, n830, n380);
xnor g1340 (n1533, n849, n445, n290, n897);
and  g1341 (n1092, n262, n579, n749, n908);
or   g1342 (n1210, n459, n687, n781, n300);
or   g1343 (n1071, n259, n557, n523, n581);
xor  g1344 (n1344, n911, n537, n368, n889);
xnor g1345 (n1317, n498, n761, n881, n827);
and  g1346 (n936, n621, n283, n371, n709);
xnor g1347 (n1051, n316, n669, n539, n357);
nand g1348 (n1423, n248, n445, n791, n886);
xor  g1349 (n1127, n887, n520, n450, n509);
xnor g1350 (n1248, n790, n563, n431, n250);
xor  g1351 (n1557, n413, n663, n652, n230);
and  g1352 (n1342, n341, n629, n570, n622);
and  g1353 (n1596, n887, n345, n885, n781);
or   g1354 (n1068, n543, n823, n804, n564);
xnor g1355 (n1208, n599, n711, n410, n537);
nand g1356 (n1432, n494, n656, n736, n411);
xor  g1357 (n1355, n397, n600, n672, n679);
nand g1358 (n1120, n840, n736, n356, n721);
or   g1359 (n1021, n793, n503, n295, n627);
or   g1360 (n1181, n623, n656, n565, n553);
and  g1361 (n1547, n881, n716, n483, n785);
xor  g1362 (n1026, n726, n734, n804, n340);
and  g1363 (n1445, n622, n861, n398, n713);
xnor g1364 (n1273, n906, n300, n308, n678);
nand g1365 (n1299, n659, n627, n471, n781);
xor  g1366 (n1053, n795, n768, n821, n440);
nand g1367 (n1221, n880, n406, n782, n762);
or   g1368 (n1359, n718, n508, n878, n690);
or   g1369 (n947, n728, n874, n710, n743);
nor  g1370 (n1293, n912, n463, n356, n533);
nor  g1371 (n1411, n763, n637, n444, n918);
xnor g1372 (n1277, n706, n528, n867, n848);
xnor g1373 (n1467, n378, n736, n835, n843);
or   g1374 (n1005, n675, n502, n324, n742);
and  g1375 (n1002, n900, n652, n874, n535);
or   g1376 (n968, n817, n255, n482, n683);
xnor g1377 (n1042, n690, n451, n914, n449);
and  g1378 (n1121, n285, n612, n853, n353);
and  g1379 (n1594, n622, n669, n458, n917);
or   g1380 (n1505, n633, n828, n817, n792);
xnor g1381 (n1192, n324, n234, n290, n812);
nand g1382 (n979, n346, n911, n882, n253);
nor  g1383 (n1353, n630, n434, n839, n826);
or   g1384 (n1465, n761, n625, n302, n805);
nor  g1385 (n1460, n244, n766, n367, n805);
nor  g1386 (n1491, n755, n511, n909, n725);
nand g1387 (n1033, n782, n379, n684, n653);
nand g1388 (n1399, n552, n442, n756, n681);
xnor g1389 (n1551, n754, n751, n521, n354);
nand g1390 (n1354, n612, n355, n771, n338);
and  g1391 (n989, n507, n916, n895, n478);
nor  g1392 (n1049, n855, n444, n241, n673);
xor  g1393 (n1325, n275, n466, n286, n917);
or   g1394 (n1086, n668, n758, n915, n674);
xnor g1395 (n1117, n505, n313, n791, n636);
or   g1396 (n1412, n624, n411, n355, n478);
nor  g1397 (n1269, n394, n270, n701, n302);
nor  g1398 (n1054, n342, n328, n845, n400);
xor  g1399 (n1251, n401, n259, n648, n308);
or   g1400 (n1407, n654, n352, n364, n889);
or   g1401 (n1292, n859, n787, n504, n873);
xnor g1402 (n1154, n384, n324, n758, n575);
xnor g1403 (n998, n741, n837, n660, n912);
xnor g1404 (n1170, n379, n540, n536, n541);
nor  g1405 (n1190, n434, n688, n430, n321);
xor  g1406 (n1153, n749, n307, n246, n612);
xnor g1407 (n1244, n252, n342, n719, n616);
or   g1408 (n1312, n576, n606, n830, n558);
xnor g1409 (n1577, n663, n558, n609, n569);
nand g1410 (n1037, n294, n446, n571, n386);
nand g1411 (n1418, n707, n521, n388, n593);
xor  g1412 (n1543, n647, n871, n893, n237);
xor  g1413 (n1442, n852, n357, n614, n860);
xnor g1414 (n1272, n885, n524, n777, n286);
xnor g1415 (n1488, n799, n356, n485, n301);
nand g1416 (n956, n331, n725, n775, n647);
and  g1417 (n1252, n883, n335, n382, n810);
nor  g1418 (n1582, n525, n332, n343, n563);
or   g1419 (n1011, n638, n271, n816, n788);
xnor g1420 (n1345, n742, n682, n887, n486);
nor  g1421 (n933, n683, n469, n863, n402);
and  g1422 (n1155, n715, n321, n623, n910);
nand g1423 (n1561, n416, n665, n879, n305);
nor  g1424 (n1047, n269, n316, n491, n836);
xor  g1425 (n1152, n411, n719, n920, n877);
xor  g1426 (n1077, n363, n804, n260, n755);
xor  g1427 (n1084, n254, n401, n322, n509);
and  g1428 (n1401, n296, n457, n786, n805);
xnor g1429 (n930, n407, n733, n879, n266);
or   g1430 (n1372, n596, n691, n707, n232);
xnor g1431 (n1394, n634, n389, n779, n450);
nand g1432 (n1303, n883, n867, n740, n651);
nand g1433 (n1373, n424, n687, n535, n384);
xnor g1434 (n1023, n570, n530, n732, n667);
xnor g1435 (n1249, n414, n239, n758, n448);
xor  g1436 (n1471, n921, n420, n496, n700);
xor  g1437 (n1078, n598, n658, n793, n811);
xnor g1438 (n1307, n653, n540, n670, n458);
and  g1439 (n1070, n828, n342, n808, n901);
xor  g1440 (n963, n613, n682, n245, n795);
nand g1441 (n1497, n583, n909, n351, n672);
nor  g1442 (n1061, n579, n621, n744, n466);
xor  g1443 (n1598, n297, n535, n845, n619);
nand g1444 (n1558, n437, n419, n433, n571);
xor  g1445 (n1302, n273, n415, n320, n903);
xnor g1446 (n1240, n574, n882, n863, n705);
nand g1447 (n1326, n743, n534, n489, n226);
or   g1448 (n1365, n594, n762, n721, n841);
and  g1449 (n1429, n372, n806, n513, n776);
or   g1450 (n1058, n708, n299, n687, n466);
xnor g1451 (n1257, n435, n602, n441, n829);
nand g1452 (n1270, n462, n369, n436, n907);
or   g1453 (n1478, n403, n593, n753, n431);
xnor g1454 (n1438, n784, n586, n915, n735);
xnor g1455 (n1450, n268, n805, n800, n505);
nand g1456 (n1531, n334, n752, n681, n757);
nor  g1457 (n961, n665, n844, n587, n729);
or   g1458 (n1100, n495, n423, n564, n901);
nor  g1459 (n1169, n447, n567, n418, n310);
or   g1460 (n1545, n796, n230, n446, n542);
xnor g1461 (n1113, n641, n892, n638, n258);
nor  g1462 (n1116, n921, n405, n397, n456);
nor  g1463 (n1479, n331, n492, n903, n439);
xnor g1464 (n1074, n888, n440, n838, n675);
and  g1465 (n1298, n839, n904, n263, n773);
or   g1466 (n1474, n766, n689, n900, n385);
nand g1467 (n1388, n477, n471, n690, n375);
and  g1468 (n1087, n715, n410, n338, n526);
nor  g1469 (n1595, n642, n324, n685, n728);
xnor g1470 (n1187, n497, n713, n809, n498);
nor  g1471 (n1226, n738, n506, n522, n417);
xor  g1472 (n1584, n514, n292, n608, n453);
xnor g1473 (n1554, n284, n275, n854, n350);
or   g1474 (n1060, n284, n310, n762, n664);
or   g1475 (n1549, n645, n487, n241, n671);
or   g1476 (n1526, n840, n770, n259, n283);
xor  g1477 (n1020, n812, n360, n669, n565);
xor  g1478 (n1449, n348, n429, n469, n681);
xor  g1479 (n1098, n364, n861, n353, n428);
nand g1480 (n1370, n577, n803, n341, n502);
xor  g1481 (n1324, n617, n606, n758, n859);
or   g1482 (n1029, n594, n520, n836, n462);
xnor g1483 (n1227, n893, n538, n336, n615);
nand g1484 (n1131, n711, n383, n676, n822);
or   g1485 (n1537, n305, n826, n869, n651);
and  g1486 (n1281, n779, n882, n318, n723);
xnor g1487 (n1176, n870, n561, n796, n304);
and  g1488 (n1284, n707, n426, n433, n789);
and  g1489 (n997, n469, n567, n818, n734);
xor  g1490 (n1088, n281, n882, n327, n736);
xnor g1491 (n1457, n803, n569, n904, n574);
and  g1492 (n1123, n721, n489, n500, n710);
xnor g1493 (n1544, n398, n243, n537, n417);
nor  g1494 (n1593, n552, n389, n531, n319);
xnor g1495 (n995, n810, n369, n619, n831);
xnor g1496 (n1309, n347, n665, n913, n416);
nand g1497 (n971, n475, n528, n433, n829);
or   g1498 (n1097, n476, n581, n387, n636);
xor  g1499 (n1233, n395, n818, n836, n287);
nand g1500 (n1036, n608, n864, n572, n568);
or   g1501 (n927, n850, n395, n248, n703);
and  g1502 (n1188, n784, n821, n278, n373);
nor  g1503 (n1540, n336, n858, n909, n450);
and  g1504 (n932, n512, n503, n616, n521);
xor  g1505 (n1334, n637, n824, n603, n547);
xnor g1506 (n1135, n740, n522, n634, n320);
nand g1507 (n1189, n746, n778, n334, n863);
xnor g1508 (n1162, n611, n724, n319, n590);
nor  g1509 (n1048, n803, n309, n515, n727);
xnor g1510 (n1506, n752, n542, n292, n772);
xnor g1511 (n1390, n371, n461, n760, n316);
xor  g1512 (n1320, n674, n899, n901, n422);
nand g1513 (n1010, n843, n738, n423, n570);
xnor g1514 (n1099, n406, n495, n904, n816);
or   g1515 (n1039, n901, n644, n646, n362);
xnor g1516 (n1306, n656, n509, n228, n916);
and  g1517 (n1571, n905, n843, n920, n712);
and  g1518 (n1397, n857, n516, n819, n368);
and  g1519 (n1546, n895, n630, n475, n727);
and  g1520 (n1535, n585, n502, n921, n602);
and  g1521 (n1351, n658, n349, n298, n873);
nor  g1522 (n1094, n598, n667, n511, n860);
nor  g1523 (n1422, n668, n329, n471, n470);
nand g1524 (n970, n603, n272, n618, n699);
nand g1525 (n1381, n800, n584, n789, n382);
nor  g1526 (n1416, n644, n365, n261, n582);
nand g1527 (n1224, n475, n543, n799, n488);
nor  g1528 (n1148, n385, n325, n334, n312);
xnor g1529 (n1161, n545, n246, n759, n534);
xnor g1530 (n1111, n644, n298, n506, n820);
or   g1531 (n1484, n742, n729, n499, n580);
xnor g1532 (n1085, n812, n486, n878, n293);
nand g1533 (n1271, n574, n422, n877, n616);
nor  g1534 (n1262, n618, n883, n396, n653);
or   g1535 (n966, n763, n480, n628, n491);
and  g1536 (n1218, n846, n413, n788, n231);
xor  g1537 (n1358, n472, n876, n769, n606);
nand g1538 (n1583, n663, n591, n791, n377);
nor  g1539 (n1073, n866, n365, n485, n723);
nor  g1540 (n1588, n703, n229, n558, n892);
nand g1541 (n1009, n620, n617, n672, n492);
xnor g1542 (n1459, n291, n794, n806, n306);
xor  g1543 (n1440, n354, n453, n504, n605);
xnor g1544 (n1444, n532, n918, n597, n238);
xnor g1545 (n1428, n829, n239, n440, n329);
or   g1546 (n1456, n650, n865, n718);
and  g1547 (n1339, n274, n730, n291, n476);
nand g1548 (n1209, n635, n492, n251, n683);
xnor g1549 (n980, n501, n505, n582, n619);
xnor g1550 (n1055, n754, n633, n777, n743);
nand g1551 (n1383, n748, n228, n364, n310);
nor  g1552 (n1310, n549, n241, n291, n502);
and  g1553 (n1590, n793, n769, n659, n830);
buf  g1554 (n1614, n944);
not  g1555 (n1615, n947);
buf  g1556 (n1606, n941);
not  g1557 (n1605, n923);
not  g1558 (n1610, n946);
buf  g1559 (n1611, n935);
not  g1560 (n1609, n928);
buf  g1561 (n1619, n939);
not  g1562 (n1608, n929);
not  g1563 (n1617, n925);
buf  g1564 (n1618, n945);
buf  g1565 (n1620, n930);
buf  g1566 (n1607, n950);
not  g1567 (n1601, n948);
or   g1568 (n1604, n936, n932);
xor  g1569 (n1612, n943, n937);
nor  g1570 (n1616, n942, n933);
nand g1571 (n1602, n927, n934);
nor  g1572 (n1603, n926, n938);
xor  g1573 (n1600, n940, n924);
and  g1574 (n1613, n931, n949);
not  g1575 (n1623, n960);
nor  g1576 (n1634, n958, n224, n1601);
and  g1577 (n1627, n965, n225, n222, n224);
xor  g1578 (n1631, n220, n222, n223);
xor  g1579 (n1624, n225, n1600, n1602, n222);
and  g1580 (n1633, n224, n961, n1602, n223);
or   g1581 (n1625, n1601, n221, n1603);
nor  g1582 (n1621, n959, n964, n1600, n962);
nor  g1583 (n1622, n952, n1601, n951, n1602);
nand g1584 (n1629, n1602, n225, n922, n1603);
nor  g1585 (n1632, n225, n954, n957, n922);
or   g1586 (n1626, n220, n1600, n1601, n221);
nand g1587 (n1635, n953, n220, n223, n963);
and  g1588 (n1628, n224, n922, n956, n223);
or   g1589 (n1630, n221, n1600, n955, n1603);
buf  g1590 (n1639, n1623);
buf  g1591 (n1640, n1621);
buf  g1592 (n1646, n1625);
not  g1593 (n1637, n1627);
not  g1594 (n1643, n1629);
buf  g1595 (n1642, n1622);
not  g1596 (n1645, n967);
not  g1597 (n1644, n1628);
not  g1598 (n1638, n1630);
not  g1599 (n1636, n1626);
and  g1600 (n1641, n1631, n966, n1624);
nand g1601 (n1650, n969, n1001, n1009, n973);
nand g1602 (n1661, n1636, n1640, n985, n974);
xnor g1603 (n1647, n979, n999, n984, n1010);
nand g1604 (n1654, n1640, n994, n1637, n1015);
or   g1605 (n1657, n986, n1636, n976, n1003);
xnor g1606 (n1648, n1012, n981, n998, n1638);
and  g1607 (n1656, n988, n1013, n1639, n1638);
or   g1608 (n1658, n972, n980, n1008, n990);
nor  g1609 (n1651, n991, n1014, n1638, n1000);
and  g1610 (n1653, n997, n1639, n992);
xor  g1611 (n1649, n1636, n970, n977, n968);
and  g1612 (n1655, n982, n983, n1007, n1638);
nor  g1613 (n1659, n996, n993, n1006, n975);
xor  g1614 (n1660, n1011, n1637, n978, n971);
nand g1615 (n1652, n1005, n1639, n1002, n987);
or   g1616 (n1662, n1637, n989, n995, n1004);
or   g1617 (n1671, n1604, n1607, n1662, n1653);
xor  g1618 (n1675, n1604, n1606, n1607, n1609);
nor  g1619 (n1670, n1604, n1612, n1655, n1654);
nand g1620 (n1676, n1608, n1614, n1610, n1615);
nand g1621 (n1672, n1611, n1604, n1609, n1613);
and  g1622 (n1677, n1611, n1658, n1657, n1608);
nor  g1623 (n1667, n1603, n1610, n1649, n1612);
or   g1624 (n1665, n1614, n1656, n1606, n1659);
nor  g1625 (n1674, n1605, n1605, n1615, n1606);
nor  g1626 (n1664, n1647, n1615, n1606, n1613);
xor  g1627 (n1669, n1608, n1648, n1612, n1651);
and  g1628 (n1668, n1607, n1605, n1610, n1652);
or   g1629 (n1663, n1611, n1609, n1612, n1661);
and  g1630 (n1673, n1610, n1609, n1613, n1608);
xor  g1631 (n1666, n1660, n1607, n1613, n1650);
nor  g1632 (n1678, n1605, n1614, n1611);
buf  g1633 (n1700, n1671);
not  g1634 (n1689, n1669);
not  g1635 (n1692, n1668);
buf  g1636 (n1701, n1670);
buf  g1637 (n1699, n1671);
not  g1638 (n1698, n1664);
buf  g1639 (n1703, n1664);
buf  g1640 (n1705, n1666);
buf  g1641 (n1691, n1669);
buf  g1642 (n1690, n1672);
not  g1643 (n1710, n1663);
not  g1644 (n1693, n1671);
buf  g1645 (n1685, n1669);
not  g1646 (n1687, n1665);
not  g1647 (n1695, n1663);
not  g1648 (n1679, n1663);
not  g1649 (n1680, n1670);
not  g1650 (n1709, n1667);
not  g1651 (n1686, n1667);
not  g1652 (n1684, n1666);
not  g1653 (n1706, n1673);
not  g1654 (n1681, n1665);
buf  g1655 (n1708, n1667);
buf  g1656 (n1702, n1672);
not  g1657 (n1688, n1664);
buf  g1658 (n1694, n1666);
buf  g1659 (n1683, n1670);
buf  g1660 (n1682, n1668);
not  g1661 (n1697, n1665);
buf  g1662 (n1696, n1672);
buf  g1663 (n1707, n1668);
not  g1664 (n1704, n1672);
buf  g1665 (n1726, n1696);
buf  g1666 (n1772, n1642);
buf  g1667 (n1792, n1644);
buf  g1668 (n1760, n1691);
buf  g1669 (n1790, n1701);
buf  g1670 (n1756, n1702);
buf  g1671 (n1725, n1645);
buf  g1672 (n1745, n1691);
buf  g1673 (n1773, n1645);
buf  g1674 (n1750, n1693);
not  g1675 (n1759, n1705);
buf  g1676 (n1793, n1692);
buf  g1677 (n1783, n1644);
buf  g1678 (n1721, n1681);
not  g1679 (n1786, n1703);
buf  g1680 (n1731, n1698);
not  g1681 (n1719, n1695);
not  g1682 (n1757, n1700);
not  g1683 (n1761, n1709);
buf  g1684 (n1768, n1642);
buf  g1685 (n1749, n1696);
not  g1686 (n1787, n1685);
not  g1687 (n1785, n1646);
buf  g1688 (n1770, n1698);
not  g1689 (n1722, n1694);
buf  g1690 (n1784, n1682);
buf  g1691 (n1724, n1690);
buf  g1692 (n1735, n1690);
not  g1693 (n1734, n1682);
not  g1694 (n1743, n1643);
buf  g1695 (n1776, n1694);
not  g1696 (n1748, n1699);
buf  g1697 (n1752, n1679);
not  g1698 (n1737, n1616);
buf  g1699 (n1712, n1701);
buf  g1700 (n1782, n1709);
not  g1701 (n1716, n1691);
not  g1702 (n1780, n1697);
not  g1703 (n1739, n1700);
not  g1704 (n1718, n1681);
buf  g1705 (n1758, n1685);
buf  g1706 (n1741, n1700);
buf  g1707 (n1764, n1701);
not  g1708 (n1714, n1702);
buf  g1709 (n1729, n1704);
buf  g1710 (n1789, n1680);
buf  g1711 (n1728, n1641);
buf  g1712 (n1747, n1700);
buf  g1713 (n1711, n1645);
buf  g1714 (n1771, n1689);
not  g1715 (n1769, n1689);
buf  g1716 (n1779, n1679);
buf  g1717 (n1713, n1690);
buf  g1718 (n1751, n1619);
buf  g1719 (n1723, n1690);
not  g1720 (n1788, n1618);
buf  g1721 (n1775, n1703);
not  g1722 (n1796, n1619);
and  g1723 (n1777, n1706, n1617);
nor  g1724 (n1738, n1707, n1685, n1646, n1643);
or   g1725 (n1754, n1704, n1705, n1692, n1695);
nand g1726 (n1732, n1705, n1699, n1706, n1681);
or   g1727 (n1744, n1705, n1617, n1707, n1645);
nand g1728 (n1733, n1680, n1689, n1684, n1691);
xor  g1729 (n1715, n1697, n1644, n1616, n1688);
and  g1730 (n1791, n1710, n1642, n1695);
or   g1731 (n1742, n1687, n1699, n1692, n1708);
nor  g1732 (n1766, n1699, n1710, n1631, n1618);
nor  g1733 (n1797, n1708, n1688, n1694, n1703);
nor  g1734 (n1767, n1646, n1683, n1685);
nor  g1735 (n1755, n1679, n1707, n1687, n1642);
nor  g1736 (n1765, n1619, n1697, n1680, n1698);
or   g1737 (n1763, n1693, n1646, n1710, n1686);
and  g1738 (n1753, n1631, n1686, n1703, n1693);
or   g1739 (n1717, n1641, n1643, n1706, n1692);
or   g1740 (n1762, n1684, n1641, n1640, n1686);
and  g1741 (n1795, n1688, n1617, n1679, n1693);
nand g1742 (n1794, n1706, n1708, n1683, n1701);
and  g1743 (n1746, n1688, n1687, n1686, n1680);
xnor g1744 (n1778, n1683, n1709, n1704, n1702);
xnor g1745 (n1727, n1643, n1641, n1644, n1696);
and  g1746 (n1720, n1618, n1694, n1702, n1687);
or   g1747 (n1781, n1681, n1684, n1708, n1640);
nor  g1748 (n1774, n1684, n1617, n1689, n1698);
or   g1749 (n1740, n1616, n1709, n1682, n1704);
nor  g1750 (n1736, n1707, n1615, n1616, n1682);
and  g1751 (n1730, n1697, n1696, n1710, n1618);
nand g1752 (n1811, n1720, n1676, n1674, n1738);
nand g1753 (n1810, n1676, n1675, n1719, n1745);
xnor g1754 (n1800, n1739, n1725, n1751, n1750);
nand g1755 (n1806, n1734, n1752, n1730, n1712);
nand g1756 (n1807, n1718, n1740, n1732, n1713);
xnor g1757 (n1812, n1711, n1744, n1749, n1727);
xnor g1758 (n1801, n1673, n1754, n1676, n1726);
nor  g1759 (n1799, n1674, n1733, n1676, n1741);
xnor g1760 (n1804, n1735, n1674, n1722, n1723);
nor  g1761 (n1803, n1673, n1717, n1746, n1742);
and  g1762 (n1802, n1674, n1743, n1721, n1753);
xor  g1763 (n1798, n1737, n1677, n1715, n1675);
xor  g1764 (n1805, n1714, n1747, n1731, n1748);
xor  g1765 (n1808, n1673, n1736, n1729, n1716);
xnor g1766 (n1809, n1728, n1724, n1675);
buf  g1767 (n1814, n1811);
not  g1768 (n1813, n1812);
xor  g1769 (n1817, n1764, n1765, n1755, n1814);
nand g1770 (n1816, n1759, n1813, n1756, n1814);
or   g1771 (n1815, n1766, n1757, n1758, n1813);
xnor g1772 (n1818, n1761, n1762, n1760, n1763);
xnor g1773 (n1822, n1775, n1777, n1770, n1768);
or   g1774 (n1823, n1818, n1779, n1815, n1774);
xor  g1775 (n1821, n1771, n1778, n1781, n1767);
nand g1776 (n1819, n1769, n1773, n1817, n1772);
and  g1777 (n1820, n1816, n1776, n1780, n1818);
buf  g1778 (n1826, n1821);
and  g1779 (n1824, n1785, n1823, n1822);
nand g1780 (n1825, n1784, n1783, n1782, n1786);
nor  g1781 (n1828, n1019, n1826, n1632, n1023);
nand g1782 (n1829, n1018, n1020, n1021, n1024);
nor  g1783 (n1827, n1825, n1826, n1016, n1025);
or   g1784 (n1830, n1824, n1017, n1022, n1632);
buf  g1785 (n1832, n1829);
nand g1786 (n1831, n1830, n1677);
not  g1787 (n1838, n1026);
buf  g1788 (n1835, n1034);
xor  g1789 (n1834, n1832, n1831, n1030, n1027);
xnor g1790 (n1837, n1831, n1032, n1036, n1029);
nand g1791 (n1833, n1037, n1832, n1033, n1831);
nor  g1792 (n1836, n1028, n1035, n1031, n1832);
not  g1793 (n1840, n1833);
not  g1794 (n1839, n1833);
or   g1795 (n1841, n1788, n1839);
or   g1796 (n1843, n1632, n1633, n1832, n1790);
xor  g1797 (n1842, n922, n1787, n1789, n1633);
buf  g1798 (n1848, n1039);
not  g1799 (n1845, n1040);
buf  g1800 (n1844, n1842);
buf  g1801 (n1846, n1841);
and  g1802 (n1847, n1038, n1843);
xnor g1803 (n1857, n1041, n1042, n1846, n1059);
nand g1804 (n1867, n1619, n1848, n1847);
nand g1805 (n1855, n1065, n1048, n1043, n1047);
and  g1806 (n1856, n1067, n1053, n1070, n1835);
nand g1807 (n1861, n1846, n1071, n1044, n1054);
or   g1808 (n1851, n1063, n1845, n1060, n1833);
or   g1809 (n1852, n1620, n1845, n1072, n1838);
xnor g1810 (n1850, n1834, n1848, n1840, n1064);
xnor g1811 (n1866, n1848, n1846, n1620, n1046);
xor  g1812 (n1862, n1068, n1844, n1837, n1836);
nor  g1813 (n1865, n1633, n1069, n1844, n1839);
xnor g1814 (n1859, n1058, n1838, n1847);
xor  g1815 (n1854, n1844, n1837, n1838);
nor  g1816 (n1853, n1845, n1061, n1837, n1049);
nor  g1817 (n1863, n1835, n1052, n1846, n1045);
xor  g1818 (n1860, n1834, n1840, n1836, n1056);
xor  g1819 (n1868, n1844, n1848, n1050, n1834);
xor  g1820 (n1849, n1057, n1835, n1836, n1062);
xnor g1821 (n1864, n1051, n1845, n1055, n1620);
nor  g1822 (n1858, n1066, n1840, n1847);
xnor g1823 (n1917, n1865, n1287, n1853, n1167);
xor  g1824 (n1923, n1246, n1860, n1267, n1281);
nor  g1825 (n1945, n1185, n1237, n1147, n1234);
or   g1826 (n1934, n1282, n1107, n1213, n1206);
and  g1827 (n1870, n1112, n1244, n1080, n1195);
or   g1828 (n1927, n1224, n1851, n1253, n1235);
or   g1829 (n1948, n1797, n1275, n1143, n1165);
nand g1830 (n1877, n1188, n1852, n1162);
xor  g1831 (n1869, n1859, n1212, n1197, n1860);
and  g1832 (n1889, n1291, n1858, n1113, n1867);
xor  g1833 (n1872, n1867, n1154, n1861, n1228);
nand g1834 (n1935, n1245, n1261, n1179, n1272);
or   g1835 (n1937, n1634, n1221, n1116, n1852);
nor  g1836 (n1926, n1238, n1172, n1229, n1248);
nand g1837 (n1896, n1201, n1163, n1297, n1233);
xnor g1838 (n1908, n1192, n1144, n1867, n1205);
nand g1839 (n1907, n1075, n1137, n1095, n1218);
or   g1840 (n1874, n1858, n1247, n1191, n1157);
xor  g1841 (n1912, n1127, n1260, n1278, n1265);
and  g1842 (n1918, n1635, n1794, n1863, n1219);
xnor g1843 (n1892, n1865, n1187, n1117, n1863);
or   g1844 (n1888, n1217, n1289, n1216, n1857);
xor  g1845 (n1876, n1850, n1128, n1171, n1796);
xor  g1846 (n1911, n1795, n1223, n1274, n1190);
xor  g1847 (n1944, n1276, n1150, n1283, n1124);
or   g1848 (n1883, n1279, n1256, n1176, n1178);
nand g1849 (n1895, n1236, n1864, n1254, n1258);
xnor g1850 (n1879, n1222, n1121, n1868, n1271);
xor  g1851 (n1936, n1851, n1270, n1864, n1853);
and  g1852 (n1897, n1791, n1249, n1277, n1858);
xnor g1853 (n1894, n1139, n1854, n1208, n1156);
nor  g1854 (n1924, n1849, n1856, n1850, n1102);
xnor g1855 (n1928, n1232, n1859, n1635, n1220);
xor  g1856 (n1919, n1136, n1131, n1852, n1298);
xnor g1857 (n1901, n1849, n1135, n1634, n1186);
xor  g1858 (n1943, n1207, n1142, n1120, n1086);
xnor g1859 (n1898, n1074, n1083, n1133, n1182);
xor  g1860 (n1939, n1082, n1097, n1856, n1862);
xnor g1861 (n1932, n1861, n1856, n1194, n1114);
xor  g1862 (n1900, n1169, n1855, n1110, n1861);
nand g1863 (n1906, n1227, n1857, n1160, n1855);
xnor g1864 (n1893, n1854, n1115, n1865, n1868);
nand g1865 (n1929, n1180, n1868, n1175, n1210);
xor  g1866 (n1880, n1090, n1849, n1093, n1105);
nor  g1867 (n1916, n1078, n1199, n1123, n1138);
or   g1868 (n1891, n1145, n1198, n1867, n1184);
xnor g1869 (n1875, n1085, n1108, n1170, n1155);
xnor g1870 (n1871, n1240, n1125, n1141, n1854);
nor  g1871 (n1922, n1087, n1111, n1293, n1865);
xor  g1872 (n1886, n1092, n1262, n1151, n1273);
nand g1873 (n1881, n1864, n1166, n1855, n1268);
xnor g1874 (n1921, n1073, n1204, n1098, n1211);
nand g1875 (n1905, n1252, n1129, n1209, n1295);
nand g1876 (n1933, n1635, n1183, n1242, n1230);
nand g1877 (n1938, n1103, n1851, n1866, n1153);
xnor g1878 (n1890, n1079, n1109, n1161, n1866);
or   g1879 (n1940, n1862, n1084, n1866, n1857);
xor  g1880 (n1913, n1850, n1088, n1859, n1101);
or   g1881 (n1947, n1854, n1286, n1266, n1132);
xnor g1882 (n1931, n1164, n1859, n1231, n1149);
or   g1883 (n1941, n1189, n1241, n1862, n1096);
xnor g1884 (n1878, n1866, n1250, n1104, n1855);
xnor g1885 (n1909, n1094, n1152, n1853, n1243);
and  g1886 (n1914, n1792, n1091, n1264, n1269);
nor  g1887 (n1942, n1119, n1081, n1292, n1076);
nor  g1888 (n1885, n1196, n1106, n1215, n1290);
xnor g1889 (n1887, n1849, n1214, n1635, n1868);
or   g1890 (n1902, n1863, n1159, n1263, n1200);
nor  g1891 (n1904, n1225, n1089, n1148, n1856);
and  g1892 (n1899, n1193, n1864, n1255, n1850);
or   g1893 (n1930, n1203, n1100, n1851, n1259);
nor  g1894 (n1873, n1146, n1860, n1158, n1173);
nand g1895 (n1946, n1239, n1130, n1294, n1860);
and  g1896 (n1925, n1861, n1140, n1181, n1077);
and  g1897 (n1882, n1251, n1226, n1634, n1122);
xor  g1898 (n1903, n1793, n1296, n1177, n1168);
nand g1899 (n1920, n1863, n1174, n1858, n1284);
or   g1900 (n1884, n1126, n1285, n1862, n1853);
and  g1901 (n1915, n1288, n1857, n1118, n1099);
or   g1902 (n1910, n1134, n1280, n1202, n1257);
not  g1903 (n2007, n1900);
not  g1904 (n2016, n1894);
not  g1905 (n1986, n1928);
not  g1906 (n2034, n1911);
not  g1907 (n2051, n1919);
not  g1908 (n2033, n1876);
not  g1909 (n2021, n1890);
not  g1910 (n1996, n1892);
buf  g1911 (n2065, n1874);
not  g1912 (n1969, n1914);
buf  g1913 (n2040, n1934);
not  g1914 (n2000, n1935);
not  g1915 (n1970, n1920);
not  g1916 (n2006, n1893);
not  g1917 (n2054, n1929);
not  g1918 (n2026, n1881);
buf  g1919 (n2036, n1942);
buf  g1920 (n2023, n1870);
buf  g1921 (n2039, n1930);
not  g1922 (n2043, n1942);
buf  g1923 (n1997, n1879);
not  g1924 (n2048, n1893);
not  g1925 (n2042, n1929);
not  g1926 (n1987, n1947);
buf  g1927 (n2047, n1878);
not  g1928 (n2035, n1896);
not  g1929 (n1957, n1917);
buf  g1930 (n2058, n1913);
buf  g1931 (n1963, n1888);
buf  g1932 (n1973, n1880);
buf  g1933 (n1985, n1892);
not  g1934 (n2068, n1899);
buf  g1935 (n1953, n1923);
not  g1936 (n2075, n1909);
not  g1937 (n2044, n1924);
buf  g1938 (n2013, n1877);
buf  g1939 (n1954, n1930);
buf  g1940 (n2009, n1919);
buf  g1941 (n2050, n1903);
not  g1942 (n2083, n1948);
not  g1943 (n1983, n1907);
not  g1944 (n2081, n1940);
buf  g1945 (n1981, n1926);
buf  g1946 (n2012, n1945);
buf  g1947 (n1989, n1904);
buf  g1948 (n2061, n1934);
buf  g1949 (n2073, n1927);
not  g1950 (n2022, n1933);
not  g1951 (n1972, n1931);
not  g1952 (n2027, n1893);
buf  g1953 (n2014, n1937);
buf  g1954 (n2017, n1933);
not  g1955 (n1977, n1941);
buf  g1956 (n2030, n1877);
not  g1957 (n2038, n1937);
buf  g1958 (n2032, n1921);
buf  g1959 (n2062, n1930);
buf  g1960 (n2045, n1882);
not  g1961 (n1955, n1881);
not  g1962 (n1962, n1914);
buf  g1963 (n2005, n1908);
buf  g1964 (n2064, n1888);
buf  g1965 (n2049, n1677);
buf  g1966 (n2037, n1936);
buf  g1967 (n2055, n1872);
not  g1968 (n1990, n1929);
not  g1969 (n1966, n1913);
buf  g1970 (n1974, n1946);
not  g1971 (n2008, n1914);
buf  g1972 (n2072, n1937);
xor  g1973 (n2052, n1911, n1912, n1931, n1678);
xnor g1974 (n2069, n1943, n1944, n1912, n1907);
nand g1975 (n2025, n1895, n1946, n1931, n1939);
nand g1976 (n1952, n1920, n1877, n1880, n1898);
nand g1977 (n2003, n1889, n1897, n1876, n1893);
nor  g1978 (n1984, n1919, n1884, n1906, n1940);
xor  g1979 (n2041, n1939, n1869, n1932, n1907);
xor  g1980 (n2078, n1915, n1940, n1920, n1883);
xor  g1981 (n2067, n1678, n1882, n1898, n1924);
xor  g1982 (n2024, n1925, n1890, n1920, n1916);
nor  g1983 (n1959, n1921, n1943, n1932, n1299);
and  g1984 (n2080, n1871, n1900, n1875, n1915);
xnor g1985 (n1978, n1926, n1678, n1948, n1941);
and  g1986 (n1999, n1620, n1892, n1891, n1871);
xor  g1987 (n2020, n1927, n1901, n1887, n1928);
nand g1988 (n2060, n1945, n1902, n1894, n1910);
nor  g1989 (n1951, n1948, n1944, n1928, n1934);
xor  g1990 (n2002, n1922, n1899, n1872, n1885);
xnor g1991 (n2053, n1890, n1902, n1891, n1871);
nand g1992 (n1960, n1925, n1921, n1932, n1872);
nor  g1993 (n1995, n1938, n1940, n1922, n1300);
xnor g1994 (n1988, n1910, n1884, n1945, n1872);
xnor g1995 (n1968, n1924, n1888, n1884, n1918);
nand g1996 (n2019, n1882, n1943, n1935, n1879);
nor  g1997 (n1993, n1910, n1886, n1678, n1301);
and  g1998 (n1979, n1947, n1938, n1927, n1897);
xnor g1999 (n2071, n1930, n1917, n1873, n1902);
and  g2000 (n2015, n1926, n1871, n1894, n1882);
or   g2001 (n1964, n1943, n1917, n1909, n1936);
nand g2002 (n2070, n1869, n1941, n1890, n1919);
xnor g2003 (n1994, n1901, n1935, n1925, n1885);
xor  g2004 (n2018, n1935, n1944, n1878, n1894);
and  g2005 (n2046, n1887, n1883, n1899, n1916);
xnor g2006 (n1998, n1887, n1900, n1895, n1921);
xor  g2007 (n2082, n1904, n1918, n1899, n1908);
and  g2008 (n1992, n1873, n1907, n1874, n1885);
and  g2009 (n2011, n1892, n1942, n1881, n1923);
nand g2010 (n2029, n1885, n1873, n1944, n1875);
nor  g2011 (n2028, n1901, n1886, n1896, n1941);
nand g2012 (n2010, n1875, n1886, n1914, n1938);
nand g2013 (n2056, n1906, n1922, n1908);
nor  g2014 (n2076, n1926, n1900, n1884, n1897);
xor  g2015 (n2077, n1874, n1909, n1876, n1916);
and  g2016 (n1958, n1928, n1905, n1906, n1873);
xnor g2017 (n2031, n1909, n1936, n1933, n1869);
nor  g2018 (n1967, n1889, n1911, n1870, n1878);
or   g2019 (n1950, n1916, n1927, n1869, n1904);
xor  g2020 (n1961, n1918, n1896, n1903, n1905);
and  g2021 (n2079, n1945, n1904, n1879, n1915);
and  g2022 (n1975, n1934, n1924, n1905, n1879);
nor  g2023 (n2074, n1929, n1946, n1915, n1876);
xnor g2024 (n2063, n1870, n1877, n1891, n1939);
and  g2025 (n2057, n1939, n1895, n1942, n1933);
and  g2026 (n1976, n1948, n1925, n1947, n1880);
xnor g2027 (n1956, n1931, n1875, n1883, n1913);
nand g2028 (n1980, n1302, n1937, n1889);
or   g2029 (n2004, n1881, n1903, n1947, n1896);
nor  g2030 (n1971, n1878, n1938, n1912, n1905);
or   g2031 (n1991, n1886, n1874, n1898, n1923);
nor  g2032 (n1949, n1901, n1932, n1891, n1936);
and  g2033 (n1982, n1908, n1880, n1888, n1870);
nor  g2034 (n2066, n1906, n1902, n1895, n1911);
xnor g2035 (n1965, n1923, n1912, n1918, n1913);
xnor g2036 (n2059, n1917, n1897, n1946, n1887);
xnor g2037 (n2001, n1898, n1910, n1883, n1903);
nor  g2038 (n2126, n1453, n1329, n1337, n1553);
or   g2039 (n2128, n2022, n2053, n2076, n1314);
and  g2040 (n2165, n2070, n1957, n1389, n1340);
nor  g2041 (n2085, n1585, n1367, n1445, n1541);
xnor g2042 (n2123, n1305, n1438, n2000, n1577);
xor  g2043 (n2162, n1400, n1960, n1545, n1403);
nor  g2044 (n2102, n2031, n1989, n1420, n1383);
and  g2045 (n2130, n2049, n2066, n1331, n1507);
nand g2046 (n2169, n1455, n1971, n1326, n1476);
xor  g2047 (n2118, n1462, n1345, n1583, n2050);
nor  g2048 (n2127, n1409, n1416, n1594, n1979);
nor  g2049 (n2172, n2041, n1408, n1479, n1562);
and  g2050 (n2101, n1961, n2017, n1518, n2037);
xor  g2051 (n2106, n1970, n1324, n1402, n1358);
nor  g2052 (n2116, n2021, n1592, n1560, n1414);
xor  g2053 (n2095, n1552, n1515, n1962, n1953);
and  g2054 (n2105, n1575, n1317, n1441, n1439);
xnor g2055 (n2142, n2002, n1352, n2026, n1558);
xor  g2056 (n2122, n1536, n1376, n1984, n1338);
xnor g2057 (n2103, n1437, n1591, n1996, n1539);
xnor g2058 (n2098, n1373, n1505, n1418, n2043);
xor  g2059 (n2147, n1374, n1313, n2030, n1956);
xor  g2060 (n2191, n1974, n2068, n1548, n1958);
xor  g2061 (n2088, n1547, n1977, n1559, n1357);
and  g2062 (n2140, n1516, n2083, n1556, n1316);
xor  g2063 (n2156, n1425, n1388, n2004, n1508);
and  g2064 (n2185, n1406, n2007, n1988, n1363);
xor  g2065 (n2158, n1955, n1514, n1482, n1963);
and  g2066 (n2178, n1571, n1386, n1472, n1387);
xor  g2067 (n2153, n2045, n1976, n1303, n1347);
nor  g2068 (n2160, n2016, n1370, n1322, n1584);
xor  g2069 (n2138, n2071, n1581, n2006, n1475);
xnor g2070 (n2129, n1336, n1982, n1465, n1521);
nor  g2071 (n2112, n1464, n2014, n1484, n1596);
or   g2072 (n2154, n1385, n1372, n1580, n1540);
nor  g2073 (n2155, n2065, n1458, n1595, n1412);
nand g2074 (n2132, n2058, n1382, n1572, n1587);
or   g2075 (n2152, n1350, n1423, n1448, n1456);
xor  g2076 (n2117, n2039, n1991, n1426, n1312);
and  g2077 (n2164, n1990, n1398, n2025, n2035);
nor  g2078 (n2121, n1306, n2013, n1494, n1546);
xnor g2079 (n2171, n1434, n1361, n1446, n2027);
xnor g2080 (n2175, n1538, n1362, n2054, n1333);
nor  g2081 (n2186, n1353, n1461, n1332, n1344);
or   g2082 (n2114, n1959, n1517, n1529, n1325);
nor  g2083 (n2131, n1429, n1474, n1483, n1371);
nand g2084 (n2148, n1304, n1579, n1492, n2080);
and  g2085 (n2157, n1404, n1566, n2061, n1466);
or   g2086 (n2137, n1993, n1341, n1401, n2073);
or   g2087 (n2150, n1318, n1951, n1535, n1574);
xnor g2088 (n2177, n1582, n1307, n1463, n2044);
xor  g2089 (n2094, n1335, n1513, n1334, n2001);
xor  g2090 (n2092, n2047, n1489, n2028, n1491);
nor  g2091 (n2167, n2060, n1987, n1557, n1319);
nor  g2092 (n2136, n1490, n1360, n1534, n1949);
xor  g2093 (n2120, n2011, n1497, n2033, n1520);
or   g2094 (n2181, n1995, n2055, n2056, n1433);
nor  g2095 (n2159, n1586, n1485, n1997, n1410);
xor  g2096 (n2168, n1365, n1509, n2009, n1502);
nor  g2097 (n2107, n2064, n1369, n1377, n2015);
nor  g2098 (n2188, n1570, n1348, n2074, n2020);
xor  g2099 (n2115, n1459, n1405, n1342, n1500);
nor  g2100 (n2124, n1522, n1442, n1597, n1569);
or   g2101 (n2119, n1328, n1496, n1486, n1506);
xor  g2102 (n2163, n2042, n2081, n1952, n1966);
xnor g2103 (n2135, n1573, n1309, n1578, n1391);
xnor g2104 (n2099, n2038, n1593, n1950, n1351);
or   g2105 (n2125, n1599, n1436, n1481, n2082);
nor  g2106 (n2183, n2063, n1395, n1537, n1551);
or   g2107 (n2134, n2069, n2048, n1381, n1498);
xor  g2108 (n2187, n2003, n1975, n1364, n1417);
or   g2109 (n2087, n1311, n1435, n1444, n1564);
xor  g2110 (n2149, n1432, n1568, n1965, n1390);
or   g2111 (n2176, n1527, n1589, n1524, n1321);
nand g2112 (n2189, n1368, n1512, n1379, n1493);
xnor g2113 (n2180, n2005, n1356, n1511, n2046);
xor  g2114 (n2184, n1549, n1588, n1983, n1470);
nor  g2115 (n2090, n1565, n1973, n1503, n1468);
or   g2116 (n2097, n1978, n1985, n2062, n1394);
xnor g2117 (n2104, n2079, n1519, n1431, n2012);
xnor g2118 (n2084, n1495, n1349, n1488, n1460);
xor  g2119 (n2161, n1378, n2023, n1422, n1427);
xor  g2120 (n2111, n2067, n2034, n1320, n1419);
and  g2121 (n2110, n1964, n1413, n1544, n2052);
nor  g2122 (n2109, n1968, n1366, n1469, n1533);
xor  g2123 (n2093, n2010, n1396, n1454, n1526);
xnor g2124 (n2190, n1561, n1473, n1504, n1994);
xor  g2125 (n2174, n2040, n1327, n1457, n1315);
xor  g2126 (n2143, n2029, n1450, n2018, n1555);
xor  g2127 (n2170, n1415, n1397, n1308, n1359);
xnor g2128 (n2173, n1449, n1375, n1530, n1339);
nand g2129 (n2096, n1501, n1999, n1543, n2059);
and  g2130 (n2166, n2077, n2057, n1384, n1330);
xor  g2131 (n2133, n1399, n2019, n2036, n1563);
or   g2132 (n2091, n1430, n1380, n2051, n1986);
and  g2133 (n2141, n2075, n1969, n1554, n1478);
xor  g2134 (n2145, n1480, n1310, n1428, n1440);
nor  g2135 (n2146, n1407, n2032, n1471, n1992);
nor  g2136 (n2139, n1411, n1523, n1499, n1528);
xnor g2137 (n2182, n1954, n1443, n1567, n1452);
nand g2138 (n2108, n1998, n1393, n1343, n1487);
and  g2139 (n2100, n1550, n1576, n1542, n1972);
xnor g2140 (n2089, n1590, n1980, n1531, n1467);
nor  g2141 (n2151, n2008, n1447, n1392, n2078);
nand g2142 (n2144, n1532, n1598, n1981, n2024);
xor  g2143 (n2179, n1424, n1525, n1354, n1355);
xor  g2144 (n2113, n2072, n1323, n1421, n1346);
xor  g2145 (n2086, n1477, n1510, n1451, n1967);
nor  g2146 (n2192, n2182, n2187, n2170, n2117);
nor  g2147 (n2218, n2177, n2085, n2137, n2159);
nand g2148 (n2200, n2119, n2088, n2166, n2148);
and  g2149 (n2205, n2171, n2106, n2143, n2162);
nor  g2150 (n2210, n2158, n2113, n2144, n2190);
and  g2151 (n2212, n2115, n2086, n2167, n2138);
or   g2152 (n2197, n2141, n2142, n2163, n2095);
nor  g2153 (n2216, n2165, n2136, n2118, n2099);
xor  g2154 (n2207, n2125, n2104, n2090, n2178);
nor  g2155 (n2202, n2120, n2109, n2147, n2128);
and  g2156 (n2193, n2091, n2152, n2145, n2174);
nand g2157 (n2206, n2130, n2134, n2151, n2172);
nand g2158 (n2196, n2189, n2129, n2168, n2179);
nor  g2159 (n2211, n2191, n2124, n2156, n2135);
or   g2160 (n2198, n2183, n2096, n2173, n2150);
xnor g2161 (n2194, n2132, n2175, n2087, n2140);
nor  g2162 (n2217, n2100, n2160, n2181, n2098);
nand g2163 (n2209, n2094, n2146, n2169, n2108);
or   g2164 (n2203, n2126, n2155, n2121, n2092);
and  g2165 (n2204, n2185, n2176, n2097, n2122);
or   g2166 (n2195, n2157, n2110, n2116, n2101);
nor  g2167 (n2214, n2114, n2093, n2111, n2149);
xor  g2168 (n2215, n2139, n2107, n2180, n2184);
nor  g2169 (n2213, n2131, n2153, n2133, n2161);
or   g2170 (n2208, n2103, n2164, n2084, n2127);
xor  g2171 (n2201, n2123, n2186, n2154, n2188);
xnor g2172 (n2199, n2112, n2105, n2102, n2089);
endmodule
