// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1425_15_11 written by SynthGen on 2021/05/24 19:45:39
module Stat_1425_15_11( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23,
 n1432, n1445, n1437, n1442, n1438, n1443, n1431, n1433,
 n1444, n1440, n1435, n1447, n1439, n1436, n1441, n1434,
 n1448, n1446);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23;

output n1432, n1445, n1437, n1442, n1438, n1443, n1431, n1433,
 n1444, n1440, n1435, n1447, n1439, n1436, n1441, n1434,
 n1448, n1446;

wire n24, n25, n26, n27, n28, n29, n30, n31,
 n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n402, n403, n404, n405, n406, n407,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n425, n426, n427, n428, n429, n430, n431,
 n432, n433, n434, n435, n436, n437, n438, n439,
 n440, n441, n442, n443, n444, n445, n446, n447,
 n448, n449, n450, n451, n452, n453, n454, n455,
 n456, n457, n458, n459, n460, n461, n462, n463,
 n464, n465, n466, n467, n468, n469, n470, n471,
 n472, n473, n474, n475, n476, n477, n478, n479,
 n480, n481, n482, n483, n484, n485, n486, n487,
 n488, n489, n490, n491, n492, n493, n494, n495,
 n496, n497, n498, n499, n500, n501, n502, n503,
 n504, n505, n506, n507, n508, n509, n510, n511,
 n512, n513, n514, n515, n516, n517, n518, n519,
 n520, n521, n522, n523, n524, n525, n526, n527,
 n528, n529, n530, n531, n532, n533, n534, n535,
 n536, n537, n538, n539, n540, n541, n542, n543,
 n544, n545, n546, n547, n548, n549, n550, n551,
 n552, n553, n554, n555, n556, n557, n558, n559,
 n560, n561, n562, n563, n564, n565, n566, n567,
 n568, n569, n570, n571, n572, n573, n574, n575,
 n576, n577, n578, n579, n580, n581, n582, n583,
 n584, n585, n586, n587, n588, n589, n590, n591,
 n592, n593, n594, n595, n596, n597, n598, n599,
 n600, n601, n602, n603, n604, n605, n606, n607,
 n608, n609, n610, n611, n612, n613, n614, n615,
 n616, n617, n618, n619, n620, n621, n622, n623,
 n624, n625, n626, n627, n628, n629, n630, n631,
 n632, n633, n634, n635, n636, n637, n638, n639,
 n640, n641, n642, n643, n644, n645, n646, n647,
 n648, n649, n650, n651, n652, n653, n654, n655,
 n656, n657, n658, n659, n660, n661, n662, n663,
 n664, n665, n666, n667, n668, n669, n670, n671,
 n672, n673, n674, n675, n676, n677, n678, n679,
 n680, n681, n682, n683, n684, n685, n686, n687,
 n688, n689, n690, n691, n692, n693, n694, n695,
 n696, n697, n698, n699, n700, n701, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735,
 n736, n737, n738, n739, n740, n741, n742, n743,
 n744, n745, n746, n747, n748, n749, n750, n751,
 n752, n753, n754, n755, n756, n757, n758, n759,
 n760, n761, n762, n763, n764, n765, n766, n767,
 n768, n769, n770, n771, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n794, n795, n796, n797, n798, n799,
 n800, n801, n802, n803, n804, n805, n806, n807,
 n808, n809, n810, n811, n812, n813, n814, n815,
 n816, n817, n818, n819, n820, n821, n822, n823,
 n824, n825, n826, n827, n828, n829, n830, n831,
 n832, n833, n834, n835, n836, n837, n838, n839,
 n840, n841, n842, n843, n844, n845, n846, n847,
 n848, n849, n850, n851, n852, n853, n854, n855,
 n856, n857, n858, n859, n860, n861, n862, n863,
 n864, n865, n866, n867, n868, n869, n870, n871,
 n872, n873, n874, n875, n876, n877, n878, n879,
 n880, n881, n882, n883, n884, n885, n886, n887,
 n888, n889, n890, n891, n892, n893, n894, n895,
 n896, n897, n898, n899, n900, n901, n902, n903,
 n904, n905, n906, n907, n908, n909, n910, n911,
 n912, n913, n914, n915, n916, n917, n918, n919,
 n920, n921, n922, n923, n924, n925, n926, n927,
 n928, n929, n930, n931, n932, n933, n934, n935,
 n936, n937, n938, n939, n940, n941, n942, n943,
 n944, n945, n946, n947, n948, n949, n950, n951,
 n952, n953, n954, n955, n956, n957, n958, n959,
 n960, n961, n962, n963, n964, n965, n966, n967,
 n968, n969, n970, n971, n972, n973, n974, n975,
 n976, n977, n978, n979, n980, n981, n982, n983,
 n984, n985, n986, n987, n988, n989, n990, n991,
 n992, n993, n994, n995, n996, n997, n998, n999,
 n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
 n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
 n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
 n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
 n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
 n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
 n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
 n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
 n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
 n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
 n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
 n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
 n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
 n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
 n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
 n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
 n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
 n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
 n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
 n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
 n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
 n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
 n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
 n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
 n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
 n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
 n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
 n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
 n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
 n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
 n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
 n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
 n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
 n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
 n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
 n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
 n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
 n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
 n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
 n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
 n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
 n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
 n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
 n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
 n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
 n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
 n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
 n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
 n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
 n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
 n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
 n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
 n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
 n1424, n1425, n1426, n1427, n1428, n1429, n1430;

buf  g0 (n52, n9);
not  g1 (n27, n14);
buf  g2 (n62, n7);
not  g3 (n25, n19);
not  g4 (n29, n7);
not  g5 (n34, n6);
not  g6 (n65, n16);
buf  g7 (n73, n21);
not  g8 (n64, n13);
buf  g9 (n66, n3);
not  g10 (n106, n15);
buf  g11 (n55, n4);
not  g12 (n95, n19);
not  g13 (n68, n22);
buf  g14 (n87, n13);
not  g15 (n32, n17);
buf  g16 (n76, n11);
buf  g17 (n94, n20);
buf  g18 (n60, n14);
not  g19 (n38, n10);
not  g20 (n77, n13);
buf  g21 (n104, n9);
buf  g22 (n49, n12);
buf  g23 (n97, n1);
not  g24 (n84, n16);
not  g25 (n69, n20);
not  g26 (n59, n18);
buf  g27 (n57, n2);
not  g28 (n91, n6);
buf  g29 (n86, n5);
buf  g30 (n24, n4);
buf  g31 (n80, n14);
not  g32 (n93, n3);
buf  g33 (n81, n1);
not  g34 (n46, n6);
buf  g35 (n92, n18);
buf  g36 (n45, n11);
buf  g37 (n102, n3);
not  g38 (n54, n6);
buf  g39 (n36, n4);
buf  g40 (n41, n11);
buf  g41 (n98, n5);
not  g42 (n82, n9);
buf  g43 (n96, n15);
not  g44 (n26, n21);
not  g45 (n39, n17);
not  g46 (n37, n15);
not  g47 (n63, n12);
buf  g48 (n61, n17);
not  g49 (n101, n15);
not  g50 (n83, n13);
buf  g51 (n89, n8);
buf  g52 (n72, n12);
buf  g53 (n33, n7);
not  g54 (n111, n2);
buf  g55 (n103, n20);
not  g56 (n67, n11);
buf  g57 (n31, n16);
buf  g58 (n51, n10);
not  g59 (n56, n8);
buf  g60 (n99, n8);
buf  g61 (n40, n5);
not  g62 (n53, n3);
not  g63 (n42, n21);
not  g64 (n75, n2);
not  g65 (n100, n16);
not  g66 (n44, n1);
buf  g67 (n43, n2);
buf  g68 (n85, n4);
buf  g69 (n90, n17);
not  g70 (n70, n21);
buf  g71 (n79, n8);
not  g72 (n71, n14);
not  g73 (n28, n19);
not  g74 (n48, n7);
buf  g75 (n50, n10);
buf  g76 (n35, n22);
not  g77 (n78, n18);
not  g78 (n58, n1);
not  g79 (n47, n10);
buf  g80 (n107, n9);
buf  g81 (n110, n22);
buf  g82 (n109, n22);
not  g83 (n105, n20);
not  g84 (n74, n5);
buf  g85 (n108, n19);
buf  g86 (n30, n18);
buf  g87 (n88, n12);
buf  g88 (n150, n66);
xor  g89 (n144, n76, n79, n89, n68);
nand g90 (n114, n57, n76, n80);
nand g91 (n134, n100, n64, n95, n104);
xor  g92 (n117, n78, n91, n73, n74);
nor  g93 (n152, n75, n46, n99, n101);
xnor g94 (n143, n26, n27, n31, n78);
or   g95 (n130, n83, n101, n96, n77);
and  g96 (n115, n71, n81, n98, n63);
and  g97 (n137, n30, n73, n59, n50);
or   g98 (n136, n25, n33, n102, n41);
and  g99 (n124, n81, n105, n90);
nand g100 (n146, n105, n49, n58, n68);
nor  g101 (n139, n73, n83, n79, n94);
and  g102 (n112, n66, n81, n105, n84);
xnor g103 (n142, n103, n92, n29, n28);
xor  g104 (n116, n98, n79, n84, n97);
nand g105 (n145, n40, n65, n75, n103);
and  g106 (n123, n96, n74, n93, n44);
and  g107 (n147, n96, n99, n85, n67);
xor  g108 (n118, n87, n70, n80, n77);
xor  g109 (n127, n100, n70, n69, n48);
nor  g110 (n138, n51, n55, n86, n91);
or   g111 (n125, n82, n37, n72, n90);
xnor g112 (n119, n92, n67, n84, n77);
xnor g113 (n140, n35, n104, n39, n32);
nand g114 (n113, n62, n98, n34, n106);
nor  g115 (n135, n82, n89, n36, n70);
and  g116 (n122, n80, n87, n56, n75);
nor  g117 (n148, n102, n74, n89, n94);
and  g118 (n149, n100, n86, n91, n52);
nand g119 (n132, n72, n42, n65, n97);
or   g120 (n133, n66, n103, n38, n93);
xor  g121 (n121, n65, n45, n102, n85);
nor  g122 (n153, n53, n68, n88, n61);
xnor g123 (n126, n88, n87, n71, n95);
nand g124 (n151, n99, n94, n67, n93);
and  g125 (n128, n43, n69, n104, n60);
nand g126 (n141, n71, n47, n78, n97);
xor  g127 (n129, n69, n95, n86, n72);
or   g128 (n120, n83, n101, n88, n24);
xnor g129 (n131, n85, n92, n82, n54);
not  g130 (n193, n146);
not  g131 (n182, n133);
not  g132 (n158, n122);
not  g133 (n172, n145);
not  g134 (n173, n116);
buf  g135 (n187, n131);
not  g136 (n164, n127);
buf  g137 (n177, n113);
buf  g138 (n186, n153);
not  g139 (n195, n134);
not  g140 (n180, n136);
not  g141 (n194, n139);
not  g142 (n190, n142);
not  g143 (n189, n151);
not  g144 (n154, n118);
buf  g145 (n181, n136);
xnor g146 (n169, n125, n119, n149, n126);
and  g147 (n170, n150, n145, n127, n114);
nor  g148 (n168, n124, n140, n134, n143);
nor  g149 (n166, n124, n131, n141, n130);
nand g150 (n156, n115, n129, n146, n140);
and  g151 (n155, n121, n148, n113);
xor  g152 (n160, n129, n119, n135, n133);
xor  g153 (n163, n140, n134, n137, n147);
xnor g154 (n176, n124, n117, n125, n131);
and  g155 (n178, n152, n137, n146, n144);
xnor g156 (n167, n128, n141, n151, n147);
nand g157 (n184, n117, n138, n139, n130);
nor  g158 (n161, n141, n135, n123);
xnor g159 (n185, n153, n126, n133, n122);
or   g160 (n159, n137, n120, n149, n123);
and  g161 (n188, n150, n139, n136, n121);
xor  g162 (n162, n126, n150, n122, n116);
xnor g163 (n175, n125, n113, n120, n117);
or   g164 (n192, n138, n114, n152, n130);
nor  g165 (n191, n129, n132, n149, n145);
and  g166 (n174, n138, n127, n144, n152);
and  g167 (n196, n132, n151, n128, n115);
xnor g168 (n183, n143, n115, n120, n142);
nand g169 (n165, n143, n147, n114, n153);
xnor g170 (n171, n144, n118, n112, n132);
and  g171 (n179, n119, n135, n148, n121);
nor  g172 (n157, n116, n128, n142, n118);
not  g173 (n208, n173);
buf  g174 (n215, n163);
not  g175 (n201, n178);
buf  g176 (n214, n157);
not  g177 (n197, n181);
buf  g178 (n210, n162);
not  g179 (n209, n170);
buf  g180 (n203, n161);
not  g181 (n216, n160);
buf  g182 (n207, n175);
buf  g183 (n202, n169);
buf  g184 (n199, n158);
buf  g185 (n205, n180);
not  g186 (n212, n174);
not  g187 (n204, n155);
buf  g188 (n217, n166);
or   g189 (n211, n156, n168);
nor  g190 (n200, n167, n154);
nor  g191 (n206, n159, n171);
or   g192 (n213, n177, n172);
nor  g193 (n218, n179, n164);
xnor g194 (n198, n176, n165);
not  g195 (n221, n205);
buf  g196 (n224, n206);
buf  g197 (n223, n202);
not  g198 (n228, n197);
buf  g199 (n222, n199);
buf  g200 (n225, n200);
buf  g201 (n227, n203);
not  g202 (n226, n201);
buf  g203 (n220, n182);
or   g204 (n219, n204, n198);
buf  g205 (n233, n228);
buf  g206 (n236, n192);
not  g207 (n247, n187);
not  g208 (n237, n219);
not  g209 (n257, n223);
not  g210 (n246, n219);
buf  g211 (n249, n227);
buf  g212 (n234, n195);
not  g213 (n238, n224);
buf  g214 (n264, n186);
not  g215 (n240, n190);
not  g216 (n258, n228);
not  g217 (n260, n110);
buf  g218 (n253, n189);
buf  g219 (n254, n23);
buf  g220 (n265, n227);
not  g221 (n239, n191);
not  g222 (n242, n220);
xor  g223 (n262, n209, n221, n194, n226);
xor  g224 (n244, n111, n227, n187, n223);
xor  g225 (n230, n219, n193, n107, n184);
nor  g226 (n256, n214, n225, n215);
nand g227 (n266, n224, n208, n192, n109);
and  g228 (n241, n207, n107, n226, n218);
nand g229 (n232, n191, n220, n108, n106);
nor  g230 (n250, n226, n108, n190, n220);
nand g231 (n231, n111, n219, n221, n227);
xor  g232 (n261, n228, n110, n23, n224);
xnor g233 (n235, n189, n226, n222, n108);
and  g234 (n255, n223, n187, n23, n210);
xnor g235 (n251, n193, n217, n225, n185);
or   g236 (n267, n190, n224, n223, n107);
xor  g237 (n245, n211, n193, n222, n183);
or   g238 (n229, n222, n23, n191, n109);
xor  g239 (n259, n221, n194, n106, n222);
xnor g240 (n252, n109, n189, n192, n110);
xor  g241 (n248, n225, n220, n195, n194);
xor  g242 (n243, n221, n188, n228, n216);
xnor g243 (n263, n188, n188, n212, n213);
not  g244 (n287, n245);
not  g245 (n270, n246);
buf  g246 (n326, n239);
buf  g247 (n292, n230);
buf  g248 (n293, n242);
not  g249 (n304, n244);
not  g250 (n298, n236);
not  g251 (n279, n236);
buf  g252 (n303, n245);
not  g253 (n341, n242);
buf  g254 (n306, n238);
buf  g255 (n334, n229);
not  g256 (n315, n229);
not  g257 (n286, n231);
buf  g258 (n312, n240);
not  g259 (n337, n248);
not  g260 (n269, n234);
not  g261 (n288, n237);
buf  g262 (n331, n241);
not  g263 (n277, n237);
not  g264 (n321, n241);
not  g265 (n319, n249);
buf  g266 (n275, n230);
buf  g267 (n285, n245);
not  g268 (n322, n244);
not  g269 (n302, n242);
buf  g270 (n273, n230);
buf  g271 (n300, n249);
buf  g272 (n325, n247);
not  g273 (n280, n239);
buf  g274 (n301, n229);
not  g275 (n289, n238);
buf  g276 (n307, n233);
buf  g277 (n308, n238);
buf  g278 (n317, n239);
buf  g279 (n305, n240);
not  g280 (n323, n247);
buf  g281 (n330, n231);
not  g282 (n335, n247);
not  g283 (n338, n248);
buf  g284 (n336, n239);
buf  g285 (n282, n233);
not  g286 (n278, n244);
buf  g287 (n268, n235);
buf  g288 (n339, n237);
not  g289 (n297, n246);
not  g290 (n320, n233);
buf  g291 (n324, n243);
not  g292 (n299, n244);
buf  g293 (n327, n248);
buf  g294 (n274, n236);
not  g295 (n332, n241);
buf  g296 (n311, n243);
not  g297 (n271, n249);
buf  g298 (n296, n235);
not  g299 (n316, n234);
not  g300 (n333, n242);
not  g301 (n328, n232);
not  g302 (n310, n232);
buf  g303 (n291, n246);
buf  g304 (n276, n243);
buf  g305 (n290, n232);
not  g306 (n329, n241);
buf  g307 (n314, n245);
not  g308 (n295, n247);
buf  g309 (n309, n243);
not  g310 (n272, n248);
buf  g311 (n313, n235);
buf  g312 (n340, n231);
not  g313 (n318, n246);
buf  g314 (n294, n240);
not  g315 (n284, n234);
not  g316 (n281, n240);
not  g317 (n283, n249);
not  g318 (n406, n254);
not  g319 (n383, n287);
buf  g320 (n384, n252);
buf  g321 (n409, n255);
not  g322 (n363, n250);
not  g323 (n379, n250);
buf  g324 (n380, n274);
buf  g325 (n366, n287);
not  g326 (n349, n280);
buf  g327 (n407, n287);
not  g328 (n344, n286);
not  g329 (n388, n285);
not  g330 (n359, n258);
buf  g331 (n351, n278);
buf  g332 (n404, n281);
not  g333 (n367, n256);
buf  g334 (n398, n253);
buf  g335 (n413, n276);
buf  g336 (n408, n281);
buf  g337 (n393, n250);
buf  g338 (n352, n281);
buf  g339 (n381, n258);
buf  g340 (n347, n279);
buf  g341 (n403, n258);
buf  g342 (n399, n284);
not  g343 (n418, n284);
not  g344 (n346, n269);
not  g345 (n354, n272);
not  g346 (n420, n279);
not  g347 (n385, n257);
buf  g348 (n356, n282);
not  g349 (n389, n283);
not  g350 (n412, n280);
not  g351 (n400, n278);
not  g352 (n405, n278);
buf  g353 (n401, n269);
buf  g354 (n396, n281);
not  g355 (n373, n259);
not  g356 (n343, n277);
buf  g357 (n345, n252);
not  g358 (n414, n250);
buf  g359 (n361, n252);
buf  g360 (n395, n259);
buf  g361 (n372, n283);
buf  g362 (n421, n272);
buf  g363 (n348, n254);
not  g364 (n370, n270);
buf  g365 (n350, n268);
buf  g366 (n410, n256);
not  g367 (n382, n286);
buf  g368 (n394, n258);
buf  g369 (n377, n257);
buf  g370 (n387, n282);
buf  g371 (n375, n272);
buf  g372 (n364, n275);
not  g373 (n419, n280);
buf  g374 (n353, n252);
buf  g375 (n374, n284);
not  g376 (n360, n268);
not  g377 (n371, n285);
not  g378 (n362, n254);
not  g379 (n417, n255);
buf  g380 (n390, n283);
not  g381 (n392, n274);
buf  g382 (n386, n256);
buf  g383 (n416, n269);
nand g384 (n358, n270, n259);
xor  g385 (n397, n275, n273, n254);
xnor g386 (n369, n251, n282, n256, n273);
nor  g387 (n342, n271, n282, n279, n285);
nor  g388 (n402, n280, n257, n255, n283);
nor  g389 (n368, n253, n251, n268, n275);
or   g390 (n376, n251, n271, n255, n277);
nand g391 (n378, n286, n270, n253);
nand g392 (n355, n251, n276, n278, n273);
or   g393 (n357, n277, n271, n274, n268);
or   g394 (n365, n277, n271, n257, n269);
and  g395 (n415, n275, n276, n287, n259);
xor  g396 (n391, n285, n279, n276, n272);
xnor g397 (n411, n274, n284, n253, n286);
not  g398 (n523, n390);
not  g399 (n526, n341);
not  g400 (n505, n315);
not  g401 (n466, n383);
buf  g402 (n554, n323);
buf  g403 (n430, n339);
not  g404 (n527, n394);
buf  g405 (n507, n365);
not  g406 (n473, n340);
not  g407 (n467, n375);
buf  g408 (n440, n350);
nand g409 (n426, n329, n293);
or   g410 (n539, n299, n366, n346, n260);
xor  g411 (n543, n302, n310, n262, n365);
nand g412 (n499, n404, n314, n297, n415);
or   g413 (n432, n311, n338, n261, n395);
and  g414 (n458, n322, n306, n399, n328);
nor  g415 (n437, n387, n395, n318, n334);
nand g416 (n427, n315, n347, n342, n379);
xnor g417 (n487, n405, n367, n368, n350);
xor  g418 (n504, n367, n331, n397, n326);
nor  g419 (n435, n336, n394, n305, n401);
or   g420 (n446, n301, n320, n339, n382);
or   g421 (n489, n291, n319, n299, n418);
or   g422 (n550, n394, n386, n260, n416);
xor  g423 (n469, n352, n421, n371, n387);
xnor g424 (n423, n335, n296, n314, n407);
or   g425 (n558, n357, n343, n310, n313);
nand g426 (n566, n297, n344, n291, n325);
or   g427 (n448, n111, n365, n305, n374);
xor  g428 (n479, n371, n289, n387, n375);
and  g429 (n534, n378, n336, n407, n261);
and  g430 (n535, n337, n356, n307, n309);
or   g431 (n444, n339, n393, n391, n400);
nand g432 (n560, n195, n416, n410, n381);
nor  g433 (n510, n316, n314, n363, n420);
and  g434 (n555, n321, n324, n289, n366);
and  g435 (n518, n389, n298, n313, n405);
xor  g436 (n447, n319, n355, n306, n301);
xnor g437 (n549, n297, n317, n420, n353);
or   g438 (n424, n325, n317, n295, n323);
nor  g439 (n517, n343, n335, n367, n361);
or   g440 (n488, n343, n348, n312, n342);
or   g441 (n438, n370, n362, n388, n378);
nand g442 (n544, n312, n361, n294, n360);
and  g443 (n500, n347, n404, n408, n368);
nor  g444 (n513, n419, n351, n359, n346);
xor  g445 (n477, n322, n294, n348, n300);
nand g446 (n509, n355, n410, n301, n288);
xnor g447 (n483, n374, n334, n386, n311);
nand g448 (n521, n348, n387, n383, n403);
and  g449 (n567, n364, n417, n346, n309);
xnor g450 (n472, n359, n421, n356, n327);
nor  g451 (n450, n343, n354, n359, n380);
or   g452 (n493, n369, n369, n301, n308);
nand g453 (n564, n345, n302, n350, n397);
or   g454 (n492, n386, n381, n421, n403);
xor  g455 (n429, n417, n353, n302);
and  g456 (n562, n352, n388, n385, n392);
xnor g457 (n553, n404, n393, n400, n351);
xnor g458 (n485, n373, n359, n361, n407);
xor  g459 (n455, n294, n381, n300, n389);
and  g460 (n512, n356, n307, n288, n355);
nor  g461 (n460, n335, n409, n318, n358);
xor  g462 (n545, n376, n358, n319, n326);
or   g463 (n542, n321, n416, n372, n326);
xnor g464 (n520, n352, n344, n378, n304);
xnor g465 (n502, n341, n344, n369, n335);
xor  g466 (n471, n377, n345, n384, n414);
xnor g467 (n552, n328, n316, n292, n318);
xor  g468 (n449, n377, n376, n332, n410);
nor  g469 (n515, n305, n358, n416, n324);
or   g470 (n494, n303, n404, n331, n317);
xor  g471 (n459, n298, n346, n299, n330);
and  g472 (n525, n337, n352, n377, n414);
xnor g473 (n461, n420, n330, n310);
xnor g474 (n425, n295, n333, n378, n393);
and  g475 (n516, n350, n261, n388, n315);
xor  g476 (n434, n398, n354, n348, n403);
nand g477 (n433, n369, n391, n384, n386);
nand g478 (n556, n417, n322, n363, n325);
nor  g479 (n561, n362, n377, n364, n349);
or   g480 (n551, n397, n357, n303, n323);
nor  g481 (n511, n357, n320, n339, n304);
xor  g482 (n490, n396, n307, n409, n384);
xnor g483 (n563, n391, n389, n406, n320);
xor  g484 (n532, n407, n289, n392, n318);
xor  g485 (n529, n368, n405, n293, n329);
and  g486 (n533, n345, n333, n327, n349);
and  g487 (n537, n329, n415, n298, n374);
xnor g488 (n522, n373, n337, n294, n323);
and  g489 (n484, n402, n296, n324, n262);
nand g490 (n546, n406, n316, n290, n379);
xnor g491 (n540, n288, n399, n332);
or   g492 (n462, n313, n392, n375, n355);
nor  g493 (n465, n327, n414, n331, n371);
nor  g494 (n475, n300, n307, n298, n370);
xor  g495 (n531, n380, n196, n309, n398);
nand g496 (n514, n398, n383, n292, n370);
and  g497 (n495, n360, n314, n336, n385);
nand g498 (n538, n351, n290, n415, n371);
nor  g499 (n454, n337, n290, n385, n400);
nor  g500 (n486, n373, n395, n295, n408);
xor  g501 (n439, n390, n379, n312, n413);
xor  g502 (n557, n296, n313, n308, n353);
nor  g503 (n496, n308, n419, n390, n364);
nor  g504 (n519, n373, n325, n411, n312);
and  g505 (n503, n415, n401, n399, n397);
nand g506 (n470, n305, n419, n341, n365);
xor  g507 (n468, n408, n322, n411, n295);
and  g508 (n524, n351, n384, n306, n410);
or   g509 (n508, n342, n389, n390, n316);
or   g510 (n456, n381, n413, n319, n328);
xor  g511 (n480, n376, n292, n347, n361);
or   g512 (n547, n372, n419, n341, n327);
xnor g513 (n498, n360, n328, n311, n379);
nand g514 (n491, n362, n414, n296, n340);
and  g515 (n478, n338, n317, n309, n383);
and  g516 (n452, n394, n392, n421, n405);
xnor g517 (n451, n310, n336, n393, n297);
and  g518 (n457, n342, n411, n261, n324);
xor  g519 (n453, n338, n396, n380, n320);
xor  g520 (n481, n388, n293, n406, n418);
xor  g521 (n443, n340, n353, n418, n326);
or   g522 (n464, n406, n315, n329, n303);
and  g523 (n428, n368, n391, n354, n363);
nor  g524 (n474, n400, n334, n288, n260);
xor  g525 (n506, n306, n347, n364, n385);
xnor g526 (n548, n418, n366, n358, n401);
and  g527 (n565, n332, n402, n412);
xnor g528 (n442, n409, n349, n299, n399);
xnor g529 (n431, n402, n338, n290, n412);
xnor g530 (n528, n291, n308, n398, n366);
xor  g531 (n476, n356, n382, n262, n380);
and  g532 (n530, n357, n413, n396, n372);
xor  g533 (n463, n344, n340, n374, n289);
nand g534 (n436, n260, n409, n345, n395);
xor  g535 (n536, n334, n408, n304, n376);
xnor g536 (n482, n413, n375, n333, n411);
and  g537 (n445, n372, n321, n330, n363);
nor  g538 (n422, n291, n321, n403, n420);
and  g539 (n541, n354, n367, n370, n396);
nand g540 (n501, n412, n331, n300, n311);
xnor g541 (n497, n401, n382, n360);
xor  g542 (n559, n349, n333, n304, n303);
nand g543 (n441, n292, n412, n417, n362);
buf  g544 (n816, n458);
not  g545 (n806, n514);
not  g546 (n913, n483);
not  g547 (n653, n496);
not  g548 (n898, n561);
not  g549 (n902, n481);
not  g550 (n929, n481);
not  g551 (n652, n534);
not  g552 (n881, n469);
not  g553 (n740, n479);
buf  g554 (n672, n483);
buf  g555 (n768, n495);
not  g556 (n885, n501);
buf  g557 (n585, n542);
buf  g558 (n646, n488);
buf  g559 (n697, n456);
buf  g560 (n640, n454);
buf  g561 (n706, n488);
not  g562 (n584, n566);
not  g563 (n804, n535);
not  g564 (n698, n480);
not  g565 (n670, n476);
not  g566 (n942, n547);
buf  g567 (n887, n427);
not  g568 (n873, n459);
not  g569 (n689, n522);
buf  g570 (n732, n559);
not  g571 (n645, n539);
not  g572 (n739, n565);
not  g573 (n759, n551);
not  g574 (n890, n540);
not  g575 (n575, n470);
not  g576 (n916, n560);
not  g577 (n907, n544);
not  g578 (n834, n545);
buf  g579 (n702, n501);
not  g580 (n909, n445);
not  g581 (n583, n552);
not  g582 (n578, n532);
not  g583 (n846, n517);
buf  g584 (n663, n546);
buf  g585 (n861, n438);
buf  g586 (n691, n519);
not  g587 (n751, n509);
buf  g588 (n860, n525);
buf  g589 (n635, n507);
buf  g590 (n744, n477);
buf  g591 (n788, n555);
not  g592 (n579, n461);
not  g593 (n918, n554);
buf  g594 (n800, n565);
not  g595 (n880, n452);
buf  g596 (n606, n500);
buf  g597 (n681, n478);
buf  g598 (n680, n549);
buf  g599 (n819, n556);
buf  g600 (n850, n486);
not  g601 (n793, n526);
buf  g602 (n827, n545);
buf  g603 (n822, n546);
buf  g604 (n883, n490);
not  g605 (n839, n462);
not  g606 (n943, n486);
buf  g607 (n667, n536);
buf  g608 (n874, n551);
buf  g609 (n664, n470);
buf  g610 (n760, n485);
buf  g611 (n758, n504);
not  g612 (n593, n522);
buf  g613 (n941, n518);
not  g614 (n684, n537);
buf  g615 (n630, n523);
not  g616 (n636, n426);
not  g617 (n810, n466);
not  g618 (n610, n437);
buf  g619 (n832, n540);
not  g620 (n725, n472);
not  g621 (n620, n530);
buf  g622 (n932, n523);
buf  g623 (n682, n496);
not  g624 (n656, n447);
buf  g625 (n794, n446);
not  g626 (n614, n514);
buf  g627 (n735, n543);
not  g628 (n651, n487);
not  g629 (n766, n560);
buf  g630 (n581, n474);
buf  g631 (n869, n516);
not  g632 (n752, n526);
not  g633 (n865, n457);
buf  g634 (n710, n498);
buf  g635 (n922, n548);
buf  g636 (n708, n507);
buf  g637 (n623, n492);
buf  g638 (n777, n530);
not  g639 (n796, n489);
not  g640 (n668, n554);
buf  g641 (n779, n511);
buf  g642 (n944, n423);
buf  g643 (n661, n520);
buf  g644 (n838, n564);
not  g645 (n780, n475);
buf  g646 (n685, n471);
not  g647 (n693, n465);
not  g648 (n848, n562);
buf  g649 (n625, n510);
buf  g650 (n650, n458);
buf  g651 (n920, n530);
not  g652 (n638, n541);
not  g653 (n836, n558);
not  g654 (n705, n567);
buf  g655 (n933, n545);
not  g656 (n809, n471);
buf  g657 (n641, n524);
buf  g658 (n703, n452);
buf  g659 (n730, n451);
buf  g660 (n724, n504);
not  g661 (n782, n500);
not  g662 (n855, n550);
not  g663 (n628, n517);
not  g664 (n720, n497);
buf  g665 (n569, n543);
not  g666 (n738, n538);
not  g667 (n683, n462);
not  g668 (n603, n527);
not  g669 (n644, n473);
buf  g670 (n715, n485);
buf  g671 (n677, n486);
buf  g672 (n755, n566);
not  g673 (n829, n547);
buf  g674 (n727, n498);
not  g675 (n891, n502);
not  g676 (n917, n521);
buf  g677 (n844, n477);
buf  g678 (n707, n505);
not  g679 (n622, n458);
not  g680 (n924, n533);
not  g681 (n787, n556);
buf  g682 (n634, n506);
buf  g683 (n927, n460);
not  g684 (n673, n559);
not  g685 (n856, n443);
not  g686 (n817, n483);
not  g687 (n925, n429);
buf  g688 (n901, n487);
buf  g689 (n778, n463);
buf  g690 (n831, n535);
buf  g691 (n807, n428);
not  g692 (n899, n562);
buf  g693 (n795, n425);
not  g694 (n769, n539);
not  g695 (n737, n454);
not  g696 (n676, n521);
buf  g697 (n826, n497);
buf  g698 (n671, n484);
buf  g699 (n776, n482);
not  g700 (n756, n502);
buf  g701 (n824, n520);
not  g702 (n658, n440);
not  g703 (n587, n460);
not  g704 (n642, n467);
not  g705 (n747, n453);
buf  g706 (n718, n509);
not  g707 (n745, n552);
not  g708 (n906, n537);
not  g709 (n763, n503);
buf  g710 (n936, n196);
buf  g711 (n892, n554);
not  g712 (n589, n464);
not  g713 (n728, n502);
not  g714 (n597, n562);
not  g715 (n701, n478);
not  g716 (n785, n548);
buf  g717 (n746, n564);
buf  g718 (n602, n494);
not  g719 (n678, n474);
not  g720 (n823, n549);
not  g721 (n815, n469);
not  g722 (n805, n472);
buf  g723 (n599, n531);
not  g724 (n731, n467);
not  g725 (n717, n436);
buf  g726 (n736, n510);
buf  g727 (n719, n476);
not  g728 (n604, n515);
not  g729 (n571, n468);
not  g730 (n875, n532);
buf  g731 (n914, n555);
not  g732 (n700, n527);
not  g733 (n821, n466);
not  g734 (n774, n474);
not  g735 (n792, n516);
buf  g736 (n611, n479);
buf  g737 (n711, n476);
not  g738 (n568, n529);
not  g739 (n862, n527);
buf  g740 (n786, n557);
buf  g741 (n757, n494);
buf  g742 (n781, n493);
buf  g743 (n930, n510);
buf  g744 (n660, n525);
not  g745 (n921, n465);
not  g746 (n905, n431);
not  g747 (n812, n473);
not  g748 (n609, n555);
not  g749 (n716, n452);
buf  g750 (n595, n524);
buf  g751 (n939, n508);
not  g752 (n935, n563);
buf  g753 (n852, n477);
buf  g754 (n940, n537);
not  g755 (n773, n435);
not  g756 (n764, n459);
not  g757 (n904, n515);
buf  g758 (n631, n433);
not  g759 (n616, n498);
buf  g760 (n798, n468);
not  g761 (n666, n457);
buf  g762 (n704, n494);
not  g763 (n864, n491);
not  g764 (n726, n455);
not  g765 (n878, n550);
not  g766 (n841, n506);
buf  g767 (n692, n567);
not  g768 (n748, n542);
not  g769 (n686, n512);
buf  g770 (n582, n424);
not  g771 (n714, n478);
buf  g772 (n910, n528);
buf  g773 (n868, n432);
not  g774 (n849, n538);
not  g775 (n833, n543);
buf  g776 (n837, n434);
not  g777 (n813, n471);
not  g778 (n879, n520);
not  g779 (n871, n519);
buf  g780 (n937, n448);
buf  g781 (n662, n485);
buf  g782 (n859, n460);
not  g783 (n742, n495);
buf  g784 (n627, n466);
not  g785 (n770, n506);
buf  g786 (n900, n557);
buf  g787 (n601, n513);
not  g788 (n863, n529);
buf  g789 (n811, n521);
buf  g790 (n655, n482);
not  g791 (n722, n512);
not  g792 (n761, n499);
buf  g793 (n851, n490);
buf  g794 (n882, n479);
buf  g795 (n590, n501);
not  g796 (n600, n469);
buf  g797 (n767, n533);
not  g798 (n699, n441);
buf  g799 (n818, n456);
not  g800 (n613, n422);
buf  g801 (n657, n529);
not  g802 (n749, n524);
buf  g803 (n753, n463);
not  g804 (n723, n511);
buf  g805 (n771, n518);
buf  g806 (n621, n511);
buf  g807 (n665, n556);
buf  g808 (n729, n531);
not  g809 (n872, n472);
not  g810 (n687, n491);
not  g811 (n743, n534);
not  g812 (n586, n455);
buf  g813 (n612, n516);
not  g814 (n574, n503);
not  g815 (n866, n558);
not  g816 (n903, n565);
buf  g817 (n842, n513);
buf  g818 (n617, n481);
not  g819 (n695, n566);
not  g820 (n934, n484);
buf  g821 (n607, n561);
not  g822 (n605, n450);
not  g823 (n931, n499);
not  g824 (n791, n430);
buf  g825 (n694, n489);
not  g826 (n802, n461);
not  g827 (n639, n454);
not  g828 (n825, n508);
not  g829 (n911, n489);
buf  g830 (n576, n509);
buf  g831 (n828, n559);
not  g832 (n928, n522);
buf  g833 (n893, n557);
buf  g834 (n884, n526);
not  g835 (n632, n505);
buf  g836 (n896, n464);
buf  g837 (n647, n544);
buf  g838 (n734, n470);
buf  g839 (n637, n439);
not  g840 (n840, n488);
buf  g841 (n762, n196);
not  g842 (n808, n525);
not  g843 (n799, n464);
not  g844 (n629, n517);
buf  g845 (n858, n550);
not  g846 (n820, n503);
buf  g847 (n675, n512);
not  g848 (n654, n535);
not  g849 (n649, n262);
not  g850 (n889, n528);
buf  g851 (n754, n533);
not  g852 (n570, n461);
not  g853 (n772, n457);
buf  g854 (n877, n519);
not  g855 (n789, n453);
buf  g856 (n573, n490);
not  g857 (n783, n442);
not  g858 (n690, n553);
not  g859 (n915, n560);
not  g860 (n857, n508);
buf  g861 (n721, n465);
not  g862 (n688, n541);
not  g863 (n912, n492);
buf  g864 (n897, n552);
buf  g865 (n596, n563);
buf  g866 (n619, n444);
buf  g867 (n867, n558);
buf  g868 (n803, n453);
not  g869 (n784, n549);
not  g870 (n712, n459);
buf  g871 (n908, n534);
not  g872 (n591, n551);
buf  g873 (n709, n480);
buf  g874 (n775, n532);
not  g875 (n919, n493);
not  g876 (n847, n561);
buf  g877 (n797, n499);
not  g878 (n835, n462);
buf  g879 (n618, n487);
buf  g880 (n801, n504);
not  g881 (n626, n455);
buf  g882 (n669, n553);
not  g883 (n830, n513);
buf  g884 (n598, n515);
not  g885 (n853, n449);
buf  g886 (n886, n500);
buf  g887 (n713, n456);
not  g888 (n845, n482);
not  g889 (n696, n505);
buf  g890 (n594, n563);
not  g891 (n814, n493);
not  g892 (n843, n548);
buf  g893 (n633, n531);
buf  g894 (n894, n546);
buf  g895 (n870, n497);
not  g896 (n741, n553);
not  g897 (n854, n492);
not  g898 (n938, n484);
not  g899 (n577, n540);
buf  g900 (n588, n514);
buf  g901 (n608, n564);
not  g902 (n888, n467);
buf  g903 (n679, n495);
not  g904 (n750, n507);
not  g905 (n643, n536);
buf  g906 (n580, n523);
not  g907 (n765, n544);
buf  g908 (n674, n473);
not  g909 (n926, n542);
not  g910 (n923, n539);
not  g911 (n733, n491);
not  g912 (n895, n538);
buf  g913 (n648, n518);
buf  g914 (n592, n480);
not  g915 (n876, n496);
buf  g916 (n659, n475);
buf  g917 (n624, n567);
not  g918 (n615, n541);
xnor g919 (n790, n475, n528);
xor  g920 (n572, n463, n468, n536, n547);
and  g921 (n1133, n913, n774, n904, n846);
xor  g922 (n1130, n872, n802, n742, n617);
xnor g923 (n985, n883, n838, n626, n698);
and  g924 (n1216, n714, n821, n710, n666);
and  g925 (n1144, n839, n623, n919, n912);
nand g926 (n1264, n758, n651, n786, n745);
xnor g927 (n1194, n635, n669, n936, n608);
nor  g928 (n1139, n832, n777, n914, n710);
nor  g929 (n1059, n827, n756, n604, n763);
and  g930 (n1225, n929, n848, n938, n811);
xnor g931 (n978, n614, n885, n613, n636);
or   g932 (n1281, n857, n877, n730, n871);
and  g933 (n1248, n644, n790, n593, n609);
xor  g934 (n1167, n857, n763, n830, n635);
nor  g935 (n1269, n888, n917, n732, n754);
nand g936 (n1169, n615, n791, n696, n576);
xnor g937 (n1190, n855, n729, n920, n737);
xor  g938 (n1249, n614, n934, n573, n697);
and  g939 (n1191, n733, n861, n634, n585);
xor  g940 (n1117, n895, n784, n776, n742);
or   g941 (n1120, n803, n597, n898, n696);
or   g942 (n1219, n678, n599, n846, n922);
xnor g943 (n1000, n908, n757, n808, n656);
and  g944 (n1220, n924, n868, n726, n878);
nor  g945 (n1231, n652, n679, n939, n676);
xor  g946 (n1273, n792, n670, n758, n892);
and  g947 (n1047, n870, n722, n784, n745);
xor  g948 (n1283, n626, n639, n691, n910);
or   g949 (n1235, n607, n737, n883, n852);
xor  g950 (n1043, n680, n896, n758, n693);
nor  g951 (n1230, n842, n783, n602, n790);
or   g952 (n1146, n716, n813, n879, n743);
xnor g953 (n1125, n721, n714, n676, n704);
and  g954 (n1013, n776, n927, n612, n926);
nor  g955 (n1166, n596, n944, n725, n786);
nor  g956 (n1062, n685, n661, n761, n766);
xor  g957 (n947, n662, n692, n654, n893);
xnor g958 (n1189, n940, n870, n900, n660);
nand g959 (n1205, n692, n925, n869, n646);
xor  g960 (n1032, n833, n718, n597, n796);
or   g961 (n1079, n632, n941, n740, n703);
xnor g962 (n991, n736, n629, n806, n852);
xnor g963 (n1042, n916, n856, n853, n748);
xor  g964 (n1008, n712, n862, n742, n593);
xor  g965 (n1050, n882, n647, n715, n826);
and  g966 (n1121, n860, n917, n823, n706);
xor  g967 (n1165, n690, n833, n805, n595);
xor  g968 (n1178, n821, n686, n605, n876);
and  g969 (n1174, n687, n851, n921, n849);
xnor g970 (n1068, n875, n817, n599, n809);
or   g971 (n1217, n794, n815, n829, n796);
xnor g972 (n1223, n920, n755, n906, n621);
or   g973 (n1029, n637, n723, n892);
nand g974 (n1019, n890, n808, n641, n787);
and  g975 (n1039, n873, n792, n938, n741);
or   g976 (n980, n653, n747, n709, n807);
xor  g977 (n1168, n884, n698, n821, n862);
or   g978 (n1212, n940, n687, n897, n664);
nand g979 (n1088, n858, n636, n926, n798);
xor  g980 (n1275, n799, n639, n666, n890);
or   g981 (n1221, n736, n929, n602, n908);
xor  g982 (n1105, n878, n666, n860, n800);
or   g983 (n1002, n798, n648, n615, n765);
xor  g984 (n1066, n747, n942, n629, n759);
xnor g985 (n1046, n590, n824, n934, n724);
xnor g986 (n1095, n666, n859, n873, n701);
and  g987 (n1017, n586, n841, n630, n750);
xnor g988 (n1015, n901, n713, n668, n886);
xor  g989 (n1090, n630, n765, n752, n732);
xor  g990 (n1285, n677, n765, n684, n905);
nor  g991 (n1234, n893, n635, n785, n611);
xor  g992 (n1010, n649, n740, n884, n699);
or   g993 (n946, n827, n700, n764, n793);
nand g994 (n961, n845, n891, n919, n691);
xnor g995 (n1024, n880, n708, n711, n717);
or   g996 (n1270, n935, n897, n810, n611);
or   g997 (n1164, n662, n724, n911, n709);
and  g998 (n1224, n711, n619, n877, n889);
and  g999 (n983, n751, n655, n714, n730);
and  g1000 (n1159, n886, n861, n654, n807);
or   g1001 (n1238, n846, n886, n720, n876);
or   g1002 (n1100, n638, n887, n603, n816);
nand g1003 (n1142, n824, n783, n938, n690);
nand g1004 (n1061, n674, n921, n713, n810);
or   g1005 (n1176, n699, n933, n826, n876);
and  g1006 (n973, n826, n750, n624, n828);
xnor g1007 (n1197, n633, n869, n596, n892);
and  g1008 (n1027, n899, n736, n768, n773);
nand g1009 (n1201, n927, n771, n765, n760);
and  g1010 (n1243, n841, n833, n737, n808);
nand g1011 (n1185, n776, n596, n914, n624);
or   g1012 (n949, n817, n745, n692, n702);
and  g1013 (n1097, n747, n836, n614, n798);
nor  g1014 (n1242, n809, n569, n856, n689);
xor  g1015 (n1034, n712, n750, n636, n935);
and  g1016 (n1161, n755, n759, n865, n682);
nand g1017 (n1056, n930, n710, n794, n901);
xnor g1018 (n1001, n943, n826, n908, n711);
xor  g1019 (n1132, n940, n615, n686, n864);
nor  g1020 (n1123, n681, n931, n659, n669);
and  g1021 (n1214, n695, n581, n899, n906);
nand g1022 (n1004, n871, n894, n632, n760);
xnor g1023 (n1158, n917, n589, n613, n631);
xnor g1024 (n1150, n858, n801, n718, n617);
xor  g1025 (n1172, n918, n739, n789, n811);
nand g1026 (n952, n891, n804, n722, n835);
nor  g1027 (n1018, n766, n802, n941, n723);
xor  g1028 (n963, n887, n813, n812, n701);
or   g1029 (n1060, n863, n888, n730, n801);
nand g1030 (n1075, n807, n658, n675, n822);
and  g1031 (n1128, n591, n755, n624, n832);
and  g1032 (n1082, n617, n901, n681, n856);
xor  g1033 (n976, n718, n893, n782, n702);
or   g1034 (n1192, n719, n902, n796, n684);
and  g1035 (n1077, n818, n931, n651, n781);
and  g1036 (n1206, n819, n697, n722, n853);
xor  g1037 (n1064, n713, n935, n737, n872);
or   g1038 (n1250, n742, n744, n935, n823);
xnor g1039 (n1202, n798, n898, n827, n625);
nand g1040 (n1003, n755, n648, n837, n689);
xor  g1041 (n1229, n788, n620, n720, n606);
or   g1042 (n1086, n683, n810, n759, n874);
nor  g1043 (n1232, n894, n932, n642, n784);
nor  g1044 (n1198, n769, n944, n835, n610);
xnor g1045 (n977, n744, n699, n836, n939);
nor  g1046 (n1246, n682, n591, n909, n713);
nand g1047 (n1259, n616, n853, n937, n942);
or   g1048 (n1129, n893, n677, n703, n812);
xnor g1049 (n1226, n688, n571, n875, n895);
xnor g1050 (n1084, n600, n926, n693, n777);
nor  g1051 (n974, n824, n793, n799, n734);
and  g1052 (n1069, n930, n921, n866, n705);
xnor g1053 (n1277, n847, n679, n657, n610);
nor  g1054 (n1089, n854, n923, n731, n841);
nor  g1055 (n1058, n900, n619, n718, n882);
and  g1056 (n1065, n793, n694, n601, n761);
xor  g1057 (n1257, n915, n670, n669, n762);
xnor g1058 (n1210, n848, n717, n704, n827);
and  g1059 (n1107, n606, n834, n930, n880);
nand g1060 (n1284, n594, n575, n693, n778);
xor  g1061 (n1119, n922, n844, n752, n835);
and  g1062 (n1151, n910, n889, n690, n683);
and  g1063 (n1126, n918, n684, n894, n867);
xor  g1064 (n1049, n929, n654, n733, n860);
and  g1065 (n1009, n905, n698, n762, n693);
or   g1066 (n1022, n744, n771, n649, n857);
xnor g1067 (n1258, n661, n849, n939, n660);
nand g1068 (n1183, n925, n782, n667, n941);
xor  g1069 (n966, n680, n717, n812, n813);
and  g1070 (n951, n795, n708, n775, n620);
or   g1071 (n975, n637, n785, n769, n779);
xor  g1072 (n954, n832, n691, n897, n804);
nor  g1073 (n1154, n944, n762, n707, n644);
xor  g1074 (n1080, n655, n943, n913, n909);
xor  g1075 (n1156, n649, n804, n640, n918);
nor  g1076 (n1237, n814, n790, n705, n904);
or   g1077 (n984, n820, n634, n684, n770);
xnor g1078 (n1140, n728, n771, n744, n797);
xor  g1079 (n997, n679, n669, n944, n735);
xor  g1080 (n1262, n761, n915, n824, n791);
nand g1081 (n998, n906, n822, n937, n899);
nand g1082 (n996, n866, n778, n867, n783);
nand g1083 (n1218, n839, n766, n867, n759);
xor  g1084 (n945, n681, n663, n773, n801);
nand g1085 (n964, n695, n792, n940, n660);
and  g1086 (n1245, n616, n597, n936, n720);
or   g1087 (n1173, n682, n631, n913, n699);
xor  g1088 (n1272, n928, n911, n820, n749);
xnor g1089 (n1005, n806, n848, n749, n677);
nand g1090 (n1033, n822, n588, n871);
or   g1091 (n982, n726, n734, n705, n708);
nand g1092 (n1180, n888, n799, n700, n685);
nor  g1093 (n987, n653, n619, n572, n899);
nand g1094 (n1247, n661, n823, n786, n785);
and  g1095 (n1261, n789, n925, n622, n629);
and  g1096 (n1112, n630, n799, n621, n672);
nor  g1097 (n948, n677, n867, n725, n878);
nor  g1098 (n1037, n725, n749, n850, n868);
nand g1099 (n1048, n855, n764, n600, n686);
nor  g1100 (n1195, n675, n820, n872, n709);
xnor g1101 (n1076, n844, n667, n748, n709);
xnor g1102 (n1260, n926, n605, n743, n770);
and  g1103 (n1203, n789, n938, n937, n643);
nor  g1104 (n1145, n668, n936, n603, n775);
and  g1105 (n1116, n639, n768, n650, n869);
xnor g1106 (n1241, n665, n891, n780, n625);
xnor g1107 (n979, n828, n828, n919, n676);
xnor g1108 (n1286, n743, n664, n777, n665);
or   g1109 (n1085, n840, n885, n829, n928);
and  g1110 (n1071, n689, n727, n767, n652);
or   g1111 (n993, n831, n875, n600, n890);
nand g1112 (n1152, n568, n620, n712, n803);
or   g1113 (n1055, n812, n888, n769, n710);
nand g1114 (n962, n687, n800, n882, n851);
nand g1115 (n1153, n928, n818, n678, n840);
or   g1116 (n1138, n838, n829, n780, n910);
xor  g1117 (n1254, n830, n663, n674, n832);
xor  g1118 (n1081, n854, n868, n797, n641);
nand g1119 (n1052, n823, n608, n838, n845);
xor  g1120 (n1098, n727, n730, n924, n579);
and  g1121 (n1115, n805, n770, n724, n657);
nand g1122 (n1073, n874, n902, n633, n820);
nor  g1123 (n989, n896, n605, n688, n920);
nand g1124 (n1256, n859, n915, n828, n734);
nand g1125 (n1016, n728, n708, n815, n818);
xnor g1126 (n1155, n725, n932, n925, n800);
nor  g1127 (n1251, n689, n942, n870, n819);
xnor g1128 (n1054, n673, n903, n907, n746);
nor  g1129 (n1026, n845, n907, n863, n795);
or   g1130 (n1175, n814, n788, n840, n914);
nand g1131 (n1108, n731, n834, n584, n582);
nor  g1132 (n1035, n807, n767, n734, n604);
nor  g1133 (n995, n733, n772, n705, n706);
and  g1134 (n1163, n704, n831, n628, n747);
xnor g1135 (n1287, n746, n645, n934, n657);
nor  g1136 (n1184, n627, n882, n941, n865);
nor  g1137 (n1110, n904, n766, n841, n788);
nor  g1138 (n1057, n774, n817, n753, n869);
nor  g1139 (n1244, n707, n864, n716, n674);
nor  g1140 (n986, n889, n690, n784, n733);
nor  g1141 (n1143, n739, n738, n775, n896);
nor  g1142 (n1147, n795, n628, n681, n738);
and  g1143 (n1091, n927, n908, n595, n738);
and  g1144 (n1072, n674, n670, n825, n796);
nor  g1145 (n1282, n900, n595, n816, n879);
nand g1146 (n953, n589, n931, n691, n701);
xnor g1147 (n1157, n658, n726, n856, n716);
nand g1148 (n1276, n753, n800, n728, n606);
and  g1149 (n970, n673, n937, n736, n740);
nor  g1150 (n1209, n808, n643, n700, n805);
nor  g1151 (n1188, n787, n599, n930, n764);
xor  g1152 (n1199, n932, n778, n763, n896);
and  g1153 (n1136, n645, n662, n761, n648);
nand g1154 (n1274, n819, n852, n727, n773);
or   g1155 (n1101, n598, n905, n777, n703);
and  g1156 (n1092, n664, n646, n621, n748);
nor  g1157 (n1177, n694, n862, n626, n644);
xnor g1158 (n1031, n884, n806, n772, n697);
nand g1159 (n1099, n697, n936, n811, n794);
xnor g1160 (n1170, n916, n787, n667, n741);
nand g1161 (n1186, n772, n667, n751, n702);
or   g1162 (n1278, n861, n916, n825, n785);
xnor g1163 (n1127, n640, n881, n750, n700);
xnor g1164 (n1213, n872, n907, n760, n642);
xnor g1165 (n1204, n868, n746, n834, n833);
and  g1166 (n971, n836, n716, n731, n881);
xor  g1167 (n1267, n721, n891, n774, n850);
nand g1168 (n1063, n701, n780, n845, n751);
xnor g1169 (n1141, n623, n837, n631, n775);
xor  g1170 (n1271, n594, n727, n781, n610);
nor  g1171 (n1040, n618, n696, n905, n756);
or   g1172 (n1122, n588, n876, n860, n842);
and  g1173 (n972, n803, n783, n607, n844);
or   g1174 (n1266, n939, n758, n735, n672);
xor  g1175 (n1279, n837, n739, n593, n583);
xnor g1176 (n1030, n570, n895, n640, n894);
xnor g1177 (n1268, n897, n612, n627, n645);
nor  g1178 (n1200, n590, n651, n818, n752);
nand g1179 (n1025, n625, n906, n789, n843);
nor  g1180 (n1211, n855, n729, n837, n741);
and  g1181 (n1131, n728, n781, n813, n729);
xor  g1182 (n1113, n776, n892, n797, n849);
nor  g1183 (n1222, n685, n866, n675, n874);
or   g1184 (n960, n858, n817, n932, n843);
or   g1185 (n1020, n769, n883, n851, n934);
xnor g1186 (n1239, n885, n767, n589, n900);
nor  g1187 (n1280, n912, n831, n756, n665);
xor  g1188 (n1148, n753, n632, n879, n857);
or   g1189 (n1007, n816, n757, n577, n743);
or   g1190 (n1041, n802, n840, n862, n902);
and  g1191 (n1215, n917, n676, n790, n695);
xnor g1192 (n1023, n904, n863, n923, n746);
and  g1193 (n1263, n830, n883, n659, n752);
xor  g1194 (n1093, n739, n608, n609, n717);
or   g1195 (n988, n751, n831, n928, n801);
xor  g1196 (n957, n943, n591, n859, n712);
nand g1197 (n1233, n682, n863, n788, n738);
xor  g1198 (n981, n819, n779, n672, n673);
xor  g1199 (n1240, n688, n748, n847, n903);
xnor g1200 (n1078, n590, n830, n672, n729);
or   g1201 (n1253, n927, n814, n911, n920);
xnor g1202 (n1070, n616, n910, n671, n756);
and  g1203 (n1187, n901, n873, n749, n779);
xnor g1204 (n1236, n922, n829, n885, n793);
xnor g1205 (n1265, n842, n587, n661, n884);
and  g1206 (n1021, n622, n668, n773, n720);
xnor g1207 (n1102, n787, n611, n647, n836);
xnor g1208 (n1053, n870, n842, n780, n843);
nand g1209 (n1006, n715, n757, n745, n864);
xnor g1210 (n1207, n850, n601, n641, n915);
nand g1211 (n1135, n839, n874, n678, n703);
nor  g1212 (n1196, n878, n865, n861, n679);
xnor g1213 (n959, n778, n844, n911, n919);
nand g1214 (n1181, n732, n923, n854, n786);
nor  g1215 (n956, n623, n603, n678, n839);
nand g1216 (n1087, n609, n574, n881, n764);
and  g1217 (n955, n754, n628, n686, n889);
nor  g1218 (n990, n791, n753, n702, n688);
nand g1219 (n1045, n921, n692, n865, n779);
and  g1220 (n1038, n722, n665, n726, n735);
and  g1221 (n1160, n594, n909, n768, n653);
and  g1222 (n1227, n795, n924, n797, n851);
nand g1223 (n1044, n854, n602, n849, n887);
and  g1224 (n1109, n815, n895, n613, n810);
nand g1225 (n1193, n771, n913, n782, n835);
nand g1226 (n1083, n754, n922, n642, n809);
nor  g1227 (n1252, n754, n803, n767, n578);
and  g1228 (n968, n719, n912, n715, n694);
nand g1229 (n1182, n659, n740, n650, n923);
nand g1230 (n1012, n723, n719, n903, n698);
nand g1231 (n1171, n770, n931, n683, n864);
nand g1232 (n999, n580, n612, n924, n943);
or   g1233 (n1028, n721, n695, n804, n652);
xnor g1234 (n1096, n656, n859, n855, n838);
and  g1235 (n1114, n664, n598, n902, n877);
nor  g1236 (n1134, n886, n706, n933, n873);
or   g1237 (n1104, n858, n662, n637, n731);
or   g1238 (n1103, n704, n871, n877, n903);
nand g1239 (n950, n601, n660, n627, n881);
or   g1240 (n1288, n805, n683, n794, n846);
xnor g1241 (n958, n671, n687, n696, n821);
or   g1242 (n1036, n918, n671, n711, n634);
and  g1243 (n1094, n806, n719, n646, n694);
and  g1244 (n1149, n822, n707, n879, n592);
nand g1245 (n1124, n735, n655, n853, n850);
and  g1246 (n965, n671, n782, n772, n914);
xnor g1247 (n992, n847, n887, n668, n791);
nand g1248 (n1137, n916, n880, n866, n741);
nand g1249 (n1179, n673, n656, n811, n658);
or   g1250 (n1208, n757, n933, n663, n638);
nor  g1251 (n969, n633, n670, n825, n912);
xor  g1252 (n1051, n875, n763, n802, n847);
nand g1253 (n1118, n768, n622, n680, n890);
xor  g1254 (n994, n760, n929, n792, n707);
xor  g1255 (n1162, n685, n942, n598, n933);
xor  g1256 (n1111, n852, n607, n834, n592);
nand g1257 (n1106, n647, n618, n762, n706);
nor  g1258 (n1067, n809, n675, n907, n848);
xnor g1259 (n967, n715, n592, n774, n880);
xor  g1260 (n1255, n816, n843, n815, n724);
xor  g1261 (n1014, n909, n643, n781, n814);
nor  g1262 (n1074, n732, n825, n680, n898);
xnor g1263 (n1228, n663, n714, n618, n604);
xor  g1264 (n1011, n721, n650, n638, n898);
buf  g1265 (n1320, n1018);
buf  g1266 (n1313, n1010);
not  g1267 (n1302, n995);
not  g1268 (n1306, n1003);
buf  g1269 (n1298, n1023);
buf  g1270 (n1307, n981);
buf  g1271 (n1319, n971);
buf  g1272 (n1301, n1034);
not  g1273 (n1300, n1008);
buf  g1274 (n1299, n961);
xnor g1275 (n1311, n1035, n1045, n1004, n1046);
nand g1276 (n1304, n1024, n954, n945, n980);
xor  g1277 (n1317, n966, n948, n969, n1031);
and  g1278 (n1295, n1013, n998, n992, n997);
nand g1279 (n1289, n978, n1039, n949, n987);
and  g1280 (n1297, n984, n1015, n985, n1030);
and  g1281 (n1310, n1025, n1032, n955, n953);
xnor g1282 (n1316, n957, n1028, n996, n1021);
and  g1283 (n1322, n988, n1026, n1043, n1040);
xnor g1284 (n1293, n1019, n970, n999, n974);
nand g1285 (n1309, n977, n958, n973, n986);
nand g1286 (n1314, n1014, n1000, n989, n1001);
nand g1287 (n1291, n960, n1011, n1038, n968);
and  g1288 (n1308, n963, n962, n1033, n967);
nor  g1289 (n1321, n1029, n1016, n1048, n975);
nor  g1290 (n1315, n1049, n982, n1006, n983);
xor  g1291 (n1290, n951, n1022, n991, n947);
xnor g1292 (n1292, n1005, n1012, n1044, n1020);
nand g1293 (n1294, n959, n979, n956, n952);
nor  g1294 (n1305, n1007, n1017, n1027, n1050);
xor  g1295 (n1312, n950, n1009, n993, n972);
xnor g1296 (n1296, n1041, n1047, n1037, n1042);
nand g1297 (n1303, n976, n990, n946, n964);
nor  g1298 (n1318, n1002, n1036, n994, n965);
nand g1299 (n1367, n1305, n1264, n1267, n1317);
nor  g1300 (n1349, n1307, n1306, n1092, n265);
xnor g1301 (n1337, n263, n1056, n1253, n1098);
nor  g1302 (n1386, n1197, n1308, n1083, n1320);
xnor g1303 (n1359, n1188, n1215, n1104, n1216);
nor  g1304 (n1358, n1189, n1126, n1294, n1124);
xnor g1305 (n1370, n1220, n1094, n1322, n263);
nor  g1306 (n1345, n1310, n1311, n1146, n1289);
xor  g1307 (n1387, n1302, n1314, n1285, n264);
xnor g1308 (n1403, n265, n1318, n1308);
and  g1309 (n1393, n1296, n1293, n1232, n1119);
xor  g1310 (n1363, n1274, n1190, n1173, n1322);
xnor g1311 (n1405, n1288, n1130, n1167, n1170);
nor  g1312 (n1380, n1224, n1141, n1247, n1316);
and  g1313 (n1347, n1313, n1191, n1118, n1282);
or   g1314 (n1418, n1066, n1062, n1054, n1321);
or   g1315 (n1333, n1193, n1128, n1278, n1292);
xnor g1316 (n1334, n1085, n1310, n1186, n1093);
xor  g1317 (n1330, n1304, n1160, n1070, n266);
xor  g1318 (n1342, n1081, n1305, n1137, n1096);
nor  g1319 (n1402, n1314, n1155, n1221, n1296);
and  g1320 (n1355, n1145, n1280, n1147, n1068);
nor  g1321 (n1408, n1303, n1231, n1300, n1222);
xnor g1322 (n1381, n1314, n1307, n1310, n1156);
xnor g1323 (n1407, n1313, n1319, n1312);
nand g1324 (n1348, n1270, n1067, n1239, n1111);
or   g1325 (n1400, n1298, n1209, n1206, n1302);
or   g1326 (n1361, n1306, n1105, n1229, n1316);
and  g1327 (n1379, n1260, n1194, n1175, n1163);
xor  g1328 (n1364, n1314, n1257, n1144, n1100);
xor  g1329 (n1325, n1198, n1072, n1245, n1291);
and  g1330 (n1395, n1205, n1311, n1182, n1090);
xor  g1331 (n1327, n1263, n1114, n1265, n1139);
xnor g1332 (n1335, n1236, n1154, n1123, n1305);
or   g1333 (n1413, n1321, n1080, n1200, n1217);
or   g1334 (n1372, n1129, n1110, n1277, n1235);
or   g1335 (n1357, n1295, n1176, n264, n1256);
nor  g1336 (n1331, n1299, n1210, n1185, n1116);
xor  g1337 (n1415, n1181, n1268, n1273, n1196);
or   g1338 (n1328, n1115, n1174, n1243, n1305);
or   g1339 (n1401, n1121, n1136, n1308, n1300);
and  g1340 (n1365, n1060, n1313, n1195, n1320);
xor  g1341 (n1362, n1180, n1259, n1089, n1234);
xor  g1342 (n1398, n1309, n1302, n1299, n1310);
or   g1343 (n1392, n1134, n1071, n266, n1228);
xor  g1344 (n1326, n1319, n1271, n263, n1254);
or   g1345 (n1324, n1286, n1148, n1317, n1058);
nor  g1346 (n1406, n1149, n1297, n1301, n1290);
nand g1347 (n1383, n1078, n1317, n1213, n1291);
xor  g1348 (n1353, n1315, n1087, n1294, n1306);
nor  g1349 (n1329, n1315, n1230, n1276, n1316);
nor  g1350 (n1368, n1287, n1289, n1075, n1103);
xor  g1351 (n1354, n1303, n1309, n1117);
xor  g1352 (n1399, n1122, n1291, n1261, n1303);
nor  g1353 (n1394, n1208, n1241, n1106, n1301);
and  g1354 (n1343, n1251, n1322, n1203, n1112);
nor  g1355 (n1411, n1294, n1171, n1097, n1113);
and  g1356 (n1417, n1292, n1293, n1211, n1237);
nand g1357 (n1391, n1281, n1315, n1275, n1138);
nor  g1358 (n1410, n1169, n1073, n1316, n1053);
nand g1359 (n1323, n1084, n1240, n1319, n1179);
and  g1360 (n1340, n1164, n1150, n1204, n1055);
xor  g1361 (n1389, n1218, n1177, n1290, n1207);
xnor g1362 (n1404, n1153, n1279, n264, n1076);
nor  g1363 (n1369, n1290, n1077, n1320, n1069);
nand g1364 (n1388, n1242, n1102, n1127, n1052);
xnor g1365 (n1378, n1079, n1312, n1225);
nor  g1366 (n1339, n1061, n1142, n1107, n1101);
or   g1367 (n1409, n1143, n1132, n1299);
xor  g1368 (n1373, n1108, n1313, n1297, n1168);
nand g1369 (n1338, n1095, n1307, n1244, n1292);
and  g1370 (n1374, n1311, n1304, n1199, n1258);
or   g1371 (n1336, n1301, n1233, n1201, n1131);
and  g1372 (n1360, n1091, n1184, n1312, n1172);
xnor g1373 (n1385, n1088, n1212, n1246, n1304);
xnor g1374 (n1332, n1255, n1269, n1082, n1162);
and  g1375 (n1414, n1300, n1183, n1214, n1289);
nor  g1376 (n1384, n1152, n1266, n1297, n1051);
xor  g1377 (n1356, n1296, n1161, n1064, n264);
nand g1378 (n1396, n1296, n1178, n1074, n1057);
or   g1379 (n1352, n1295, n1192, n1318, n1283);
xor  g1380 (n1346, n1059, n1300, n1238, n1135);
and  g1381 (n1397, n1272, n1140, n1248, n263);
xor  g1382 (n1371, n1252, n1298, n1304, n1307);
nand g1383 (n1390, n1301, n1250, n1227, n265);
or   g1384 (n1382, n1294, n1125, n1309, n1159);
and  g1385 (n1412, n1187, n1320, n1293, n1157);
or   g1386 (n1416, n1295, n1311, n1249, n1165);
or   g1387 (n1377, n1086, n1321, n1223, n1120);
and  g1388 (n1350, n1306, n1321, n1317, n1226);
and  g1389 (n1341, n1166, n265, n1133, n1303);
xnor g1390 (n1344, n1293, n1318, n1298, n1099);
nor  g1391 (n1351, n1315, n1158, n1151, n1109);
or   g1392 (n1366, n1308, n1295, n1219, n1202);
or   g1393 (n1375, n1065, n1297, n1302, n1284);
or   g1394 (n1376, n1298, n1262, n1063, n1322);
and  g1395 (n1430, n1344, n1362, n1358, n1331);
nand g1396 (n1420, n1330, n1364, n1328, n1329);
xor  g1397 (n1426, n1342, n1323, n1333, n1335);
nor  g1398 (n1425, n1351, n1363, n1332, n1334);
or   g1399 (n1422, n1359, n266, n1354, n267);
and  g1400 (n1421, n1356, n1339, n267, n1352);
nand g1401 (n1423, n267, n1343, n1353, n1345);
and  g1402 (n1419, n1341, n1326, n1325, n267);
nor  g1403 (n1428, n1336, n1327, n1349, n1357);
xor  g1404 (n1424, n1347, n1350, n1355, n1337);
nand g1405 (n1427, n1360, n1340, n1361, n1338);
nand g1406 (n1429, n1346, n266, n1348, n1324);
xnor g1407 (n1439, n1411, n1385, n1428);
or   g1408 (n1440, n1400, n1381, n1391, n1412);
xor  g1409 (n1441, n1430, n1417, n1365, n1427);
or   g1410 (n1433, n1392, n1407, n1398, n1409);
and  g1411 (n1444, n1374, n1415, n1423, n1424);
nand g1412 (n1438, n1373, n1394, n1428, n1429);
xnor g1413 (n1435, n1426, n1429, n1393, n1383);
nor  g1414 (n1436, n1378, n1413, n1382, n1414);
and  g1415 (n1442, n1366, n1404, n1401, n1375);
nand g1416 (n1445, n1369, n1420, n1377, n1416);
nand g1417 (n1432, n1390, n1380, n1410, n1399);
xnor g1418 (n1448, n1397, n1405, n1371, n1379);
xnor g1419 (n1447, n1403, n1386, n1421, n1425);
xor  g1420 (n1434, n1430, n1406, n1387, n1372);
or   g1421 (n1437, n1402, n1376, n1389, n1422);
nor  g1422 (n1443, n1429, n1396, n1430, n1419);
xor  g1423 (n1431, n1384, n1368, n1367, n1408);
xnor g1424 (n1446, n1395, n1370, n1418, n1388);
endmodule
