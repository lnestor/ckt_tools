

module Stat_100_63
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n43,
  n115,
  n88,
  n103,
  n96,
  n97,
  n80,
  n100,
  n66,
  n77,
  n102,
  n75,
  n65,
  n111,
  n78,
  n95,
  n82,
  n106,
  n129,
  n123,
  n121,
  n119,
  n124,
  n125,
  n120,
  n122,
  n127,
  n126,
  n128,
  n132,
  n131,
  n130,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n43;
  output n115;
  output n88;
  output n103;
  output n96;
  output n97;
  output n80;
  output n100;
  output n66;
  output n77;
  output n102;
  output n75;
  output n65;
  output n111;
  output n78;
  output n95;
  output n82;
  output n106;
  output n129;
  output n123;
  output n121;
  output n119;
  output n124;
  output n125;
  output n120;
  output n122;
  output n127;
  output n126;
  output n128;
  output n132;
  output n131;
  output n130;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n76;
  wire n79;
  wire n81;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n98;
  wire n99;
  wire n101;
  wire n104;
  wire n105;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n112;
  wire n113;
  wire n114;
  wire n116;
  wire n117;
  wire n118;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n35,
    n1
  );


  buf
  g1
  (
    KeyWire_0_37,
    n2
  );


  buf
  g2
  (
    KeyWire_0_48,
    n1
  );


  not
  g3
  (
    n37,
    n1
  );


  buf
  g4
  (
    KeyWire_0_55,
    n1
  );


  not
  g5
  (
    n34,
    n2
  );


  not
  g6
  (
    KeyWire_0_53,
    n37
  );


  not
  g7
  (
    KeyWire_0_56,
    n37
  );


  buf
  g8
  (
    KeyWire_0_3,
    n2
  );


  buf
  g9
  (
    n43,
    n3
  );


  nand
  g10
  (
    KeyWire_0_8,
    n2,
    n36
  );


  not
  g11
  (
    KeyWire_0_20,
    n43
  );


  buf
  g12
  (
    n46,
    n40
  );


  buf
  g13
  (
    KeyWire_0_29,
    n41
  );


  not
  g14
  (
    KeyWire_0_7,
    n42
  );


  buf
  g15
  (
    KeyWire_0_13,
    n44
  );


  buf
  g16
  (
    n58,
    n44
  );


  buf
  g17
  (
    KeyWire_0_25,
    n4
  );


  not
  g18
  (
    KeyWire_0_0,
    n5
  );


  buf
  g19
  (
    KeyWire_0_61,
    n47
  );


  buf
  g20
  (
    KeyWire_0_42,
    n45
  );


  buf
  g21
  (
    KeyWire_0_11,
    n4
  );


  buf
  g22
  (
    n63,
    n46
  );


  buf
  g23
  (
    n55,
    n6
  );


  buf
  g24
  (
    n62,
    n3
  );


  buf
  g25
  (
    KeyWire_0_63,
    n46
  );


  buf
  g26
  (
    n53,
    n46
  );


  nor
  g27
  (
    KeyWire_0_16,
    n45,
    n4,
    n5,
    n46
  );


  nor
  g28
  (
    KeyWire_0_59,
    n45,
    n47,
    n44
  );


  xnor
  g29
  (
    KeyWire_0_58,
    n44,
    n5,
    n3,
    n4
  );


  or
  g30
  (
    KeyWire_0_15,
    n47,
    n45,
    n5,
    n3
  );


  not
  g31
  (
    KeyWire_0_31,
    n9
  );


  buf
  g32
  (
    KeyWire_0_40,
    n7
  );


  buf
  g33
  (
    KeyWire_0_22,
    n59
  );


  buf
  g34
  (
    KeyWire_0_62,
    n52
  );


  not
  g35
  (
    n117,
    n26
  );


  not
  g36
  (
    KeyWire_0_6,
    n23
  );


  buf
  g37
  (
    KeyWire_0_5,
    n19
  );


  not
  g38
  (
    n86,
    n50
  );


  buf
  g39
  (
    KeyWire_0_38,
    n38
  );


  not
  g40
  (
    KeyWire_0_28,
    n20
  );


  not
  g41
  (
    n107,
    n60
  );


  not
  g42
  (
    KeyWire_0_27,
    n6
  );


  not
  g43
  (
    KeyWire_0_26,
    n9
  );


  buf
  g44
  (
    KeyWire_0_50,
    n8
  );


  not
  g45
  (
    KeyWire_0_30,
    n28
  );


  xor
  g46
  (
    KeyWire_0_45,
    n20,
    n61,
    n10
  );


  xnor
  g47
  (
    KeyWire_0_34,
    n8,
    n14,
    n18,
    n28
  );


  nor
  g48
  (
    n88,
    n57,
    n56,
    n58,
    n31
  );


  xnor
  g49
  (
    n67,
    n51,
    n56,
    n11,
    n13
  );


  xnor
  g50
  (
    n84,
    n18,
    n61,
    n27,
    n60
  );


  nand
  g51
  (
    KeyWire_0_32,
    n53,
    n18,
    n62
  );


  and
  g52
  (
    n79,
    n14,
    n48,
    n31,
    n7
  );


  xor
  g53
  (
    n89,
    n28,
    n57,
    n60,
    n49
  );


  nor
  g54
  (
    KeyWire_0_41,
    n16,
    n32,
    n15,
    n57
  );


  nor
  g55
  (
    KeyWire_0_1,
    n26,
    n12,
    n31,
    n27
  );


  xnor
  g56
  (
    KeyWire_0_54,
    n21,
    n12,
    n49,
    n32
  );


  nor
  g57
  (
    n102,
    n28,
    n30,
    n14,
    n16
  );


  xnor
  g58
  (
    n78,
    n32,
    n11,
    n15,
    n54
  );


  or
  g59
  (
    n71,
    n16,
    n63,
    n18,
    n25
  );


  nor
  g60
  (
    KeyWire_0_43,
    n53,
    n14,
    n51,
    n57
  );


  nand
  g61
  (
    KeyWire_0_33,
    n22,
    n30,
    n63,
    n58
  );


  xor
  g62
  (
    n74,
    n23,
    n10,
    n37,
    n27
  );


  xor
  g63
  (
    n85,
    n60,
    n29,
    n6,
    n27
  );


  xor
  g64
  (
    KeyWire_0_9,
    n55,
    n53,
    n12,
    n13
  );


  xnor
  g65
  (
    KeyWire_0_36,
    n52,
    n52,
    n21,
    n16
  );


  and
  g66
  (
    n106,
    n25,
    n19,
    n23,
    n55
  );


  or
  g67
  (
    KeyWire_0_19,
    n26,
    n55,
    n63,
    n29
  );


  xnor
  g68
  (
    KeyWire_0_57,
    n59,
    n52,
    n50,
    n13
  );


  or
  g69
  (
    n91,
    n53,
    n15,
    n19,
    n24
  );


  or
  g70
  (
    n116,
    n58,
    n29,
    n56,
    n62
  );


  and
  g71
  (
    KeyWire_0_60,
    n21,
    n38,
    n22,
    n17
  );


  nand
  g72
  (
    n82,
    n23,
    n10,
    n48,
    n51
  );


  xnor
  g73
  (
    KeyWire_0_49,
    n20,
    n48,
    n9,
    n13
  );


  and
  g74
  (
    KeyWire_0_12,
    n6,
    n63,
    n49,
    n10
  );


  and
  g75
  (
    KeyWire_0_14,
    n24,
    n50,
    n7,
    n59
  );


  nor
  g76
  (
    n83,
    n21,
    n24,
    n30
  );


  nand
  g77
  (
    n112,
    n51,
    n54,
    n8,
    n56
  );


  xnor
  g78
  (
    n98,
    n8,
    n22,
    n9,
    n26
  );


  nand
  g79
  (
    KeyWire_0_46,
    n20,
    n59,
    n54,
    n17
  );


  nand
  g80
  (
    n77,
    n49,
    n25,
    n29,
    n61
  );


  nor
  g81
  (
    KeyWire_0_47,
    n15,
    n31,
    n19,
    n12
  );


  and
  g82
  (
    n90,
    n38,
    n58,
    n22,
    n11
  );


  and
  g83
  (
    KeyWire_0_51,
    n55,
    n32,
    n62,
    n48
  );


  nand
  g84
  (
    KeyWire_0_18,
    n7,
    n50,
    n25,
    n54
  );


  or
  g85
  (
    n70,
    n11,
    n30,
    n17
  );


  xnor
  g86
  (
    KeyWire_0_2,
    n118,
    n101,
    n107,
    n115
  );


  xnor
  g87
  (
    KeyWire_0_39,
    n95,
    n110,
    n113,
    n103
  );


  xor
  g88
  (
    KeyWire_0_52,
    n115,
    n111,
    n116,
    n118
  );


  xnor
  g89
  (
    KeyWire_0_44,
    n86,
    n106,
    n100,
    n84
  );


  nor
  g90
  (
    KeyWire_0_23,
    n112,
    n99,
    n94,
    n82
  );


  xnor
  g91
  (
    n120,
    n80,
    n77,
    n117,
    n93
  );


  and
  g92
  (
    KeyWire_0_24,
    n117,
    n97,
    n116,
    n115
  );


  or
  g93
  (
    KeyWire_0_21,
    n117,
    n89,
    n104,
    n98
  );


  and
  g94
  (
    KeyWire_0_35,
    n114,
    n116,
    n88,
    n87
  );


  nand
  g95
  (
    KeyWire_0_10,
    n105,
    n113,
    n96,
    n92
  );


  nor
  g96
  (
    KeyWire_0_17,
    n85,
    n109,
    n102,
    n78
  );


  nand
  g97
  (
    KeyWire_0_4,
    n112,
    n114,
    n90,
    n113
  );


  and
  g98
  (
    n123,
    n79,
    n108,
    n114,
    n112
  );


  and
  g99
  (
    n121,
    n83,
    n118,
    n81,
    n91
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n50,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n118,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n130,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n42,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n129,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n94,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n73,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n45,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n39,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n69,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n125,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n49,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n76,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n61,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n113,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n51,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n60,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n127,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n114,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n64,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n44,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n128,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n80,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n132,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n124,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n59,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n68,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n72,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n97,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n47,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n81,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n110,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n103,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n93,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n105,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n126,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n99,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n36,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n75,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n122,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n100,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n95,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n54,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n96,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n119,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n66,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n101,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n111,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n33,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n65,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n115,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n92,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n131,
    KeyNOTWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n40,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n109,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n38,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n41,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n87,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n48,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n57,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n104,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n56,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n108,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n52,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

