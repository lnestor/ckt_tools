

module Stat_387_1118
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n175,
  n170,
  n167,
  n159,
  n166,
  n151,
  n174,
  n160,
  n157,
  n152,
  n173,
  n182,
  n162,
  n169,
  n406,
  n408,
  n407,
  n409,
  n411,
  n410,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n175;
  output n170;
  output n167;
  output n159;
  output n166;
  output n151;
  output n174;
  output n160;
  output n157;
  output n152;
  output n173;
  output n182;
  output n162;
  output n169;
  output n406;
  output n408;
  output n407;
  output n409;
  output n411;
  output n410;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n158;
  wire n161;
  wire n163;
  wire n164;
  wire n165;
  wire n168;
  wire n171;
  wire n172;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n66,
    n9
  );


  buf
  g1
  (
    n41,
    n11
  );


  not
  g2
  (
    n43,
    n16
  );


  not
  g3
  (
    n45,
    n20
  );


  not
  g4
  (
    n62,
    n14
  );


  buf
  g5
  (
    n35,
    n15
  );


  not
  g6
  (
    n61,
    n4
  );


  not
  g7
  (
    n69,
    n4
  );


  not
  g8
  (
    KeyWire_0_18,
    n17
  );


  not
  g9
  (
    n96,
    n11
  );


  buf
  g10
  (
    KeyWire_0_10,
    n22
  );


  buf
  g11
  (
    n57,
    n6
  );


  buf
  g12
  (
    n91,
    n18
  );


  buf
  g13
  (
    n30,
    n5
  );


  not
  g14
  (
    n67,
    n10
  );


  buf
  g15
  (
    n38,
    n16
  );


  not
  g16
  (
    n25,
    n8
  );


  not
  g17
  (
    n60,
    n17
  );


  buf
  g18
  (
    n74,
    n19
  );


  buf
  g19
  (
    n100,
    n13
  );


  not
  g20
  (
    n83,
    n14
  );


  not
  g21
  (
    n98,
    n23
  );


  not
  g22
  (
    n32,
    n20
  );


  not
  g23
  (
    n99,
    n6
  );


  not
  g24
  (
    n85,
    n15
  );


  not
  g25
  (
    n54,
    n7
  );


  buf
  g26
  (
    n75,
    n8
  );


  not
  g27
  (
    n48,
    n10
  );


  not
  g28
  (
    n49,
    n23
  );


  buf
  g29
  (
    n97,
    n10
  );


  not
  g30
  (
    n87,
    n6
  );


  not
  g31
  (
    n81,
    n20
  );


  buf
  g32
  (
    n70,
    n13
  );


  not
  g33
  (
    n28,
    n18
  );


  buf
  g34
  (
    n36,
    n5
  );


  buf
  g35
  (
    n42,
    n12
  );


  not
  g36
  (
    n92,
    n9
  );


  not
  g37
  (
    n89,
    n8
  );


  buf
  g38
  (
    n47,
    n23
  );


  buf
  g39
  (
    n40,
    n9
  );


  not
  g40
  (
    n84,
    n20
  );


  not
  g41
  (
    n55,
    n15
  );


  not
  g42
  (
    n26,
    n19
  );


  buf
  g43
  (
    n72,
    n21
  );


  not
  g44
  (
    n63,
    n11
  );


  not
  g45
  (
    n39,
    n21
  );


  not
  g46
  (
    n46,
    n16
  );


  not
  g47
  (
    n102,
    n19
  );


  not
  g48
  (
    n37,
    n13
  );


  not
  g49
  (
    n65,
    n18
  );


  not
  g50
  (
    n44,
    n17
  );


  not
  g51
  (
    KeyWire_0_22,
    n22
  );


  not
  g52
  (
    n27,
    n1
  );


  buf
  g53
  (
    KeyWire_0_14,
    n14
  );


  buf
  g54
  (
    n68,
    n2
  );


  buf
  g55
  (
    n86,
    n19
  );


  buf
  g56
  (
    n95,
    n18
  );


  not
  g57
  (
    n56,
    n11
  );


  not
  g58
  (
    n73,
    n7
  );


  buf
  g59
  (
    n31,
    n7
  );


  buf
  g60
  (
    n64,
    n22
  );


  buf
  g61
  (
    n29,
    n7
  );


  not
  g62
  (
    n78,
    n21
  );


  buf
  g63
  (
    n76,
    n14
  );


  buf
  g64
  (
    n79,
    n3
  );


  not
  g65
  (
    KeyWire_0_19,
    n12
  );


  not
  g66
  (
    n88,
    n9
  );


  buf
  g67
  (
    n34,
    n13
  );


  not
  g68
  (
    n50,
    n12
  );


  not
  g69
  (
    n53,
    n10
  );


  buf
  g70
  (
    n52,
    n21
  );


  not
  g71
  (
    n71,
    n12
  );


  not
  g72
  (
    n77,
    n15
  );


  not
  g73
  (
    n51,
    n6
  );


  not
  g74
  (
    n33,
    n16
  );


  not
  g75
  (
    n59,
    n8
  );


  not
  g76
  (
    n94,
    n17
  );


  not
  g77
  (
    n93,
    n22
  );


  buf
  g78
  (
    n143,
    n28
  );


  not
  g79
  (
    n147,
    n61
  );


  not
  g80
  (
    n113,
    n67
  );


  buf
  g81
  (
    n132,
    n44
  );


  not
  g82
  (
    KeyWire_0_12,
    n32
  );


  buf
  g83
  (
    n140,
    n27
  );


  buf
  g84
  (
    n130,
    n43
  );


  not
  g85
  (
    n137,
    n56
  );


  not
  g86
  (
    KeyWire_0_5,
    n70
  );


  not
  g87
  (
    n114,
    n58
  );


  buf
  g88
  (
    n127,
    n64
  );


  not
  g89
  (
    n112,
    n39
  );


  not
  g90
  (
    n104,
    n55
  );


  buf
  g91
  (
    KeyWire_0_1,
    n59
  );


  not
  g92
  (
    n111,
    n36
  );


  buf
  g93
  (
    n148,
    n71
  );


  buf
  g94
  (
    n146,
    n42
  );


  buf
  g95
  (
    n118,
    n30
  );


  buf
  g96
  (
    KeyWire_0_24,
    n34
  );


  not
  g97
  (
    n124,
    n50
  );


  buf
  g98
  (
    n109,
    n48
  );


  not
  g99
  (
    n106,
    n54
  );


  buf
  g100
  (
    n149,
    n33
  );


  not
  g101
  (
    n122,
    n60
  );


  buf
  g102
  (
    n131,
    n35
  );


  not
  g103
  (
    n117,
    n49
  );


  buf
  g104
  (
    n134,
    n46
  );


  not
  g105
  (
    n121,
    n69
  );


  buf
  g106
  (
    n136,
    n37
  );


  not
  g107
  (
    n128,
    n38
  );


  buf
  g108
  (
    n115,
    n29
  );


  buf
  g109
  (
    n150,
    n51
  );


  buf
  g110
  (
    n120,
    n63
  );


  buf
  g111
  (
    n103,
    n68
  );


  buf
  g112
  (
    n116,
    n40
  );


  not
  g113
  (
    n144,
    n31
  );


  buf
  g114
  (
    n142,
    n62
  );


  not
  g115
  (
    n119,
    n52
  );


  not
  g116
  (
    n138,
    n72
  );


  not
  g117
  (
    n139,
    n41
  );


  not
  g118
  (
    n108,
    n26
  );


  buf
  g119
  (
    n141,
    n53
  );


  not
  g120
  (
    n125,
    n65
  );


  buf
  g121
  (
    n133,
    n57
  );


  not
  g122
  (
    n145,
    n25
  );


  not
  g123
  (
    n110,
    n47
  );


  not
  g124
  (
    n129,
    n66
  );


  buf
  g125
  (
    n126,
    n45
  );


  not
  g126
  (
    n153,
    n116
  );


  buf
  g127
  (
    n155,
    n146
  );


  not
  g128
  (
    n172,
    n135
  );


  not
  g129
  (
    n163,
    n124
  );


  not
  g130
  (
    n177,
    n138
  );


  buf
  g131
  (
    n168,
    n137
  );


  buf
  g132
  (
    n179,
    n121
  );


  not
  g133
  (
    n161,
    n148
  );


  not
  g134
  (
    n167,
    n145
  );


  not
  g135
  (
    n176,
    n141
  );


  not
  g136
  (
    KeyWire_0_29,
    n143
  );


  not
  g137
  (
    n152,
    n108
  );


  not
  g138
  (
    n165,
    n139
  );


  not
  g139
  (
    n166,
    n149
  );


  buf
  g140
  (
    n178,
    n127
  );


  buf
  g141
  (
    KeyWire_0_30,
    n128
  );


  not
  g142
  (
    n169,
    n150
  );


  buf
  g143
  (
    n170,
    n133
  );


  not
  g144
  (
    n173,
    n118
  );


  not
  g145
  (
    n159,
    n103
  );


  buf
  g146
  (
    n180,
    n136
  );


  buf
  g147
  (
    n181,
    n140
  );


  buf
  g148
  (
    n156,
    n114
  );


  buf
  g149
  (
    n154,
    n110
  );


  not
  g150
  (
    n164,
    n104
  );


  buf
  g151
  (
    n162,
    n130
  );


  and
  g152
  (
    n160,
    n117,
    n105
  );


  xnor
  g153
  (
    n158,
    n142,
    n144,
    n113,
    n106
  );


  xnor
  g154
  (
    n174,
    n131,
    n123,
    n129,
    n115
  );


  or
  g155
  (
    n171,
    n119,
    n107,
    n125,
    n111
  );


  and
  g156
  (
    n157,
    n126,
    n132,
    n120,
    n147
  );


  and
  g157
  (
    n182,
    n134,
    n109,
    n112,
    n122
  );


  not
  g158
  (
    n197,
    n81
  );


  not
  g159
  (
    n189,
    n175
  );


  buf
  g160
  (
    n192,
    n165
  );


  not
  g161
  (
    n198,
    n172
  );


  not
  g162
  (
    n186,
    n77
  );


  buf
  g163
  (
    n184,
    n75
  );


  buf
  g164
  (
    n195,
    n170
  );


  buf
  g165
  (
    n200,
    n173
  );


  buf
  g166
  (
    n199,
    n171
  );


  buf
  g167
  (
    n193,
    n169
  );


  not
  g168
  (
    n191,
    n174
  );


  not
  g169
  (
    KeyWire_0_28,
    n179
  );


  buf
  g170
  (
    n183,
    n176
  );


  buf
  g171
  (
    n187,
    n167
  );


  nand
  g172
  (
    n196,
    n80,
    n168
  );


  or
  g173
  (
    n188,
    n177,
    n74,
    n79,
    n178
  );


  xnor
  g174
  (
    n185,
    n78,
    n180,
    n76,
    n73
  );


  xor
  g175
  (
    n194,
    n182,
    n166,
    n181,
    n150
  );


  buf
  g176
  (
    n202,
    n188
  );


  buf
  g177
  (
    n210,
    n186
  );


  not
  g178
  (
    n209,
    n189
  );


  buf
  g179
  (
    n203,
    n193
  );


  not
  g180
  (
    n211,
    n192
  );


  buf
  g181
  (
    n205,
    n183
  );


  buf
  g182
  (
    n201,
    n187
  );


  buf
  g183
  (
    KeyWire_0_16,
    n185
  );


  buf
  g184
  (
    n208,
    n191
  );


  not
  g185
  (
    n206,
    n190
  );


  buf
  g186
  (
    n207,
    n184
  );


  buf
  g187
  (
    n222,
    n205
  );


  not
  g188
  (
    n246,
    n201
  );


  buf
  g189
  (
    n252,
    n202
  );


  not
  g190
  (
    n234,
    n209
  );


  buf
  g191
  (
    n244,
    n207
  );


  buf
  g192
  (
    n245,
    n202
  );


  buf
  g193
  (
    n214,
    n202
  );


  not
  g194
  (
    n248,
    n211
  );


  not
  g195
  (
    n243,
    n207
  );


  buf
  g196
  (
    KeyWire_0_31,
    n209
  );


  not
  g197
  (
    n216,
    n194
  );


  not
  g198
  (
    n213,
    n205
  );


  not
  g199
  (
    n219,
    n206
  );


  buf
  g200
  (
    n229,
    n206
  );


  not
  g201
  (
    n237,
    n203
  );


  buf
  g202
  (
    n227,
    n205
  );


  buf
  g203
  (
    n225,
    n207
  );


  not
  g204
  (
    n233,
    n205
  );


  not
  g205
  (
    n242,
    n204
  );


  not
  g206
  (
    n241,
    n206
  );


  not
  g207
  (
    n228,
    n204
  );


  not
  g208
  (
    n236,
    n204
  );


  buf
  g209
  (
    n232,
    n203
  );


  not
  g210
  (
    n253,
    n209
  );


  buf
  g211
  (
    KeyWire_0_23,
    n210
  );


  not
  g212
  (
    n247,
    n207
  );


  not
  g213
  (
    n238,
    n209
  );


  not
  g214
  (
    n239,
    n203
  );


  buf
  g215
  (
    n226,
    n203
  );


  buf
  g216
  (
    n224,
    n206
  );


  not
  g217
  (
    n249,
    n201
  );


  not
  g218
  (
    n212,
    n210
  );


  not
  g219
  (
    n217,
    n208
  );


  buf
  g220
  (
    n230,
    n202
  );


  buf
  g221
  (
    n231,
    n211
  );


  buf
  g222
  (
    n221,
    n208
  );


  not
  g223
  (
    KeyWire_0_7,
    n194
  );


  not
  g224
  (
    n218,
    n208
  );


  not
  g225
  (
    n251,
    n201
  );


  not
  g226
  (
    KeyWire_0_15,
    n204
  );


  not
  g227
  (
    n235,
    n210
  );


  buf
  g228
  (
    n223,
    n210
  );


  buf
  g229
  (
    n240,
    n201
  );


  nor
  g230
  (
    n254,
    n208,
    n211
  );


  buf
  g231
  (
    n260,
    n231
  );


  buf
  g232
  (
    n264,
    n215
  );


  buf
  g233
  (
    n268,
    n224
  );


  not
  g234
  (
    n256,
    n212
  );


  not
  g235
  (
    KeyWire_0_11,
    n226
  );


  buf
  g236
  (
    n262,
    n228
  );


  buf
  g237
  (
    n270,
    n218
  );


  not
  g238
  (
    n257,
    n230
  );


  buf
  g239
  (
    n273,
    n229
  );


  not
  g240
  (
    n272,
    n223
  );


  not
  g241
  (
    KeyWire_0_17,
    n222
  );


  buf
  g242
  (
    n267,
    n225
  );


  not
  g243
  (
    n269,
    n217
  );


  not
  g244
  (
    n271,
    n213
  );


  buf
  g245
  (
    n259,
    n216
  );


  buf
  g246
  (
    n275,
    n221
  );


  buf
  g247
  (
    n261,
    n227
  );


  not
  g248
  (
    KeyWire_0_4,
    n219
  );


  not
  g249
  (
    n263,
    n214
  );


  buf
  g250
  (
    KeyWire_0_9,
    n220
  );


  not
  g251
  (
    n314,
    n263
  );


  buf
  g252
  (
    n288,
    n247
  );


  buf
  g253
  (
    n309,
    n264
  );


  not
  g254
  (
    n319,
    n266
  );


  not
  g255
  (
    n330,
    n253
  );


  buf
  g256
  (
    n303,
    n238
  );


  buf
  g257
  (
    n287,
    n97
  );


  buf
  g258
  (
    n285,
    n264
  );


  not
  g259
  (
    n276,
    n195
  );


  buf
  g260
  (
    n304,
    n83
  );


  buf
  g261
  (
    n298,
    n241
  );


  not
  g262
  (
    KeyWire_0_27,
    n260
  );


  not
  g263
  (
    KeyWire_0_13,
    n244
  );


  buf
  g264
  (
    n317,
    n263
  );


  not
  g265
  (
    n310,
    n254
  );


  buf
  g266
  (
    n333,
    n195
  );


  not
  g267
  (
    n295,
    n246
  );


  buf
  g268
  (
    n318,
    n236
  );


  buf
  g269
  (
    n292,
    n92
  );


  buf
  g270
  (
    n301,
    n265
  );


  buf
  g271
  (
    n323,
    n82
  );


  not
  g272
  (
    n300,
    n196
  );


  buf
  g273
  (
    n279,
    n268
  );


  not
  g274
  (
    n296,
    n263
  );


  not
  g275
  (
    n302,
    n253
  );


  buf
  g276
  (
    n313,
    n253
  );


  not
  g277
  (
    n328,
    n270
  );


  buf
  g278
  (
    n307,
    n259
  );


  buf
  g279
  (
    n311,
    n251
  );


  not
  g280
  (
    n334,
    n271
  );


  buf
  g281
  (
    n327,
    n271
  );


  not
  g282
  (
    n299,
    n245
  );


  not
  g283
  (
    n297,
    n256
  );


  not
  g284
  (
    n290,
    n249
  );


  nor
  g285
  (
    KeyWire_0_6,
    n240,
    n250,
    n272
  );


  xnor
  g286
  (
    n329,
    n266,
    n270,
    n275,
    n249
  );


  nor
  g287
  (
    n332,
    n89,
    n274,
    n242,
    n233
  );


  and
  g288
  (
    n293,
    n272,
    n267,
    n268
  );


  xnor
  g289
  (
    n286,
    n269,
    n252,
    n262,
    n99
  );


  and
  g290
  (
    n322,
    n273,
    n101,
    n196,
    n237
  );


  xnor
  g291
  (
    n321,
    n98,
    n272,
    n95,
    n250
  );


  xor
  g292
  (
    n324,
    n266,
    n264,
    n250,
    n195
  );


  xnor
  g293
  (
    n278,
    n96,
    n274,
    n253
  );


  or
  g294
  (
    n284,
    n197,
    n243,
    n102,
    n195
  );


  xnor
  g295
  (
    n335,
    n271,
    n232,
    n248,
    n252
  );


  nand
  g296
  (
    n289,
    n254,
    n251,
    n258,
    n273
  );


  nor
  g297
  (
    n325,
    n251,
    n100,
    n235,
    n271
  );


  and
  g298
  (
    n316,
    n197,
    n275,
    n250,
    n270
  );


  and
  g299
  (
    n281,
    n265,
    n197,
    n252,
    n251
  );


  nand
  g300
  (
    n312,
    n86,
    n268,
    n267,
    n94
  );


  nor
  g301
  (
    n306,
    n198,
    n196,
    n254,
    n267
  );


  nor
  g302
  (
    KeyWire_0_0,
    n257,
    n249,
    n93
  );


  xor
  g303
  (
    n305,
    n269,
    n263,
    n90,
    n275
  );


  xor
  g304
  (
    n331,
    n88,
    n265,
    n274,
    n239
  );


  or
  g305
  (
    n282,
    n262,
    n84,
    n85,
    n273
  );


  and
  g306
  (
    n326,
    n194,
    n261,
    n197,
    n264
  );


  nor
  g307
  (
    n294,
    n254,
    n196,
    n267,
    n265
  );


  xnor
  g308
  (
    n291,
    n275,
    n273,
    n252,
    n87
  );


  and
  g309
  (
    n280,
    n91,
    n266,
    n198,
    n270
  );


  nor
  g310
  (
    n308,
    n234,
    n194,
    n269
  );


  nor
  g311
  (
    n368,
    n330,
    n306,
    n326,
    n329
  );


  nor
  g312
  (
    n362,
    n295,
    n317,
    n298,
    n324
  );


  and
  g313
  (
    n364,
    n276,
    n286,
    n298,
    n310
  );


  nor
  g314
  (
    n386,
    n333,
    n288,
    n311,
    n322
  );


  xor
  g315
  (
    n338,
    n303,
    n286,
    n294
  );


  xnor
  g316
  (
    KeyWire_0_20,
    n312,
    n329,
    n299,
    n327
  );


  nand
  g317
  (
    n346,
    n323,
    n291,
    n320,
    n328
  );


  xnor
  g318
  (
    n347,
    n279,
    n296,
    n331,
    n310
  );


  and
  g319
  (
    n383,
    n321,
    n302,
    n255,
    n287
  );


  nor
  g320
  (
    n337,
    n305,
    n291,
    n328,
    n325
  );


  xor
  g321
  (
    n387,
    n327,
    n287,
    n295,
    n302
  );


  and
  g322
  (
    KeyWire_0_3,
    n295,
    n332,
    n322,
    n282
  );


  nor
  g323
  (
    KeyWire_0_21,
    n312,
    n285,
    n280,
    n325
  );


  xnor
  g324
  (
    n372,
    n323,
    n320,
    n307,
    n335
  );


  xor
  g325
  (
    n370,
    n324,
    n319,
    n301,
    n289
  );


  or
  g326
  (
    n391,
    n314,
    n299,
    n305,
    n278
  );


  nor
  g327
  (
    KeyWire_0_2,
    n286,
    n317,
    n303,
    n324
  );


  nand
  g328
  (
    n361,
    n306,
    n290,
    n281
  );


  and
  g329
  (
    n341,
    n284,
    n325,
    n301,
    n320
  );


  xnor
  g330
  (
    n376,
    n311,
    n314,
    n302,
    n307
  );


  nand
  g331
  (
    n379,
    n304,
    n329,
    n293,
    n294
  );


  xnor
  g332
  (
    n351,
    n321,
    n292,
    n313,
    n332
  );


  xnor
  g333
  (
    n373,
    n335,
    n308,
    n333,
    n316
  );


  xnor
  g334
  (
    n381,
    n324,
    n289,
    n316,
    n293
  );


  nand
  g335
  (
    n336,
    n327,
    n305,
    n283,
    n322
  );


  xor
  g336
  (
    n390,
    n307,
    n299,
    n301,
    n288
  );


  xor
  g337
  (
    n354,
    n334,
    n255,
    n294,
    n331
  );


  and
  g338
  (
    n340,
    n298,
    n300,
    n332,
    n296
  );


  nand
  g339
  (
    n343,
    n335,
    n331,
    n297,
    n289
  );


  nand
  g340
  (
    n350,
    n317,
    n24,
    n286,
    n314
  );


  nor
  g341
  (
    n366,
    n284,
    n313,
    n307,
    n323
  );


  nand
  g342
  (
    n382,
    n317,
    n326,
    n303,
    n318
  );


  xnor
  g343
  (
    n344,
    n297,
    n296,
    n283,
    n295
  );


  xor
  g344
  (
    n380,
    n292,
    n309,
    n308,
    n24
  );


  xor
  g345
  (
    n357,
    n288,
    n291,
    n293,
    n304
  );


  nor
  g346
  (
    n359,
    n312,
    n318,
    n292,
    n255
  );


  xnor
  g347
  (
    KeyWire_0_25,
    n311,
    n316,
    n321
  );


  xnor
  g348
  (
    n375,
    n285,
    n315,
    n319,
    n331
  );


  nand
  g349
  (
    n339,
    n304,
    n313,
    n287,
    n308
  );


  xor
  g350
  (
    n367,
    n326,
    n292,
    n330,
    n300
  );


  xor
  g351
  (
    n358,
    n332,
    n309,
    n306,
    n334
  );


  nor
  g352
  (
    n374,
    n319,
    n300,
    n310,
    n277
  );


  nand
  g353
  (
    n352,
    n334,
    n297,
    n301,
    n325
  );


  and
  g354
  (
    n389,
    n24,
    n318,
    n315,
    n291
  );


  or
  g355
  (
    n384,
    n308,
    n288,
    n289,
    n328
  );


  xnor
  g356
  (
    n353,
    n297,
    n330,
    n309,
    n290
  );


  nand
  g357
  (
    n355,
    n296,
    n305,
    n309,
    n313
  );


  and
  g358
  (
    n369,
    n328,
    n300,
    n24,
    n326
  );


  and
  g359
  (
    n388,
    n303,
    n285,
    n333,
    n293
  );


  and
  g360
  (
    n371,
    n323,
    n23,
    n298,
    n304
  );


  xor
  g361
  (
    n356,
    n299,
    n334,
    n318,
    n330
  );


  and
  g362
  (
    n377,
    n320,
    n333,
    n287,
    n329
  );


  nand
  g363
  (
    n385,
    n335,
    n255,
    n312,
    n315
  );


  and
  g364
  (
    n349,
    n322,
    n314,
    n310,
    n315
  );


  xor
  g365
  (
    n365,
    n302,
    n290,
    n327,
    n306
  );


  xor
  g366
  (
    n345,
    n319,
    n311,
    n316,
    n285
  );


  or
  g367
  (
    n399,
    n345,
    n364,
    n360,
    n377
  );


  or
  g368
  (
    n392,
    n337,
    n378,
    n340,
    n344
  );


  nand
  g369
  (
    n401,
    n356,
    n341,
    n389,
    n384
  );


  xnor
  g370
  (
    n405,
    n370,
    n348,
    n358,
    n373
  );


  nor
  g371
  (
    n403,
    n379,
    n359,
    n390,
    n363
  );


  xnor
  g372
  (
    n398,
    n346,
    n380,
    n342,
    n367
  );


  nand
  g373
  (
    n397,
    n355,
    n374,
    n383,
    n369
  );


  nor
  g374
  (
    n393,
    n339,
    n354,
    n361,
    n382
  );


  nand
  g375
  (
    KeyWire_0_8,
    n388,
    n347,
    n357,
    n336
  );


  and
  g376
  (
    KeyWire_0_26,
    n385,
    n343,
    n349,
    n387
  );


  nand
  g377
  (
    n402,
    n368,
    n352,
    n350,
    n386
  );


  nand
  g378
  (
    n396,
    n372,
    n375,
    n366,
    n353
  );


  or
  g379
  (
    n400,
    n338,
    n362,
    n351,
    n365
  );


  xnor
  g380
  (
    n395,
    n371,
    n376,
    n381,
    n391
  );


  and
  g381
  (
    n409,
    n394,
    n402,
    n200,
    n395
  );


  or
  g382
  (
    n408,
    n401,
    n200,
    n199,
    n403
  );


  and
  g383
  (
    n411,
    n397,
    n393,
    n392,
    n198
  );


  nor
  g384
  (
    n407,
    n200,
    n396,
    n199,
    n404
  );


  and
  g385
  (
    n410,
    n198,
    n199,
    n200,
    n398
  );


  nor
  g386
  (
    n406,
    n199,
    n399,
    n405,
    n400
  );


  xor
  KeyGate_0_0
  (
    n283,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n105,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n363,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n378,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n258,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n135,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n277,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n250,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n404,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n274,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n80,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n266,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n107,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n315,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n90,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n220,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n204,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n265,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n58,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n101,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n348,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n342,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n82,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n255,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n123,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n360,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n394,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n320,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n190,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n175,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n151,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n215,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

