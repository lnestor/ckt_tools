// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1071_333 written by SynthGen on 2021/05/24 19:42:16
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1071_333 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52,
 n358, n361, n340, n360, n355, n345, n338, n362,
 n356, n335, n353, n359, n354, n1004, n1070, n1059,
 n1056, n1053, n1060, n1062, n1057, n1052, n1071, n1072,
 n1058, n1055, n1073, n1065, n1061, n1074, n1063, n1114,
 n1092, n1093, n1107, n1102, n1113, n1105, n1120, n1094,
 n1121, n1098, n1104, n1116, n1101, n1112, n1119, n1097,
 n1118, n1110, n1103, n1095, n1123, n1100, n1117, n1111,
 n1109, n1099, n1096, n1106, n1115, n1108, n1122);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52;

output n358, n361, n340, n360, n355, n345, n338, n362,
 n356, n335, n353, n359, n354, n1004, n1070, n1059,
 n1056, n1053, n1060, n1062, n1057, n1052, n1071, n1072,
 n1058, n1055, n1073, n1065, n1061, n1074, n1063, n1114,
 n1092, n1093, n1107, n1102, n1113, n1105, n1120, n1094,
 n1121, n1098, n1104, n1116, n1101, n1112, n1119, n1097,
 n1118, n1110, n1103, n1095, n1123, n1100, n1117, n1111,
 n1109, n1099, n1096, n1106, n1115, n1108, n1122;

wire n53, n54, n55, n56, n57, n58, n59, n60,
 n61, n62, n63, n64, n65, n66, n67, n68,
 n69, n70, n71, n72, n73, n74, n75, n76,
 n77, n78, n79, n80, n81, n82, n83, n84,
 n85, n86, n87, n88, n89, n90, n91, n92,
 n93, n94, n95, n96, n97, n98, n99, n100,
 n101, n102, n103, n104, n105, n106, n107, n108,
 n109, n110, n111, n112, n113, n114, n115, n116,
 n117, n118, n119, n120, n121, n122, n123, n124,
 n125, n126, n127, n128, n129, n130, n131, n132,
 n133, n134, n135, n136, n137, n138, n139, n140,
 n141, n142, n143, n144, n145, n146, n147, n148,
 n149, n150, n151, n152, n153, n154, n155, n156,
 n157, n158, n159, n160, n161, n162, n163, n164,
 n165, n166, n167, n168, n169, n170, n171, n172,
 n173, n174, n175, n176, n177, n178, n179, n180,
 n181, n182, n183, n184, n185, n186, n187, n188,
 n189, n190, n191, n192, n193, n194, n195, n196,
 n197, n198, n199, n200, n201, n202, n203, n204,
 n205, n206, n207, n208, n209, n210, n211, n212,
 n213, n214, n215, n216, n217, n218, n219, n220,
 n221, n222, n223, n224, n225, n226, n227, n228,
 n229, n230, n231, n232, n233, n234, n235, n236,
 n237, n238, n239, n240, n241, n242, n243, n244,
 n245, n246, n247, n248, n249, n250, n251, n252,
 n253, n254, n255, n256, n257, n258, n259, n260,
 n261, n262, n263, n264, n265, n266, n267, n268,
 n269, n270, n271, n272, n273, n274, n275, n276,
 n277, n278, n279, n280, n281, n282, n283, n284,
 n285, n286, n287, n288, n289, n290, n291, n292,
 n293, n294, n295, n296, n297, n298, n299, n300,
 n301, n302, n303, n304, n305, n306, n307, n308,
 n309, n310, n311, n312, n313, n314, n315, n316,
 n317, n318, n319, n320, n321, n322, n323, n324,
 n325, n326, n327, n328, n329, n330, n331, n332,
 n333, n334, n336, n337, n339, n341, n342, n343,
 n344, n346, n347, n348, n349, n350, n351, n352,
 n357, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1054, n1064, n1066, n1067, n1068, n1069, n1075,
 n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
 n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091;

not  g0 (n81, n21);
buf  g1 (n90, n34);
not  g2 (n186, n17);
not  g3 (n131, n27);
not  g4 (n86, n43);
buf  g5 (n75, n35);
buf  g6 (n165, n23);
not  g7 (n118, n37);
buf  g8 (n132, n7);
not  g9 (n217, n41);
buf  g10 (n91, n12);
buf  g11 (n202, n15);
buf  g12 (n181, n33);
buf  g13 (n155, n38);
not  g14 (n211, n17);
buf  g15 (n56, n9);
not  g16 (n218, n46);
not  g17 (n92, n28);
not  g18 (n177, n20);
not  g19 (n68, n27);
not  g20 (n224, n22);
not  g21 (n144, n31);
not  g22 (n72, n16);
not  g23 (n191, n12);
not  g24 (n120, n41);
not  g25 (n114, n17);
not  g26 (n125, n22);
not  g27 (n149, n16);
not  g28 (n195, n41);
buf  g29 (n167, n28);
not  g30 (n89, n34);
not  g31 (n99, n9);
buf  g32 (n200, n42);
buf  g33 (n94, n12);
buf  g34 (n219, n29);
not  g35 (n112, n30);
buf  g36 (n123, n13);
buf  g37 (n192, n31);
not  g38 (n142, n4);
not  g39 (n166, n19);
not  g40 (n203, n4);
not  g41 (n110, n5);
not  g42 (n184, n13);
buf  g43 (n170, n23);
buf  g44 (n182, n18);
not  g45 (n204, n32);
not  g46 (n162, n22);
buf  g47 (n158, n40);
not  g48 (n199, n45);
buf  g49 (n117, n23);
not  g50 (n226, n14);
not  g51 (n212, n42);
buf  g52 (n65, n44);
not  g53 (n220, n35);
buf  g54 (n208, n28);
not  g55 (n95, n47);
not  g56 (n221, n39);
not  g57 (n126, n46);
buf  g58 (n135, n26);
buf  g59 (n215, n18);
buf  g60 (n105, n35);
buf  g61 (n97, n1);
not  g62 (n148, n33);
buf  g63 (n57, n7);
not  g64 (n156, n3);
buf  g65 (n185, n43);
not  g66 (n160, n7);
buf  g67 (n150, n11);
not  g68 (n139, n38);
not  g69 (n198, n25);
not  g70 (n61, n27);
not  g71 (n84, n46);
buf  g72 (n128, n23);
not  g73 (n79, n31);
not  g74 (n176, n9);
not  g75 (n67, n26);
not  g76 (n141, n14);
buf  g77 (n136, n36);
buf  g78 (n80, n1);
buf  g79 (n146, n22);
not  g80 (n213, n24);
not  g81 (n122, n10);
buf  g82 (n71, n6);
not  g83 (n133, n5);
buf  g84 (n147, n34);
buf  g85 (n164, n40);
buf  g86 (n154, n15);
not  g87 (n109, n39);
buf  g88 (n77, n44);
buf  g89 (n159, n33);
buf  g90 (n207, n16);
not  g91 (n223, n18);
buf  g92 (n174, n40);
buf  g93 (n124, n24);
not  g94 (n87, n36);
buf  g95 (n60, n42);
buf  g96 (n134, n39);
not  g97 (n111, n15);
not  g98 (n169, n3);
buf  g99 (n93, n10);
not  g100 (n188, n18);
not  g101 (n103, n19);
buf  g102 (n121, n20);
not  g103 (n171, n32);
buf  g104 (n113, n29);
buf  g105 (n64, n20);
not  g106 (n145, n6);
buf  g107 (n173, n20);
buf  g108 (n175, n33);
buf  g109 (n54, n8);
buf  g110 (n201, n32);
not  g111 (n225, n10);
not  g112 (n190, n8);
not  g113 (n197, n36);
not  g114 (n107, n37);
buf  g115 (n62, n7);
buf  g116 (n161, n25);
buf  g117 (n116, n44);
buf  g118 (n83, n43);
not  g119 (n108, n40);
not  g120 (n187, n21);
not  g121 (n88, n47);
not  g122 (n63, n31);
not  g123 (n209, n38);
buf  g124 (n193, n45);
buf  g125 (n101, n28);
buf  g126 (n102, n43);
not  g127 (n82, n30);
not  g128 (n196, n11);
buf  g129 (n153, n14);
buf  g130 (n168, n24);
buf  g131 (n106, n16);
not  g132 (n73, n30);
buf  g133 (n127, n45);
buf  g134 (n157, n12);
buf  g135 (n137, n32);
not  g136 (n172, n19);
not  g137 (n189, n13);
buf  g138 (n138, n36);
not  g139 (n98, n21);
buf  g140 (n163, n46);
buf  g141 (n70, n26);
buf  g142 (n222, n25);
not  g143 (n151, n29);
buf  g144 (n74, n41);
buf  g145 (n69, n24);
not  g146 (n104, n2);
buf  g147 (n119, n9);
not  g148 (n85, n10);
not  g149 (n115, n15);
buf  g150 (n55, n2);
buf  g151 (n205, n26);
buf  g152 (n58, n39);
buf  g153 (n78, n14);
not  g154 (n129, n44);
buf  g155 (n214, n8);
buf  g156 (n53, n37);
buf  g157 (n76, n29);
buf  g158 (n100, n11);
buf  g159 (n210, n35);
not  g160 (n194, n19);
buf  g161 (n66, n42);
not  g162 (n206, n25);
not  g163 (n143, n11);
not  g164 (n152, n45);
buf  g165 (n178, n38);
buf  g166 (n183, n8);
buf  g167 (n216, n13);
buf  g168 (n130, n34);
not  g169 (n180, n37);
not  g170 (n96, n30);
not  g171 (n59, n21);
buf  g172 (n140, n27);
not  g173 (n179, n17);
buf  g174 (n314, n124);
not  g175 (n301, n121);
buf  g176 (n229, n115);
not  g177 (n275, n71);
buf  g178 (n296, n72);
buf  g179 (n298, n92);
buf  g180 (n260, n106);
buf  g181 (n268, n90);
not  g182 (n321, n110);
buf  g183 (n323, n95);
not  g184 (n262, n120);
not  g185 (n292, n65);
buf  g186 (n289, n87);
buf  g187 (n315, n68);
buf  g188 (n249, n56);
not  g189 (n228, n91);
buf  g190 (n310, n74);
buf  g191 (n328, n83);
buf  g192 (n251, n89);
buf  g193 (n320, n113);
not  g194 (n239, n91);
buf  g195 (n243, n95);
not  g196 (n317, n63);
not  g197 (n327, n92);
buf  g198 (n253, n55);
buf  g199 (n306, n58);
buf  g200 (n265, n103);
buf  g201 (n311, n98);
not  g202 (n264, n122);
not  g203 (n333, n66);
buf  g204 (n303, n79);
not  g205 (n281, n104);
not  g206 (n242, n107);
buf  g207 (n330, n57);
not  g208 (n284, n105);
buf  g209 (n259, n100);
not  g210 (n304, n96);
not  g211 (n232, n111);
not  g212 (n250, n119);
not  g213 (n270, n60);
not  g214 (n247, n125);
not  g215 (n231, n93);
buf  g216 (n300, n73);
not  g217 (n322, n102);
not  g218 (n291, n64);
buf  g219 (n316, n116);
not  g220 (n263, n90);
buf  g221 (n278, n89);
buf  g222 (n283, n107);
buf  g223 (n288, n87);
buf  g224 (n332, n76);
not  g225 (n257, n114);
not  g226 (n307, n67);
not  g227 (n318, n93);
buf  g228 (n258, n112);
not  g229 (n240, n80);
buf  g230 (n234, n99);
not  g231 (n256, n84);
buf  g232 (n241, n113);
not  g233 (n293, n88);
not  g234 (n227, n88);
not  g235 (n271, n105);
not  g236 (n277, n81);
buf  g237 (n269, n69);
not  g238 (n309, n59);
not  g239 (n313, n94);
buf  g240 (n329, n75);
buf  g241 (n245, n77);
buf  g242 (n308, n125);
buf  g243 (n286, n101);
not  g244 (n324, n122);
buf  g245 (n236, n121);
buf  g246 (n279, n61);
not  g247 (n266, n123);
not  g248 (n326, n114);
not  g249 (n261, n70);
buf  g250 (n312, n96);
not  g251 (n287, n62);
buf  g252 (n297, n117);
not  g253 (n280, n119);
buf  g254 (n274, n94);
not  g255 (n267, n106);
not  g256 (n273, n110);
buf  g257 (n255, n116);
not  g258 (n299, n126);
not  g259 (n325, n54);
buf  g260 (n248, n120);
buf  g261 (n331, n97);
not  g262 (n302, n98);
buf  g263 (n246, n118);
buf  g264 (n238, n109);
not  g265 (n334, n53);
buf  g266 (n254, n78);
not  g267 (n285, n123);
buf  g268 (n295, n102);
not  g269 (n244, n101);
buf  g270 (n272, n111);
buf  g271 (n252, n109);
not  g272 (n230, n100);
buf  g273 (n305, n117);
not  g274 (n290, n124);
not  g275 (n282, n97);
not  g276 (n237, n86);
not  g277 (n235, n115);
not  g278 (n294, n99);
buf  g279 (n276, n85);
xnor g280 (n233, n108, n118, n112);
nand g281 (n319, n103, n104, n108, n82);
nor  g282 (n353, n230, n127);
nand g283 (n359, n289, n257, n240, n275);
nor  g284 (n339, n251, n273, n242, n255);
nor  g285 (n362, n303, n295, n282, n228);
or   g286 (n340, n262, n235, n284, n247);
nor  g287 (n360, n241, n298, n261, n297);
nor  g288 (n355, n266, n290, n319, n278);
nor  g289 (n337, n129, n271, n128, n311);
and  g290 (n348, n283, n329, n310, n236);
and  g291 (n346, n245, n127, n288, n231);
xnor g292 (n357, n299, n321, n291, n252);
nor  g293 (n352, n307, n277, n269, n272);
xor  g294 (n341, n315, n300, n265, n246);
nor  g295 (n344, n227, n332, n293, n243);
and  g296 (n350, n233, n308, n260, n232);
and  g297 (n356, n274, n287, n258, n314);
xnor g298 (n361, n254, n267, n305, n244);
nor  g299 (n354, n229, n280, n325, n238);
xor  g300 (n349, n126, n323, n302, n306);
or   g301 (n342, n322, n237, n256, n263);
xor  g302 (n338, n320, n264, n253, n285);
and  g303 (n336, n249, n309, n270, n331);
xor  g304 (n358, n334, n318, n276, n286);
nor  g305 (n347, n326, n301, n294, n328);
or   g306 (n363, n248, n317, n279, n312);
or   g307 (n343, n313, n330, n259, n268);
nor  g308 (n335, n234, n333, n128, n296);
xnor g309 (n345, n250, n292, n316, n239);
xor  g310 (n351, n281, n304, n327, n324);
buf  g311 (n368, n49);
not  g312 (n372, n51);
not  g313 (n370, n358);
not  g314 (n365, n356);
buf  g315 (n367, n50);
xor  g316 (n375, n50, n351);
xnor g317 (n374, n48, n49);
xnor g318 (n364, n48, n47, n348);
nor  g319 (n376, n48, n360, n359);
nand g320 (n371, n354, n50);
xor  g321 (n369, n350, n355, n352);
xnor g322 (n366, n357, n47, n353);
and  g323 (n373, n49, n349, n48);
xnor g324 (n387, n140, n366, n365);
or   g325 (n385, n144, n140, n143, n137);
nor  g326 (n388, n133, n132, n135, n367);
and  g327 (n383, n132, n142, n143, n366);
nor  g328 (n379, n365, n136, n129, n146);
nor  g329 (n386, n145, n364, n131);
and  g330 (n380, n144, n146, n138, n133);
nand g331 (n382, n139, n134, n366, n135);
nand g332 (n381, n130, n139, n142, n136);
or   g333 (n378, n147, n131, n366, n367);
and  g334 (n384, n134, n145, n137, n130);
or   g335 (n377, n365, n141, n138);
buf  g336 (n391, n379);
not  g337 (n393, n380);
not  g338 (n398, n377);
not  g339 (n397, n378);
not  g340 (n392, n378);
buf  g341 (n396, n381);
not  g342 (n390, n379);
not  g343 (n395, n381);
not  g344 (n389, n380);
buf  g345 (n394, n377);
buf  g346 (n400, n362);
not  g347 (n401, n392);
buf  g348 (n402, n361);
and  g349 (n399, n389, n390, n391);
buf  g350 (n406, n400);
not  g351 (n408, n399);
not  g352 (n409, n400);
buf  g353 (n404, n401);
not  g354 (n405, n400);
not  g355 (n407, n399);
not  g356 (n412, n399);
not  g357 (n403, n400);
buf  g358 (n411, n401);
buf  g359 (n410, n399);
not  g360 (n414, n406);
buf  g361 (n422, n404);
buf  g362 (n418, n385);
not  g363 (n417, n404);
buf  g364 (n425, n403);
not  g365 (n427, n403);
not  g366 (n419, n403);
buf  g367 (n426, n383);
not  g368 (n415, n405);
buf  g369 (n421, n403);
buf  g370 (n420, n406);
not  g371 (n413, n404);
nand g372 (n424, n404, n386, n384, n382);
xnor g373 (n416, n385, n405, n406);
nor  g374 (n423, n383, n382, n405, n384);
nor  g375 (n436, n163, n157, n156, n153);
and  g376 (n428, n151, n164, n152, n158);
nand g377 (n431, n150, n155, n413, n152);
xnor g378 (n435, n396, n166, n162);
xor  g379 (n434, n163, n150, n414, n147);
nand g380 (n432, n416, n413, n414, n167);
nor  g381 (n444, n161, n168, n169, n413);
nand g382 (n430, n393, n168, n416, n414);
nand g383 (n440, n154, n157, n415);
and  g384 (n443, n415, n149, n395);
xnor g385 (n439, n165, n161, n414, n167);
xor  g386 (n442, n159, n166, n160, n154);
xnor g387 (n429, n148, n151, n413, n165);
nor  g388 (n437, n416, n155, n160, n417);
xor  g389 (n433, n394, n415, n153, n416);
nand g390 (n441, n398, n148, n164, n158);
nand g391 (n438, n159, n156, n169, n397);
buf  g392 (n446, n433);
buf  g393 (n475, n428);
buf  g394 (n470, n429);
not  g395 (n458, n436);
buf  g396 (n467, n429);
not  g397 (n468, n433);
not  g398 (n478, n435);
not  g399 (n469, n431);
not  g400 (n454, n429);
buf  g401 (n471, n430);
not  g402 (n453, n430);
buf  g403 (n449, n434);
buf  g404 (n477, n434);
buf  g405 (n474, n432);
buf  g406 (n447, n435);
not  g407 (n462, n434);
buf  g408 (n455, n433);
buf  g409 (n459, n430);
not  g410 (n460, n431);
buf  g411 (n451, n401);
buf  g412 (n448, n437);
not  g413 (n464, n432);
buf  g414 (n476, n436);
buf  g415 (n473, n432);
buf  g416 (n456, n431);
not  g417 (n457, n401);
buf  g418 (n465, n402);
buf  g419 (n445, n431);
not  g420 (n472, n436);
not  g421 (n463, n402);
buf  g422 (n452, n429);
not  g423 (n466, n402);
xnor g424 (n461, n430, n435, n433, n402);
nand g425 (n450, n435, n436, n432, n434);
not  g426 (n492, n460);
buf  g427 (n527, n472);
not  g428 (n522, n453);
not  g429 (n520, n462);
not  g430 (n521, n412);
buf  g431 (n496, n477);
buf  g432 (n533, n476);
buf  g433 (n497, n452);
buf  g434 (n498, n463);
buf  g435 (n529, n412);
buf  g436 (n495, n475);
buf  g437 (n547, n474);
not  g438 (n534, n412);
not  g439 (n523, n410);
not  g440 (n516, n455);
not  g441 (n532, n463);
buf  g442 (n511, n466);
buf  g443 (n528, n451);
not  g444 (n526, n451);
buf  g445 (n517, n464);
buf  g446 (n513, n458);
not  g447 (n536, n409);
buf  g448 (n530, n412);
buf  g449 (n524, n407);
not  g450 (n509, n467);
buf  g451 (n518, n445);
not  g452 (n546, n454);
not  g453 (n541, n407);
not  g454 (n525, n448);
buf  g455 (n499, n457);
not  g456 (n484, n478);
buf  g457 (n551, n462);
buf  g458 (n481, n447);
buf  g459 (n488, n468);
not  g460 (n543, n453);
buf  g461 (n480, n409);
buf  g462 (n519, n408);
not  g463 (n505, n469);
not  g464 (n504, n473);
buf  g465 (n507, n446);
buf  g466 (n514, n471);
not  g467 (n539, n410);
not  g468 (n549, n470);
not  g469 (n537, n410);
buf  g470 (n502, n410);
not  g471 (n506, n458);
buf  g472 (n500, n469);
buf  g473 (n487, n457);
not  g474 (n503, n472);
buf  g475 (n508, n452);
not  g476 (n485, n411);
buf  g477 (n512, n411);
not  g478 (n479, n467);
not  g479 (n542, n406);
not  g480 (n515, n476);
buf  g481 (n548, n459);
buf  g482 (n491, n465);
buf  g483 (n540, n408);
not  g484 (n486, n468);
buf  g485 (n494, n461);
not  g486 (n531, n409);
not  g487 (n483, n477);
buf  g488 (n510, n476);
not  g489 (n482, n475);
nor  g490 (n490, n409, n478);
xor  g491 (n489, n408, n454, n411, n456);
xnor g492 (n493, n466, n464, n407, n470);
or   g493 (n535, n477, n447, n411, n449);
nor  g494 (n550, n460, n474, n450);
nand g495 (n538, n478, n465, n473, n477);
nand g496 (n545, n476, n445, n446, n459);
and  g497 (n544, n407, n449, n461, n455);
xor  g498 (n501, n408, n456, n471, n448);
buf  g499 (n679, n374);
not  g500 (n583, n525);
not  g501 (n556, n506);
buf  g502 (n736, n504);
buf  g503 (n669, n371);
not  g504 (n690, n488);
not  g505 (n732, n502);
not  g506 (n589, n372);
buf  g507 (n705, n424);
not  g508 (n668, n421);
not  g509 (n594, n522);
buf  g510 (n597, n419);
not  g511 (n622, n486);
buf  g512 (n579, n489);
not  g513 (n581, n512);
not  g514 (n719, n523);
not  g515 (n708, n518);
buf  g516 (n649, n370);
not  g517 (n704, n417);
buf  g518 (n738, n523);
buf  g519 (n667, n367);
not  g520 (n695, n524);
buf  g521 (n559, n486);
buf  g522 (n701, n425);
buf  g523 (n682, n482);
buf  g524 (n663, n498);
not  g525 (n716, n369);
buf  g526 (n595, n516);
buf  g527 (n647, n485);
buf  g528 (n602, n482);
buf  g529 (n606, n525);
not  g530 (n684, n51);
not  g531 (n591, n514);
not  g532 (n554, n515);
buf  g533 (n672, n484);
not  g534 (n697, n499);
buf  g535 (n648, n483);
not  g536 (n607, n507);
buf  g537 (n747, n508);
not  g538 (n592, n521);
buf  g539 (n702, n514);
not  g540 (n557, n512);
not  g541 (n715, n485);
buf  g542 (n694, n507);
not  g543 (n641, n375);
not  g544 (n588, n523);
buf  g545 (n689, n505);
buf  g546 (n656, n500);
not  g547 (n565, n526);
buf  g548 (n662, n503);
not  g549 (n564, n525);
not  g550 (n692, n505);
not  g551 (n745, n370);
not  g552 (n660, n495);
buf  g553 (n568, n483);
buf  g554 (n670, n504);
buf  g555 (n737, n513);
not  g556 (n561, n513);
not  g557 (n643, n374);
buf  g558 (n610, n427);
buf  g559 (n553, n482);
buf  g560 (n612, n519);
not  g561 (n666, n512);
not  g562 (n638, n526);
not  g563 (n603, n417);
not  g564 (n575, n487);
not  g565 (n582, n371);
not  g566 (n664, n519);
not  g567 (n744, n506);
buf  g568 (n584, n512);
not  g569 (n593, n495);
buf  g570 (n713, n523);
buf  g571 (n628, n424);
not  g572 (n632, n510);
not  g573 (n640, n524);
not  g574 (n609, n494);
buf  g575 (n634, n370);
not  g576 (n650, n514);
not  g577 (n717, n521);
not  g578 (n600, n527);
not  g579 (n636, n422);
not  g580 (n631, n492);
not  g581 (n651, n486);
buf  g582 (n611, n374);
buf  g583 (n659, n479);
buf  g584 (n567, n479);
buf  g585 (n635, n368);
not  g586 (n637, n420);
not  g587 (n680, n484);
not  g588 (n729, n423);
not  g589 (n639, n484);
not  g590 (n574, n503);
not  g591 (n566, n491);
not  g592 (n655, n524);
not  g593 (n723, n498);
buf  g594 (n601, n499);
buf  g595 (n552, n424);
not  g596 (n710, n490);
buf  g597 (n709, n425);
buf  g598 (n590, n487);
buf  g599 (n735, n480);
not  g600 (n731, n518);
not  g601 (n645, n517);
buf  g602 (n742, n498);
not  g603 (n586, n481);
not  g604 (n711, n502);
buf  g605 (n569, n368);
buf  g606 (n617, n373);
not  g607 (n573, n421);
buf  g608 (n726, n491);
not  g609 (n571, n496);
buf  g610 (n703, n480);
buf  g611 (n721, n485);
buf  g612 (n707, n423);
buf  g613 (n678, n375);
buf  g614 (n706, n490);
not  g615 (n741, n504);
not  g616 (n728, n511);
not  g617 (n677, n501);
buf  g618 (n654, n488);
not  g619 (n714, n499);
buf  g620 (n691, n422);
not  g621 (n587, n516);
not  g622 (n646, n521);
not  g623 (n657, n518);
not  g624 (n661, n418);
buf  g625 (n696, n418);
not  g626 (n621, n506);
not  g627 (n577, n500);
buf  g628 (n722, n509);
not  g629 (n739, n503);
buf  g630 (n720, n527);
buf  g631 (n683, n498);
buf  g632 (n674, n490);
buf  g633 (n626, n516);
not  g634 (n743, n419);
buf  g635 (n576, n522);
buf  g636 (n693, n509);
buf  g637 (n700, n481);
buf  g638 (n653, n495);
not  g639 (n624, n497);
not  g640 (n676, n501);
not  g641 (n604, n426);
not  g642 (n681, n526);
buf  g643 (n699, n369);
buf  g644 (n608, n525);
buf  g645 (n652, n519);
not  g646 (n630, n504);
not  g647 (n614, n492);
not  g648 (n616, n516);
not  g649 (n740, n502);
not  g650 (n688, n491);
buf  g651 (n633, n493);
not  g652 (n727, n426);
not  g653 (n733, n509);
buf  g654 (n725, n519);
buf  g655 (n734, n421);
buf  g656 (n730, n427);
buf  g657 (n686, n483);
buf  g658 (n665, n510);
not  g659 (n599, n511);
not  g660 (n625, n493);
buf  g661 (n555, n499);
buf  g662 (n558, n375);
buf  g663 (n642, n508);
buf  g664 (n658, n488);
buf  g665 (n580, n372);
not  g666 (n629, n495);
not  g667 (n644, n368);
buf  g668 (n578, n522);
nor  g669 (n746, n487, n487, n505, n501);
xor  g670 (n675, n518, n421, n493, n484);
nand g671 (n619, n419, n520, n508, n506);
nor  g672 (n687, n372, n427, n502, n492);
and  g673 (n718, n481, n522, n427, n510);
xnor g674 (n724, n486, n520, n524, n420);
xnor g675 (n671, n493, n371, n425, n419);
xor  g676 (n605, n526, n510, n485, n491);
nor  g677 (n623, n511, n511, n501, n517);
xor  g678 (n615, n503, n515, n423, n418);
xor  g679 (n712, n497, n521, n368, n492);
nand g680 (n618, n508, n370, n488, n509);
and  g681 (n620, n424, n373, n507, n482);
xnor g682 (n563, n517, n496, n515, n373);
xor  g683 (n585, n423, n514, n479, n494);
xnor g684 (n685, n520, n527, n417, n422);
xor  g685 (n698, n489, n372, n527, n497);
xnor g686 (n570, n373, n418, n479, n481);
nor  g687 (n596, n489, n515, n500, n367);
and  g688 (n562, n513, n507, n489, n490);
nand g689 (n572, n480, n420, n425, n375);
nor  g690 (n673, n494, n497, n369, n420);
or   g691 (n560, n513, n422, n505, n426);
and  g692 (n598, n520, n496, n500);
xor  g693 (n627, n369, n517, n494, n426);
nand g694 (n613, n374, n480, n371, n483);
buf  g695 (n748, n556);
not  g696 (n753, n552);
not  g697 (n749, n555);
not  g698 (n751, n557);
not  g699 (n754, n553);
and  g700 (n750, n552, n554, n556);
nor  g701 (n752, n557, n555, n553, n554);
not  g702 (n761, n561);
nor  g703 (n762, n564, n748, n562);
or   g704 (n755, n558, n753, n566, n750);
nand g705 (n757, n752, n478, n564, n565);
nor  g706 (n759, n563, n559, n562, n565);
xor  g707 (n756, n560, n563, n754, n561);
and  g708 (n760, n170, n560, n559, n558);
nor  g709 (n758, n566, n751, n749, n754);
xnor g710 (n791, n538, n541, n551, n542);
xor  g711 (n780, n544, n543, n529, n539);
nor  g712 (n764, n759, n755, n533, n535);
xnor g713 (n766, n758, n539, n550, n551);
nand g714 (n786, n761, n534, n536, n539);
xor  g715 (n788, n755, n757, n529, n538);
xor  g716 (n768, n760, n550, n545, n759);
xnor g717 (n785, n548, n545, n536, n538);
xnor g718 (n763, n547, n755, n530, n535);
nand g719 (n772, n534, n546, n544, n759);
or   g720 (n783, n548, n756, n541);
and  g721 (n767, n543, n756, n544, n530);
and  g722 (n787, n543, n528, n760, n762);
or   g723 (n776, n757, n540, n543, n551);
nor  g724 (n765, n535, n540, n545, n528);
xor  g725 (n774, n529, n549, n542, n537);
or   g726 (n770, n762, n548, n547, n758);
nor  g727 (n781, n531, n762, n542, n540);
and  g728 (n775, n761, n756, n528, n546);
and  g729 (n784, n547, n544, n755, n546);
and  g730 (n779, n550, n528, n761);
xor  g731 (n773, n538, n530, n535, n551);
nand g732 (n794, n760, n757, n541, n547);
and  g733 (n771, n529, n534, n542, n545);
xnor g734 (n793, n536, n537, n532, n533);
or   g735 (n778, n533, n762, n758, n757);
xnor g736 (n782, n532, n534, n531);
xor  g737 (n792, n531, n530, n760, n532);
xnor g738 (n789, n537, n541, n549, n536);
nand g739 (n790, n550, n759, n532, n533);
or   g740 (n777, n758, n539, n546, n549);
nor  g741 (n769, n537, n549, n548, n540);
not  g742 (n810, n780);
buf  g743 (n801, n570);
buf  g744 (n814, n568);
not  g745 (n804, n569);
buf  g746 (n796, n766);
not  g747 (n809, n773);
buf  g748 (n808, n764);
buf  g749 (n813, n779);
not  g750 (n795, n780);
not  g751 (n798, n778);
not  g752 (n812, n765);
not  g753 (n797, n569);
not  g754 (n802, n567);
not  g755 (n803, n567);
not  g756 (n811, n568);
not  g757 (n805, n767);
buf  g758 (n799, n781);
not  g759 (n806, n768);
xor  g760 (n800, n777, n770);
nor  g761 (n807, n763, n771, n769, n772);
nor  g762 (n815, n774, n775, n776, n779);
xnor g763 (n820, n171, n212, n196, n800);
xnor g764 (n853, n797, n796, n191);
and  g765 (n847, n215, n193, n206);
xor  g766 (n838, n174, n203, n216, n795);
xor  g767 (n842, n799, n575, n800, n796);
nand g768 (n849, n216, n185, n173, n573);
nor  g769 (n827, n217, n804, n226, n225);
nor  g770 (n817, n207, n191, n209, n176);
nand g771 (n856, n571, n795, n192, n179);
xor  g772 (n816, n223, n204, n209, n193);
xor  g773 (n852, n183, n201, n204, n197);
or   g774 (n846, n184, n210, n219, n187);
xor  g775 (n841, n182, n798, n217, n223);
nor  g776 (n843, n179, n576, n186, n220);
and  g777 (n833, n180, n805, n226, n804);
and  g778 (n826, n800, n207, n225, n574);
nor  g779 (n857, n796, n214, n181, n196);
nand g780 (n854, n577, n214, n799, n194);
nor  g781 (n850, n213, n186, n202, n578);
nor  g782 (n819, n195, n208, n804, n220);
nand g783 (n845, n570, n195, n221, n175);
and  g784 (n823, n218, n575, n572, n221);
or   g785 (n839, n797, n571, n218, n574);
xor  g786 (n822, n205, n801, n188);
and  g787 (n837, n198, n177, n170, n224);
nor  g788 (n818, n181, n212, n172, n798);
xnor g789 (n825, n798, n222, n803, n573);
and  g790 (n832, n802, n205, n219, n190);
or   g791 (n831, n199, n189, n187, n201);
nand g792 (n844, n199, n211, n215, n801);
xor  g793 (n855, n178, n224, n797, n184);
and  g794 (n828, n176, n222, n572, n194);
or   g795 (n858, n211, n797, n803, n802);
xnor g796 (n829, n175, n171, n182, n801);
and  g797 (n840, n803, n197, n208, n189);
or   g798 (n821, n210, n803, n576, n795);
nor  g799 (n836, n802, n190, n178, n577);
or   g800 (n835, n798, n200, n802);
nor  g801 (n834, n174, n173, n801, n198);
or   g802 (n848, n795, n800, n172, n799);
xnor g803 (n824, n202, n192, n177, n180);
nand g804 (n851, n185, n805, n183, n203);
xor  g805 (n830, n213, n805, n804, n799);
buf  g806 (n863, n819);
buf  g807 (n859, n828);
not  g808 (n861, n822);
buf  g809 (n862, n817);
buf  g810 (n860, n51);
xnor g811 (n866, n827, n52, n826);
nor  g812 (n864, n818, n816, n825, n821);
xnor g813 (n865, n824, n823, n51, n820);
and  g814 (n871, n579, n860, n863, n792);
xnor g815 (n874, n794, n861, n782);
nor  g816 (n873, n794, n792, n793, n784);
nor  g817 (n870, n785, n783, n790, n863);
xor  g818 (n872, n862, n859, n788, n789);
xor  g819 (n869, n786, n793, n781, n784);
or   g820 (n875, n860, n859, n791, n787);
or   g821 (n867, n788, n791, n862, n789);
nor  g822 (n868, n787, n785, n861, n578);
and  g823 (n876, n579, n790, n786, n783);
xnor g824 (n888, n814, n870, n583, n875);
nor  g825 (n887, n806, n585, n813, n808);
nand g826 (n878, n809, n876, n807, n814);
nor  g827 (n893, n873, n811, n812, n809);
and  g828 (n882, n584, n586, n815);
nor  g829 (n889, n585, n868, n813);
xnor g830 (n883, n580, n807, n869, n876);
nand g831 (n886, n815, n811, n874, n867);
nor  g832 (n881, n810, n810, n815, n808);
xor  g833 (n890, n809, n875, n874, n807);
or   g834 (n880, n810, n814, n582, n807);
xor  g835 (n885, n872, n580, n805, n871);
and  g836 (n879, n806, n873, n581, n871);
nor  g837 (n892, n808, n808, n582, n869);
nand g838 (n877, n583, n812, n810);
or   g839 (n891, n811, n581, n806, n813);
and  g840 (n884, n870, n584, n809, n814);
xnor g841 (n894, n872, n812, n811, n806);
nor  g842 (n921, n882, n598, n596, n884);
or   g843 (n943, n656, n879, n659);
nand g844 (n932, n847, n625, n631, n637);
xor  g845 (n896, n620, n609, n832, n660);
and  g846 (n942, n625, n888, n635, n894);
nand g847 (n908, n617, n663, n590, n636);
xnor g848 (n945, n650, n892, n669, n656);
nor  g849 (n963, n889, n884, n586, n599);
xnor g850 (n901, n631, n661, n880, n842);
and  g851 (n922, n880, n657, n605, n626);
xnor g852 (n931, n632, n882, n619, n603);
xnor g853 (n937, n587, n649, n668, n597);
and  g854 (n903, n597, n890, n637, n883);
or   g855 (n965, n604, n880, n611, n881);
and  g856 (n899, n670, n851, n622, n882);
xor  g857 (n957, n830, n659, n652, n878);
xor  g858 (n898, n881, n651, n878, n890);
or   g859 (n920, n894, n837, n600, n886);
and  g860 (n948, n833, n593, n849, n630);
nand g861 (n952, n849, n642, n622, n893);
nand g862 (n918, n601, n885, n612, n610);
nand g863 (n900, n846, n852, n626, n666);
nor  g864 (n964, n606, n592, n588, n621);
xor  g865 (n905, n884, n891, n646, n605);
xnor g866 (n930, n891, n665, n877, n842);
nand g867 (n923, n623, n669, n643, n640);
nor  g868 (n949, n654, n604, n594, n613);
and  g869 (n958, n607, n628, n632, n655);
xnor g870 (n929, n840, n846, n589, n606);
or   g871 (n961, n608, n848, n850, n645);
nand g872 (n924, n589, n641, n613, n834);
xor  g873 (n928, n841, n829, n616, n591);
and  g874 (n950, n599, n612, n661, n630);
nand g875 (n960, n835, n670, n624, n843);
or   g876 (n966, n633, n884, n878, n837);
or   g877 (n935, n590, n840, n648, n608);
xor  g878 (n944, n888, n634, n838, n835);
xnor g879 (n959, n614, n883, n587, n888);
xor  g880 (n940, n880, n618, n892);
nor  g881 (n946, n651, n894, n889, n847);
xnor g882 (n912, n883, n643, n641, n607);
or   g883 (n926, n595, n889, n891, n666);
nand g884 (n915, n640, n636, n893, n885);
and  g885 (n925, n662, n883, n600, n592);
nand g886 (n910, n639, n644, n629, n619);
or   g887 (n941, n888, n617, n658, n645);
and  g888 (n916, n646, n634, n653, n844);
or   g889 (n954, n887, n594, n662, n881);
and  g890 (n953, n664, n660, n596, n879);
nand g891 (n936, n602, n887, n663, n603);
or   g892 (n927, n839, n650, n892, n618);
or   g893 (n938, n602, n621, n639, n889);
xor  g894 (n933, n610, n667, n629);
xor  g895 (n895, n886, n839, n593, n668);
nor  g896 (n934, n615, n638, n623, n614);
nand g897 (n939, n653, n893, n624, n894);
nand g898 (n907, n655, n627, n595, n845);
nand g899 (n897, n834, n890, n844, n601);
xor  g900 (n955, n620, n628, n654, n881);
nor  g901 (n962, n588, n887, n879, n882);
nor  g902 (n902, n836, n635, n886, n831);
xor  g903 (n919, n885, n838, n831, n609);
nor  g904 (n956, n648, n833, n611, n843);
nor  g905 (n917, n633, n845, n644, n591);
and  g906 (n947, n598, n878, n830, n638);
nand g907 (n951, n848, n657, n649, n877);
xnor g908 (n906, n851, n665, n877, n829);
and  g909 (n909, n658, n647, n885, n615);
nand g910 (n913, n877, n647, n891, n850);
and  g911 (n914, n616, n890, n832, n841);
xor  g912 (n904, n836, n627, n887, n652);
xnor g913 (n911, n664, n893, n642, n886);
buf  g914 (n990, n898);
not  g915 (n972, n900);
not  g916 (n967, n918);
buf  g917 (n974, n916);
buf  g918 (n975, n912);
not  g919 (n991, n917);
not  g920 (n988, n922);
buf  g921 (n977, n914);
buf  g922 (n982, n906);
not  g923 (n968, n903);
buf  g924 (n978, n899);
buf  g925 (n970, n919);
buf  g926 (n969, n897);
buf  g927 (n987, n907);
not  g928 (n994, n913);
not  g929 (n980, n910);
not  g930 (n986, n904);
not  g931 (n973, n908);
buf  g932 (n983, n901);
buf  g933 (n976, n902);
buf  g934 (n985, n896);
buf  g935 (n984, n915);
buf  g936 (n981, n905);
not  g937 (n993, n895);
not  g938 (n989, n909);
buf  g939 (n971, n911);
buf  g940 (n979, n920);
buf  g941 (n992, n921);
xor  g942 (n1004, n970, n982, n441, n437);
or   g943 (n1007, n387, n438, n439, n437);
or   g944 (n1002, n441, n443, n967, n439);
xor  g945 (n1009, n438, n994, n442);
nor  g946 (n997, n440, n439, n443, n444);
xor  g947 (n1012, n974, n989, n986, n981);
xor  g948 (n999, n993, n972, n439, n437);
and  g949 (n1003, n991, n442, n976, n444);
or   g950 (n1005, n442, n968, n388, n985);
nor  g951 (n1006, n988, n991, n984, n388);
xnor g952 (n996, n438, n441, n977, n993);
xnor g953 (n995, n992, n969, n443, n990);
nor  g954 (n998, n973, n978, n983, n438);
or   g955 (n1001, n992, n979, n987, n923);
nor  g956 (n1011, n440, n994, n989, n386);
xnor g957 (n1010, n387, n975, n443, n671);
nor  g958 (n1000, n671, n444, n980, n440);
xor  g959 (n1008, n440, n971, n441, n990);
xor  g960 (n1023, n1006, n855, n1001, n376);
or   g961 (n1013, n856, n855, n927, n940);
xnor g962 (n1016, n933, n376, n931, n924);
xnor g963 (n1025, n998, n997, n852, n1008);
nand g964 (n1015, n1003, n929, n376);
and  g965 (n1021, n935, n853, n363, n947);
nand g966 (n1020, n856, n925, n936, n854);
and  g967 (n1022, n1007, n943, n854, n1002);
or   g968 (n1018, n937, n945, n672, n996);
or   g969 (n1024, n942, n939, n1009, n1000);
nor  g970 (n1017, n938, n932, n672, n946);
nand g971 (n1026, n857, n999, n944, n928);
nand g972 (n1014, n941, n1004, n948, n1005);
nand g973 (n1019, n930, n934, n853, n926);
xnor g974 (n1027, n959, n1014, n960, n954);
xnor g975 (n1030, n1013, n956, n950, n1014);
xor  g976 (n1028, n952, n1013, n949, n953);
xor  g977 (n1029, n951, n955, n957, n958);
not  g978 (n1034, n1028);
buf  g979 (n1033, n673);
xnor g980 (n1031, n674, n673);
nor  g981 (n1032, n674, n1027);
not  g982 (n1045, n866);
buf  g983 (n1050, n52);
buf  g984 (n1038, n388);
buf  g985 (n1037, n1033);
buf  g986 (n1035, n858);
and  g987 (n1046, n866, n961, n1033);
and  g988 (n1041, n866, n1032, n388, n1034);
xnor g989 (n1047, n1031, n865, n1010);
xnor g990 (n1040, n963, n858, n864, n1012);
xnor g991 (n1048, n1031, n865, n864, n52);
nor  g992 (n1044, n1034, n965, n1032, n864);
xor  g993 (n1042, n863, n1033, n964);
xor  g994 (n1036, n1034, n857, n962, n1031);
nand g995 (n1043, n444, n1031, n1032, n1011);
or   g996 (n1049, n1032, n52, n1034, n863);
nor  g997 (n1039, n866, n865, n966, n864);
or   g998 (n1061, n1043, n690, n682);
xor  g999 (n1074, n1035, n1018, n1026, n1022);
xor  g1000 (n1054, n676, n1042, n1020, n677);
xnor g1001 (n1053, n1025, n685, n1021, n1044);
nand g1002 (n1057, n1019, n1044, n1049, n1020);
nand g1003 (n1051, n680, n1050, n682);
nor  g1004 (n1065, n681, n1018, n1025, n1047);
xnor g1005 (n1058, n1020, n683, n686, n1024);
xnor g1006 (n1067, n1020, n676, n686, n1017);
or   g1007 (n1068, n689, n1017, n1025, n675);
or   g1008 (n1066, n679, n1026, n1023, n1038);
nand g1009 (n1052, n1025, n1046, n1048, n1024);
nand g1010 (n1060, n1024, n1021, n1022);
and  g1011 (n1064, n1015, n683, n1023, n1049);
xnor g1012 (n1070, n687, n1019, n1015, n1023);
or   g1013 (n1062, n1037, n1021, n689, n688);
or   g1014 (n1072, n1040, n1047, n1023, n679);
or   g1015 (n1056, n677, n1043, n1016, n1045);
nor  g1016 (n1055, n691, n1026, n684, n688);
or   g1017 (n1069, n1048, n685, n1026, n678);
nand g1018 (n1059, n684, n1021, n1022, n1036);
nand g1019 (n1063, n691, n681, n687, n675);
xnor g1020 (n1071, n1041, n1016, n1024, n1039);
and  g1021 (n1073, n1046, n678, n1045, n680);
nand g1022 (n1075, n693, n695, n1029, n1028);
nand g1023 (n1077, n1072, n1030, n1028, n696);
xor  g1024 (n1076, n693, n1074, n1030, n1071);
xnor g1025 (n1081, n1073, n694, n692, n695);
or   g1026 (n1080, n1069, n694, n692, n1028);
nor  g1027 (n1079, n1030, n1030, n1070, n696);
xnor g1028 (n1078, n1068, n1029);
not  g1029 (n1083, n1075);
not  g1030 (n1082, n1075);
xor  g1031 (n1091, n702, n707, n1082, n705);
nor  g1032 (n1087, n700, n1083, n701, n704);
or   g1033 (n1088, n698, n704, n701, n699);
and  g1034 (n1086, n1083, n1082, n706);
nand g1035 (n1085, n700, n707, n697, n699);
nand g1036 (n1084, n708, n703, n697);
and  g1037 (n1089, n702, n1082, n708, n705);
or   g1038 (n1090, n698, n706, n1083);
xnor g1039 (n1110, n1085, n712, n741, n1090);
and  g1040 (n1103, n729, n718, n736, n745);
nand g1041 (n1092, n1085, n732, n731, n1076);
xnor g1042 (n1111, n745, n719, n1081, n1078);
xor  g1043 (n1100, n1078, n746, n747, n1091);
nor  g1044 (n1112, n746, n1081, n727, n738);
nor  g1045 (n1105, n712, n735, n1085, n1077);
xnor g1046 (n1114, n711, n711, n1086, n729);
or   g1047 (n1119, n1088, n715, n1084);
xnor g1048 (n1106, n717, n740, n1089, n731);
nand g1049 (n1104, n1087, n1091, n1089, n1084);
or   g1050 (n1120, n1086, n1080, n737, n747);
xnor g1051 (n1109, n718, n710, n744);
or   g1052 (n1122, n728, n733, n1086);
xor  g1053 (n1097, n742, n713, n734, n730);
xnor g1054 (n1101, n717, n1091, n716, n724);
xnor g1055 (n1094, n1091, n726, n734, n1077);
nand g1056 (n1116, n1076, n742, n730, n728);
xor  g1057 (n1115, n1089, n741, n721, n1090);
xnor g1058 (n1118, n1088, n716, n723, n714);
xor  g1059 (n1095, n1087, n1086, n1081, n710);
and  g1060 (n1096, n721, n713, n738, n1090);
and  g1061 (n1098, n719, n743, n1079);
or   g1062 (n1108, n709, n714, n720, n1085);
nor  g1063 (n1107, n746, n724, n723, n737);
or   g1064 (n1123, n722, n740, n735, n732);
or   g1065 (n1113, n722, n1084, n746, n747);
or   g1066 (n1102, n1080, n743, n747, n720);
and  g1067 (n1121, n1087, n736, n1089, n1090);
xnor g1068 (n1099, n715, n739, n1087, n725);
xor  g1069 (n1093, n1088, n727, n726, n709);
xnor g1070 (n1117, n1088, n725, n739, n1081);
endmodule
