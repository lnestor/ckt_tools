

module Stat_2000_203
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1036,
  n1038,
  n1043,
  n1030,
  n1033,
  n1048,
  n1045,
  n1047,
  n1035,
  n1039,
  n1032,
  n1044,
  n1031,
  n1040,
  n1046,
  n1041,
  n1109,
  n1097,
  n1105,
  n1087,
  n1084,
  n1100,
  n1094,
  n1107,
  n1083,
  n2026,
  n2032,
  n2031,
  n2029,
  n2027,
  n2030,
  n2028
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1036;output n1038;output n1043;output n1030;output n1033;output n1048;output n1045;output n1047;output n1035;output n1039;output n1032;output n1044;output n1031;output n1040;output n1046;output n1041;output n1109;output n1097;output n1105;output n1087;output n1084;output n1100;output n1094;output n1107;output n1083;output n2026;output n2032;output n2031;output n2029;output n2027;output n2030;output n2028;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1034;wire n1037;wire n1042;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1085;wire n1086;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1095;wire n1096;wire n1098;wire n1099;wire n1101;wire n1102;wire n1103;wire n1104;wire n1106;wire n1108;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;wire KeyWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyNOTWire_0_35;wire KeyWire_0_36;wire KeyNOTWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyNOTWire_0_57;wire KeyWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyNOTWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    n68,
    n14
  );


  not
  g1
  (
    n114,
    n27
  );


  buf
  g2
  (
    n67,
    n25
  );


  buf
  g3
  (
    n88,
    n31
  );


  buf
  g4
  (
    n36,
    n30
  );


  not
  g5
  (
    n43,
    n28
  );


  buf
  g6
  (
    n78,
    n16
  );


  buf
  g7
  (
    n46,
    n1
  );


  not
  g8
  (
    n83,
    n25
  );


  not
  g9
  (
    n142,
    n6
  );


  buf
  g10
  (
    n94,
    n3
  );


  buf
  g11
  (
    n77,
    n2
  );


  buf
  g12
  (
    n150,
    n6
  );


  not
  g13
  (
    n121,
    n23
  );


  not
  g14
  (
    n47,
    n31
  );


  buf
  g15
  (
    n37,
    n12
  );


  not
  g16
  (
    n74,
    n12
  );


  buf
  g17
  (
    n60,
    n24
  );


  not
  g18
  (
    n117,
    n21
  );


  not
  g19
  (
    n127,
    n24
  );


  buf
  g20
  (
    n58,
    n8
  );


  buf
  g21
  (
    n56,
    n17
  );


  not
  g22
  (
    n124,
    n22
  );


  not
  g23
  (
    KeyWire_0_38,
    n20
  );


  buf
  g24
  (
    n120,
    n22
  );


  buf
  g25
  (
    n138,
    n19
  );


  not
  g26
  (
    n81,
    n27
  );


  buf
  g27
  (
    n84,
    n2
  );


  buf
  g28
  (
    n91,
    n18
  );


  not
  g29
  (
    n133,
    n16
  );


  not
  g30
  (
    n69,
    n12
  );


  not
  g31
  (
    n66,
    n23
  );


  buf
  g32
  (
    n50,
    n9
  );


  buf
  g33
  (
    n100,
    n28
  );


  buf
  g34
  (
    n49,
    n26
  );


  buf
  g35
  (
    n63,
    n23
  );


  buf
  g36
  (
    n147,
    n10
  );


  not
  g37
  (
    n129,
    n5
  );


  not
  g38
  (
    n85,
    n16
  );


  buf
  g39
  (
    n119,
    n6
  );


  not
  g40
  (
    n80,
    n26
  );


  not
  g41
  (
    n72,
    n2
  );


  not
  g42
  (
    n54,
    n20
  );


  buf
  g43
  (
    n86,
    n14
  );


  not
  g44
  (
    n44,
    n3
  );


  buf
  g45
  (
    n134,
    n7
  );


  not
  g46
  (
    n135,
    n6
  );


  not
  g47
  (
    n89,
    n13
  );


  buf
  g48
  (
    n57,
    n5
  );


  buf
  g49
  (
    n33,
    n15
  );


  not
  g50
  (
    n141,
    n13
  );


  not
  g51
  (
    n82,
    n10
  );


  not
  g52
  (
    n149,
    n14
  );


  not
  g53
  (
    n108,
    n4
  );


  not
  g54
  (
    n41,
    n10
  );


  not
  g55
  (
    n35,
    n18
  );


  not
  g56
  (
    n128,
    n13
  );


  not
  g57
  (
    n145,
    n9
  );


  buf
  g58
  (
    n111,
    n29
  );


  buf
  g59
  (
    KeyWire_0_62,
    n31
  );


  not
  g60
  (
    n151,
    n29
  );


  buf
  g61
  (
    n92,
    n1
  );


  not
  g62
  (
    n156,
    n24
  );


  not
  g63
  (
    n146,
    n3
  );


  buf
  g64
  (
    n112,
    n15
  );


  not
  g65
  (
    n93,
    n19
  );


  buf
  g66
  (
    n115,
    n22
  );


  not
  g67
  (
    n87,
    n1
  );


  not
  g68
  (
    n118,
    n4
  );


  buf
  g69
  (
    n122,
    n27
  );


  not
  g70
  (
    n64,
    n11
  );


  buf
  g71
  (
    n132,
    n8
  );


  buf
  g72
  (
    n70,
    n19
  );


  not
  g73
  (
    n104,
    n25
  );


  not
  g74
  (
    n73,
    n24
  );


  buf
  g75
  (
    n155,
    n9
  );


  not
  g76
  (
    n103,
    n25
  );


  not
  g77
  (
    n125,
    n8
  );


  not
  g78
  (
    n79,
    n11
  );


  buf
  g79
  (
    KeyWire_0_23,
    n4
  );


  buf
  g80
  (
    n116,
    n31
  );


  buf
  g81
  (
    n61,
    n10
  );


  buf
  g82
  (
    n53,
    n11
  );


  buf
  g83
  (
    n99,
    n28
  );


  buf
  g84
  (
    n90,
    n15
  );


  not
  g85
  (
    n144,
    n17
  );


  not
  g86
  (
    n113,
    n26
  );


  buf
  g87
  (
    n136,
    n16
  );


  buf
  g88
  (
    n62,
    n13
  );


  not
  g89
  (
    n34,
    n18
  );


  not
  g90
  (
    n45,
    n12
  );


  buf
  g91
  (
    n71,
    n27
  );


  not
  g92
  (
    n105,
    n26
  );


  buf
  g93
  (
    n153,
    n20
  );


  buf
  g94
  (
    n109,
    n23
  );


  buf
  g95
  (
    n126,
    n17
  );


  not
  g96
  (
    n130,
    n5
  );


  not
  g97
  (
    n123,
    n8
  );


  not
  g98
  (
    n76,
    n1
  );


  not
  g99
  (
    n52,
    n7
  );


  buf
  g100
  (
    n39,
    n22
  );


  buf
  g101
  (
    n48,
    n29
  );


  not
  g102
  (
    n40,
    n15
  );


  buf
  g103
  (
    n101,
    n30
  );


  buf
  g104
  (
    n143,
    n4
  );


  not
  g105
  (
    n107,
    n21
  );


  not
  g106
  (
    n139,
    n30
  );


  buf
  g107
  (
    n97,
    n7
  );


  buf
  g108
  (
    n106,
    n3
  );


  not
  g109
  (
    n140,
    n30
  );


  not
  g110
  (
    n95,
    n2
  );


  buf
  g111
  (
    n137,
    n21
  );


  not
  g112
  (
    n55,
    n28
  );


  not
  g113
  (
    n96,
    n20
  );


  not
  g114
  (
    n152,
    n9
  );


  not
  g115
  (
    n42,
    n5
  );


  not
  g116
  (
    n98,
    n21
  );


  not
  g117
  (
    n131,
    n7
  );


  not
  g118
  (
    n65,
    n14
  );


  not
  g119
  (
    n38,
    n17
  );


  not
  g120
  (
    n154,
    n29
  );


  not
  g121
  (
    KeyWire_0_40,
    n11
  );


  buf
  g122
  (
    n110,
    n19
  );


  not
  g123
  (
    n51,
    n18
  );


  not
  g124
  (
    n561,
    n48
  );


  buf
  g125
  (
    n326,
    n47
  );


  buf
  g126
  (
    n570,
    n92
  );


  buf
  g127
  (
    n271,
    n95
  );


  buf
  g128
  (
    n559,
    n85
  );


  buf
  g129
  (
    n285,
    n124
  );


  not
  g130
  (
    n241,
    n81
  );


  not
  g131
  (
    n424,
    n66
  );


  not
  g132
  (
    n236,
    n55
  );


  buf
  g133
  (
    n164,
    n131
  );


  buf
  g134
  (
    n518,
    n78
  );


  buf
  g135
  (
    n458,
    n89
  );


  buf
  g136
  (
    n306,
    n50
  );


  not
  g137
  (
    n293,
    n87
  );


  not
  g138
  (
    n477,
    n41
  );


  not
  g139
  (
    n340,
    n66
  );


  not
  g140
  (
    n507,
    n70
  );


  not
  g141
  (
    n339,
    n78
  );


  buf
  g142
  (
    n425,
    n72
  );


  buf
  g143
  (
    n262,
    n65
  );


  not
  g144
  (
    n302,
    n105
  );


  not
  g145
  (
    n544,
    n82
  );


  buf
  g146
  (
    n439,
    n53
  );


  not
  g147
  (
    n299,
    n110
  );


  not
  g148
  (
    n167,
    n113
  );


  not
  g149
  (
    n207,
    n34
  );


  buf
  g150
  (
    n432,
    n103
  );


  not
  g151
  (
    n443,
    n118
  );


  not
  g152
  (
    n185,
    n110
  );


  buf
  g153
  (
    n500,
    n98
  );


  not
  g154
  (
    n400,
    n47
  );


  buf
  g155
  (
    n158,
    n127
  );


  not
  g156
  (
    n170,
    n127
  );


  buf
  g157
  (
    n358,
    n46
  );


  buf
  g158
  (
    n305,
    n66
  );


  buf
  g159
  (
    n498,
    n88
  );


  buf
  g160
  (
    n516,
    n76
  );


  buf
  g161
  (
    n321,
    n49
  );


  buf
  g162
  (
    n213,
    n125
  );


  not
  g163
  (
    n403,
    n106
  );


  not
  g164
  (
    n275,
    n46
  );


  not
  g165
  (
    n379,
    n50
  );


  buf
  g166
  (
    n292,
    n70
  );


  not
  g167
  (
    n368,
    n138
  );


  buf
  g168
  (
    n511,
    n64
  );


  not
  g169
  (
    n261,
    n135
  );


  buf
  g170
  (
    n573,
    n44
  );


  buf
  g171
  (
    n401,
    n41
  );


  not
  g172
  (
    n260,
    n67
  );


  buf
  g173
  (
    n374,
    n79
  );


  not
  g174
  (
    n469,
    n108
  );


  buf
  g175
  (
    n256,
    n36
  );


  buf
  g176
  (
    n535,
    n122
  );


  buf
  g177
  (
    n233,
    n55
  );


  not
  g178
  (
    n253,
    n132
  );


  not
  g179
  (
    n376,
    n115
  );


  buf
  g180
  (
    n471,
    n69
  );


  not
  g181
  (
    n472,
    n84
  );


  not
  g182
  (
    n397,
    n65
  );


  not
  g183
  (
    n291,
    n71
  );


  not
  g184
  (
    n485,
    n95
  );


  not
  g185
  (
    n332,
    n107
  );


  not
  g186
  (
    n230,
    n73
  );


  not
  g187
  (
    n398,
    n76
  );


  buf
  g188
  (
    n240,
    n133
  );


  not
  g189
  (
    n457,
    n68
  );


  not
  g190
  (
    n418,
    n133
  );


  buf
  g191
  (
    n541,
    n72
  );


  buf
  g192
  (
    n248,
    n128
  );


  buf
  g193
  (
    n337,
    n51
  );


  buf
  g194
  (
    n545,
    n99
  );


  not
  g195
  (
    n204,
    n75
  );


  not
  g196
  (
    n197,
    n85
  );


  not
  g197
  (
    n459,
    n80
  );


  not
  g198
  (
    n557,
    n113
  );


  not
  g199
  (
    n529,
    n86
  );


  buf
  g200
  (
    n222,
    n124
  );


  not
  g201
  (
    n389,
    n110
  );


  buf
  g202
  (
    n243,
    n45
  );


  buf
  g203
  (
    n417,
    n114
  );


  not
  g204
  (
    n325,
    n132
  );


  not
  g205
  (
    n440,
    n104
  );


  not
  g206
  (
    n497,
    n120
  );


  buf
  g207
  (
    n411,
    n41
  );


  not
  g208
  (
    KeyWire_0_54,
    n73
  );


  buf
  g209
  (
    n329,
    n115
  );


  not
  g210
  (
    n504,
    n63
  );


  buf
  g211
  (
    n377,
    n52
  );


  not
  g212
  (
    KeyWire_0_61,
    n134
  );


  buf
  g213
  (
    n426,
    n106
  );


  not
  g214
  (
    n528,
    n56
  );


  not
  g215
  (
    n202,
    n77
  );


  buf
  g216
  (
    n514,
    n120
  );


  not
  g217
  (
    n546,
    n112
  );


  not
  g218
  (
    n433,
    n68
  );


  not
  g219
  (
    n567,
    n96
  );


  buf
  g220
  (
    n238,
    n52
  );


  buf
  g221
  (
    n381,
    n62
  );


  buf
  g222
  (
    n183,
    n131
  );


  buf
  g223
  (
    n198,
    n105
  );


  buf
  g224
  (
    n552,
    n83
  );


  not
  g225
  (
    n218,
    n36
  );


  not
  g226
  (
    n454,
    n97
  );


  not
  g227
  (
    n569,
    n84
  );


  buf
  g228
  (
    n476,
    n57
  );


  buf
  g229
  (
    n408,
    n62
  );


  buf
  g230
  (
    n563,
    n128
  );


  not
  g231
  (
    n444,
    n135
  );


  not
  g232
  (
    n406,
    n115
  );


  not
  g233
  (
    n527,
    n38
  );


  buf
  g234
  (
    n282,
    n46
  );


  not
  g235
  (
    n239,
    n77
  );


  not
  g236
  (
    n520,
    n54
  );


  not
  g237
  (
    n348,
    n137
  );


  not
  g238
  (
    n226,
    n55
  );


  not
  g239
  (
    n189,
    n54
  );


  buf
  g240
  (
    n547,
    n84
  );


  buf
  g241
  (
    n255,
    n109
  );


  buf
  g242
  (
    n375,
    n90
  );


  not
  g243
  (
    n493,
    n130
  );


  buf
  g244
  (
    n468,
    n61
  );


  not
  g245
  (
    n521,
    n100
  );


  not
  g246
  (
    n482,
    n33
  );


  not
  g247
  (
    n412,
    n93
  );


  buf
  g248
  (
    n531,
    n78
  );


  not
  g249
  (
    n200,
    n92
  );


  buf
  g250
  (
    n180,
    n69
  );


  buf
  g251
  (
    n553,
    n81
  );


  buf
  g252
  (
    n451,
    n128
  );


  not
  g253
  (
    n437,
    n103
  );


  not
  g254
  (
    n539,
    n36
  );


  buf
  g255
  (
    n249,
    n77
  );


  not
  g256
  (
    n172,
    n129
  );


  not
  g257
  (
    n429,
    n42
  );


  buf
  g258
  (
    n259,
    n37
  );


  not
  g259
  (
    n483,
    n90
  );


  not
  g260
  (
    n228,
    n74
  );


  buf
  g261
  (
    n346,
    n138
  );


  not
  g262
  (
    n351,
    n113
  );


  buf
  g263
  (
    KeyWire_0_58,
    n105
  );


  not
  g264
  (
    n176,
    n112
  );


  buf
  g265
  (
    n513,
    n59
  );


  not
  g266
  (
    n434,
    n138
  );


  buf
  g267
  (
    n157,
    n43
  );


  buf
  g268
  (
    n281,
    n35
  );


  not
  g269
  (
    n267,
    n38
  );


  buf
  g270
  (
    n499,
    n88
  );


  buf
  g271
  (
    n347,
    n82
  );


  not
  g272
  (
    n519,
    n79
  );


  not
  g273
  (
    n314,
    n40
  );


  buf
  g274
  (
    n582,
    n118
  );


  not
  g275
  (
    n201,
    n94
  );


  buf
  g276
  (
    n273,
    n104
  );


  not
  g277
  (
    n254,
    n102
  );


  not
  g278
  (
    KeyWire_0_29,
    n33
  );


  buf
  g279
  (
    n268,
    n61
  );


  buf
  g280
  (
    n336,
    n48
  );


  not
  g281
  (
    n536,
    n90
  );


  buf
  g282
  (
    n423,
    n101
  );


  buf
  g283
  (
    n533,
    n124
  );


  buf
  g284
  (
    n246,
    n56
  );


  not
  g285
  (
    n331,
    n75
  );


  buf
  g286
  (
    n288,
    n97
  );


  not
  g287
  (
    n396,
    n43
  );


  buf
  g288
  (
    n328,
    n43
  );


  buf
  g289
  (
    n280,
    n111
  );


  buf
  g290
  (
    n470,
    n122
  );


  not
  g291
  (
    n462,
    n44
  );


  buf
  g292
  (
    n502,
    n93
  );


  not
  g293
  (
    n359,
    n91
  );


  buf
  g294
  (
    n307,
    n37
  );


  not
  g295
  (
    n242,
    n57
  );


  not
  g296
  (
    n510,
    n80
  );


  buf
  g297
  (
    n436,
    n116
  );


  buf
  g298
  (
    n577,
    n56
  );


  not
  g299
  (
    n304,
    n129
  );


  buf
  g300
  (
    n385,
    n108
  );


  not
  g301
  (
    n205,
    n91
  );


  buf
  g302
  (
    n534,
    n82
  );


  buf
  g303
  (
    n495,
    n94
  );


  buf
  g304
  (
    KeyWire_0_48,
    n116
  );


  not
  g305
  (
    n298,
    n40
  );


  buf
  g306
  (
    n555,
    n38
  );


  buf
  g307
  (
    n214,
    n67
  );


  not
  g308
  (
    n435,
    n132
  );


  buf
  g309
  (
    n225,
    n75
  );


  buf
  g310
  (
    n327,
    n127
  );


  buf
  g311
  (
    n479,
    n39
  );


  buf
  g312
  (
    n522,
    n137
  );


  not
  g313
  (
    n447,
    n62
  );


  buf
  g314
  (
    n491,
    n72
  );


  not
  g315
  (
    n341,
    n136
  );


  buf
  g316
  (
    n380,
    n90
  );


  not
  g317
  (
    n313,
    n83
  );


  buf
  g318
  (
    n461,
    n136
  );


  buf
  g319
  (
    n301,
    n68
  );


  buf
  g320
  (
    n442,
    n134
  );


  buf
  g321
  (
    n187,
    n118
  );


  buf
  g322
  (
    n182,
    n49
  );


  buf
  g323
  (
    n463,
    n71
  );


  buf
  g324
  (
    n466,
    n59
  );


  buf
  g325
  (
    n496,
    n104
  );


  buf
  g326
  (
    n196,
    n34
  );


  not
  g327
  (
    n524,
    n100
  );


  buf
  g328
  (
    n245,
    n52
  );


  buf
  g329
  (
    n428,
    n95
  );


  not
  g330
  (
    n574,
    n69
  );


  not
  g331
  (
    n550,
    n63
  );


  not
  g332
  (
    n490,
    n133
  );


  buf
  g333
  (
    n251,
    n109
  );


  buf
  g334
  (
    n395,
    n81
  );


  buf
  g335
  (
    n272,
    n139
  );


  buf
  g336
  (
    n320,
    n70
  );


  buf
  g337
  (
    n160,
    n89
  );


  buf
  g338
  (
    n274,
    n103
  );


  buf
  g339
  (
    KeyWire_0_8,
    n64
  );


  buf
  g340
  (
    n515,
    n116
  );


  buf
  g341
  (
    n478,
    n125
  );


  buf
  g342
  (
    n334,
    n54
  );


  not
  g343
  (
    n391,
    n99
  );


  buf
  g344
  (
    n364,
    n117
  );


  buf
  g345
  (
    n413,
    n120
  );


  not
  g346
  (
    n441,
    n118
  );


  not
  g347
  (
    n363,
    n86
  );


  buf
  g348
  (
    n343,
    n58
  );


  not
  g349
  (
    n366,
    n42
  );


  buf
  g350
  (
    n265,
    n60
  );


  buf
  g351
  (
    n309,
    n36
  );


  buf
  g352
  (
    n315,
    n60
  );


  not
  g353
  (
    n316,
    n88
  );


  not
  g354
  (
    n162,
    n54
  );


  buf
  g355
  (
    n300,
    n126
  );


  not
  g356
  (
    n512,
    n126
  );


  not
  g357
  (
    n386,
    n78
  );


  buf
  g358
  (
    n173,
    n77
  );


  buf
  g359
  (
    n486,
    n76
  );


  buf
  g360
  (
    n453,
    n137
  );


  buf
  g361
  (
    n576,
    n87
  );


  not
  g362
  (
    n501,
    n139
  );


  not
  g363
  (
    n171,
    n105
  );


  buf
  g364
  (
    n450,
    n102
  );


  not
  g365
  (
    n191,
    n80
  );


  buf
  g366
  (
    n221,
    n40
  );


  buf
  g367
  (
    n549,
    n57
  );


  not
  g368
  (
    n455,
    n96
  );


  buf
  g369
  (
    n538,
    n133
  );


  buf
  g370
  (
    n410,
    n98
  );


  not
  g371
  (
    n258,
    n107
  );


  not
  g372
  (
    n247,
    n44
  );


  buf
  g373
  (
    n209,
    n40
  );


  buf
  g374
  (
    n556,
    n39
  );


  not
  g375
  (
    n324,
    n58
  );


  buf
  g376
  (
    n388,
    n121
  );


  buf
  g377
  (
    n168,
    n39
  );


  buf
  g378
  (
    n421,
    n76
  );


  buf
  g379
  (
    n223,
    n107
  );


  buf
  g380
  (
    n357,
    n136
  );


  buf
  g381
  (
    n542,
    n59
  );


  not
  g382
  (
    n390,
    n112
  );


  buf
  g383
  (
    n480,
    n43
  );


  buf
  g384
  (
    n188,
    n111
  );


  buf
  g385
  (
    n407,
    n126
  );


  buf
  g386
  (
    n430,
    n86
  );


  buf
  g387
  (
    n445,
    n86
  );


  not
  g388
  (
    n393,
    n125
  );


  not
  g389
  (
    n427,
    n112
  );


  not
  g390
  (
    n572,
    n61
  );


  not
  g391
  (
    n179,
    n96
  );


  buf
  g392
  (
    n193,
    n33
  );


  not
  g393
  (
    n409,
    n135
  );


  buf
  g394
  (
    n530,
    n35
  );


  not
  g395
  (
    n270,
    n92
  );


  buf
  g396
  (
    n311,
    n134
  );


  buf
  g397
  (
    n250,
    n130
  );


  buf
  g398
  (
    n192,
    n71
  );


  buf
  g399
  (
    n489,
    n75
  );


  not
  g400
  (
    n165,
    n82
  );


  not
  g401
  (
    n558,
    n63
  );


  buf
  g402
  (
    n562,
    n115
  );


  not
  g403
  (
    n231,
    n89
  );


  buf
  g404
  (
    n355,
    n34
  );


  buf
  g405
  (
    n276,
    n129
  );


  buf
  g406
  (
    n571,
    n89
  );


  not
  g407
  (
    n540,
    n84
  );


  not
  g408
  (
    n487,
    n39
  );


  not
  g409
  (
    n295,
    n131
  );


  buf
  g410
  (
    n372,
    n73
  );


  not
  g411
  (
    n194,
    n123
  );


  buf
  g412
  (
    n517,
    n60
  );


  buf
  g413
  (
    n551,
    n58
  );


  buf
  g414
  (
    n575,
    n33
  );


  not
  g415
  (
    n523,
    n56
  );


  not
  g416
  (
    n237,
    n38
  );


  buf
  g417
  (
    n289,
    n94
  );


  not
  g418
  (
    n473,
    n65
  );


  not
  g419
  (
    n215,
    n119
  );


  buf
  g420
  (
    n580,
    n47
  );


  not
  g421
  (
    n446,
    n53
  );


  buf
  g422
  (
    n405,
    n79
  );


  not
  g423
  (
    n349,
    n64
  );


  not
  g424
  (
    n322,
    n61
  );


  not
  g425
  (
    n220,
    n123
  );


  not
  g426
  (
    n548,
    n60
  );


  not
  g427
  (
    n373,
    n117
  );


  buf
  g428
  (
    n465,
    n102
  );


  not
  g429
  (
    n352,
    n124
  );


  buf
  g430
  (
    n216,
    n138
  );


  buf
  g431
  (
    n186,
    n101
  );


  not
  g432
  (
    n277,
    n96
  );


  not
  g433
  (
    n537,
    n121
  );


  buf
  g434
  (
    n219,
    n101
  );


  buf
  g435
  (
    n229,
    n45
  );


  not
  g436
  (
    n257,
    n80
  );


  buf
  g437
  (
    n392,
    n45
  );


  buf
  g438
  (
    n422,
    n104
  );


  buf
  g439
  (
    n506,
    n48
  );


  not
  g440
  (
    n212,
    n127
  );


  buf
  g441
  (
    n365,
    n34
  );


  buf
  g442
  (
    n323,
    n121
  );


  not
  g443
  (
    n382,
    n128
  );


  not
  g444
  (
    n278,
    n117
  );


  not
  g445
  (
    n161,
    n35
  );


  not
  g446
  (
    n367,
    n126
  );


  buf
  g447
  (
    n448,
    n132
  );


  buf
  g448
  (
    n252,
    n130
  );


  buf
  g449
  (
    n294,
    n53
  );


  not
  g450
  (
    n361,
    n63
  );


  not
  g451
  (
    n206,
    n46
  );


  not
  g452
  (
    n370,
    n42
  );


  buf
  g453
  (
    n177,
    n83
  );


  not
  g454
  (
    n360,
    n88
  );


  not
  g455
  (
    n159,
    n73
  );


  not
  g456
  (
    n554,
    n107
  );


  buf
  g457
  (
    n308,
    n51
  );


  buf
  g458
  (
    n356,
    n101
  );


  not
  g459
  (
    n286,
    n119
  );


  not
  g460
  (
    n452,
    n74
  );


  buf
  g461
  (
    n526,
    n92
  );


  buf
  g462
  (
    n419,
    n123
  );


  not
  g463
  (
    n344,
    n37
  );


  buf
  g464
  (
    n383,
    n122
  );


  buf
  g465
  (
    n431,
    n59
  );


  buf
  g466
  (
    n195,
    n117
  );


  buf
  g467
  (
    n353,
    n51
  );


  not
  g468
  (
    n467,
    n98
  );


  not
  g469
  (
    n224,
    n49
  );


  not
  g470
  (
    n369,
    n68
  );


  buf
  g471
  (
    n509,
    n66
  );


  not
  g472
  (
    n203,
    n109
  );


  buf
  g473
  (
    n508,
    n62
  );


  buf
  g474
  (
    n568,
    n64
  );


  buf
  g475
  (
    n414,
    n114
  );


  not
  g476
  (
    n371,
    n113
  );


  not
  g477
  (
    n345,
    n45
  );


  buf
  g478
  (
    n264,
    n108
  );


  not
  g479
  (
    n211,
    n85
  );


  not
  g480
  (
    n416,
    n47
  );


  buf
  g481
  (
    n235,
    n114
  );


  not
  g482
  (
    n210,
    n57
  );


  not
  g483
  (
    n169,
    n49
  );


  not
  g484
  (
    n399,
    n125
  );


  buf
  g485
  (
    n505,
    n97
  );


  not
  g486
  (
    n338,
    n111
  );


  buf
  g487
  (
    n199,
    n119
  );


  buf
  g488
  (
    n163,
    n58
  );


  buf
  g489
  (
    n378,
    n106
  );


  buf
  g490
  (
    n464,
    n69
  );


  buf
  g491
  (
    n208,
    n123
  );


  not
  g492
  (
    n263,
    n72
  );


  buf
  g493
  (
    n342,
    n129
  );


  buf
  g494
  (
    n456,
    n120
  );


  buf
  g495
  (
    n579,
    n91
  );


  buf
  g496
  (
    n296,
    n97
  );


  not
  g497
  (
    n312,
    n50
  );


  not
  g498
  (
    n384,
    n137
  );


  buf
  g499
  (
    n394,
    n44
  );


  buf
  g500
  (
    n387,
    n71
  );


  not
  g501
  (
    n335,
    n99
  );


  not
  g502
  (
    n525,
    n48
  );


  not
  g503
  (
    n420,
    n121
  );


  not
  g504
  (
    n350,
    n42
  );


  not
  g505
  (
    n484,
    n108
  );


  not
  g506
  (
    n234,
    n70
  );


  buf
  g507
  (
    n319,
    n85
  );


  buf
  g508
  (
    n317,
    n93
  );


  buf
  g509
  (
    n532,
    n50
  );


  not
  g510
  (
    n488,
    n130
  );


  buf
  g511
  (
    n279,
    n41
  );


  not
  g512
  (
    n474,
    n52
  );


  not
  g513
  (
    n178,
    n83
  );


  buf
  g514
  (
    n244,
    n53
  );


  not
  g515
  (
    n492,
    n79
  );


  not
  g516
  (
    n578,
    n114
  );


  not
  g517
  (
    n438,
    n93
  );


  not
  g518
  (
    KeyWire_0_60,
    n111
  );


  not
  g519
  (
    n460,
    n131
  );


  buf
  g520
  (
    n404,
    n81
  );


  not
  g521
  (
    n449,
    n94
  );


  not
  g522
  (
    n581,
    n51
  );


  not
  g523
  (
    n290,
    n106
  );


  buf
  g524
  (
    n415,
    n119
  );


  not
  g525
  (
    n402,
    n67
  );


  buf
  g526
  (
    n175,
    n100
  );


  buf
  g527
  (
    n564,
    n37
  );


  not
  g528
  (
    n184,
    n102
  );


  not
  g529
  (
    n303,
    n95
  );


  not
  g530
  (
    n543,
    n87
  );


  not
  g531
  (
    n297,
    n136
  );


  not
  g532
  (
    n475,
    n74
  );


  not
  g533
  (
    n503,
    n110
  );


  buf
  g534
  (
    n318,
    n74
  );


  buf
  g535
  (
    n232,
    n35
  );


  buf
  g536
  (
    n217,
    n65
  );


  buf
  g537
  (
    n565,
    n99
  );


  buf
  g538
  (
    n227,
    n103
  );


  not
  g539
  (
    n287,
    n100
  );


  not
  g540
  (
    n284,
    n109
  );


  not
  g541
  (
    n333,
    n55
  );


  buf
  g542
  (
    n330,
    n116
  );


  buf
  g543
  (
    n494,
    n98
  );


  not
  g544
  (
    n560,
    n134
  );


  buf
  g545
  (
    n266,
    n67
  );


  buf
  g546
  (
    n166,
    n135
  );


  not
  g547
  (
    n269,
    n87
  );


  buf
  g548
  (
    n310,
    n122
  );


  not
  g549
  (
    n354,
    n91
  );


  and
  g550
  (
    n602,
    n337,
    n357,
    n342,
    n321
  );


  nor
  g551
  (
    n623,
    n282,
    n234,
    n205,
    n383
  );


  or
  g552
  (
    n590,
    n244,
    n364,
    n238,
    n166
  );


  xor
  g553
  (
    n609,
    n344,
    n356,
    n263,
    n362
  );


  xor
  g554
  (
    n601,
    n349,
    n232,
    n377,
    n176
  );


  nand
  g555
  (
    n603,
    n308,
    n348,
    n223,
    n256
  );


  nand
  g556
  (
    n608,
    n301,
    n233,
    n253,
    n312
  );


  nor
  g557
  (
    n620,
    n363,
    n216,
    n274,
    n339
  );


  or
  g558
  (
    n615,
    n252,
    n251,
    n317,
    n376
  );


  nand
  g559
  (
    n625,
    n273,
    n313,
    n323,
    n316
  );


  nand
  g560
  (
    n604,
    n219,
    n236,
    n359,
    n199
  );


  nand
  g561
  (
    n626,
    n172,
    n217,
    n335,
    n206
  );


  and
  g562
  (
    n618,
    n358,
    n182,
    n343,
    n369
  );


  and
  g563
  (
    n624,
    n331,
    n367,
    n379,
    n299
  );


  and
  g564
  (
    n614,
    n355,
    n157,
    n277,
    n178
  );


  nor
  g565
  (
    n585,
    n300,
    n283,
    n187,
    n332
  );


  or
  g566
  (
    n600,
    n288,
    n180,
    n162,
    n272
  );


  xnor
  g567
  (
    n639,
    n249,
    n202,
    n280,
    n188
  );


  nor
  g568
  (
    n593,
    n198,
    n354,
    n250,
    n302
  );


  and
  g569
  (
    n632,
    n171,
    n245,
    n315,
    n380
  );


  xor
  g570
  (
    n583,
    n220,
    n345,
    n292,
    n381
  );


  and
  g571
  (
    n622,
    n164,
    n254,
    n211,
    n196
  );


  or
  g572
  (
    n610,
    n371,
    n372,
    n241,
    n258
  );


  or
  g573
  (
    n616,
    n210,
    n351,
    n384,
    n341
  );


  nor
  g574
  (
    n598,
    n226,
    n324,
    n290,
    n262
  );


  xnor
  g575
  (
    n613,
    n294,
    n237,
    n231,
    n304
  );


  or
  g576
  (
    n599,
    n201,
    n230,
    n183,
    n271
  );


  xor
  g577
  (
    n633,
    n158,
    n375,
    n320,
    n336
  );


  nor
  g578
  (
    KeyWire_0_42,
    n235,
    n267,
    n209,
    n305
  );


  xnor
  g579
  (
    n627,
    n228,
    n378,
    n189,
    n260
  );


  xor
  g580
  (
    n597,
    n338,
    n327,
    n309,
    n311
  );


  xnor
  g581
  (
    n596,
    n179,
    n177,
    n303,
    n194
  );


  nand
  g582
  (
    n636,
    n373,
    n319,
    n265,
    n185
  );


  xor
  g583
  (
    n612,
    n255,
    n248,
    n186,
    n382
  );


  nand
  g584
  (
    KeyWire_0_33,
    n257,
    n213,
    n276,
    n246
  );


  nor
  g585
  (
    n589,
    n229,
    n275,
    n322,
    n287
  );


  xor
  g586
  (
    n588,
    n306,
    n240,
    n168,
    n184
  );


  nor
  g587
  (
    n617,
    n318,
    n374,
    n286,
    n352
  );


  xnor
  g588
  (
    n606,
    n270,
    n350,
    n243,
    n297
  );


  xnor
  g589
  (
    n621,
    n366,
    n208,
    n247,
    n329
  );


  or
  g590
  (
    n635,
    n190,
    n218,
    n191,
    n325
  );


  or
  g591
  (
    n605,
    n328,
    n298,
    n224,
    n307
  );


  nand
  g592
  (
    n587,
    n242,
    n163,
    n370,
    n269
  );


  xor
  g593
  (
    n586,
    n281,
    n340,
    n361,
    n326
  );


  nor
  g594
  (
    n594,
    n261,
    n259,
    n310,
    n207
  );


  xor
  g595
  (
    n595,
    n215,
    n365,
    n353,
    n330
  );


  nor
  g596
  (
    n584,
    n295,
    n204,
    n181,
    n170
  );


  nand
  g597
  (
    n631,
    n268,
    n346,
    n203,
    n212
  );


  xnor
  g598
  (
    n607,
    n214,
    n197,
    n159,
    n285
  );


  or
  g599
  (
    n611,
    n284,
    n314,
    n167,
    n165
  );


  and
  g600
  (
    n592,
    n227,
    n266,
    n291,
    n225
  );


  and
  g601
  (
    n629,
    n161,
    n173,
    n160,
    n360
  );


  nand
  g602
  (
    n591,
    n296,
    n193,
    n264,
    n175
  );


  xnor
  g603
  (
    n638,
    n192,
    n293,
    n279,
    n278
  );


  nand
  g604
  (
    n619,
    n222,
    n239,
    n333,
    n200
  );


  or
  g605
  (
    n634,
    n221,
    n334,
    n174,
    n169
  );


  and
  g606
  (
    n628,
    n195,
    n289,
    n347,
    n368
  );


  not
  g607
  (
    n686,
    n615
  );


  buf
  g608
  (
    KeyWire_0_45,
    n623
  );


  not
  g609
  (
    n675,
    n625
  );


  buf
  g610
  (
    n692,
    n593
  );


  buf
  g611
  (
    n682,
    n610
  );


  buf
  g612
  (
    n660,
    n619
  );


  buf
  g613
  (
    KeyWire_0_47,
    n595
  );


  not
  g614
  (
    n643,
    n141
  );


  buf
  g615
  (
    n640,
    n636
  );


  buf
  g616
  (
    n680,
    n586
  );


  buf
  g617
  (
    n690,
    n612
  );


  not
  g618
  (
    KeyWire_0_39,
    n587
  );


  not
  g619
  (
    n691,
    n141
  );


  not
  g620
  (
    n681,
    n617
  );


  not
  g621
  (
    n684,
    n608
  );


  not
  g622
  (
    n644,
    n632
  );


  buf
  g623
  (
    n673,
    n596
  );


  not
  g624
  (
    n659,
    n589
  );


  buf
  g625
  (
    n651,
    n627
  );


  not
  g626
  (
    n654,
    n616
  );


  buf
  g627
  (
    n669,
    n583
  );


  buf
  g628
  (
    n661,
    n630
  );


  buf
  g629
  (
    KeyWire_0_28,
    n624
  );


  buf
  g630
  (
    n662,
    n591
  );


  buf
  g631
  (
    n676,
    n585
  );


  not
  g632
  (
    n648,
    n611
  );


  not
  g633
  (
    n641,
    n622
  );


  buf
  g634
  (
    n670,
    n141
  );


  buf
  g635
  (
    n693,
    n598
  );


  buf
  g636
  (
    n656,
    n609
  );


  not
  g637
  (
    n671,
    n592
  );


  not
  g638
  (
    n642,
    n613
  );


  buf
  g639
  (
    n647,
    n607
  );


  buf
  g640
  (
    n679,
    n621
  );


  buf
  g641
  (
    n652,
    n597
  );


  not
  g642
  (
    n677,
    n140
  );


  not
  g643
  (
    n667,
    n140
  );


  not
  g644
  (
    n688,
    n629
  );


  buf
  g645
  (
    n668,
    n606
  );


  buf
  g646
  (
    n663,
    n139
  );


  buf
  g647
  (
    n674,
    n594
  );


  buf
  g648
  (
    n678,
    n604
  );


  buf
  g649
  (
    n687,
    n603
  );


  buf
  g650
  (
    n657,
    n631
  );


  not
  g651
  (
    n683,
    n601
  );


  buf
  g652
  (
    n649,
    n599
  );


  not
  g653
  (
    n672,
    n634
  );


  buf
  g654
  (
    n646,
    n140
  );


  not
  g655
  (
    n653,
    n584
  );


  not
  g656
  (
    n665,
    n614
  );


  nand
  g657
  (
    n664,
    n600,
    n141
  );


  and
  g658
  (
    n650,
    n628,
    n618,
    n626,
    n140
  );


  nand
  g659
  (
    n645,
    n635,
    n633,
    n588,
    n602
  );


  or
  g660
  (
    n655,
    n139,
    n620,
    n590,
    n605
  );


  not
  g661
  (
    n714,
    n641
  );


  buf
  g662
  (
    n731,
    n687
  );


  not
  g663
  (
    n886,
    n673
  );


  not
  g664
  (
    n786,
    n152
  );


  not
  g665
  (
    n709,
    n654
  );


  not
  g666
  (
    KeyWire_0_18,
    n144
  );


  buf
  g667
  (
    n862,
    n663
  );


  not
  g668
  (
    n739,
    n667
  );


  not
  g669
  (
    n790,
    n645
  );


  buf
  g670
  (
    n764,
    n684
  );


  not
  g671
  (
    n809,
    n144
  );


  not
  g672
  (
    n779,
    n147
  );


  buf
  g673
  (
    n840,
    n660
  );


  not
  g674
  (
    n889,
    n671
  );


  buf
  g675
  (
    n825,
    n648
  );


  buf
  g676
  (
    n706,
    n662
  );


  buf
  g677
  (
    n870,
    n656
  );


  not
  g678
  (
    n838,
    n150
  );


  not
  g679
  (
    n888,
    n661
  );


  buf
  g680
  (
    n784,
    n658
  );


  not
  g681
  (
    n874,
    n145
  );


  not
  g682
  (
    n720,
    n652
  );


  not
  g683
  (
    n780,
    n677
  );


  buf
  g684
  (
    n831,
    n686
  );


  not
  g685
  (
    n799,
    n146
  );


  buf
  g686
  (
    n702,
    n651
  );


  not
  g687
  (
    KeyWire_0_51,
    n648
  );


  buf
  g688
  (
    n844,
    n674
  );


  buf
  g689
  (
    n859,
    n151
  );


  not
  g690
  (
    n819,
    n669
  );


  not
  g691
  (
    KeyWire_0_34,
    n654
  );


  buf
  g692
  (
    n716,
    n647
  );


  not
  g693
  (
    n881,
    n152
  );


  buf
  g694
  (
    n726,
    n652
  );


  buf
  g695
  (
    n807,
    n642
  );


  buf
  g696
  (
    n757,
    n649
  );


  buf
  g697
  (
    n877,
    n684
  );


  not
  g698
  (
    n800,
    n648
  );


  not
  g699
  (
    n861,
    n650
  );


  not
  g700
  (
    n697,
    n688
  );


  not
  g701
  (
    n738,
    n662
  );


  buf
  g702
  (
    n772,
    n661
  );


  buf
  g703
  (
    n759,
    n643
  );


  not
  g704
  (
    n884,
    n655
  );


  not
  g705
  (
    n715,
    n149
  );


  not
  g706
  (
    n857,
    n673
  );


  buf
  g707
  (
    n815,
    n145
  );


  not
  g708
  (
    n745,
    n658
  );


  buf
  g709
  (
    n754,
    n656
  );


  not
  g710
  (
    n843,
    n674
  );


  not
  g711
  (
    n871,
    n666
  );


  not
  g712
  (
    n851,
    n649
  );


  buf
  g713
  (
    n725,
    n669
  );


  buf
  g714
  (
    n782,
    n678
  );


  not
  g715
  (
    n766,
    n151
  );


  not
  g716
  (
    n719,
    n682
  );


  buf
  g717
  (
    n763,
    n685
  );


  buf
  g718
  (
    n873,
    n675
  );


  not
  g719
  (
    n867,
    n684
  );


  not
  g720
  (
    n748,
    n661
  );


  not
  g721
  (
    n841,
    n653
  );


  buf
  g722
  (
    n860,
    n663
  );


  not
  g723
  (
    n864,
    n640
  );


  not
  g724
  (
    n769,
    n147
  );


  buf
  g725
  (
    n774,
    n647
  );


  not
  g726
  (
    KeyWire_0_16,
    n150
  );


  buf
  g727
  (
    n821,
    n658
  );


  not
  g728
  (
    n750,
    n149
  );


  not
  g729
  (
    n768,
    n659
  );


  buf
  g730
  (
    n848,
    n657
  );


  not
  g731
  (
    n741,
    n643
  );


  not
  g732
  (
    n744,
    n148
  );


  not
  g733
  (
    n736,
    n681
  );


  buf
  g734
  (
    n858,
    n641
  );


  buf
  g735
  (
    n802,
    n676
  );


  not
  g736
  (
    n883,
    n646
  );


  buf
  g737
  (
    n836,
    n145
  );


  not
  g738
  (
    n710,
    n659
  );


  not
  g739
  (
    n876,
    n662
  );


  not
  g740
  (
    n696,
    n670
  );


  not
  g741
  (
    n747,
    n646
  );


  buf
  g742
  (
    KeyWire_0_43,
    n673
  );


  not
  g743
  (
    n855,
    n659
  );


  buf
  g744
  (
    n712,
    n151
  );


  buf
  g745
  (
    n824,
    n666
  );


  not
  g746
  (
    n869,
    n657
  );


  not
  g747
  (
    n701,
    n653
  );


  not
  g748
  (
    KeyWire_0_52,
    n662
  );


  not
  g749
  (
    n775,
    n688
  );


  buf
  g750
  (
    n791,
    n675
  );


  buf
  g751
  (
    n845,
    n660
  );


  not
  g752
  (
    n827,
    n687
  );


  not
  g753
  (
    n723,
    n658
  );


  not
  g754
  (
    n765,
    n641
  );


  not
  g755
  (
    n789,
    n142
  );


  not
  g756
  (
    n850,
    n685
  );


  not
  g757
  (
    n835,
    n683
  );


  buf
  g758
  (
    n794,
    n665
  );


  buf
  g759
  (
    n797,
    n659
  );


  buf
  g760
  (
    n879,
    n672
  );


  not
  g761
  (
    n760,
    n642
  );


  not
  g762
  (
    n770,
    n672
  );


  buf
  g763
  (
    n756,
    n150
  );


  buf
  g764
  (
    n853,
    n677
  );


  not
  g765
  (
    n808,
    n645
  );


  buf
  g766
  (
    n793,
    n681
  );


  buf
  g767
  (
    n762,
    n686
  );


  not
  g768
  (
    n730,
    n142
  );


  not
  g769
  (
    n818,
    n647
  );


  not
  g770
  (
    n713,
    n143
  );


  buf
  g771
  (
    n755,
    n667
  );


  not
  g772
  (
    n734,
    n679
  );


  not
  g773
  (
    n761,
    n672
  );


  not
  g774
  (
    n866,
    n642
  );


  buf
  g775
  (
    n842,
    n651
  );


  not
  g776
  (
    n875,
    n645
  );


  buf
  g777
  (
    n834,
    n644
  );


  buf
  g778
  (
    n854,
    n664
  );


  buf
  g779
  (
    n694,
    n687
  );


  buf
  g780
  (
    n865,
    n657
  );


  not
  g781
  (
    n826,
    n150
  );


  buf
  g782
  (
    n724,
    n640
  );


  not
  g783
  (
    n721,
    n688
  );


  not
  g784
  (
    n828,
    n679
  );


  not
  g785
  (
    n746,
    n680
  );


  buf
  g786
  (
    n717,
    n668
  );


  not
  g787
  (
    n796,
    n143
  );


  not
  g788
  (
    n722,
    n669
  );


  not
  g789
  (
    n711,
    n686
  );


  buf
  g790
  (
    n887,
    n149
  );


  not
  g791
  (
    n820,
    n678
  );


  not
  g792
  (
    n695,
    n675
  );


  buf
  g793
  (
    n823,
    n661
  );


  not
  g794
  (
    n735,
    n657
  );


  buf
  g795
  (
    n810,
    n666
  );


  not
  g796
  (
    n878,
    n681
  );


  not
  g797
  (
    n773,
    n650
  );


  not
  g798
  (
    KeyWire_0_26,
    n680
  );


  buf
  g799
  (
    n872,
    n649
  );


  not
  g800
  (
    n792,
    n648
  );


  not
  g801
  (
    n707,
    n642
  );


  not
  g802
  (
    n856,
    n664
  );


  buf
  g803
  (
    n829,
    n144
  );


  not
  g804
  (
    n846,
    n668
  );


  not
  g805
  (
    n718,
    n686
  );


  not
  g806
  (
    n785,
    n647
  );


  not
  g807
  (
    n727,
    n146
  );


  not
  g808
  (
    n813,
    n146
  );


  not
  g809
  (
    n811,
    n678
  );


  buf
  g810
  (
    n863,
    n143
  );


  buf
  g811
  (
    n822,
    n147
  );


  not
  g812
  (
    n728,
    n142
  );


  not
  g813
  (
    n804,
    n665
  );


  not
  g814
  (
    n806,
    n646
  );


  buf
  g815
  (
    n852,
    n142
  );


  buf
  g816
  (
    n778,
    n656
  );


  not
  g817
  (
    n812,
    n143
  );


  not
  g818
  (
    n729,
    n671
  );


  buf
  g819
  (
    n742,
    n147
  );


  buf
  g820
  (
    KeyWire_0_1,
    n643
  );


  buf
  g821
  (
    n733,
    n148
  );


  buf
  g822
  (
    n880,
    n679
  );


  not
  g823
  (
    n832,
    n675
  );


  buf
  g824
  (
    n788,
    n678
  );


  not
  g825
  (
    n704,
    n649
  );


  buf
  g826
  (
    n805,
    n665
  );


  not
  g827
  (
    n698,
    n680
  );


  not
  g828
  (
    n708,
    n674
  );


  not
  g829
  (
    n740,
    n654
  );


  buf
  g830
  (
    n781,
    n152
  );


  buf
  g831
  (
    n833,
    n667
  );


  buf
  g832
  (
    n795,
    n688
  );


  buf
  g833
  (
    n776,
    n654
  );


  buf
  g834
  (
    n839,
    n672
  );


  buf
  g835
  (
    n837,
    n644
  );


  buf
  g836
  (
    n798,
    n683
  );


  not
  g837
  (
    n753,
    n646
  );


  not
  g838
  (
    n737,
    n655
  );


  not
  g839
  (
    n749,
    n684
  );


  buf
  g840
  (
    n699,
    n148
  );


  or
  g841
  (
    n817,
    n676,
    n667
  );


  nor
  g842
  (
    n703,
    n144,
    n685
  );


  and
  g843
  (
    n752,
    n650,
    n652,
    n677,
    n145
  );


  xor
  g844
  (
    n816,
    n663,
    n683,
    n640,
    n682
  );


  xnor
  g845
  (
    n771,
    n671,
    n668,
    n670,
    n665
  );


  xor
  g846
  (
    n801,
    n676,
    n663,
    n655,
    n640
  );


  nand
  g847
  (
    n700,
    n676,
    n677,
    n651,
    n670
  );


  or
  g848
  (
    n767,
    n664,
    n666,
    n644,
    n679
  );


  and
  g849
  (
    n787,
    n664,
    n671,
    n146,
    n660
  );


  nor
  g850
  (
    n732,
    n682,
    n653,
    n655
  );


  xor
  g851
  (
    n803,
    n668,
    n660,
    n650,
    n683
  );


  and
  g852
  (
    n814,
    n152,
    n645,
    n680,
    n643
  );


  xor
  g853
  (
    n705,
    n644,
    n670,
    n669,
    n148
  );


  xor
  g854
  (
    n777,
    n673,
    n652,
    n151,
    n656
  );


  and
  g855
  (
    n849,
    n674,
    n685,
    n149,
    n651
  );


  xor
  g856
  (
    n751,
    n687,
    n681,
    n682,
    n641
  );


  xor
  g857
  (
    n1028,
    n571,
    n478,
    n504,
    n827
  );


  or
  g858
  (
    n976,
    n794,
    n812,
    n715,
    n765
  );


  xor
  g859
  (
    n908,
    n700,
    n517,
    n770,
    n537
  );


  and
  g860
  (
    n927,
    n718,
    n774,
    n445,
    n567
  );


  nor
  g861
  (
    n989,
    n711,
    n516,
    n509,
    n830
  );


  nor
  g862
  (
    KeyWire_0_21,
    n552,
    n772,
    n714,
    n544
  );


  xor
  g863
  (
    n1013,
    n836,
    n556,
    n515,
    n492
  );


  xnor
  g864
  (
    n936,
    n750,
    n727,
    n436,
    n449
  );


  xnor
  g865
  (
    n975,
    n565,
    n569,
    n441,
    n564
  );


  xnor
  g866
  (
    n960,
    n726,
    n564,
    n430,
    n546
  );


  or
  g867
  (
    n963,
    n833,
    n769,
    n808,
    n507
  );


  and
  g868
  (
    n980,
    n555,
    n734,
    n709,
    n735
  );


  nor
  g869
  (
    n947,
    n698,
    n815,
    n786,
    n501
  );


  and
  g870
  (
    n946,
    n568,
    n554,
    n455,
    n548
  );


  or
  g871
  (
    n1021,
    n559,
    n749,
    n731,
    n785
  );


  or
  g872
  (
    n952,
    n820,
    n788,
    n519,
    n762
  );


  nor
  g873
  (
    n921,
    n825,
    n570,
    n526,
    n450
  );


  xnor
  g874
  (
    n979,
    n837,
    n563,
    n468,
    n516
  );


  xor
  g875
  (
    n977,
    n560,
    n824,
    n409,
    n523
  );


  and
  g876
  (
    n961,
    n469,
    n435,
    n764,
    n485
  );


  nor
  g877
  (
    n926,
    n550,
    n730,
    n708,
    n466
  );


  xor
  g878
  (
    n899,
    n795,
    n695,
    n525,
    n754
  );


  nor
  g879
  (
    n900,
    n520,
    n710,
    n555,
    n524
  );


  nand
  g880
  (
    n992,
    n801,
    n545,
    n700,
    n829
  );


  and
  g881
  (
    n974,
    n431,
    n790,
    n749,
    n813
  );


  xnor
  g882
  (
    n928,
    n807,
    n793,
    n560,
    n410
  );


  nand
  g883
  (
    n933,
    n823,
    n538,
    n727,
    n758
  );


  xor
  g884
  (
    n965,
    n407,
    n811,
    n558,
    n773
  );


  xor
  g885
  (
    n994,
    n824,
    n459,
    n735,
    n718
  );


  nor
  g886
  (
    n1024,
    n443,
    n408,
    n780,
    n838
  );


  nand
  g887
  (
    n895,
    n780,
    n712,
    n433,
    n756
  );


  or
  g888
  (
    n905,
    n422,
    n391,
    n759,
    n713
  );


  nor
  g889
  (
    n983,
    n439,
    n522,
    n471,
    n543
  );


  xor
  g890
  (
    n1020,
    n781,
    n527,
    n766,
    n519
  );


  nand
  g891
  (
    n914,
    n804,
    n771,
    n551,
    n719
  );


  nand
  g892
  (
    n892,
    n406,
    n529,
    n545,
    n794
  );


  and
  g893
  (
    n950,
    n518,
    n534,
    n787,
    n568
  );


  and
  g894
  (
    n918,
    n820,
    n544,
    n782,
    n696
  );


  nand
  g895
  (
    n920,
    n779,
    n553,
    n501,
    n523
  );


  and
  g896
  (
    n909,
    n807,
    n739,
    n387,
    n771
  );


  nor
  g897
  (
    n923,
    n415,
    n751,
    n446,
    n831
  );


  xor
  g898
  (
    n982,
    n509,
    n474,
    n806,
    n536
  );


  xnor
  g899
  (
    n1000,
    n764,
    n529,
    n801,
    n708
  );


  xnor
  g900
  (
    n1015,
    n743,
    n760,
    n514,
    n778
  );


  and
  g901
  (
    n938,
    n453,
    n800,
    n833,
    n746
  );


  nor
  g902
  (
    n1001,
    n748,
    n806,
    n442,
    n702
  );


  nor
  g903
  (
    n1025,
    n569,
    n405,
    n740,
    n793
  );


  and
  g904
  (
    KeyWire_0_19,
    n479,
    n805,
    n840,
    n429
  );


  nor
  g905
  (
    n897,
    n723,
    n738,
    n543,
    n799
  );


  nand
  g906
  (
    n1027,
    n828,
    n808,
    n426,
    n530
  );


  and
  g907
  (
    n949,
    n819,
    n497,
    n508,
    n502
  );


  nor
  g908
  (
    n1016,
    n491,
    n798,
    n573,
    n540
  );


  nor
  g909
  (
    n1012,
    n412,
    n456,
    n777,
    n417
  );


  nor
  g910
  (
    n1005,
    n505,
    n716,
    n755,
    n398
  );


  xnor
  g911
  (
    n894,
    n802,
    n757,
    n719,
    n753
  );


  nand
  g912
  (
    n934,
    n490,
    n835,
    n473,
    n448
  );


  and
  g913
  (
    n987,
    n752,
    n486,
    n452,
    n488
  );


  xor
  g914
  (
    n890,
    n528,
    n495,
    n472,
    n724
  );


  xor
  g915
  (
    KeyWire_0_27,
    n517,
    n732,
    n783,
    n461
  );


  nand
  g916
  (
    KeyWire_0_5,
    n394,
    n504,
    n553,
    n829
  );


  or
  g917
  (
    n925,
    n776,
    n521,
    n742,
    n520
  );


  xor
  g918
  (
    n998,
    n470,
    n538,
    n481,
    n744
  );


  or
  g919
  (
    n919,
    n798,
    n542,
    n707,
    n482
  );


  xor
  g920
  (
    n1023,
    n728,
    n532,
    n546,
    n725
  );


  nand
  g921
  (
    n893,
    n571,
    n745,
    n710,
    n532
  );


  or
  g922
  (
    n944,
    n549,
    n411,
    n542,
    n775
  );


  nand
  g923
  (
    n990,
    n721,
    n558,
    n424,
    n722
  );


  xor
  g924
  (
    n922,
    n772,
    n760,
    n751,
    n502
  );


  or
  g925
  (
    n967,
    n460,
    n561,
    n528,
    n511
  );


  and
  g926
  (
    n917,
    n434,
    n804,
    n717,
    n789
  );


  nor
  g927
  (
    n913,
    n723,
    n755,
    n747,
    n694
  );


  xnor
  g928
  (
    n981,
    n818,
    n761,
    n438,
    n769
  );


  xor
  g929
  (
    n1022,
    n796,
    n420,
    n770,
    n822
  );


  nand
  g930
  (
    n1003,
    n716,
    n416,
    n540,
    n821
  );


  xnor
  g931
  (
    n932,
    n728,
    n554,
    n499,
    n739
  );


  nor
  g932
  (
    n988,
    n697,
    n813,
    n809,
    n839
  );


  xnor
  g933
  (
    n930,
    n548,
    n530,
    n779,
    n547
  );


  nand
  g934
  (
    n903,
    n791,
    n714,
    n782,
    n831
  );


  and
  g935
  (
    n995,
    n786,
    n803,
    n699,
    n552
  );


  nand
  g936
  (
    n939,
    n707,
    n752,
    n503,
    n774
  );


  and
  g937
  (
    n953,
    n514,
    n572,
    n531,
    n521
  );


  and
  g938
  (
    n1002,
    n512,
    n389,
    n834,
    n561
  );


  nor
  g939
  (
    n1014,
    n392,
    n536,
    n787,
    n464
  );


  or
  g940
  (
    n1017,
    n432,
    n822,
    n814,
    n753
  );


  xor
  g941
  (
    n901,
    n508,
    n777,
    n788,
    n451
  );


  and
  g942
  (
    n902,
    n698,
    n830,
    n697,
    n447
  );


  nand
  g943
  (
    n907,
    n393,
    n518,
    n525,
    n737
  );


  nor
  g944
  (
    n942,
    n732,
    n722,
    n494,
    n513
  );


  or
  g945
  (
    n959,
    n701,
    n388,
    n733,
    n730
  );


  or
  g946
  (
    n941,
    n816,
    n818,
    n505,
    n427
  );


  nor
  g947
  (
    n1018,
    n773,
    n531,
    n810,
    n791
  );


  and
  g948
  (
    n896,
    n498,
    n792,
    n385,
    n535
  );


  nor
  g949
  (
    n940,
    n704,
    n784,
    n712,
    n480
  );


  nand
  g950
  (
    n958,
    n566,
    n766,
    n817,
    n699
  );


  or
  g951
  (
    n912,
    n738,
    n703,
    n510,
    n487
  );


  and
  g952
  (
    n931,
    n454,
    n709,
    n399,
    n832
  );


  xnor
  g953
  (
    n943,
    n507,
    n547,
    n503,
    n397
  );


  nand
  g954
  (
    n945,
    n767,
    n781,
    n828,
    n396
  );


  nor
  g955
  (
    n972,
    n506,
    n795,
    n476,
    n836
  );


  nand
  g956
  (
    KeyWire_0_4,
    n562,
    n541,
    n563,
    n499
  );


  or
  g957
  (
    n999,
    n694,
    n425,
    n784,
    n811
  );


  nor
  g958
  (
    KeyWire_0_6,
    n827,
    n562,
    n759,
    n783
  );


  or
  g959
  (
    n915,
    n403,
    n741,
    n803,
    n423
  );


  nand
  g960
  (
    n966,
    n725,
    n825,
    n513,
    n720
  );


  nor
  g961
  (
    n955,
    n744,
    n437,
    n826,
    n386
  );


  xnor
  g962
  (
    n985,
    n535,
    n810,
    n785,
    n823
  );


  xor
  g963
  (
    n929,
    n701,
    n762,
    n834,
    n489
  );


  and
  g964
  (
    n1019,
    n706,
    n467,
    n705,
    n741
  );


  nand
  g965
  (
    n970,
    n500,
    n734,
    n413,
    n715
  );


  and
  g966
  (
    n1009,
    n567,
    n477,
    n748,
    n726
  );


  xnor
  g967
  (
    n935,
    n565,
    n835,
    n706,
    n465
  );


  and
  g968
  (
    n1007,
    n703,
    n541,
    n717,
    n839
  );


  xor
  g969
  (
    n968,
    n400,
    n705,
    n792,
    n566
  );


  xnor
  g970
  (
    n986,
    n826,
    n729,
    n570,
    n402
  );


  nor
  g971
  (
    n910,
    n736,
    n522,
    n534,
    n790
  );


  xor
  g972
  (
    n898,
    n526,
    n837,
    n539,
    n756
  );


  xor
  g973
  (
    n891,
    n390,
    n572,
    n747,
    n419
  );


  and
  g974
  (
    n1006,
    n832,
    n696,
    n440,
    n797
  );


  xor
  g975
  (
    n973,
    n733,
    n702,
    n800,
    n713
  );


  or
  g976
  (
    n1026,
    n720,
    n737,
    n421,
    n731
  );


  or
  g977
  (
    n904,
    n483,
    n821,
    n484,
    n695
  );


  xor
  g978
  (
    n1008,
    n750,
    n458,
    n496,
    n736
  );


  or
  g979
  (
    n993,
    n493,
    n817,
    n533,
    n506
  );


  xnor
  g980
  (
    KeyWire_0_50,
    n768,
    n557,
    n814,
    n812
  );


  xnor
  g981
  (
    n969,
    n768,
    n512,
    n724,
    n789
  );


  nor
  g982
  (
    n911,
    n796,
    n763,
    n711,
    n418
  );


  and
  g983
  (
    n978,
    n704,
    n550,
    n757,
    n475
  );


  nor
  g984
  (
    n948,
    n533,
    n758,
    n462,
    n799
  );


  and
  g985
  (
    n957,
    n767,
    n395,
    n775,
    n743
  );


  xnor
  g986
  (
    n991,
    n537,
    n463,
    n511,
    n556
  );


  xnor
  g987
  (
    n996,
    n539,
    n809,
    n778,
    n797
  );


  or
  g988
  (
    n954,
    n729,
    n515,
    n524,
    n802
  );


  nand
  g989
  (
    n924,
    n428,
    n404,
    n549,
    n457
  );


  nor
  g990
  (
    n984,
    n746,
    n444,
    n776,
    n816
  );


  nor
  g991
  (
    n997,
    n742,
    n740,
    n765,
    n838
  );


  xor
  g992
  (
    n956,
    n745,
    n815,
    n500,
    n721
  );


  xnor
  g993
  (
    KeyWire_0_17,
    n559,
    n551,
    n819,
    n754
  );


  or
  g994
  (
    n1011,
    n401,
    n527,
    n510,
    n805
  );


  and
  g995
  (
    n916,
    n557,
    n763,
    n414,
    n761
  );


  not
  g996
  (
    n1042,
    n899
  );


  not
  g997
  (
    n1035,
    n903
  );


  not
  g998
  (
    n1030,
    n905
  );


  not
  g999
  (
    n1033,
    n890
  );


  buf
  g1000
  (
    KeyWire_0_22,
    n904
  );


  not
  g1001
  (
    n1047,
    n907
  );


  buf
  g1002
  (
    n1031,
    n900
  );


  buf
  g1003
  (
    n1048,
    n901
  );


  not
  g1004
  (
    n1037,
    n908
  );


  not
  g1005
  (
    n1032,
    n898
  );


  not
  g1006
  (
    n1029,
    n895
  );


  not
  g1007
  (
    n1043,
    n894
  );


  not
  g1008
  (
    n1034,
    n909
  );


  buf
  g1009
  (
    n1040,
    n892
  );


  not
  g1010
  (
    n1041,
    n902
  );


  buf
  g1011
  (
    KeyWire_0_35,
    n891
  );


  not
  g1012
  (
    n1044,
    n897
  );


  not
  g1013
  (
    n1039,
    n906
  );


  buf
  g1014
  (
    n1036,
    n896
  );


  not
  g1015
  (
    n1038,
    n893
  );


  and
  g1016
  (
    n1062,
    n850,
    n914,
    n1035,
    n1032
  );


  and
  g1017
  (
    n1053,
    n1036,
    n844,
    n855,
    n858
  );


  nor
  g1018
  (
    n1051,
    n842,
    n1031,
    n856,
    n843
  );


  xor
  g1019
  (
    n1055,
    n850,
    n841,
    n1034,
    n855
  );


  nor
  g1020
  (
    n1065,
    n843,
    n853,
    n911,
    n916
  );


  xor
  g1021
  (
    n1050,
    n857,
    n1031,
    n846,
    n1029
  );


  or
  g1022
  (
    n1052,
    n850,
    n847,
    n851,
    n857
  );


  or
  g1023
  (
    n1056,
    n848,
    n1037,
    n849,
    n915
  );


  or
  g1024
  (
    n1058,
    n853,
    n1030,
    n848
  );


  xnor
  g1025
  (
    n1064,
    n848,
    n1038,
    n847,
    n858
  );


  and
  g1026
  (
    n1061,
    n849,
    n856,
    n689,
    n1033
  );


  or
  g1027
  (
    KeyWire_0_13,
    n849,
    n852,
    n857,
    n913
  );


  xor
  g1028
  (
    n1049,
    n858,
    n854,
    n852,
    n1037
  );


  xor
  g1029
  (
    n1054,
    n1038,
    n852,
    n1037,
    n1029
  );


  nor
  g1030
  (
    n1057,
    n847,
    n844,
    n854,
    n840
  );


  and
  g1031
  (
    n1067,
    n854,
    n1038,
    n842,
    n845
  );


  nand
  g1032
  (
    n1068,
    n850,
    n689,
    n848,
    n856
  );


  or
  g1033
  (
    n1070,
    n910,
    n849,
    n853,
    n851
  );


  nor
  g1034
  (
    n1069,
    n851,
    n853,
    n1035,
    n1032
  );


  or
  g1035
  (
    KeyWire_0_41,
    n847,
    n852,
    n689,
    n1033
  );


  xor
  g1036
  (
    n1072,
    n851,
    n846,
    n856,
    n845
  );


  xnor
  g1037
  (
    n1071,
    n912,
    n689,
    n1034,
    n1036
  );


  xnor
  g1038
  (
    n1063,
    n1038,
    n841,
    n1037,
    n855
  );


  and
  g1039
  (
    n1060,
    n917,
    n854,
    n857,
    n855
  );


  xor
  g1040
  (
    n1091,
    n865,
    n878,
    n1066,
    n858
  );


  xnor
  g1041
  (
    n1109,
    n880,
    n1063,
    n883,
    n862
  );


  and
  g1042
  (
    n1105,
    n874,
    n1067,
    n919,
    n864
  );


  xnor
  g1043
  (
    n1099,
    n881,
    n1068,
    n1055,
    n884
  );


  xnor
  g1044
  (
    n1092,
    n874,
    n870,
    n866,
    n861
  );


  or
  g1045
  (
    n1075,
    n866,
    n1062,
    n861,
    n868
  );


  xor
  g1046
  (
    n1097,
    n877,
    n918,
    n1049,
    n861
  );


  nand
  g1047
  (
    n1084,
    n881,
    n859,
    n884,
    n871
  );


  nand
  g1048
  (
    n1080,
    n867,
    n883,
    n875,
    n868
  );


  nand
  g1049
  (
    n1082,
    n880,
    n1069,
    n1070,
    n866
  );


  or
  g1050
  (
    n1085,
    n872,
    n859,
    n1068,
    n873
  );


  xnor
  g1051
  (
    KeyWire_0_37,
    n1058,
    n863,
    n869,
    n864
  );


  nand
  g1052
  (
    n1087,
    n864,
    n1071,
    n885,
    n881
  );


  or
  g1053
  (
    n1083,
    n879,
    n862,
    n878,
    n876
  );


  xnor
  g1054
  (
    n1103,
    n877,
    n875,
    n1071,
    n882
  );


  xor
  g1055
  (
    n1098,
    n883,
    n872,
    n1064,
    n863
  );


  xor
  g1056
  (
    n1078,
    n884,
    n865,
    n869,
    n859
  );


  xor
  g1057
  (
    n1088,
    n870,
    n1070,
    n864,
    n869
  );


  or
  g1058
  (
    n1086,
    n1061,
    n1070,
    n867,
    n1071
  );


  xor
  g1059
  (
    KeyWire_0_25,
    n865,
    n885,
    n882,
    n860
  );


  xor
  g1060
  (
    n1096,
    n862,
    n1056,
    n875,
    n1052
  );


  or
  g1061
  (
    n1077,
    n876,
    n861,
    n870,
    n871
  );


  nand
  g1062
  (
    n1090,
    n873,
    n878,
    n1069
  );


  xor
  g1063
  (
    n1107,
    n871,
    n875,
    n862,
    n885
  );


  and
  g1064
  (
    n1100,
    n1067,
    n871,
    n882,
    n872
  );


  nor
  g1065
  (
    n1104,
    n882,
    n880,
    n1053,
    n868
  );


  xnor
  g1066
  (
    n1106,
    n869,
    n874,
    n867,
    n870
  );


  nand
  g1067
  (
    n1076,
    n878,
    n866,
    n1060,
    n1069
  );


  nand
  g1068
  (
    n1073,
    n1057,
    n1051,
    n865,
    n1068
  );


  and
  g1069
  (
    n1101,
    n877,
    n879,
    n873
  );


  xor
  g1070
  (
    n1102,
    n1054,
    n1067,
    n872,
    n863
  );


  and
  g1071
  (
    n1094,
    n885,
    n860,
    n873,
    n868
  );


  and
  g1072
  (
    n1079,
    n877,
    n876,
    n1059,
    n860
  );


  nand
  g1073
  (
    n1095,
    n1068,
    n881,
    n874,
    n859
  );


  nor
  g1074
  (
    n1074,
    n1065,
    n879,
    n876,
    n883
  );


  or
  g1075
  (
    n1089,
    n863,
    n860,
    n1070,
    n1050
  );


  xnor
  g1076
  (
    n1108,
    n880,
    n1067,
    n884,
    n867
  );


  not
  g1077
  (
    n1110,
    n930
  );


  not
  g1078
  (
    n1124,
    n922
  );


  buf
  g1079
  (
    n1125,
    n1102
  );


  buf
  g1080
  (
    n1114,
    n1083
  );


  buf
  g1081
  (
    n1111,
    n928
  );


  not
  g1082
  (
    n1120,
    n931
  );


  buf
  g1083
  (
    n1133,
    n1091
  );


  not
  g1084
  (
    n1127,
    n1084
  );


  not
  g1085
  (
    n1123,
    n1101
  );


  buf
  g1086
  (
    n1118,
    n1092
  );


  buf
  g1087
  (
    n1131,
    n925
  );


  buf
  g1088
  (
    n1116,
    n1100
  );


  buf
  g1089
  (
    n1119,
    n920
  );


  not
  g1090
  (
    n1112,
    n1093
  );


  buf
  g1091
  (
    n1113,
    n1088
  );


  not
  g1092
  (
    n1122,
    n923
  );


  buf
  g1093
  (
    n1126,
    n1095
  );


  buf
  g1094
  (
    n1117,
    n924
  );


  buf
  g1095
  (
    n1132,
    n929
  );


  buf
  g1096
  (
    n1128,
    n1105
  );


  nand
  g1097
  (
    n1115,
    n1082,
    n1096,
    n1087,
    n1094
  );


  nand
  g1098
  (
    n1130,
    n1085,
    n1086,
    n1090,
    n1089
  );


  nand
  g1099
  (
    n1129,
    n926,
    n1099,
    n1098,
    n1104
  );


  xor
  g1100
  (
    n1121,
    n1097,
    n927,
    n921,
    n1103
  );


  xnor
  g1101
  (
    n1135,
    n1117,
    n886,
    n1114
  );


  nor
  g1102
  (
    n1204,
    n1121,
    n1128,
    n943
  );


  or
  g1103
  (
    n1164,
    n638,
    n1132,
    n154
  );


  xnor
  g1104
  (
    n1165,
    n886,
    n1123
  );


  or
  g1105
  (
    n1207,
    n954,
    n933,
    n969
  );


  xor
  g1106
  (
    n1181,
    n1109,
    n1111,
    n32
  );


  nand
  g1107
  (
    n1195,
    n949,
    n1045,
    n1123
  );


  or
  g1108
  (
    n1213,
    n1122,
    n691,
    n1048
  );


  xnor
  g1109
  (
    KeyWire_0_2,
    n1130,
    n1004,
    n1114
  );


  and
  g1110
  (
    n1194,
    n984,
    n993,
    n959
  );


  xor
  g1111
  (
    n1171,
    n1007,
    n1046,
    n982
  );


  nand
  g1112
  (
    n1177,
    n1117,
    n963,
    n1130
  );


  nor
  g1113
  (
    n1139,
    n1132,
    n1005,
    n980
  );


  xor
  g1114
  (
    n1174,
    n1108,
    n1016,
    n1041
  );


  or
  g1115
  (
    n1217,
    n888,
    n981,
    n968
  );


  xnor
  g1116
  (
    n1144,
    n690,
    n952,
    n965
  );


  nor
  g1117
  (
    n1169,
    n946,
    n887,
    n1047
  );


  xnor
  g1118
  (
    n1211,
    n888,
    n1041,
    n991
  );


  nand
  g1119
  (
    n1209,
    n955,
    n889,
    n1048
  );


  nor
  g1120
  (
    n1153,
    n1125,
    n950,
    n1048
  );


  and
  g1121
  (
    n1145,
    n1124,
    n1045,
    n1046
  );


  or
  g1122
  (
    n1200,
    n939,
    n1115,
    n1132
  );


  xor
  g1123
  (
    n1140,
    n1113,
    n1124,
    n1048
  );


  and
  g1124
  (
    n1191,
    n889,
    n575,
    n886
  );


  nor
  g1125
  (
    n1206,
    n1121,
    n956,
    n935
  );


  nand
  g1126
  (
    n1188,
    n153,
    n691,
    n577
  );


  xnor
  g1127
  (
    n1214,
    n966,
    n972,
    n975
  );


  xor
  g1128
  (
    n1143,
    n690,
    n1041,
    n1116
  );


  nand
  g1129
  (
    n1157,
    n1042,
    n1046
  );


  xnor
  g1130
  (
    n1199,
    n1001,
    n1112,
    n887
  );


  nor
  g1131
  (
    n1180,
    n154,
    n970,
    n1117
  );


  xor
  g1132
  (
    n1189,
    n1122,
    n887,
    n1040
  );


  xor
  g1133
  (
    n1193,
    n934,
    n1133,
    n32
  );


  nand
  g1134
  (
    n1212,
    n957,
    n1119,
    n999
  );


  nand
  g1135
  (
    n1141,
    n1111,
    n1072,
    n1129
  );


  xnor
  g1136
  (
    n1203,
    n889,
    n1129
  );


  nor
  g1137
  (
    n1182,
    n691,
    n967,
    n1119
  );


  nand
  g1138
  (
    n1196,
    n1039,
    n1131,
    n983
  );


  xnor
  g1139
  (
    n1161,
    n692,
    n1039,
    n1128
  );


  xnor
  g1140
  (
    n1137,
    n1118,
    n1121,
    n153
  );


  xnor
  g1141
  (
    n1152,
    n1132,
    n1120,
    n1041
  );


  or
  g1142
  (
    n1210,
    n973,
    n958,
    n637
  );


  or
  g1143
  (
    n1147,
    n1000,
    n1107,
    n577
  );


  nand
  g1144
  (
    n1154,
    n1120,
    n1042,
    n945
  );


  and
  g1145
  (
    n1172,
    n1043,
    n1128,
    n888
  );


  or
  g1146
  (
    n1156,
    n1006,
    n1110,
    n1116
  );


  nor
  g1147
  (
    n1192,
    n1043,
    n888,
    n1113
  );


  nor
  g1148
  (
    n1218,
    n1130,
    n692,
    n998
  );


  nor
  g1149
  (
    n1149,
    n1124,
    n576,
    n938
  );


  xor
  g1150
  (
    n1168,
    n1013,
    n1039,
    n1119
  );


  or
  g1151
  (
    n1197,
    n971,
    n573,
    n994
  );


  or
  g1152
  (
    n1160,
    n987,
    n974,
    n1071
  );


  nand
  g1153
  (
    n1148,
    n1011,
    n1126,
    n1117
  );


  nor
  g1154
  (
    n1183,
    n1045,
    n1119,
    n1040
  );


  nor
  g1155
  (
    n1175,
    n577,
    n1118,
    n1131
  );


  xor
  g1156
  (
    n1163,
    n1116,
    n1115,
    n577
  );


  or
  g1157
  (
    n1159,
    n960,
    n1044,
    n154
  );


  xnor
  g1158
  (
    n1208,
    n692,
    n992,
    n1120
  );


  nand
  g1159
  (
    n1173,
    n886,
    n1131,
    n693
  );


  xor
  g1160
  (
    n1155,
    n1112,
    n1128,
    n1115
  );


  xor
  g1161
  (
    n1146,
    n1106,
    n1047,
    n941
  );


  xnor
  g1162
  (
    n1178,
    n1043,
    n1118,
    n997
  );


  nand
  g1163
  (
    n1150,
    n574,
    n1002,
    n1008
  );


  xor
  g1164
  (
    n1186,
    n1126,
    n1042,
    n1122
  );


  nand
  g1165
  (
    n1219,
    n1127,
    n576,
    n1112,
    n1120
  );


  xnor
  g1166
  (
    n1184,
    n639,
    n575,
    n1124,
    n1121
  );


  or
  g1167
  (
    n1221,
    n940,
    n1040,
    n691,
    n692
  );


  nand
  g1168
  (
    n1138,
    n889,
    n951,
    n1072,
    n996
  );


  nor
  g1169
  (
    n1162,
    n978,
    n1047,
    n944,
    n1072
  );


  nor
  g1170
  (
    n1187,
    n1003,
    n153,
    n932,
    n1116
  );


  nor
  g1171
  (
    n1201,
    n1125,
    n1039,
    n1110,
    n575
  );


  xnor
  g1172
  (
    n1142,
    n153,
    n953,
    n936,
    n1111
  );


  xnor
  g1173
  (
    n1220,
    n947,
    n1133,
    n990,
    n1127
  );


  xnor
  g1174
  (
    n1158,
    n1113,
    n961,
    n1009,
    n937
  );


  xnor
  g1175
  (
    n1151,
    n1125,
    n964,
    n1126,
    n576
  );


  or
  g1176
  (
    n1176,
    n1015,
    n1111,
    n948,
    n1113
  );


  nand
  g1177
  (
    n1190,
    n690,
    n887,
    n995,
    n988
  );


  nor
  g1178
  (
    n1222,
    n1040,
    n154,
    n1133,
    n1012
  );


  nor
  g1179
  (
    n1134,
    n1044,
    n1129,
    n1127,
    n962
  );


  or
  g1180
  (
    n1215,
    n32,
    n1115,
    n693,
    n942
  );


  nor
  g1181
  (
    n1136,
    n639,
    n1044,
    n1043,
    n976
  );


  xnor
  g1182
  (
    n1205,
    n977,
    n690,
    n1125,
    n985
  );


  nand
  g1183
  (
    n1202,
    n979,
    n1042,
    n693,
    n1122
  );


  nor
  g1184
  (
    n1166,
    n1114,
    n1045,
    n1126,
    n1010
  );


  and
  g1185
  (
    KeyWire_0_24,
    n1044,
    n574,
    n1131,
    n1118
  );


  or
  g1186
  (
    KeyWire_0_49,
    n1047,
    n1130,
    n1072,
    n986
  );


  and
  g1187
  (
    n1198,
    n1112,
    n1133,
    n1123,
    n1114
  );


  and
  g1188
  (
    n1167,
    n578,
    n1127,
    n1014,
    n576
  );


  xor
  g1189
  (
    n1170,
    n693,
    n989,
    n32,
    n575
  );


  buf
  g1190
  (
    n1246,
    n1136
  );


  buf
  g1191
  (
    n1255,
    n1134
  );


  not
  g1192
  (
    n1225,
    n1166
  );


  not
  g1193
  (
    n1237,
    n1152
  );


  not
  g1194
  (
    n1234,
    n1138
  );


  not
  g1195
  (
    n1244,
    n1149
  );


  buf
  g1196
  (
    n1228,
    n1162
  );


  buf
  g1197
  (
    n1235,
    n1165
  );


  buf
  g1198
  (
    n1229,
    n1167
  );


  buf
  g1199
  (
    n1241,
    n1139
  );


  buf
  g1200
  (
    n1238,
    n1150
  );


  not
  g1201
  (
    n1231,
    n1158
  );


  not
  g1202
  (
    n1247,
    n1164
  );


  not
  g1203
  (
    n1232,
    n1163
  );


  buf
  g1204
  (
    n1251,
    n1137
  );


  not
  g1205
  (
    n1245,
    n1154
  );


  not
  g1206
  (
    n1250,
    n1151
  );


  buf
  g1207
  (
    n1236,
    n1156
  );


  buf
  g1208
  (
    n1249,
    n1155
  );


  buf
  g1209
  (
    n1252,
    n1135
  );


  not
  g1210
  (
    n1224,
    n1144
  );


  buf
  g1211
  (
    n1242,
    n1140
  );


  not
  g1212
  (
    n1230,
    n1145
  );


  not
  g1213
  (
    n1253,
    n1159
  );


  buf
  g1214
  (
    n1233,
    n1148
  );


  not
  g1215
  (
    n1226,
    n1161
  );


  buf
  g1216
  (
    n1239,
    n1160
  );


  buf
  g1217
  (
    n1227,
    n1153
  );


  not
  g1218
  (
    n1223,
    n1142
  );


  buf
  g1219
  (
    n1248,
    n1146
  );


  not
  g1220
  (
    n1240,
    n1157
  );


  not
  g1221
  (
    n1254,
    n1141
  );


  not
  g1222
  (
    n1256,
    n1147
  );


  not
  g1223
  (
    n1243,
    n1143
  );


  not
  g1224
  (
    n1264,
    n1225
  );


  buf
  g1225
  (
    n1268,
    n1223
  );


  not
  g1226
  (
    n1261,
    n1225
  );


  buf
  g1227
  (
    n1258,
    n1225
  );


  buf
  g1228
  (
    n1267,
    n1223
  );


  not
  g1229
  (
    n1257,
    n1223
  );


  not
  g1230
  (
    n1263,
    n1224
  );


  not
  g1231
  (
    n1259,
    n1224
  );


  buf
  g1232
  (
    n1260,
    n1224
  );


  buf
  g1233
  (
    n1266,
    n1225
  );


  buf
  g1234
  (
    n1265,
    n1224
  );


  not
  g1235
  (
    n1262,
    n1223
  );


  buf
  g1236
  (
    n1296,
    n1263
  );


  buf
  g1237
  (
    n1273,
    n1268
  );


  not
  g1238
  (
    n1270,
    n1267
  );


  buf
  g1239
  (
    n1295,
    n156
  );


  not
  g1240
  (
    n1274,
    n1027
  );


  not
  g1241
  (
    n1293,
    n1258
  );


  or
  g1242
  (
    n1281,
    n1261,
    n1188,
    n578,
    n1260
  );


  nand
  g1243
  (
    n1272,
    n1257,
    n1263,
    n1259
  );


  nand
  g1244
  (
    n1278,
    n1191,
    n1265,
    n1190,
    n1189
  );


  or
  g1245
  (
    n1269,
    n1261,
    n1258,
    n1184,
    n155
  );


  xor
  g1246
  (
    n1286,
    n579,
    n578,
    n1263,
    n1028
  );


  xor
  g1247
  (
    n1297,
    n1187,
    n1264,
    n1174,
    n156
  );


  nor
  g1248
  (
    n1294,
    n1182,
    n579,
    n156,
    n1019
  );


  nor
  g1249
  (
    n1289,
    n1266,
    n1259,
    n155,
    n1258
  );


  or
  g1250
  (
    n1298,
    n580,
    n1260,
    n1262,
    n1169
  );


  nor
  g1251
  (
    n1277,
    n1025,
    n1178,
    n1181,
    n1268
  );


  xnor
  g1252
  (
    n1271,
    n1257,
    n1020,
    n1265,
    n1260
  );


  xor
  g1253
  (
    n1288,
    n1179,
    n1266,
    n1177,
    n1257
  );


  nand
  g1254
  (
    n1275,
    n1176,
    n1261,
    n580,
    n155
  );


  or
  g1255
  (
    n1285,
    n1265,
    n579,
    n1017,
    n1185
  );


  nand
  g1256
  (
    n1290,
    n1024,
    n1172,
    n1186,
    n1259
  );


  nor
  g1257
  (
    n1279,
    n1266,
    n1023,
    n156,
    n1170
  );


  nand
  g1258
  (
    n1292,
    n1263,
    n1266,
    n1264,
    n1018
  );


  or
  g1259
  (
    n1283,
    n1268,
    n1175,
    n1267,
    n1262
  );


  xnor
  g1260
  (
    n1291,
    n1262,
    n1021,
    n1264,
    n580
  );


  and
  g1261
  (
    n1284,
    n1173,
    n1262,
    n1265,
    n155
  );


  and
  g1262
  (
    n1276,
    n1267,
    n1168,
    n1268,
    n1171
  );


  or
  g1263
  (
    n1287,
    n578,
    n1257,
    n1180,
    n1026
  );


  xnor
  g1264
  (
    n1280,
    n1267,
    n1264,
    n1183,
    n1258
  );


  or
  g1265
  (
    n1282,
    n1261,
    n1022,
    n579,
    n1260
  );


  buf
  g1266
  (
    n1320,
    n1283
  );


  not
  g1267
  (
    n1310,
    n1295
  );


  not
  g1268
  (
    n1326,
    n1288
  );


  not
  g1269
  (
    n1306,
    n1205
  );


  not
  g1270
  (
    n1311,
    n1212
  );


  buf
  g1271
  (
    n1299,
    n1204
  );


  buf
  g1272
  (
    n1309,
    n1291
  );


  not
  g1273
  (
    n1300,
    n1294
  );


  buf
  g1274
  (
    n1301,
    n1220
  );


  not
  g1275
  (
    n1313,
    n1218
  );


  buf
  g1276
  (
    n1305,
    n1284
  );


  not
  g1277
  (
    n1302,
    n1193
  );


  buf
  g1278
  (
    n1322,
    n1210
  );


  buf
  g1279
  (
    n1325,
    n1287
  );


  buf
  g1280
  (
    n1316,
    n1272
  );


  not
  g1281
  (
    n1319,
    n1270
  );


  or
  g1282
  (
    n1321,
    n1200,
    n1285,
    n1297,
    n1194
  );


  and
  g1283
  (
    n1303,
    n1296,
    n1271,
    n1279,
    n1192
  );


  or
  g1284
  (
    n1324,
    n1207,
    n1208,
    n1216,
    n1211
  );


  xor
  g1285
  (
    KeyWire_0_0,
    n1201,
    n1202,
    n1273,
    n1209
  );


  xnor
  g1286
  (
    n1312,
    n1197,
    n1277,
    n1276,
    n1293
  );


  nand
  g1287
  (
    n1323,
    n1215,
    n1199,
    n1280,
    n1198
  );


  xnor
  g1288
  (
    n1304,
    n1275,
    n1290,
    n1217,
    n1292
  );


  or
  g1289
  (
    n1314,
    n1281,
    n1214,
    n1282,
    n1206
  );


  and
  g1290
  (
    n1315,
    n1289,
    n1296,
    n1269,
    n1286
  );


  or
  g1291
  (
    n1318,
    n1203,
    n1274,
    n1222,
    n1298
  );


  or
  g1292
  (
    n1317,
    n1221,
    n1298,
    n1195,
    n1213
  );


  nand
  g1293
  (
    n1307,
    n1278,
    n1297,
    n1196,
    n1219
  );


  buf
  g1294
  (
    n1416,
    n1254
  );


  buf
  g1295
  (
    n1372,
    n1310
  );


  buf
  g1296
  (
    n1379,
    n581
  );


  not
  g1297
  (
    n1392,
    n1303
  );


  not
  g1298
  (
    n1334,
    n1240
  );


  not
  g1299
  (
    n1432,
    n1244
  );


  not
  g1300
  (
    n1419,
    n1230
  );


  not
  g1301
  (
    n1421,
    n1245
  );


  not
  g1302
  (
    n1409,
    n1319
  );


  not
  g1303
  (
    n1433,
    n1323
  );


  not
  g1304
  (
    n1339,
    n1248
  );


  not
  g1305
  (
    n1393,
    n1245
  );


  not
  g1306
  (
    n1400,
    n1227
  );


  buf
  g1307
  (
    n1420,
    n1234
  );


  not
  g1308
  (
    n1345,
    n1243
  );


  not
  g1309
  (
    n1394,
    n1304
  );


  buf
  g1310
  (
    n1351,
    n1302
  );


  not
  g1311
  (
    n1357,
    n1319
  );


  not
  g1312
  (
    n1367,
    n1230
  );


  buf
  g1313
  (
    n1335,
    n1235
  );


  buf
  g1314
  (
    n1386,
    n1236
  );


  not
  g1315
  (
    KeyWire_0_36,
    n1302
  );


  not
  g1316
  (
    n1333,
    n1313
  );


  not
  g1317
  (
    n1346,
    n1243
  );


  not
  g1318
  (
    n1430,
    n1251
  );


  buf
  g1319
  (
    n1354,
    n1228
  );


  not
  g1320
  (
    n1329,
    n1229
  );


  not
  g1321
  (
    n1383,
    n1241
  );


  buf
  g1322
  (
    n1426,
    n1239
  );


  buf
  g1323
  (
    n1434,
    n1325
  );


  buf
  g1324
  (
    n1401,
    n1310
  );


  buf
  g1325
  (
    n1381,
    n1248
  );


  not
  g1326
  (
    n1418,
    n1244
  );


  buf
  g1327
  (
    n1413,
    n1250
  );


  buf
  g1328
  (
    n1427,
    n1311
  );


  not
  g1329
  (
    n1328,
    n1235
  );


  buf
  g1330
  (
    n1368,
    n1303
  );


  not
  g1331
  (
    n1388,
    n1324
  );


  not
  g1332
  (
    n1382,
    n1238
  );


  not
  g1333
  (
    n1438,
    n1313
  );


  not
  g1334
  (
    n1404,
    n1317
  );


  not
  g1335
  (
    n1340,
    n1228
  );


  buf
  g1336
  (
    n1391,
    n1250
  );


  buf
  g1337
  (
    n1407,
    n1308
  );


  buf
  g1338
  (
    n1402,
    n1232
  );


  not
  g1339
  (
    KeyWire_0_11,
    n1238
  );


  buf
  g1340
  (
    n1385,
    n1249
  );


  not
  g1341
  (
    n1347,
    n1239
  );


  buf
  g1342
  (
    n1437,
    n1253
  );


  buf
  g1343
  (
    n1341,
    n1325
  );


  buf
  g1344
  (
    n1355,
    n1326
  );


  buf
  g1345
  (
    n1344,
    n1301
  );


  not
  g1346
  (
    n1411,
    n1304
  );


  not
  g1347
  (
    n1406,
    n1302
  );


  buf
  g1348
  (
    n1389,
    n1321
  );


  not
  g1349
  (
    n1366,
    n1228
  );


  buf
  g1350
  (
    n1362,
    n1226
  );


  buf
  g1351
  (
    n1331,
    n1303
  );


  not
  g1352
  (
    n1364,
    n1317
  );


  not
  g1353
  (
    n1377,
    n1302
  );


  buf
  g1354
  (
    KeyWire_0_9,
    n1237
  );


  buf
  g1355
  (
    n1359,
    n1250
  );


  not
  g1356
  (
    n1425,
    n1306
  );


  not
  g1357
  (
    n1410,
    n1324
  );


  buf
  g1358
  (
    n1343,
    n1299
  );


  not
  g1359
  (
    n1374,
    n1324
  );


  not
  g1360
  (
    n1384,
    n1315
  );


  not
  g1361
  (
    n1435,
    n1309
  );


  nand
  g1362
  (
    n1405,
    n1246,
    n1307
  );


  or
  g1363
  (
    n1370,
    n1226,
    n1234,
    n582,
    n1299
  );


  xnor
  g1364
  (
    n1363,
    n1244,
    n1255,
    n1229,
    n1248
  );


  and
  g1365
  (
    n1332,
    n1247,
    n1312,
    n1311,
    n1246
  );


  and
  g1366
  (
    n1436,
    n1237,
    n1326,
    n1242,
    n1251
  );


  nor
  g1367
  (
    n1338,
    n1315,
    n1322,
    n1313,
    n1229
  );


  or
  g1368
  (
    n1376,
    n1243,
    n1243,
    n1236,
    n1308
  );


  nor
  g1369
  (
    n1412,
    n1323,
    n1256,
    n1249,
    n1232
  );


  xnor
  g1370
  (
    n1431,
    n1311,
    n1325,
    n1318,
    n1321
  );


  and
  g1371
  (
    n1336,
    n1248,
    n1239,
    n1320,
    n1315
  );


  or
  g1372
  (
    n1387,
    n1227,
    n1233,
    n1241,
    n1316
  );


  nand
  g1373
  (
    n1399,
    n1255,
    n1326,
    n1300,
    n1320
  );


  nand
  g1374
  (
    n1361,
    n1232,
    n1320,
    n1319,
    n1227
  );


  and
  g1375
  (
    n1423,
    n1229,
    n1318,
    n1252,
    n1239
  );


  xor
  g1376
  (
    n1414,
    n1301,
    n1299,
    n1305,
    n1306
  );


  xnor
  g1377
  (
    n1378,
    n1307,
    n1227,
    n1237,
    n1301
  );


  nor
  g1378
  (
    n1356,
    n1228,
    n1306,
    n1253,
    n1305
  );


  xor
  g1379
  (
    n1365,
    n1233,
    n1310,
    n1246,
    n1305
  );


  xnor
  g1380
  (
    n1360,
    n1252,
    n1310,
    n1241,
    n1251
  );


  and
  g1381
  (
    n1380,
    n581,
    n580,
    n1322,
    n1231
  );


  and
  g1382
  (
    n1337,
    n1323,
    n1326,
    n1234,
    n1230
  );


  nor
  g1383
  (
    n1403,
    n1247,
    n1315,
    n1235,
    n1249
  );


  xor
  g1384
  (
    n1408,
    n1300,
    n1254,
    n1242
  );


  xnor
  g1385
  (
    n1350,
    n1256,
    n1304,
    n1317,
    n1236
  );


  xnor
  g1386
  (
    n1390,
    n1316,
    n1247,
    n1242,
    n1231
  );


  and
  g1387
  (
    n1353,
    n1312,
    n1305,
    n581,
    n1317
  );


  xnor
  g1388
  (
    n1396,
    n1226,
    n1249,
    n1316,
    n1233
  );


  xnor
  g1389
  (
    n1397,
    n1226,
    n1256,
    n1230,
    n1240
  );


  and
  g1390
  (
    n1327,
    n1236,
    n1250,
    n1307,
    n1322
  );


  xor
  g1391
  (
    n1424,
    n1314,
    n1309,
    n1247,
    n1253
  );


  and
  g1392
  (
    n1429,
    n1318,
    n1308,
    n1231,
    n1238
  );


  or
  g1393
  (
    n1358,
    n1325,
    n1300,
    n1244,
    n1314
  );


  xnor
  g1394
  (
    n1398,
    n1241,
    n1256,
    n1309,
    n1312
  );


  xnor
  g1395
  (
    n1342,
    n1254,
    n1308,
    n1307,
    n1245
  );


  xnor
  g1396
  (
    n1349,
    n1313,
    n1231,
    n1311,
    n1237
  );


  or
  g1397
  (
    n1369,
    n1324,
    n1245,
    n1253,
    n1319
  );


  xor
  g1398
  (
    n1371,
    n1238,
    n1316,
    n1314,
    n1240
  );


  xnor
  g1399
  (
    n1428,
    n1301,
    n581,
    n1309,
    n1321
  );


  xor
  g1400
  (
    n1422,
    n1242,
    n1252,
    n1321,
    n1240
  );


  xnor
  g1401
  (
    n1373,
    n1312,
    n1300,
    n1232,
    n1314
  );


  xor
  g1402
  (
    n1415,
    n1322,
    n1252,
    n1320,
    n1233
  );


  or
  g1403
  (
    n1330,
    n1234,
    n1323,
    n1306,
    n1251
  );


  or
  g1404
  (
    n1395,
    n1299,
    n1235,
    n1303,
    n1255
  );


  or
  g1405
  (
    n1352,
    n1255,
    n1318,
    n1246,
    n1304
  );


  not
  g1406
  (
    n1834,
    n1406
  );


  buf
  g1407
  (
    n1538,
    n1417
  );


  not
  g1408
  (
    KeyWire_0_14,
    n1409
  );


  not
  g1409
  (
    n1526,
    n1366
  );


  not
  g1410
  (
    n1811,
    n1343
  );


  not
  g1411
  (
    n1780,
    n1421
  );


  buf
  g1412
  (
    n1553,
    n1333
  );


  buf
  g1413
  (
    n1674,
    n1405
  );


  buf
  g1414
  (
    n1852,
    n1431
  );


  not
  g1415
  (
    n1699,
    n1413
  );


  not
  g1416
  (
    n1530,
    n1401
  );


  not
  g1417
  (
    n1762,
    n1383
  );


  buf
  g1418
  (
    n1872,
    n1367
  );


  buf
  g1419
  (
    n1703,
    n1369
  );


  buf
  g1420
  (
    n1623,
    n1391
  );


  not
  g1421
  (
    n1876,
    n1364
  );


  buf
  g1422
  (
    n1575,
    n1352
  );


  buf
  g1423
  (
    n1464,
    n1395
  );


  buf
  g1424
  (
    n1452,
    n1431
  );


  not
  g1425
  (
    n1719,
    n1368
  );


  not
  g1426
  (
    n1552,
    n1383
  );


  buf
  g1427
  (
    n1794,
    n1358
  );


  not
  g1428
  (
    n1616,
    n1372
  );


  not
  g1429
  (
    n1563,
    n1432
  );


  not
  g1430
  (
    n1607,
    n1336
  );


  buf
  g1431
  (
    n1457,
    n1406
  );


  not
  g1432
  (
    n1493,
    n1379
  );


  buf
  g1433
  (
    n1841,
    n1426
  );


  buf
  g1434
  (
    n1716,
    n1413
  );


  not
  g1435
  (
    n1519,
    n1414
  );


  buf
  g1436
  (
    n1637,
    n1343
  );


  not
  g1437
  (
    n1684,
    n1376
  );


  not
  g1438
  (
    n1524,
    n1349
  );


  not
  g1439
  (
    n1879,
    n1428
  );


  not
  g1440
  (
    n1827,
    n582
  );


  not
  g1441
  (
    n1695,
    n1350
  );


  not
  g1442
  (
    n1448,
    n1410
  );


  buf
  g1443
  (
    KeyWire_0_56,
    n1427
  );


  not
  g1444
  (
    n1500,
    n1374
  );


  buf
  g1445
  (
    n1700,
    n1416
  );


  not
  g1446
  (
    n1686,
    n1373
  );


  not
  g1447
  (
    n1735,
    n1400
  );


  not
  g1448
  (
    n1820,
    n1404
  );


  not
  g1449
  (
    n1506,
    n1400
  );


  not
  g1450
  (
    n1786,
    n1328
  );


  buf
  g1451
  (
    n1865,
    n1361
  );


  not
  g1452
  (
    n1511,
    n1357
  );


  buf
  g1453
  (
    n1828,
    n1364
  );


  not
  g1454
  (
    n1785,
    n1397
  );


  not
  g1455
  (
    n1815,
    n1435
  );


  buf
  g1456
  (
    n1845,
    n1392
  );


  buf
  g1457
  (
    n1835,
    n1406
  );


  not
  g1458
  (
    n1647,
    n1348
  );


  not
  g1459
  (
    n1534,
    n1357
  );


  not
  g1460
  (
    n1729,
    n1347
  );


  not
  g1461
  (
    n1788,
    n1386
  );


  not
  g1462
  (
    n1471,
    n1367
  );


  not
  g1463
  (
    n1777,
    n1335
  );


  not
  g1464
  (
    n1672,
    n1341
  );


  buf
  g1465
  (
    KeyWire_0_63,
    n1386
  );


  not
  g1466
  (
    n1614,
    n1437
  );


  not
  g1467
  (
    n1767,
    n1437
  );


  buf
  g1468
  (
    n1573,
    n1396
  );


  not
  g1469
  (
    n1856,
    n1393
  );


  buf
  g1470
  (
    n1628,
    n1429
  );


  buf
  g1471
  (
    n1714,
    n1352
  );


  not
  g1472
  (
    n1510,
    n1351
  );


  buf
  g1473
  (
    n1503,
    n1336
  );


  buf
  g1474
  (
    n1861,
    n1382
  );


  not
  g1475
  (
    n1665,
    n1438
  );


  buf
  g1476
  (
    n1681,
    n1410
  );


  buf
  g1477
  (
    n1544,
    n1374
  );


  buf
  g1478
  (
    n1508,
    n1425
  );


  buf
  g1479
  (
    n1807,
    n1380
  );


  not
  g1480
  (
    n1697,
    n1346
  );


  buf
  g1481
  (
    n1869,
    n1382
  );


  not
  g1482
  (
    n1643,
    n1374
  );


  buf
  g1483
  (
    n1825,
    n1366
  );


  not
  g1484
  (
    n1504,
    n1378
  );


  buf
  g1485
  (
    n1769,
    n1393
  );


  buf
  g1486
  (
    n1758,
    n1400
  );


  buf
  g1487
  (
    n1779,
    n1369
  );


  buf
  g1488
  (
    n1617,
    n1434
  );


  not
  g1489
  (
    n1768,
    n1336
  );


  not
  g1490
  (
    n1666,
    n1404
  );


  not
  g1491
  (
    n1860,
    n1408
  );


  buf
  g1492
  (
    n1585,
    n1378
  );


  not
  g1493
  (
    n1644,
    n1333
  );


  buf
  g1494
  (
    n1596,
    n1329
  );


  buf
  g1495
  (
    n1696,
    n1357
  );


  not
  g1496
  (
    n1746,
    n1389
  );


  buf
  g1497
  (
    n1738,
    n1423
  );


  not
  g1498
  (
    n1507,
    n1397
  );


  buf
  g1499
  (
    n1718,
    n1356
  );


  buf
  g1500
  (
    n1560,
    n1434
  );


  buf
  g1501
  (
    n1734,
    n1386
  );


  not
  g1502
  (
    n1839,
    n1390
  );


  not
  g1503
  (
    n1749,
    n1338
  );


  buf
  g1504
  (
    n1489,
    n1335
  );


  not
  g1505
  (
    n1747,
    n1353
  );


  not
  g1506
  (
    n1583,
    n1385
  );


  not
  g1507
  (
    n1648,
    n1334
  );


  buf
  g1508
  (
    n1635,
    n1363
  );


  not
  g1509
  (
    n1754,
    n1429
  );


  not
  g1510
  (
    n1466,
    n1371
  );


  buf
  g1511
  (
    n1629,
    n1388
  );


  buf
  g1512
  (
    n1773,
    n1433
  );


  buf
  g1513
  (
    n1586,
    n1399
  );


  buf
  g1514
  (
    n1441,
    n1348
  );


  not
  g1515
  (
    n1578,
    n1415
  );


  buf
  g1516
  (
    n1639,
    n1378
  );


  not
  g1517
  (
    n1447,
    n1370
  );


  not
  g1518
  (
    n1883,
    n1350
  );


  buf
  g1519
  (
    n1630,
    n1365
  );


  buf
  g1520
  (
    n1606,
    n1355
  );


  not
  g1521
  (
    KeyWire_0_57,
    n1342
  );


  buf
  g1522
  (
    n1701,
    n1378
  );


  not
  g1523
  (
    n1725,
    n1385
  );


  buf
  g1524
  (
    n1540,
    n1403
  );


  not
  g1525
  (
    n1581,
    n1375
  );


  buf
  g1526
  (
    n1481,
    n1393
  );


  not
  g1527
  (
    n1821,
    n582
  );


  buf
  g1528
  (
    n1531,
    n1339
  );


  buf
  g1529
  (
    n1631,
    n1425
  );


  not
  g1530
  (
    n1473,
    n1366
  );


  buf
  g1531
  (
    n1659,
    n1337
  );


  not
  g1532
  (
    n1536,
    n1364
  );


  buf
  g1533
  (
    n1576,
    n1433
  );


  buf
  g1534
  (
    n1474,
    n1415
  );


  not
  g1535
  (
    n1569,
    n1338
  );


  buf
  g1536
  (
    n1812,
    n1379
  );


  not
  g1537
  (
    n1771,
    n1422
  );


  buf
  g1538
  (
    n1626,
    n1380
  );


  not
  g1539
  (
    n1634,
    n1360
  );


  not
  g1540
  (
    n1527,
    n1391
  );


  not
  g1541
  (
    n1761,
    n1330
  );


  buf
  g1542
  (
    KeyWire_0_31,
    n1411
  );


  not
  g1543
  (
    KeyWire_0_59,
    n1377
  );


  buf
  g1544
  (
    n1671,
    n1342
  );


  buf
  g1545
  (
    n1525,
    n1346
  );


  buf
  g1546
  (
    n1817,
    n1406
  );


  buf
  g1547
  (
    n1810,
    n1412
  );


  buf
  g1548
  (
    n1662,
    n1387
  );


  not
  g1549
  (
    n1599,
    n1375
  );


  not
  g1550
  (
    n1642,
    n1436
  );


  buf
  g1551
  (
    n1833,
    n1332
  );


  buf
  g1552
  (
    n1698,
    n1338
  );


  not
  g1553
  (
    n1756,
    n1377
  );


  not
  g1554
  (
    n1819,
    n1343
  );


  buf
  g1555
  (
    n1477,
    n1438
  );


  not
  g1556
  (
    n1640,
    n1375
  );


  buf
  g1557
  (
    n1783,
    n1341
  );


  buf
  g1558
  (
    n1522,
    n1379
  );


  buf
  g1559
  (
    n1866,
    n1376
  );


  not
  g1560
  (
    n1731,
    n1430
  );


  buf
  g1561
  (
    n1801,
    n1368
  );


  buf
  g1562
  (
    n1562,
    n1408
  );


  not
  g1563
  (
    n1479,
    n1423
  );


  buf
  g1564
  (
    n1533,
    n1412
  );


  buf
  g1565
  (
    n1615,
    n1438
  );


  buf
  g1566
  (
    n1791,
    n1347
  );


  buf
  g1567
  (
    n1789,
    n1388
  );


  not
  g1568
  (
    n1884,
    n1427
  );


  not
  g1569
  (
    n1470,
    n1384
  );


  buf
  g1570
  (
    n1882,
    n1353
  );


  buf
  g1571
  (
    n1649,
    n1404
  );


  not
  g1572
  (
    n1655,
    n1392
  );


  buf
  g1573
  (
    n1458,
    n1434
  );


  buf
  g1574
  (
    n1676,
    n1349
  );


  not
  g1575
  (
    n1838,
    n1404
  );


  not
  g1576
  (
    n1497,
    n1354
  );


  not
  g1577
  (
    n1487,
    n1423
  );


  buf
  g1578
  (
    n1751,
    n1365
  );


  buf
  g1579
  (
    n1546,
    n1425
  );


  buf
  g1580
  (
    n1822,
    n1381
  );


  not
  g1581
  (
    n1814,
    n1387
  );


  not
  g1582
  (
    n1736,
    n1360
  );


  not
  g1583
  (
    n1483,
    n1420
  );


  not
  g1584
  (
    n1502,
    n1374
  );


  buf
  g1585
  (
    n1661,
    n1424
  );


  not
  g1586
  (
    n1439,
    n1363
  );


  buf
  g1587
  (
    n1803,
    n1432
  );


  not
  g1588
  (
    n1664,
    n1410
  );


  not
  g1589
  (
    n1455,
    n1419
  );


  not
  g1590
  (
    n1463,
    n1335
  );


  not
  g1591
  (
    n1728,
    n1345
  );


  not
  g1592
  (
    n1885,
    n1426
  );


  buf
  g1593
  (
    n1873,
    n1420
  );


  not
  g1594
  (
    n1867,
    n1409
  );


  not
  g1595
  (
    n1543,
    n1399
  );


  buf
  g1596
  (
    n1831,
    n1401
  );


  not
  g1597
  (
    n1516,
    n1362
  );


  not
  g1598
  (
    n1495,
    n1428
  );


  not
  g1599
  (
    n1529,
    n1422
  );


  not
  g1600
  (
    n1793,
    n1409
  );


  buf
  g1601
  (
    n1491,
    n1422
  );


  buf
  g1602
  (
    n1485,
    n1424
  );


  not
  g1603
  (
    n1750,
    n1418
  );


  not
  g1604
  (
    n1871,
    n1395
  );


  not
  g1605
  (
    n1778,
    n1398
  );


  buf
  g1606
  (
    n1826,
    n1424
  );


  buf
  g1607
  (
    n1624,
    n1389
  );


  not
  g1608
  (
    n1702,
    n1329
  );


  buf
  g1609
  (
    n1796,
    n1349
  );


  buf
  g1610
  (
    n1570,
    n1417
  );


  not
  g1611
  (
    n1480,
    n1383
  );


  not
  g1612
  (
    n1737,
    n1412
  );


  buf
  g1613
  (
    n1782,
    n1387
  );


  buf
  g1614
  (
    n1490,
    n1392
  );


  not
  g1615
  (
    n1757,
    n1368
  );


  not
  g1616
  (
    n1805,
    n1344
  );


  not
  g1617
  (
    n1446,
    n1384
  );


  not
  g1618
  (
    KeyWire_0_55,
    n1411
  );


  not
  g1619
  (
    n1741,
    n1429
  );


  buf
  g1620
  (
    n1707,
    n1387
  );


  not
  g1621
  (
    n1870,
    n1358
  );


  not
  g1622
  (
    n1775,
    n1412
  );


  not
  g1623
  (
    n1680,
    n1428
  );


  buf
  g1624
  (
    n1848,
    n1334
  );


  not
  g1625
  (
    n1611,
    n1395
  );


  not
  g1626
  (
    KeyWire_0_3,
    n1436
  );


  not
  g1627
  (
    n1462,
    n1438
  );


  buf
  g1628
  (
    n1613,
    n1411
  );


  not
  g1629
  (
    n1740,
    n1356
  );


  not
  g1630
  (
    n1465,
    n1328
  );


  not
  g1631
  (
    n1857,
    n1336
  );


  not
  g1632
  (
    n1565,
    n1376
  );


  buf
  g1633
  (
    n1598,
    n1390
  );


  buf
  g1634
  (
    n1484,
    n1339
  );


  buf
  g1635
  (
    n1597,
    n1390
  );


  buf
  g1636
  (
    n1693,
    n1373
  );


  not
  g1637
  (
    n1830,
    n1337
  );


  not
  g1638
  (
    n1667,
    n1382
  );


  buf
  g1639
  (
    n1668,
    n1417
  );


  buf
  g1640
  (
    n1711,
    n1409
  );


  buf
  g1641
  (
    n1787,
    n1373
  );


  not
  g1642
  (
    n1733,
    n1411
  );


  not
  g1643
  (
    n1498,
    n1432
  );


  buf
  g1644
  (
    n1774,
    n1399
  );


  not
  g1645
  (
    n1475,
    n1418
  );


  buf
  g1646
  (
    n1704,
    n1342
  );


  not
  g1647
  (
    KeyWire_0_30,
    n1365
  );


  not
  g1648
  (
    n1878,
    n1431
  );


  buf
  g1649
  (
    n1853,
    n1390
  );


  not
  g1650
  (
    n1460,
    n1349
  );


  buf
  g1651
  (
    n1548,
    n1405
  );


  buf
  g1652
  (
    n1632,
    n1354
  );


  not
  g1653
  (
    n1843,
    n1331
  );


  buf
  g1654
  (
    n1713,
    n1413
  );


  not
  g1655
  (
    n1712,
    n1396
  );


  not
  g1656
  (
    n1658,
    n1328
  );


  buf
  g1657
  (
    n1881,
    n1421
  );


  buf
  g1658
  (
    n1646,
    n1407
  );


  not
  g1659
  (
    n1772,
    n1350
  );


  buf
  g1660
  (
    n1654,
    n1428
  );


  buf
  g1661
  (
    n1603,
    n1340
  );


  buf
  g1662
  (
    n1641,
    n1424
  );


  not
  g1663
  (
    n1804,
    n1379
  );


  not
  g1664
  (
    n1673,
    n1334
  );


  not
  g1665
  (
    n1625,
    n1430
  );


  not
  g1666
  (
    n1610,
    n1353
  );


  buf
  g1667
  (
    n1561,
    n1430
  );


  buf
  g1668
  (
    n1663,
    n1418
  );


  buf
  g1669
  (
    n1816,
    n1344
  );


  buf
  g1670
  (
    n1842,
    n1392
  );


  buf
  g1671
  (
    n1584,
    n1415
  );


  buf
  g1672
  (
    n1592,
    n1350
  );


  buf
  g1673
  (
    n1564,
    n1382
  );


  not
  g1674
  (
    KeyWire_0_12,
    n582
  );


  buf
  g1675
  (
    n1795,
    n1352
  );


  not
  g1676
  (
    n1743,
    n1398
  );


  buf
  g1677
  (
    n1809,
    n1344
  );


  buf
  g1678
  (
    n1798,
    n1369
  );


  buf
  g1679
  (
    n1579,
    n1351
  );


  not
  g1680
  (
    n1720,
    n1344
  );


  not
  g1681
  (
    n1679,
    n1436
  );


  buf
  g1682
  (
    n1567,
    n1361
  );


  buf
  g1683
  (
    n1745,
    n1357
  );


  not
  g1684
  (
    n1566,
    n1397
  );


  not
  g1685
  (
    n1532,
    n1348
  );


  not
  g1686
  (
    n1727,
    n1414
  );


  buf
  g1687
  (
    n1453,
    n1363
  );


  not
  g1688
  (
    n1687,
    n1407
  );


  not
  g1689
  (
    n1513,
    n1340
  );


  not
  g1690
  (
    n1515,
    n1337
  );


  buf
  g1691
  (
    n1808,
    n1327
  );


  buf
  g1692
  (
    n1823,
    n1333
  );


  buf
  g1693
  (
    n1709,
    n1347
  );


  not
  g1694
  (
    n1850,
    n1419
  );


  not
  g1695
  (
    n1549,
    n1359
  );


  buf
  g1696
  (
    n1660,
    n1365
  );


  buf
  g1697
  (
    n1724,
    n1381
  );


  buf
  g1698
  (
    n1656,
    n1346
  );


  buf
  g1699
  (
    n1689,
    n1354
  );


  not
  g1700
  (
    n1442,
    n1396
  );


  not
  g1701
  (
    n1645,
    n1407
  );


  buf
  g1702
  (
    n1691,
    n1345
  );


  not
  g1703
  (
    n1550,
    n1327
  );


  not
  g1704
  (
    n1554,
    n1360
  );


  buf
  g1705
  (
    n1517,
    n1394
  );


  not
  g1706
  (
    n1717,
    n1394
  );


  not
  g1707
  (
    n1675,
    n1384
  );


  buf
  g1708
  (
    n1682,
    n1435
  );


  not
  g1709
  (
    KeyWire_0_32,
    n1370
  );


  not
  g1710
  (
    n1705,
    n1372
  );


  not
  g1711
  (
    n1595,
    n1389
  );


  buf
  g1712
  (
    n1467,
    n1394
  );


  not
  g1713
  (
    n1764,
    n1422
  );


  buf
  g1714
  (
    n1440,
    n1369
  );


  not
  g1715
  (
    n1708,
    n1435
  );


  not
  g1716
  (
    n1763,
    n1391
  );


  buf
  g1717
  (
    n1582,
    n1335
  );


  buf
  g1718
  (
    n1706,
    n1398
  );


  not
  g1719
  (
    n1577,
    n1381
  );


  not
  g1720
  (
    n1753,
    n1381
  );


  buf
  g1721
  (
    n1685,
    n1327
  );


  buf
  g1722
  (
    n1723,
    n1414
  );


  not
  g1723
  (
    n1557,
    n1356
  );


  buf
  g1724
  (
    n1818,
    n1343
  );


  not
  g1725
  (
    n1730,
    n1435
  );


  not
  g1726
  (
    n1692,
    n1434
  );


  buf
  g1727
  (
    n1690,
    n1332
  );


  not
  g1728
  (
    n1555,
    n1426
  );


  buf
  g1729
  (
    n1744,
    n1415
  );


  buf
  g1730
  (
    n1609,
    n1345
  );


  not
  g1731
  (
    n1461,
    n1380
  );


  not
  g1732
  (
    n1478,
    n1341
  );


  buf
  g1733
  (
    n1541,
    n1416
  );


  not
  g1734
  (
    n1784,
    n1358
  );


  not
  g1735
  (
    n1636,
    n1403
  );


  buf
  g1736
  (
    n1499,
    n1427
  );


  not
  g1737
  (
    KeyWire_0_15,
    n1361
  );


  not
  g1738
  (
    n1612,
    n1385
  );


  not
  g1739
  (
    n1688,
    n1345
  );


  not
  g1740
  (
    n1605,
    n1433
  );


  not
  g1741
  (
    n1792,
    n1391
  );


  not
  g1742
  (
    n1755,
    n1383
  );


  not
  g1743
  (
    n1851,
    n1405
  );


  buf
  g1744
  (
    n1523,
    n1388
  );


  buf
  g1745
  (
    n1694,
    n1416
  );


  buf
  g1746
  (
    n1622,
    n1340
  );


  buf
  g1747
  (
    n1670,
    n1359
  );


  not
  g1748
  (
    n1608,
    n1396
  );


  not
  g1749
  (
    n1618,
    n1333
  );


  not
  g1750
  (
    n1535,
    n1362
  );


  buf
  g1751
  (
    n1486,
    n1376
  );


  buf
  g1752
  (
    n1571,
    n1351
  );


  buf
  g1753
  (
    n1514,
    n1370
  );


  buf
  g1754
  (
    n1501,
    n1355
  );


  not
  g1755
  (
    n1594,
    n1360
  );


  not
  g1756
  (
    n1589,
    n1332
  );


  buf
  g1757
  (
    n1837,
    n1371
  );


  not
  g1758
  (
    n1859,
    n1366
  );


  not
  g1759
  (
    n1726,
    n1359
  );


  not
  g1760
  (
    n1602,
    n1354
  );


  not
  g1761
  (
    n1651,
    n1359
  );


  buf
  g1762
  (
    n1669,
    n1364
  );


  not
  g1763
  (
    n1844,
    n1358
  );


  not
  g1764
  (
    n1721,
    n1339
  );


  not
  g1765
  (
    n1505,
    n1423
  );


  not
  g1766
  (
    n1568,
    n1384
  );


  not
  g1767
  (
    n1829,
    n1371
  );


  not
  g1768
  (
    n1677,
    n1397
  );


  buf
  g1769
  (
    n1528,
    n1429
  );


  buf
  g1770
  (
    n1864,
    n1401
  );


  not
  g1771
  (
    n1551,
    n1405
  );


  not
  g1772
  (
    n1824,
    n1421
  );


  not
  g1773
  (
    KeyWire_0_53,
    n1408
  );


  not
  g1774
  (
    n1765,
    n1371
  );


  not
  g1775
  (
    n1542,
    n1330
  );


  buf
  g1776
  (
    n1444,
    n1418
  );


  buf
  g1777
  (
    n1521,
    n1419
  );


  not
  g1778
  (
    n1619,
    n1402
  );


  not
  g1779
  (
    n1877,
    n1377
  );


  buf
  g1780
  (
    n1678,
    n1337
  );


  buf
  g1781
  (
    n1862,
    n1340
  );


  not
  g1782
  (
    n1715,
    n1375
  );


  not
  g1783
  (
    n1847,
    n1386
  );


  not
  g1784
  (
    n1512,
    n1372
  );


  not
  g1785
  (
    n1509,
    n1413
  );


  buf
  g1786
  (
    n1806,
    n1329
  );


  not
  g1787
  (
    n1638,
    n1367
  );


  not
  g1788
  (
    n1593,
    n1332
  );


  not
  g1789
  (
    n1621,
    n1426
  );


  not
  g1790
  (
    n1496,
    n1420
  );


  not
  g1791
  (
    n1781,
    n1433
  );


  not
  g1792
  (
    n1802,
    n1402
  );


  not
  g1793
  (
    n1836,
    n1377
  );


  not
  g1794
  (
    n1739,
    n1427
  );


  not
  g1795
  (
    n1732,
    n1399
  );


  not
  g1796
  (
    n1652,
    n1334
  );


  buf
  g1797
  (
    n1492,
    n1400
  );


  not
  g1798
  (
    n1875,
    n1437
  );


  buf
  g1799
  (
    n1683,
    n1394
  );


  buf
  g1800
  (
    n1574,
    n1356
  );


  buf
  g1801
  (
    n1601,
    n1432
  );


  buf
  g1802
  (
    n1547,
    n1408
  );


  not
  g1803
  (
    n1545,
    n1351
  );


  not
  g1804
  (
    n1494,
    n1327
  );


  buf
  g1805
  (
    n1874,
    n1361
  );


  not
  g1806
  (
    n1760,
    n1430
  );


  buf
  g1807
  (
    n1854,
    n1330
  );


  not
  g1808
  (
    n1587,
    n1355
  );


  buf
  g1809
  (
    n1443,
    n1431
  );


  buf
  g1810
  (
    n1742,
    n1437
  );


  buf
  g1811
  (
    n1858,
    n1407
  );


  not
  g1812
  (
    n1653,
    n1398
  );


  buf
  g1813
  (
    n1539,
    n1425
  );


  buf
  g1814
  (
    n1520,
    n1393
  );


  buf
  g1815
  (
    n1759,
    n1372
  );


  not
  g1816
  (
    n1620,
    n1331
  );


  buf
  g1817
  (
    n1600,
    n1373
  );


  not
  g1818
  (
    n1770,
    n1331
  );


  not
  g1819
  (
    n1482,
    n1388
  );


  buf
  g1820
  (
    n1445,
    n1380
  );


  buf
  g1821
  (
    n1748,
    n1385
  );


  not
  g1822
  (
    n1450,
    n1403
  );


  not
  g1823
  (
    n1832,
    n1402
  );


  not
  g1824
  (
    n1558,
    n1353
  );


  buf
  g1825
  (
    n1799,
    n1414
  );


  buf
  g1826
  (
    n1868,
    n1368
  );


  not
  g1827
  (
    n1572,
    n1420
  );


  buf
  g1828
  (
    n1556,
    n1395
  );


  not
  g1829
  (
    n1488,
    n1339
  );


  not
  g1830
  (
    n1468,
    n1342
  );


  not
  g1831
  (
    n1604,
    n1330
  );


  buf
  g1832
  (
    n1590,
    n1352
  );


  buf
  g1833
  (
    n1454,
    n1417
  );


  buf
  g1834
  (
    n1650,
    n1416
  );


  buf
  g1835
  (
    n1518,
    n1341
  );


  not
  g1836
  (
    n1846,
    n1346
  );


  buf
  g1837
  (
    n1456,
    n1401
  );


  buf
  g1838
  (
    KeyWire_0_20,
    n1403
  );


  buf
  g1839
  (
    n1840,
    n1421
  );


  buf
  g1840
  (
    n1591,
    n1367
  );


  buf
  g1841
  (
    n1588,
    n1410
  );


  buf
  g1842
  (
    n1710,
    n1328
  );


  buf
  g1843
  (
    n1537,
    n1389
  );


  not
  g1844
  (
    n1722,
    n1436
  );


  buf
  g1845
  (
    n1776,
    n1347
  );


  buf
  g1846
  (
    n1559,
    n1362
  );


  buf
  g1847
  (
    n1797,
    n1355
  );


  buf
  g1848
  (
    n1657,
    n1338
  );


  buf
  g1849
  (
    n1627,
    n1329
  );


  buf
  g1850
  (
    n1476,
    n1362
  );


  nand
  g1851
  (
    n1880,
    n1402,
    n1419
  );


  xnor
  g1852
  (
    n1863,
    n1370,
    n1331,
    n1363,
    n1348
  );


  nor
  g1853
  (
    KeyWire_0_10,
    n1699,
    n1471,
    n1509,
    n1607
  );


  nand
  g1854
  (
    n1968,
    n1756,
    n1750,
    n1870,
    n1741
  );


  xnor
  g1855
  (
    n1914,
    n1794,
    n1589,
    n1723,
    n1580
  );


  xnor
  g1856
  (
    n1900,
    n1582,
    n1641,
    n1883,
    n1553
  );


  or
  g1857
  (
    n1997,
    n1830,
    n1653,
    n1876,
    n1591
  );


  xor
  g1858
  (
    n1910,
    n1604,
    n1490,
    n1752,
    n1686
  );


  or
  g1859
  (
    n1896,
    n1640,
    n1719,
    n1611,
    n1491
  );


  xnor
  g1860
  (
    n1886,
    n1487,
    n1687,
    n1838,
    n1868
  );


  xnor
  g1861
  (
    n1993,
    n1709,
    n1803,
    n1694,
    n1657
  );


  and
  g1862
  (
    n1911,
    n1871,
    n1873,
    n1726,
    n1579
  );


  xnor
  g1863
  (
    n1972,
    n1880,
    n1691,
    n1720,
    n1677
  );


  and
  g1864
  (
    n1925,
    n1557,
    n1674,
    n1618,
    n1525
  );


  or
  g1865
  (
    n1929,
    n1476,
    n1587,
    n1474,
    n1764
  );


  nand
  g1866
  (
    n1894,
    n1624,
    n1465,
    n1682,
    n1565
  );


  nor
  g1867
  (
    n1985,
    n1548,
    n1777,
    n1533,
    n1772
  );


  or
  g1868
  (
    n1967,
    n1608,
    n1658,
    n1762,
    n1732
  );


  nand
  g1869
  (
    n1978,
    n1669,
    n1737,
    n1483,
    n1600
  );


  and
  g1870
  (
    n1928,
    n1603,
    n1859,
    n1526,
    n1494
  );


  nor
  g1871
  (
    n1952,
    n1828,
    n1638,
    n1824,
    n1452
  );


  or
  g1872
  (
    n1927,
    n1552,
    n1554,
    n1724,
    n1633
  );


  or
  g1873
  (
    n1913,
    n1754,
    n1708,
    n1831,
    n1662
  );


  nand
  g1874
  (
    n1956,
    n1468,
    n1462,
    n1853,
    n1498
  );


  nand
  g1875
  (
    n1909,
    n1747,
    n1761,
    n1558,
    n1793
  );


  nand
  g1876
  (
    n1986,
    n1703,
    n1775,
    n1728,
    n1593
  );


  nor
  g1877
  (
    n1970,
    n1616,
    n1501,
    n1517,
    n1855
  );


  xnor
  g1878
  (
    n1976,
    n1632,
    n1734,
    n1510,
    n1837
  );


  nor
  g1879
  (
    n1938,
    n1845,
    n1518,
    n1820,
    n1811
  );


  xnor
  g1880
  (
    n1994,
    n1527,
    n1697,
    n1626,
    n1701
  );


  nor
  g1881
  (
    n1947,
    n1692,
    n1778,
    n1693,
    n1759
  );


  xnor
  g1882
  (
    n1966,
    n1573,
    n1666,
    n1808,
    n1874
  );


  xor
  g1883
  (
    n1901,
    n1758,
    n1696,
    n1451,
    n1771
  );


  and
  g1884
  (
    n1948,
    n1672,
    n1800,
    n1722,
    n1541
  );


  nand
  g1885
  (
    n1954,
    n1536,
    n1877,
    n1664,
    n1866
  );


  xnor
  g1886
  (
    n1916,
    n1520,
    n1839,
    n1738,
    n1574
  );


  xnor
  g1887
  (
    n1899,
    n1826,
    n1569,
    n1576,
    n1715
  );


  nand
  g1888
  (
    n1971,
    n1822,
    n1727,
    n1511,
    n1757
  );


  nand
  g1889
  (
    n1939,
    n1702,
    n1862,
    n1856,
    n1879
  );


  nor
  g1890
  (
    n1962,
    n1571,
    n1532,
    n1622,
    n1537
  );


  xnor
  g1891
  (
    n1991,
    n1502,
    n1599,
    n1755,
    n1524
  );


  xor
  g1892
  (
    n1919,
    n1647,
    n1543,
    n1790,
    n1765
  );


  and
  g1893
  (
    n1924,
    n1883,
    n1463,
    n1514,
    n1745
  );


  or
  g1894
  (
    KeyWire_0_46,
    n1516,
    n1884,
    n1551,
    n1780
  );


  and
  g1895
  (
    n1958,
    n1566,
    n1508,
    n1560,
    n1546
  );


  nor
  g1896
  (
    n1969,
    n1817,
    n1807,
    n1716,
    n1717
  );


  xor
  g1897
  (
    n1979,
    n1482,
    n1739,
    n1766,
    n1467
  );


  xor
  g1898
  (
    n1964,
    n1875,
    n1815,
    n1583,
    n1749
  );


  or
  g1899
  (
    n1988,
    n1499,
    n1595,
    n1504,
    n1735
  );


  or
  g1900
  (
    n1935,
    n1818,
    n1782,
    n1473,
    n1631
  );


  and
  g1901
  (
    n1918,
    n1788,
    n1547,
    n1821,
    n1832
  );


  or
  g1902
  (
    KeyWire_0_44,
    n1481,
    n1833,
    n1492,
    n1522
  );


  xnor
  g1903
  (
    n1960,
    n1614,
    n1721,
    n1661,
    n1835
  );


  nand
  g1904
  (
    n1921,
    n1515,
    n1671,
    n1834,
    n1564
  );


  nor
  g1905
  (
    n1892,
    n1455,
    n1884,
    n1464,
    n1812
  );


  or
  g1906
  (
    n1915,
    n1779,
    n1549,
    n1531,
    n1851
  );


  nand
  g1907
  (
    n1905,
    n1823,
    n1848,
    n1729,
    n1810
  );


  and
  g1908
  (
    n1961,
    n1841,
    n1581,
    n1705,
    n1470
  );


  xnor
  g1909
  (
    n1973,
    n1654,
    n1453,
    n1500,
    n1883
  );


  nand
  g1910
  (
    n1941,
    n1519,
    n1733,
    n1506,
    n1784
  );


  xor
  g1911
  (
    n1995,
    n1769,
    n1836,
    n1594,
    n1450
  );


  nor
  g1912
  (
    n1917,
    n1539,
    n1740,
    n1863,
    n1528
  );


  xnor
  g1913
  (
    n1946,
    n1459,
    n1707,
    n1885,
    n1458
  );


  or
  g1914
  (
    n1982,
    n1713,
    n1454,
    n1685,
    n1477
  );


  nand
  g1915
  (
    n1907,
    n1665,
    n1645,
    n1844,
    n1760
  );


  nor
  g1916
  (
    n1898,
    n1663,
    n1885,
    n1773,
    n1563
  );


  or
  g1917
  (
    n1992,
    n1601,
    n1646,
    n1598,
    n1688
  );


  xor
  g1918
  (
    n1951,
    n1489,
    n1689,
    n1829,
    n1783
  );


  or
  g1919
  (
    n1904,
    n1683,
    n1753,
    n1725,
    n1639
  );


  xor
  g1920
  (
    n1959,
    n1858,
    n1860,
    n1854,
    n1555
  );


  or
  g1921
  (
    n1932,
    n1449,
    n1628,
    n1781,
    n1636
  );


  nand
  g1922
  (
    n1981,
    n1675,
    n1610,
    n1710,
    n1776
  );


  nand
  g1923
  (
    n1944,
    n1602,
    n1751,
    n1568,
    n1488
  );


  and
  g1924
  (
    n1950,
    n1679,
    n1774,
    n1670,
    n1617
  );


  xor
  g1925
  (
    n1903,
    n1507,
    n1621,
    n1486,
    n1570
  );


  nand
  g1926
  (
    n1888,
    n1649,
    n1630,
    n1872,
    n1544
  );


  or
  g1927
  (
    n1983,
    n1612,
    n1770,
    n1850,
    n1840
  );


  xor
  g1928
  (
    n1963,
    n1609,
    n1816,
    n1586,
    n1673
  );


  and
  g1929
  (
    n1955,
    n1534,
    n1575,
    n1786,
    n1503
  );


  xnor
  g1930
  (
    n1920,
    n1648,
    n1561,
    n1643,
    n1712
  );


  xor
  g1931
  (
    n1922,
    n1495,
    n1825,
    n1796,
    n1843
  );


  or
  g1932
  (
    n1934,
    n1813,
    n1513,
    n1852,
    n1613
  );


  and
  g1933
  (
    n1953,
    n1698,
    n1572,
    n1521,
    n1731
  );


  xor
  g1934
  (
    n1937,
    n1883,
    n1791,
    n1676,
    n1884
  );


  xnor
  g1935
  (
    n1931,
    n1809,
    n1655,
    n1744,
    n1827
  );


  or
  g1936
  (
    n1942,
    n1885,
    n1512,
    n1627,
    n1785
  );


  xor
  g1937
  (
    n1984,
    n1885,
    n1804,
    n1606,
    n1882
  );


  or
  g1938
  (
    n1945,
    n1681,
    n1478,
    n1448,
    n1730
  );


  nor
  g1939
  (
    n1980,
    n1629,
    n1846,
    n1805,
    n1748
  );


  xnor
  g1940
  (
    n1940,
    n1615,
    n1475,
    n1801,
    n1585
  );


  and
  g1941
  (
    n1974,
    n1667,
    n1484,
    n1461,
    n1651
  );


  nor
  g1942
  (
    n1895,
    n1590,
    n1619,
    n1540,
    n1718
  );


  xnor
  g1943
  (
    n1906,
    n1704,
    n1559,
    n1881,
    n1861
  );


  xor
  g1944
  (
    n1975,
    n1789,
    n1695,
    n1625,
    n1869
  );


  xnor
  g1945
  (
    n1930,
    n1597,
    n1497,
    n1798,
    n1634
  );


  and
  g1946
  (
    n1908,
    n1523,
    n1678,
    n1592,
    n1819
  );


  nor
  g1947
  (
    n1923,
    n1469,
    n1652,
    n1605,
    n1711
  );


  or
  g1948
  (
    n1887,
    n1797,
    n1505,
    n1865,
    n1644
  );


  nor
  g1949
  (
    n1891,
    n1746,
    n1690,
    n1457,
    n1496
  );


  xnor
  g1950
  (
    n1926,
    n1562,
    n1700,
    n1787,
    n1806
  );


  xnor
  g1951
  (
    n1989,
    n1447,
    n1656,
    n1706,
    n1642
  );


  xor
  g1952
  (
    n1889,
    n1795,
    n1479,
    n1714,
    n1736
  );


  xnor
  g1953
  (
    n1890,
    n1542,
    n1842,
    n1460,
    n1680
  );


  and
  g1954
  (
    n1902,
    n1635,
    n1485,
    n1660,
    n1847
  );


  nor
  g1955
  (
    n1936,
    n1743,
    n1637,
    n1867,
    n1814
  );


  xor
  g1956
  (
    n1949,
    n1456,
    n1567,
    n1742,
    n1668
  );


  nand
  g1957
  (
    n1897,
    n1623,
    n1857,
    n1556,
    n1472
  );


  xor
  g1958
  (
    n1893,
    n1650,
    n1545,
    n1466,
    n1529
  );


  or
  g1959
  (
    n1912,
    n1577,
    n1659,
    n1767,
    n1493
  );


  nand
  g1960
  (
    KeyWire_0_7,
    n1535,
    n1768,
    n1849,
    n1620
  );


  nand
  g1961
  (
    n1987,
    n1802,
    n1864,
    n1799,
    n1480
  );


  xor
  g1962
  (
    n1977,
    n1588,
    n1538,
    n1584,
    n1550
  );


  or
  g1963
  (
    n1965,
    n1878,
    n1578,
    n1763,
    n1596
  );


  xor
  g1964
  (
    n1996,
    n1792,
    n1884,
    n1684,
    n1530
  );


  or
  g1965
  (
    n1998,
    n1899,
    n1938,
    n1948,
    n1963
  );


  xor
  g1966
  (
    n1999,
    n1940,
    n1901,
    n1945,
    n1993
  );


  or
  g1967
  (
    n2002,
    n1928,
    n1966,
    n1990,
    n1905
  );


  nand
  g1968
  (
    n2020,
    n1922,
    n1958,
    n1918,
    n1925
  );


  xor
  g1969
  (
    n2022,
    n1906,
    n1950,
    n1980,
    n1991
  );


  xnor
  g1970
  (
    n2024,
    n1944,
    n1894,
    n1976,
    n1939
  );


  and
  g1971
  (
    n2017,
    n1974,
    n1971,
    n1888,
    n1926
  );


  nor
  g1972
  (
    n2005,
    n1979,
    n1962,
    n1947,
    n1912
  );


  or
  g1973
  (
    n2021,
    n1931,
    n1903,
    n1985,
    n1916
  );


  xnor
  g1974
  (
    n2025,
    n1951,
    n1890,
    n1933,
    n1970
  );


  nor
  g1975
  (
    n2000,
    n1967,
    n1889,
    n1913,
    n1937
  );


  nor
  g1976
  (
    n2001,
    n1992,
    n1989,
    n1911,
    n1914
  );


  or
  g1977
  (
    n2018,
    n1952,
    n1981,
    n1886,
    n1900
  );


  nand
  g1978
  (
    n2003,
    n1920,
    n1978,
    n1996,
    n1935
  );


  nand
  g1979
  (
    n2004,
    n1910,
    n1904,
    n1960,
    n1927
  );


  nor
  g1980
  (
    n2015,
    n1924,
    n1892,
    n1994,
    n1983
  );


  and
  g1981
  (
    n2010,
    n1984,
    n1929,
    n1977,
    n1915
  );


  and
  g1982
  (
    n2007,
    n1988,
    n1995,
    n1955,
    n1923
  );


  xor
  g1983
  (
    n2006,
    n1941,
    n1987,
    n1954,
    n1896
  );


  nor
  g1984
  (
    n2019,
    n1893,
    n1997,
    n1959,
    n1897
  );


  nor
  g1985
  (
    n2023,
    n1953,
    n1930,
    n1895,
    n1956
  );


  or
  g1986
  (
    n2011,
    n1908,
    n1934,
    n1887,
    n1949
  );


  nand
  g1987
  (
    n2013,
    n1936,
    n1921,
    n1902,
    n1973
  );


  nand
  g1988
  (
    n2016,
    n1986,
    n1907,
    n1946,
    n1961
  );


  and
  g1989
  (
    n2009,
    n1972,
    n1969,
    n1957,
    n1919
  );


  and
  g1990
  (
    n2008,
    n1968,
    n1943,
    n1917,
    n1965
  );


  nor
  g1991
  (
    n2012,
    n1932,
    n1898,
    n1942,
    n1891
  );


  xnor
  g1992
  (
    n2014,
    n1982,
    n1964,
    n1909,
    n1975
  );


  or
  g1993
  (
    n2027,
    n2008,
    n2019,
    n2004,
    n2003
  );


  nand
  g1994
  (
    n2030,
    n2013,
    n2020,
    n2006,
    n2015
  );


  and
  g1995
  (
    n2032,
    n2018,
    n1999,
    n2001,
    n2010
  );


  and
  g1996
  (
    n2029,
    n2016,
    n2011,
    n2023,
    n2021
  );


  xor
  g1997
  (
    n2026,
    n2000,
    n2022,
    n1998,
    n2014
  );


  or
  g1998
  (
    n2031,
    n2005,
    n2012,
    n2025,
    n2017
  );


  nor
  g1999
  (
    n2028,
    n2024,
    n2002,
    n2009,
    n2007
  );


  xor
  KeyGate_0_0
  (
    n1308,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n758,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1185,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1451,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n964,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n962,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1004,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1957,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n362,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1348,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1990,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1417,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n1459,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n1059,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1849,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1813,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n882,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n906,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n885,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1010,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1752,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n971,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1046,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n148,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n1179,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n1081,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n743,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n937,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n689,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n181,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1800,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n1790,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n1766,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n630,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n868,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n1045,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n1375,
    KeyNOTWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n1093,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n75,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n685,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n102,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n1066,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n637,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n830,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n1933,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n666,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n1943,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n658,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n190,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n1216,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n951,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n847,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n783,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n1469,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n283,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n1633,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n1855,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n1449,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n174,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n1580,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n566,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n481,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n59,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n1472,
    KeyNOTWire_0_63
  );


endmodule


