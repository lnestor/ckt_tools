// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_47 written by SynthGen on 2021/04/05 11:08:37
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_47 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n110, n132, n126, n125, n102, n121, n127, n112,
 n115, n129, n119, n109, n107, n108, n128, n131,
 n114, n103, n104, n113, n111, n122, n105, n117,
 n118, n124, n101, n120, n116, n123, n106, n130);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n110, n132, n126, n125, n102, n121, n127, n112,
 n115, n129, n119, n109, n107, n108, n128, n131,
 n114, n103, n104, n113, n111, n122, n105, n117,
 n118, n124, n101, n120, n116, n123, n106, n130;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

not  g0 (n33, n1);
buf  g1 (n37, n1);
buf  g2 (n34, n1);
not  g3 (n36, n2);
not  g4 (n35, n1);
buf  g5 (n45, n34);
buf  g6 (n46, n35);
not  g7 (n40, n34);
buf  g8 (n48, n34);
buf  g9 (n56, n33);
buf  g10 (n42, n35);
buf  g11 (n53, n33);
not  g12 (n44, n37);
buf  g13 (n47, n36);
buf  g14 (n52, n33);
buf  g15 (n38, n34);
buf  g16 (n41, n37);
buf  g17 (n55, n36);
not  g18 (n54, n37);
buf  g19 (n43, n33);
buf  g20 (n50, n36);
buf  g21 (n51, n35);
not  g22 (n49, n35);
buf  g23 (n39, n36);
not  g24 (n79, n28);
buf  g25 (n75, n9);
and  g26 (n65, n47, n18, n8, n29);
nor  g27 (n70, n26, n8, n55, n20);
or   g28 (n91, n48, n11, n56, n6);
xnor g29 (n63, n31, n42, n45, n29);
xor  g30 (n82, n7, n2, n50);
xnor g31 (n78, n22, n25, n13, n26);
xor  g32 (n92, n52, n5, n7, n40);
nand g33 (n67, n52, n10, n7, n21);
nor  g34 (n94, n14, n11, n32, n21);
or   g35 (n60, n12, n17, n28, n21);
nor  g36 (n85, n6, n48, n41, n4);
xor  g37 (n58, n30, n16, n51, n27);
nand g38 (n71, n12, n4, n31, n27);
nor  g39 (n93, n53, n14, n17, n23);
nor  g40 (n66, n11, n15, n4, n25);
or   g41 (n89, n54, n26, n25, n3);
and  g42 (n72, n24, n31, n9, n18);
or   g43 (n97, n27, n22, n6, n24);
or   g44 (n83, n49, n43, n56, n39);
and  g45 (n98, n12, n52, n23, n51);
nand g46 (n61, n19, n50, n9);
and  g47 (n73, n22, n56, n28, n20);
or   g48 (n84, n15, n19, n17, n47);
xnor g49 (n100, n14, n19, n54, n16);
or   g50 (n81, n10, n13, n52, n51);
xnor g51 (n57, n46, n55, n18, n38);
or   g52 (n69, n29, n6, n48, n54);
nand g53 (n62, n16, n15, n12, n14);
and  g54 (n88, n51, n23, n47, n3);
xor  g55 (n74, n19, n30, n56, n47);
or   g56 (n86, n3, n55, n15, n18);
nor  g57 (n76, n2, n13, n5, n10);
and  g58 (n68, n13, n32, n48, n11);
and  g59 (n80, n23, n44, n7, n55);
nor  g60 (n64, n49, n20, n5, n54);
or   g61 (n59, n10, n8, n28, n26);
or   g62 (n87, n17, n20, n2, n5);
and  g63 (n99, n4, n53, n49, n3);
xnor g64 (n77, n31, n24, n27);
xnor g65 (n95, n16, n29, n22, n50);
xor  g66 (n96, n49, n53, n8);
xnor g67 (n90, n21, n30, n25);
nor  g68 (n119, n79, n94, n64, n58);
xor  g69 (n115, n100, n79, n81, n87);
xnor g70 (n123, n85, n98, n92, n91);
nand g71 (n132, n78, n76, n95, n83);
or   g72 (n101, n67, n76, n92, n77);
or   g73 (n105, n92, n95, n79, n68);
nor  g74 (n108, n95, n93, n80, n79);
xor  g75 (n118, n94, n94, n81, n90);
xnor g76 (n128, n61, n77, n87, n82);
and  g77 (n121, n63, n72, n87, n78);
or   g78 (n131, n73, n96, n84, n80);
xnor g79 (n127, n96, n97, n81, n74);
and  g80 (n116, n84, n96, n71, n83);
nor  g81 (n129, n85, n88, n84, n98);
and  g82 (n111, n65, n100, n97, n94);
and  g83 (n124, n88, n59, n76, n99);
or   g84 (n130, n75, n60, n97, n57);
or   g85 (n112, n74, n66, n77, n93);
xor  g86 (n109, n77, n99, n93, n74);
xor  g87 (n102, n89, n86, n90, n82);
nor  g88 (n113, n82, n90, n76, n78);
nor  g89 (n122, n89, n82, n88, n100);
xor  g90 (n120, n83, n88, n86, n91);
nand g91 (n125, n100, n99, n32, n75);
xor  g92 (n103, n93, n92, n74, n98);
xnor g93 (n106, n99, n70, n80);
or   g94 (n114, n90, n87, n91, n69);
xnor g95 (n104, n86, n78, n98, n83);
and  g96 (n126, n95, n62, n85, n89);
xor  g97 (n117, n84, n37, n91, n97);
and  g98 (n110, n86, n85, n75);
and  g99 (n107, n32, n89, n81, n96);
endmodule
