

module Stat_1905_21_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n1530,
  n1551,
  n1559,
  n1562,
  n1548,
  n1549,
  n1556,
  n1560,
  n1547,
  n1552,
  n1543,
  n1564,
  n1545,
  n1919,
  n1921,
  n1911,
  n1915,
  n1918,
  n1916,
  n1925,
  n1914,
  n1926,
  n1924,
  n1913,
  n1920,
  n1917,
  n1923,
  n1922,
  n1912,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n1530;
  output n1551;
  output n1559;
  output n1562;
  output n1548;
  output n1549;
  output n1556;
  output n1560;
  output n1547;
  output n1552;
  output n1543;
  output n1564;
  output n1545;
  output n1919;
  output n1921;
  output n1911;
  output n1915;
  output n1918;
  output n1916;
  output n1925;
  output n1914;
  output n1926;
  output n1924;
  output n1913;
  output n1920;
  output n1917;
  output n1923;
  output n1922;
  output n1912;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1544;
  wire n1546;
  wire n1550;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1557;
  wire n1558;
  wire n1561;
  wire n1563;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    n93,
    n9
  );


  buf
  g1
  (
    n99,
    n11
  );


  not
  g2
  (
    n59,
    n8
  );


  not
  g3
  (
    n84,
    n10
  );


  not
  g4
  (
    n53,
    n7
  );


  not
  g5
  (
    n102,
    n10
  );


  buf
  g6
  (
    n40,
    n11
  );


  not
  g7
  (
    n75,
    n5
  );


  buf
  g8
  (
    n46,
    n6
  );


  not
  g9
  (
    n88,
    n13
  );


  not
  g10
  (
    n54,
    n17
  );


  not
  g11
  (
    n72,
    n15
  );


  not
  g12
  (
    n87,
    n17
  );


  buf
  g13
  (
    n91,
    n15
  );


  buf
  g14
  (
    n43,
    n4
  );


  not
  g15
  (
    n81,
    n5
  );


  buf
  g16
  (
    n67,
    n4
  );


  not
  g17
  (
    n63,
    n14
  );


  not
  g18
  (
    n52,
    n14
  );


  buf
  g19
  (
    n80,
    n4
  );


  not
  g20
  (
    n73,
    n16
  );


  buf
  g21
  (
    n69,
    n15
  );


  not
  g22
  (
    n83,
    n21
  );


  buf
  g23
  (
    n23,
    n4
  );


  buf
  g24
  (
    n105,
    n3
  );


  not
  g25
  (
    n97,
    n21
  );


  not
  g26
  (
    n35,
    n5
  );


  not
  g27
  (
    n68,
    n10
  );


  buf
  g28
  (
    n28,
    n16
  );


  buf
  g29
  (
    n30,
    n2
  );


  not
  g30
  (
    n70,
    n18
  );


  buf
  g31
  (
    n45,
    n20
  );


  not
  g32
  (
    n62,
    n12
  );


  not
  g33
  (
    n29,
    n10
  );


  not
  g34
  (
    n96,
    n1
  );


  buf
  g35
  (
    n86,
    n19
  );


  buf
  g36
  (
    n89,
    n3
  );


  not
  g37
  (
    KeyWire_0_6,
    n9
  );


  not
  g38
  (
    n26,
    n7
  );


  not
  g39
  (
    n32,
    n19
  );


  buf
  g40
  (
    n65,
    n3
  );


  not
  g41
  (
    n24,
    n13
  );


  buf
  g42
  (
    n33,
    n1
  );


  not
  g43
  (
    n44,
    n14
  );


  buf
  g44
  (
    n79,
    n7
  );


  not
  g45
  (
    n103,
    n13
  );


  not
  g46
  (
    n34,
    n9
  );


  buf
  g47
  (
    n49,
    n9
  );


  buf
  g48
  (
    n36,
    n14
  );


  buf
  g49
  (
    n48,
    n19
  );


  not
  g50
  (
    n78,
    n1
  );


  not
  g51
  (
    n57,
    n6
  );


  buf
  g52
  (
    n98,
    n6
  );


  not
  g53
  (
    n90,
    n20
  );


  buf
  g54
  (
    n64,
    n20
  );


  buf
  g55
  (
    n77,
    n18
  );


  not
  g56
  (
    n76,
    n8
  );


  buf
  g57
  (
    KeyWire_0_0,
    n7
  );


  not
  g58
  (
    n60,
    n21
  );


  not
  g59
  (
    n100,
    n11
  );


  not
  g60
  (
    n22,
    n2
  );


  buf
  g61
  (
    n71,
    n2
  );


  not
  g62
  (
    n37,
    n19
  );


  buf
  g63
  (
    n94,
    n1
  );


  not
  g64
  (
    n58,
    n17
  );


  buf
  g65
  (
    KeyWire_0_4,
    n6
  );


  buf
  g66
  (
    n74,
    n12
  );


  not
  g67
  (
    n56,
    n8
  );


  buf
  g68
  (
    n55,
    n16
  );


  not
  g69
  (
    n39,
    n3
  );


  buf
  g70
  (
    n66,
    n18
  );


  not
  g71
  (
    n38,
    n16
  );


  buf
  g72
  (
    n51,
    n21
  );


  not
  g73
  (
    n50,
    n15
  );


  not
  g74
  (
    n85,
    n12
  );


  not
  g75
  (
    n42,
    n11
  );


  not
  g76
  (
    n95,
    n13
  );


  buf
  g77
  (
    n41,
    n2
  );


  buf
  g78
  (
    n61,
    n5
  );


  not
  g79
  (
    n104,
    n12
  );


  buf
  g80
  (
    n47,
    n18
  );


  not
  g81
  (
    n25,
    n20
  );


  buf
  g82
  (
    n101,
    n8
  );


  not
  g83
  (
    n82,
    n17
  );


  not
  g84
  (
    n329,
    n46
  );


  not
  g85
  (
    n362,
    n69
  );


  buf
  g86
  (
    n293,
    n54
  );


  not
  g87
  (
    n201,
    n77
  );


  buf
  g88
  (
    n397,
    n62
  );


  buf
  g89
  (
    n413,
    n91
  );


  not
  g90
  (
    n230,
    n74
  );


  buf
  g91
  (
    n303,
    n46
  );


  not
  g92
  (
    n106,
    n95
  );


  buf
  g93
  (
    n437,
    n26
  );


  not
  g94
  (
    n147,
    n87
  );


  not
  g95
  (
    n138,
    n35
  );


  buf
  g96
  (
    n321,
    n54
  );


  not
  g97
  (
    n337,
    n68
  );


  buf
  g98
  (
    n237,
    n26
  );


  buf
  g99
  (
    n262,
    n38
  );


  not
  g100
  (
    n364,
    n63
  );


  not
  g101
  (
    n108,
    n60
  );


  not
  g102
  (
    n388,
    n65
  );


  not
  g103
  (
    n291,
    n85
  );


  buf
  g104
  (
    n405,
    n59
  );


  not
  g105
  (
    n122,
    n105
  );


  not
  g106
  (
    n307,
    n80
  );


  not
  g107
  (
    n112,
    n66
  );


  not
  g108
  (
    n164,
    n40
  );


  not
  g109
  (
    n171,
    n90
  );


  not
  g110
  (
    n238,
    n30
  );


  not
  g111
  (
    n415,
    n37
  );


  buf
  g112
  (
    n257,
    n80
  );


  not
  g113
  (
    n156,
    n87
  );


  not
  g114
  (
    n380,
    n25
  );


  buf
  g115
  (
    n139,
    n60
  );


  buf
  g116
  (
    n382,
    n42
  );


  not
  g117
  (
    n183,
    n54
  );


  not
  g118
  (
    n114,
    n26
  );


  buf
  g119
  (
    n166,
    n103
  );


  buf
  g120
  (
    n280,
    n81
  );


  not
  g121
  (
    n423,
    n60
  );


  not
  g122
  (
    n181,
    n48
  );


  not
  g123
  (
    n130,
    n96
  );


  buf
  g124
  (
    n246,
    n38
  );


  not
  g125
  (
    n353,
    n50
  );


  buf
  g126
  (
    n211,
    n30
  );


  not
  g127
  (
    n304,
    n62
  );


  buf
  g128
  (
    n207,
    n85
  );


  not
  g129
  (
    n232,
    n43
  );


  not
  g130
  (
    n187,
    n41
  );


  buf
  g131
  (
    n319,
    n100
  );


  not
  g132
  (
    n158,
    n98
  );


  not
  g133
  (
    n289,
    n55
  );


  buf
  g134
  (
    n137,
    n103
  );


  not
  g135
  (
    n368,
    n53
  );


  buf
  g136
  (
    n123,
    n55
  );


  buf
  g137
  (
    KeyWire_0_2,
    n55
  );


  buf
  g138
  (
    n345,
    n62
  );


  not
  g139
  (
    n435,
    n85
  );


  buf
  g140
  (
    n386,
    n70
  );


  not
  g141
  (
    n340,
    n83
  );


  not
  g142
  (
    n326,
    n96
  );


  buf
  g143
  (
    n261,
    n57
  );


  buf
  g144
  (
    n430,
    n104
  );


  not
  g145
  (
    n401,
    n30
  );


  buf
  g146
  (
    n378,
    n59
  );


  not
  g147
  (
    n408,
    n62
  );


  buf
  g148
  (
    n195,
    n90
  );


  buf
  g149
  (
    n283,
    n91
  );


  buf
  g150
  (
    n119,
    n81
  );


  buf
  g151
  (
    n323,
    n25
  );


  not
  g152
  (
    n421,
    n22
  );


  not
  g153
  (
    n190,
    n35
  );


  not
  g154
  (
    n285,
    n56
  );


  buf
  g155
  (
    n431,
    n28
  );


  buf
  g156
  (
    n165,
    n71
  );


  buf
  g157
  (
    n126,
    n42
  );


  not
  g158
  (
    n243,
    n49
  );


  buf
  g159
  (
    n167,
    n81
  );


  buf
  g160
  (
    n360,
    n33
  );


  not
  g161
  (
    n361,
    n97
  );


  buf
  g162
  (
    n152,
    n37
  );


  not
  g163
  (
    n159,
    n43
  );


  not
  g164
  (
    n197,
    n68
  );


  not
  g165
  (
    n301,
    n58
  );


  buf
  g166
  (
    n172,
    n46
  );


  buf
  g167
  (
    n127,
    n49
  );


  buf
  g168
  (
    n244,
    n95
  );


  not
  g169
  (
    n409,
    n89
  );


  not
  g170
  (
    n271,
    n73
  );


  not
  g171
  (
    n286,
    n47
  );


  buf
  g172
  (
    n330,
    n91
  );


  buf
  g173
  (
    n233,
    n70
  );


  not
  g174
  (
    n315,
    n87
  );


  buf
  g175
  (
    n325,
    n35
  );


  buf
  g176
  (
    n418,
    n26
  );


  buf
  g177
  (
    n436,
    n84
  );


  not
  g178
  (
    n297,
    n63
  );


  buf
  g179
  (
    n118,
    n36
  );


  not
  g180
  (
    KeyWire_0_29,
    n28
  );


  not
  g181
  (
    n375,
    n95
  );


  buf
  g182
  (
    n347,
    n82
  );


  buf
  g183
  (
    n221,
    n99
  );


  not
  g184
  (
    n427,
    n42
  );


  not
  g185
  (
    n426,
    n52
  );


  buf
  g186
  (
    n205,
    n49
  );


  not
  g187
  (
    n210,
    n101
  );


  buf
  g188
  (
    n163,
    n53
  );


  not
  g189
  (
    n214,
    n27
  );


  buf
  g190
  (
    n270,
    n100
  );


  not
  g191
  (
    n202,
    n22
  );


  buf
  g192
  (
    n140,
    n24
  );


  not
  g193
  (
    n384,
    n41
  );


  buf
  g194
  (
    n281,
    n78
  );


  buf
  g195
  (
    n393,
    n104
  );


  buf
  g196
  (
    n157,
    n79
  );


  buf
  g197
  (
    n107,
    n70
  );


  not
  g198
  (
    n222,
    n76
  );


  not
  g199
  (
    n363,
    n74
  );


  not
  g200
  (
    n178,
    n103
  );


  buf
  g201
  (
    n357,
    n41
  );


  not
  g202
  (
    n400,
    n78
  );


  not
  g203
  (
    n115,
    n24
  );


  buf
  g204
  (
    n160,
    n80
  );


  not
  g205
  (
    n407,
    n73
  );


  buf
  g206
  (
    n179,
    n98
  );


  not
  g207
  (
    n255,
    n38
  );


  not
  g208
  (
    n193,
    n84
  );


  buf
  g209
  (
    n367,
    n30
  );


  buf
  g210
  (
    n116,
    n77
  );


  buf
  g211
  (
    n219,
    n101
  );


  not
  g212
  (
    n296,
    n39
  );


  buf
  g213
  (
    n204,
    n94
  );


  buf
  g214
  (
    n206,
    n27
  );


  not
  g215
  (
    n429,
    n58
  );


  buf
  g216
  (
    n161,
    n32
  );


  not
  g217
  (
    n273,
    n34
  );


  buf
  g218
  (
    n334,
    n47
  );


  not
  g219
  (
    n333,
    n23
  );


  not
  g220
  (
    n250,
    n65
  );


  buf
  g221
  (
    n133,
    n28
  );


  not
  g222
  (
    n410,
    n67
  );


  not
  g223
  (
    n151,
    n44
  );


  not
  g224
  (
    n175,
    n65
  );


  buf
  g225
  (
    n194,
    n92
  );


  buf
  g226
  (
    n241,
    n45
  );


  not
  g227
  (
    n290,
    n45
  );


  buf
  g228
  (
    n298,
    n101
  );


  buf
  g229
  (
    n125,
    n105
  );


  not
  g230
  (
    n381,
    n86
  );


  not
  g231
  (
    n268,
    n79
  );


  buf
  g232
  (
    n314,
    n76
  );


  buf
  g233
  (
    n128,
    n93
  );


  not
  g234
  (
    n121,
    n53
  );


  not
  g235
  (
    n234,
    n71
  );


  not
  g236
  (
    n328,
    n102
  );


  not
  g237
  (
    n282,
    n88
  );


  not
  g238
  (
    n336,
    n86
  );


  not
  g239
  (
    n327,
    n22
  );


  buf
  g240
  (
    n343,
    n64
  );


  not
  g241
  (
    n110,
    n89
  );


  buf
  g242
  (
    n352,
    n81
  );


  buf
  g243
  (
    n226,
    n82
  );


  not
  g244
  (
    n189,
    n75
  );


  buf
  g245
  (
    n335,
    n25
  );


  not
  g246
  (
    n253,
    n47
  );


  not
  g247
  (
    n144,
    n66
  );


  not
  g248
  (
    n168,
    n84
  );


  buf
  g249
  (
    n320,
    n75
  );


  not
  g250
  (
    n331,
    n64
  );


  buf
  g251
  (
    n287,
    n50
  );


  not
  g252
  (
    n176,
    n61
  );


  not
  g253
  (
    n182,
    n34
  );


  buf
  g254
  (
    n389,
    n56
  );


  buf
  g255
  (
    n228,
    n50
  );


  not
  g256
  (
    n371,
    n72
  );


  not
  g257
  (
    n213,
    n29
  );


  not
  g258
  (
    n428,
    n93
  );


  buf
  g259
  (
    n425,
    n29
  );


  buf
  g260
  (
    n383,
    n35
  );


  buf
  g261
  (
    n373,
    n71
  );


  buf
  g262
  (
    n424,
    n101
  );


  buf
  g263
  (
    n146,
    n94
  );


  not
  g264
  (
    n249,
    n61
  );


  buf
  g265
  (
    n220,
    n25
  );


  not
  g266
  (
    n145,
    n57
  );


  buf
  g267
  (
    n369,
    n32
  );


  not
  g268
  (
    n153,
    n31
  );


  not
  g269
  (
    n258,
    n74
  );


  buf
  g270
  (
    n306,
    n38
  );


  not
  g271
  (
    n177,
    n102
  );


  not
  g272
  (
    n131,
    n56
  );


  buf
  g273
  (
    n142,
    n92
  );


  buf
  g274
  (
    n208,
    n56
  );


  buf
  g275
  (
    n366,
    n34
  );


  buf
  g276
  (
    n251,
    n39
  );


  not
  g277
  (
    n284,
    n58
  );


  buf
  g278
  (
    n196,
    n67
  );


  not
  g279
  (
    n239,
    n37
  );


  not
  g280
  (
    n376,
    n90
  );


  buf
  g281
  (
    n439,
    n48
  );


  buf
  g282
  (
    n235,
    n79
  );


  not
  g283
  (
    n344,
    n45
  );


  not
  g284
  (
    n200,
    n44
  );


  buf
  g285
  (
    n186,
    n67
  );


  buf
  g286
  (
    n385,
    n44
  );


  buf
  g287
  (
    n318,
    n77
  );


  not
  g288
  (
    KeyWire_0_21,
    n59
  );


  buf
  g289
  (
    n229,
    n94
  );


  not
  g290
  (
    n227,
    n52
  );


  not
  g291
  (
    n170,
    n51
  );


  buf
  g292
  (
    n419,
    n83
  );


  buf
  g293
  (
    n154,
    n48
  );


  not
  g294
  (
    n402,
    n48
  );


  not
  g295
  (
    n120,
    n33
  );


  not
  g296
  (
    n254,
    n103
  );


  not
  g297
  (
    n379,
    n73
  );


  not
  g298
  (
    n300,
    n72
  );


  buf
  g299
  (
    n416,
    n31
  );


  not
  g300
  (
    n274,
    n70
  );


  not
  g301
  (
    n414,
    n39
  );


  buf
  g302
  (
    n387,
    n33
  );


  not
  g303
  (
    n422,
    n45
  );


  buf
  g304
  (
    KeyWire_0_14,
    n88
  );


  buf
  g305
  (
    n174,
    n82
  );


  buf
  g306
  (
    n180,
    n36
  );


  not
  g307
  (
    n148,
    n104
  );


  buf
  g308
  (
    n256,
    n60
  );


  buf
  g309
  (
    n399,
    n79
  );


  buf
  g310
  (
    n267,
    n24
  );


  not
  g311
  (
    n316,
    n40
  );


  buf
  g312
  (
    n348,
    n61
  );


  not
  g313
  (
    n404,
    n95
  );


  buf
  g314
  (
    n312,
    n86
  );


  not
  g315
  (
    n370,
    n29
  );


  buf
  g316
  (
    n278,
    n68
  );


  buf
  g317
  (
    n433,
    n78
  );


  buf
  g318
  (
    n292,
    n29
  );


  not
  g319
  (
    n149,
    n97
  );


  not
  g320
  (
    n231,
    n75
  );


  not
  g321
  (
    n136,
    n31
  );


  not
  g322
  (
    n275,
    n102
  );


  buf
  g323
  (
    n338,
    n76
  );


  buf
  g324
  (
    n403,
    n105
  );


  not
  g325
  (
    n398,
    n24
  );


  buf
  g326
  (
    n217,
    n28
  );


  buf
  g327
  (
    n218,
    n57
  );


  buf
  g328
  (
    n311,
    n80
  );


  not
  g329
  (
    n132,
    n86
  );


  buf
  g330
  (
    n134,
    n32
  );


  not
  g331
  (
    n247,
    n99
  );


  buf
  g332
  (
    n143,
    n32
  );


  buf
  g333
  (
    n272,
    n39
  );


  buf
  g334
  (
    n391,
    n73
  );


  buf
  g335
  (
    n309,
    n58
  );


  not
  g336
  (
    n264,
    n64
  );


  buf
  g337
  (
    n223,
    n69
  );


  not
  g338
  (
    n350,
    n67
  );


  not
  g339
  (
    n109,
    n99
  );


  buf
  g340
  (
    n295,
    n100
  );


  buf
  g341
  (
    n169,
    n36
  );


  not
  g342
  (
    n215,
    n66
  );


  not
  g343
  (
    n276,
    n43
  );


  buf
  g344
  (
    n240,
    n34
  );


  buf
  g345
  (
    n259,
    n51
  );


  buf
  g346
  (
    n317,
    n44
  );


  not
  g347
  (
    n339,
    n57
  );


  not
  g348
  (
    n341,
    n65
  );


  buf
  g349
  (
    n199,
    n68
  );


  buf
  g350
  (
    n417,
    n54
  );


  buf
  g351
  (
    n302,
    n96
  );


  buf
  g352
  (
    n162,
    n102
  );


  not
  g353
  (
    KeyWire_0_3,
    n43
  );


  not
  g354
  (
    n117,
    n92
  );


  not
  g355
  (
    n198,
    n36
  );


  not
  g356
  (
    n394,
    n72
  );


  buf
  g357
  (
    n356,
    n92
  );


  not
  g358
  (
    n150,
    n59
  );


  buf
  g359
  (
    n358,
    n97
  );


  buf
  g360
  (
    n440,
    n87
  );


  not
  g361
  (
    n288,
    n83
  );


  not
  g362
  (
    n432,
    n69
  );


  not
  g363
  (
    n396,
    n52
  );


  not
  g364
  (
    n355,
    n41
  );


  buf
  g365
  (
    n266,
    n49
  );


  not
  g366
  (
    n185,
    n33
  );


  buf
  g367
  (
    n392,
    n51
  );


  buf
  g368
  (
    n342,
    n82
  );


  buf
  g369
  (
    n310,
    n69
  );


  not
  g370
  (
    n372,
    n27
  );


  not
  g371
  (
    n260,
    n31
  );


  buf
  g372
  (
    n351,
    n71
  );


  buf
  g373
  (
    n191,
    n63
  );


  buf
  g374
  (
    n269,
    n63
  );


  buf
  g375
  (
    n365,
    n89
  );


  buf
  g376
  (
    n277,
    n91
  );


  not
  g377
  (
    n390,
    n98
  );


  not
  g378
  (
    n113,
    n77
  );


  not
  g379
  (
    n225,
    n27
  );


  buf
  g380
  (
    n209,
    n83
  );


  buf
  g381
  (
    n245,
    n61
  );


  not
  g382
  (
    n294,
    n84
  );


  buf
  g383
  (
    n252,
    n74
  );


  buf
  g384
  (
    n305,
    n23
  );


  not
  g385
  (
    n406,
    n42
  );


  not
  g386
  (
    n322,
    n98
  );


  not
  g387
  (
    n299,
    n88
  );


  buf
  g388
  (
    n184,
    n97
  );


  not
  g389
  (
    n308,
    n88
  );


  buf
  g390
  (
    n155,
    n85
  );


  not
  g391
  (
    n236,
    n40
  );


  buf
  g392
  (
    n346,
    n55
  );


  buf
  g393
  (
    n374,
    n47
  );


  not
  g394
  (
    n349,
    n93
  );


  not
  g395
  (
    n377,
    n94
  );


  not
  g396
  (
    n438,
    n100
  );


  not
  g397
  (
    n412,
    n72
  );


  not
  g398
  (
    n141,
    n104
  );


  not
  g399
  (
    n224,
    n23
  );


  not
  g400
  (
    n248,
    n40
  );


  buf
  g401
  (
    n324,
    n93
  );


  buf
  g402
  (
    n332,
    n37
  );


  buf
  g403
  (
    n313,
    n51
  );


  not
  g404
  (
    n188,
    n46
  );


  not
  g405
  (
    n359,
    n52
  );


  buf
  g406
  (
    n265,
    n89
  );


  buf
  g407
  (
    n111,
    n22
  );


  not
  g408
  (
    n124,
    n99
  );


  not
  g409
  (
    n434,
    n78
  );


  buf
  g410
  (
    n203,
    n90
  );


  buf
  g411
  (
    n135,
    n75
  );


  buf
  g412
  (
    n395,
    n50
  );


  buf
  g413
  (
    n354,
    n96
  );


  not
  g414
  (
    n411,
    n23
  );


  buf
  g415
  (
    n212,
    n64
  );


  not
  g416
  (
    n192,
    n66
  );


  buf
  g417
  (
    n129,
    n53
  );


  buf
  g418
  (
    n242,
    n76
  );


  not
  g419
  (
    n676,
    n317
  );


  buf
  g420
  (
    n699,
    n187
  );


  buf
  g421
  (
    n824,
    n112
  );


  buf
  g422
  (
    n941,
    n354
  );


  not
  g423
  (
    n961,
    n324
  );


  not
  g424
  (
    n570,
    n212
  );


  buf
  g425
  (
    n753,
    n243
  );


  not
  g426
  (
    n1116,
    n362
  );


  not
  g427
  (
    n611,
    n220
  );


  buf
  g428
  (
    n475,
    n210
  );


  buf
  g429
  (
    n1074,
    n340
  );


  not
  g430
  (
    n510,
    n309
  );


  not
  g431
  (
    n913,
    n192
  );


  not
  g432
  (
    n1021,
    n314
  );


  buf
  g433
  (
    n872,
    n198
  );


  buf
  g434
  (
    n701,
    n210
  );


  not
  g435
  (
    n444,
    n222
  );


  not
  g436
  (
    n932,
    n134
  );


  not
  g437
  (
    n1119,
    n257
  );


  not
  g438
  (
    n1041,
    n174
  );


  buf
  g439
  (
    n1069,
    n270
  );


  buf
  g440
  (
    n471,
    n158
  );


  not
  g441
  (
    n1170,
    n269
  );


  not
  g442
  (
    n454,
    n161
  );


  not
  g443
  (
    n876,
    n246
  );


  buf
  g444
  (
    n456,
    n198
  );


  not
  g445
  (
    n746,
    n233
  );


  not
  g446
  (
    n739,
    n154
  );


  not
  g447
  (
    n1096,
    n147
  );


  not
  g448
  (
    n639,
    n344
  );


  not
  g449
  (
    n590,
    n182
  );


  not
  g450
  (
    n787,
    n336
  );


  not
  g451
  (
    n582,
    n232
  );


  not
  g452
  (
    n925,
    n256
  );


  not
  g453
  (
    n804,
    n128
  );


  buf
  g454
  (
    n664,
    n312
  );


  not
  g455
  (
    n720,
    n304
  );


  buf
  g456
  (
    n886,
    n350
  );


  not
  g457
  (
    n596,
    n335
  );


  buf
  g458
  (
    n1164,
    n125
  );


  not
  g459
  (
    n813,
    n328
  );


  buf
  g460
  (
    n920,
    n157
  );


  not
  g461
  (
    n1017,
    n294
  );


  buf
  g462
  (
    n856,
    n291
  );


  buf
  g463
  (
    n934,
    n262
  );


  not
  g464
  (
    n995,
    n264
  );


  not
  g465
  (
    n738,
    n226
  );


  not
  g466
  (
    n839,
    n134
  );


  not
  g467
  (
    n484,
    n229
  );


  buf
  g468
  (
    n852,
    n149
  );


  buf
  g469
  (
    n773,
    n190
  );


  buf
  g470
  (
    n761,
    n355
  );


  buf
  g471
  (
    n1043,
    n174
  );


  buf
  g472
  (
    n662,
    n363
  );


  not
  g473
  (
    n1048,
    n128
  );


  buf
  g474
  (
    n1095,
    n374
  );


  not
  g475
  (
    n819,
    n363
  );


  not
  g476
  (
    n693,
    n317
  );


  buf
  g477
  (
    n731,
    n195
  );


  buf
  g478
  (
    n1015,
    n285
  );


  not
  g479
  (
    n732,
    n366
  );


  not
  g480
  (
    n548,
    n107
  );


  buf
  g481
  (
    n851,
    n248
  );


  buf
  g482
  (
    n816,
    n196
  );


  not
  g483
  (
    n626,
    n143
  );


  buf
  g484
  (
    n985,
    n217
  );


  not
  g485
  (
    n1137,
    n252
  );


  buf
  g486
  (
    n975,
    n314
  );


  not
  g487
  (
    n750,
    n161
  );


  not
  g488
  (
    n757,
    n351
  );


  buf
  g489
  (
    n531,
    n383
  );


  not
  g490
  (
    n478,
    n336
  );


  not
  g491
  (
    n631,
    n138
  );


  buf
  g492
  (
    n997,
    n325
  );


  not
  g493
  (
    n690,
    n126
  );


  not
  g494
  (
    n508,
    n107
  );


  buf
  g495
  (
    n1161,
    n109
  );


  not
  g496
  (
    n809,
    n316
  );


  buf
  g497
  (
    n1030,
    n236
  );


  not
  g498
  (
    n1169,
    n357
  );


  buf
  g499
  (
    n465,
    n373
  );


  buf
  g500
  (
    n542,
    n357
  );


  buf
  g501
  (
    n891,
    n115
  );


  buf
  g502
  (
    n496,
    n352
  );


  not
  g503
  (
    n1040,
    n363
  );


  not
  g504
  (
    n501,
    n386
  );


  not
  g505
  (
    n1025,
    n163
  );


  not
  g506
  (
    n989,
    n153
  );


  buf
  g507
  (
    n747,
    n201
  );


  not
  g508
  (
    n726,
    n124
  );


  buf
  g509
  (
    KeyWire_0_23,
    n310
  );


  not
  g510
  (
    n1072,
    n242
  );


  buf
  g511
  (
    n649,
    n342
  );


  buf
  g512
  (
    n794,
    n192
  );


  not
  g513
  (
    n874,
    n353
  );


  not
  g514
  (
    n767,
    n328
  );


  not
  g515
  (
    n777,
    n359
  );


  buf
  g516
  (
    n957,
    n258
  );


  buf
  g517
  (
    n620,
    n174
  );


  not
  g518
  (
    n530,
    n251
  );


  buf
  g519
  (
    n778,
    n136
  );


  buf
  g520
  (
    n566,
    n123
  );


  buf
  g521
  (
    n1122,
    n261
  );


  not
  g522
  (
    n855,
    n144
  );


  buf
  g523
  (
    n1088,
    n206
  );


  buf
  g524
  (
    n771,
    n356
  );


  buf
  g525
  (
    n513,
    n197
  );


  buf
  g526
  (
    n1118,
    n150
  );


  not
  g527
  (
    n1127,
    n301
  );


  not
  g528
  (
    n618,
    n257
  );


  not
  g529
  (
    n953,
    n304
  );


  buf
  g530
  (
    n905,
    n111
  );


  not
  g531
  (
    n1054,
    n327
  );


  buf
  g532
  (
    n752,
    n342
  );


  buf
  g533
  (
    n1110,
    n380
  );


  not
  g534
  (
    n546,
    n299
  );


  not
  g535
  (
    n1151,
    n267
  );


  not
  g536
  (
    n987,
    n262
  );


  buf
  g537
  (
    n741,
    n323
  );


  not
  g538
  (
    n758,
    n377
  );


  not
  g539
  (
    n955,
    n320
  );


  not
  g540
  (
    n719,
    n110
  );


  not
  g541
  (
    n922,
    n246
  );


  buf
  g542
  (
    n1132,
    n193
  );


  buf
  g543
  (
    n674,
    n234
  );


  buf
  g544
  (
    n1128,
    n285
  );


  not
  g545
  (
    n635,
    n182
  );


  buf
  g546
  (
    n994,
    n246
  );


  buf
  g547
  (
    n877,
    n207
  );


  not
  g548
  (
    n799,
    n340
  );


  not
  g549
  (
    n715,
    n371
  );


  not
  g550
  (
    n939,
    n253
  );


  buf
  g551
  (
    n580,
    n219
  );


  buf
  g552
  (
    n469,
    n241
  );


  not
  g553
  (
    n560,
    n231
  );


  buf
  g554
  (
    n462,
    n123
  );


  buf
  g555
  (
    n1022,
    n229
  );


  buf
  g556
  (
    n768,
    n237
  );


  buf
  g557
  (
    n770,
    n261
  );


  buf
  g558
  (
    n935,
    n231
  );


  not
  g559
  (
    n883,
    n167
  );


  not
  g560
  (
    n453,
    n152
  );


  buf
  g561
  (
    n900,
    n226
  );


  buf
  g562
  (
    n571,
    n276
  );


  buf
  g563
  (
    n788,
    n292
  );


  not
  g564
  (
    n1065,
    n215
  );


  buf
  g565
  (
    n822,
    n303
  );


  not
  g566
  (
    n871,
    n251
  );


  not
  g567
  (
    n1131,
    n346
  );


  buf
  g568
  (
    n873,
    n167
  );


  buf
  g569
  (
    n928,
    n249
  );


  not
  g570
  (
    n583,
    n288
  );


  not
  g571
  (
    n775,
    n154
  );


  not
  g572
  (
    n599,
    n312
  );


  not
  g573
  (
    n1007,
    n229
  );


  not
  g574
  (
    n898,
    n346
  );


  buf
  g575
  (
    n536,
    n372
  );


  not
  g576
  (
    n556,
    n129
  );


  buf
  g577
  (
    n575,
    n375
  );


  buf
  g578
  (
    n1155,
    n161
  );


  buf
  g579
  (
    n659,
    n238
  );


  buf
  g580
  (
    n979,
    n369
  );


  buf
  g581
  (
    n742,
    n311
  );


  buf
  g582
  (
    n616,
    n216
  );


  not
  g583
  (
    n554,
    n376
  );


  buf
  g584
  (
    n517,
    n288
  );


  not
  g585
  (
    n466,
    n313
  );


  not
  g586
  (
    n1093,
    n261
  );


  buf
  g587
  (
    n756,
    n184
  );


  not
  g588
  (
    n1044,
    n346
  );


  not
  g589
  (
    n704,
    n149
  );


  not
  g590
  (
    n1001,
    n284
  );


  not
  g591
  (
    n880,
    n272
  );


  buf
  g592
  (
    n780,
    n271
  );


  not
  g593
  (
    n769,
    n371
  );


  not
  g594
  (
    n1109,
    n341
  );


  buf
  g595
  (
    n1016,
    n107
  );


  buf
  g596
  (
    n667,
    n113
  );


  not
  g597
  (
    n1111,
    n211
  );


  buf
  g598
  (
    n765,
    n326
  );


  buf
  g599
  (
    n544,
    n371
  );


  not
  g600
  (
    n827,
    n292
  );


  buf
  g601
  (
    n656,
    n296
  );


  not
  g602
  (
    n723,
    n131
  );


  buf
  g603
  (
    n579,
    n213
  );


  not
  g604
  (
    n1010,
    n190
  );


  buf
  g605
  (
    n993,
    n119
  );


  not
  g606
  (
    n1121,
    n166
  );


  buf
  g607
  (
    n672,
    n123
  );


  buf
  g608
  (
    n606,
    n161
  );


  not
  g609
  (
    n792,
    n269
  );


  buf
  g610
  (
    n832,
    n292
  );


  not
  g611
  (
    n550,
    n157
  );


  buf
  g612
  (
    n485,
    n115
  );


  not
  g613
  (
    n705,
    n368
  );


  not
  g614
  (
    n464,
    n359
  );


  not
  g615
  (
    n535,
    n254
  );


  not
  g616
  (
    n1050,
    n283
  );


  buf
  g617
  (
    n1087,
    n373
  );


  not
  g618
  (
    n791,
    n191
  );


  not
  g619
  (
    n1157,
    n310
  );


  not
  g620
  (
    n947,
    n334
  );


  buf
  g621
  (
    n807,
    n352
  );


  not
  g622
  (
    n966,
    n288
  );


  buf
  g623
  (
    n729,
    n262
  );


  buf
  g624
  (
    n492,
    n350
  );


  not
  g625
  (
    n673,
    n318
  );


  buf
  g626
  (
    n1032,
    n248
  );


  not
  g627
  (
    n645,
    n289
  );


  buf
  g628
  (
    n1113,
    n351
  );


  not
  g629
  (
    n609,
    n112
  );


  not
  g630
  (
    n936,
    n131
  );


  buf
  g631
  (
    n521,
    n311
  );


  not
  g632
  (
    n481,
    n130
  );


  not
  g633
  (
    n823,
    n204
  );


  not
  g634
  (
    n1100,
    n178
  );


  buf
  g635
  (
    n915,
    n244
  );


  buf
  g636
  (
    n1173,
    n210
  );


  buf
  g637
  (
    n868,
    n162
  );


  not
  g638
  (
    n1163,
    n148
  );


  not
  g639
  (
    n793,
    n115
  );


  buf
  g640
  (
    n1150,
    n295
  );


  buf
  g641
  (
    n474,
    n245
  );


  not
  g642
  (
    n952,
    n143
  );


  buf
  g643
  (
    n1052,
    n223
  );


  not
  g644
  (
    n1012,
    n145
  );


  not
  g645
  (
    n808,
    n143
  );


  buf
  g646
  (
    n786,
    n364
  );


  buf
  g647
  (
    n721,
    n383
  );


  buf
  g648
  (
    n789,
    n206
  );


  not
  g649
  (
    n614,
    n249
  );


  not
  g650
  (
    n971,
    n302
  );


  not
  g651
  (
    n986,
    n243
  );


  buf
  g652
  (
    n930,
    n235
  );


  buf
  g653
  (
    n815,
    n319
  );


  buf
  g654
  (
    n684,
    n279
  );


  not
  g655
  (
    n516,
    n305
  );


  buf
  g656
  (
    n885,
    n207
  );


  buf
  g657
  (
    n826,
    n249
  );


  buf
  g658
  (
    n725,
    n275
  );


  buf
  g659
  (
    n929,
    n341
  );


  not
  g660
  (
    n447,
    n289
  );


  not
  g661
  (
    n901,
    n376
  );


  not
  g662
  (
    n895,
    n230
  );


  buf
  g663
  (
    n472,
    n133
  );


  buf
  g664
  (
    n702,
    n107
  );


  not
  g665
  (
    n569,
    n329
  );


  buf
  g666
  (
    n653,
    n214
  );


  buf
  g667
  (
    n722,
    n200
  );


  buf
  g668
  (
    n1075,
    n268
  );


  buf
  g669
  (
    n1056,
    n127
  );


  not
  g670
  (
    n759,
    n178
  );


  not
  g671
  (
    n563,
    n360
  );


  not
  g672
  (
    n489,
    n211
  );


  not
  g673
  (
    n592,
    n152
  );


  buf
  g674
  (
    n845,
    n300
  );


  not
  g675
  (
    n992,
    n329
  );


  not
  g676
  (
    n1160,
    n290
  );


  not
  g677
  (
    n1174,
    n320
  );


  not
  g678
  (
    n538,
    n152
  );


  buf
  g679
  (
    n710,
    n385
  );


  not
  g680
  (
    n628,
    n356
  );


  not
  g681
  (
    n743,
    n188
  );


  not
  g682
  (
    n1147,
    n139
  );


  not
  g683
  (
    n545,
    n227
  );


  buf
  g684
  (
    n479,
    n116
  );


  not
  g685
  (
    n1049,
    n359
  );


  not
  g686
  (
    n760,
    n377
  );


  not
  g687
  (
    n679,
    n315
  );


  buf
  g688
  (
    n1108,
    n186
  );


  not
  g689
  (
    n652,
    n203
  );


  buf
  g690
  (
    n526,
    n372
  );


  buf
  g691
  (
    n970,
    n121
  );


  buf
  g692
  (
    n1144,
    n218
  );


  buf
  g693
  (
    n641,
    n108
  );


  not
  g694
  (
    n1059,
    n208
  );


  buf
  g695
  (
    n613,
    n127
  );


  not
  g696
  (
    n842,
    n336
  );


  not
  g697
  (
    n605,
    n259
  );


  buf
  g698
  (
    n960,
    n296
  );


  buf
  g699
  (
    n703,
    n233
  );


  buf
  g700
  (
    n578,
    n172
  );


  not
  g701
  (
    n996,
    n162
  );


  buf
  g702
  (
    n984,
    n349
  );


  not
  g703
  (
    n849,
    n384
  );


  not
  g704
  (
    n1179,
    n313
  );


  not
  g705
  (
    n1020,
    n261
  );


  not
  g706
  (
    KeyWire_0_25,
    n201
  );


  not
  g707
  (
    n740,
    n327
  );


  buf
  g708
  (
    n1104,
    n147
  );


  not
  g709
  (
    n1076,
    n287
  );


  buf
  g710
  (
    n646,
    n240
  );


  not
  g711
  (
    n918,
    n304
  );


  not
  g712
  (
    n625,
    n155
  );


  buf
  g713
  (
    n998,
    n324
  );


  not
  g714
  (
    n840,
    n181
  );


  buf
  g715
  (
    n924,
    n369
  );


  not
  g716
  (
    n745,
    n211
  );


  buf
  g717
  (
    n983,
    n354
  );


  not
  g718
  (
    n734,
    n258
  );


  buf
  g719
  (
    KeyWire_0_10,
    n231
  );


  buf
  g720
  (
    n495,
    n266
  );


  buf
  g721
  (
    n473,
    n118
  );


  buf
  g722
  (
    n593,
    n178
  );


  not
  g723
  (
    n834,
    n240
  );


  buf
  g724
  (
    n749,
    n318
  );


  buf
  g725
  (
    n817,
    n247
  );


  not
  g726
  (
    n946,
    n185
  );


  not
  g727
  (
    n1046,
    n120
  );


  buf
  g728
  (
    n527,
    n198
  );


  buf
  g729
  (
    n627,
    n260
  );


  buf
  g730
  (
    n505,
    n191
  );


  buf
  g731
  (
    n547,
    n349
  );


  buf
  g732
  (
    n451,
    n190
  );


  buf
  g733
  (
    n712,
    n330
  );


  buf
  g734
  (
    n798,
    n311
  );


  buf
  g735
  (
    n608,
    n146
  );


  buf
  g736
  (
    n532,
    n140
  );


  buf
  g737
  (
    n1117,
    n289
  );


  buf
  g738
  (
    n498,
    n176
  );


  not
  g739
  (
    n561,
    n307
  );


  buf
  g740
  (
    n982,
    n164
  );


  not
  g741
  (
    n763,
    n256
  );


  not
  g742
  (
    n642,
    n229
  );


  not
  g743
  (
    n663,
    n239
  );


  buf
  g744
  (
    n728,
    n128
  );


  buf
  g745
  (
    n643,
    n374
  );


  not
  g746
  (
    n638,
    n156
  );


  buf
  g747
  (
    n717,
    n206
  );


  buf
  g748
  (
    n458,
    n385
  );


  buf
  g749
  (
    n460,
    n186
  );


  buf
  g750
  (
    n540,
    n187
  );


  not
  g751
  (
    n452,
    n352
  );


  buf
  g752
  (
    n706,
    n314
  );


  buf
  g753
  (
    n612,
    n140
  );


  buf
  g754
  (
    n991,
    n300
  );


  not
  g755
  (
    n682,
    n384
  );


  buf
  g756
  (
    n1133,
    n322
  );


  buf
  g757
  (
    n1003,
    n177
  );


  not
  g758
  (
    n647,
    n296
  );


  not
  g759
  (
    n711,
    n132
  );


  not
  g760
  (
    n607,
    n116
  );


  buf
  g761
  (
    n669,
    n241
  );


  buf
  g762
  (
    n621,
    n374
  );


  buf
  g763
  (
    n718,
    n306
  );


  not
  g764
  (
    n1057,
    n116
  );


  buf
  g765
  (
    n630,
    n340
  );


  not
  g766
  (
    n1038,
    n143
  );


  not
  g767
  (
    n1162,
    n289
  );


  not
  g768
  (
    n797,
    n153
  );


  buf
  g769
  (
    n1071,
    n122
  );


  buf
  g770
  (
    n1002,
    n150
  );


  buf
  g771
  (
    n867,
    n334
  );


  buf
  g772
  (
    n904,
    n163
  );


  not
  g773
  (
    n1094,
    n207
  );


  not
  g774
  (
    n506,
    n273
  );


  not
  g775
  (
    n782,
    n254
  );


  buf
  g776
  (
    n1168,
    n176
  );


  buf
  g777
  (
    n724,
    n222
  );


  buf
  g778
  (
    n879,
    n204
  );


  buf
  g779
  (
    n1060,
    n284
  );


  buf
  g780
  (
    n829,
    n353
  );


  not
  g781
  (
    n1097,
    n130
  );


  buf
  g782
  (
    n655,
    n306
  );


  not
  g783
  (
    n755,
    n121
  );


  not
  g784
  (
    n1084,
    n138
  );


  or
  g785
  (
    n1145,
    n226,
    n142
  );


  nand
  g786
  (
    n549,
    n308,
    n345
  );


  xnor
  g787
  (
    n1148,
    n290,
    n317
  );


  and
  g788
  (
    n565,
    n108,
    n227
  );


  xor
  g789
  (
    n1172,
    n284,
    n167
  );


  nand
  g790
  (
    n818,
    n300,
    n148
  );


  nand
  g791
  (
    n927,
    n312,
    n147
  );


  xor
  g792
  (
    n528,
    n313,
    n137
  );


  nand
  g793
  (
    n785,
    n158,
    n320
  );


  nand
  g794
  (
    n801,
    n106,
    n159
  );


  nor
  g795
  (
    n1114,
    n370,
    n266
  );


  or
  g796
  (
    n1042,
    n113,
    n276
  );


  xor
  g797
  (
    n1035,
    n141,
    n142
  );


  and
  g798
  (
    n636,
    n225,
    n245
  );


  nand
  g799
  (
    n658,
    n214,
    n381
  );


  xor
  g800
  (
    n633,
    n346,
    n149
  );


  and
  g801
  (
    n1167,
    n302,
    n184
  );


  xnor
  g802
  (
    n515,
    n247,
    n294
  );


  xor
  g803
  (
    n455,
    n263,
    n297
  );


  nor
  g804
  (
    n468,
    n358,
    n270
  );


  nor
  g805
  (
    n1178,
    n114,
    n117
  );


  nor
  g806
  (
    n899,
    n177,
    n151
  );


  nand
  g807
  (
    n480,
    n168,
    n115
  );


  nand
  g808
  (
    n958,
    n182,
    n323
  );


  xnor
  g809
  (
    n486,
    n320,
    n234
  );


  nor
  g810
  (
    KeyWire_0_7,
    n264,
    n216
  );


  nand
  g811
  (
    n1083,
    n208,
    n165
  );


  and
  g812
  (
    n1053,
    n240,
    n370
  );


  xnor
  g813
  (
    n1140,
    n378,
    n205
  );


  or
  g814
  (
    n795,
    n177,
    n109
  );


  nand
  g815
  (
    n461,
    n348,
    n108
  );


  nor
  g816
  (
    n963,
    n378,
    n218
  );


  xor
  g817
  (
    n796,
    n277,
    n330
  );


  and
  g818
  (
    n892,
    n384,
    n203
  );


  xnor
  g819
  (
    n919,
    n287,
    n355
  );


  nor
  g820
  (
    n1103,
    n146,
    n212
  );


  nor
  g821
  (
    n783,
    n343,
    n249
  );


  xor
  g822
  (
    n965,
    n254,
    n355
  );


  xnor
  g823
  (
    n727,
    n203,
    n300
  );


  and
  g824
  (
    n843,
    n338,
    n123
  );


  xor
  g825
  (
    n803,
    n243,
    n163
  );


  and
  g826
  (
    KeyWire_0_18,
    n347,
    n307
  );


  xnor
  g827
  (
    n716,
    n278,
    n209
  );


  or
  g828
  (
    n476,
    n217,
    n189
  );


  xor
  g829
  (
    n602,
    n194,
    n268
  );


  xnor
  g830
  (
    n1181,
    n295,
    n140
  );


  and
  g831
  (
    n1051,
    n332,
    n257
  );


  xor
  g832
  (
    n903,
    n188,
    n122
  );


  or
  g833
  (
    n854,
    n369,
    n324
  );


  xnor
  g834
  (
    n520,
    n194,
    n277
  );


  and
  g835
  (
    n776,
    n379,
    n305
  );


  xor
  g836
  (
    n604,
    n281,
    n178
  );


  nand
  g837
  (
    n990,
    n136,
    n151
  );


  xor
  g838
  (
    n564,
    n134,
    n272
  );


  or
  g839
  (
    n944,
    n309,
    n303
  );


  nor
  g840
  (
    n1154,
    n171,
    n190
  );


  or
  g841
  (
    n574,
    n306,
    n360
  );


  xor
  g842
  (
    n812,
    n272,
    n230
  );


  and
  g843
  (
    n847,
    n341,
    n185
  );


  xor
  g844
  (
    n503,
    n132,
    n377
  );


  nand
  g845
  (
    n1098,
    n151,
    n120
  );


  nand
  g846
  (
    n499,
    n335,
    n307
  );


  xnor
  g847
  (
    KeyWire_0_11,
    n295,
    n302
  );


  nand
  g848
  (
    n736,
    n239,
    n172
  );


  nor
  g849
  (
    n831,
    n318,
    n270
  );


  xnor
  g850
  (
    n977,
    n113,
    n321
  );


  xor
  g851
  (
    n698,
    n288,
    n279
  );


  and
  g852
  (
    KeyWire_0_28,
    n182,
    n137
  );


  nor
  g853
  (
    n677,
    n339,
    n296
  );


  nand
  g854
  (
    n594,
    n283,
    n174
  );


  nor
  g855
  (
    n909,
    n330,
    n213
  );


  xnor
  g856
  (
    n1171,
    n248,
    n209
  );


  xor
  g857
  (
    n666,
    n160,
    n364
  );


  nand
  g858
  (
    n695,
    n227,
    n183
  );


  or
  g859
  (
    n619,
    n299,
    n375
  );


  nor
  g860
  (
    n1085,
    n135,
    n224
  );


  xnor
  g861
  (
    n1149,
    n186,
    n335
  );


  nand
  g862
  (
    n890,
    n256,
    n211
  );


  or
  g863
  (
    n576,
    n166,
    n165
  );


  nand
  g864
  (
    n543,
    n148,
    n335
  );


  xor
  g865
  (
    n587,
    n361,
    n285
  );


  xor
  g866
  (
    n833,
    n133,
    n160
  );


  xnor
  g867
  (
    KeyWire_0_13,
    n341,
    n331
  );


  nand
  g868
  (
    n691,
    n181,
    n294
  );


  xor
  g869
  (
    n1024,
    n325,
    n326
  );


  nand
  g870
  (
    KeyWire_0_12,
    n331,
    n233
  );


  or
  g871
  (
    n1165,
    n308,
    n349
  );


  nand
  g872
  (
    n916,
    n282,
    n299
  );


  xor
  g873
  (
    n1102,
    n375,
    n348
  );


  nor
  g874
  (
    n533,
    n192,
    n257
  );


  nand
  g875
  (
    n683,
    n347,
    n120
  );


  xor
  g876
  (
    n629,
    n118,
    n147
  );


  nor
  g877
  (
    n1009,
    n180,
    n364
  );


  nand
  g878
  (
    n519,
    n265,
    n130
  );


  and
  g879
  (
    n591,
    n274,
    n225
  );


  nand
  g880
  (
    n811,
    n127,
    n365
  );


  xnor
  g881
  (
    n509,
    n128,
    n259
  );


  xnor
  g882
  (
    n800,
    n291,
    n177
  );


  and
  g883
  (
    n493,
    n160,
    n365
  );


  nand
  g884
  (
    n1055,
    n331,
    n170
  );


  xnor
  g885
  (
    n821,
    n153,
    n263
  );


  or
  g886
  (
    n889,
    n171,
    n228
  );


  xnor
  g887
  (
    n640,
    n225,
    n189
  );


  xor
  g888
  (
    n730,
    n153,
    n110
  );


  xnor
  g889
  (
    n881,
    n151,
    n232
  );


  xor
  g890
  (
    n700,
    n145,
    n167
  );


  or
  g891
  (
    n457,
    n271,
    n129
  );


  xor
  g892
  (
    n491,
    n344,
    n319
  );


  xor
  g893
  (
    n846,
    n163,
    n193
  );


  xor
  g894
  (
    n624,
    n199,
    n334
  );


  xor
  g895
  (
    n954,
    n186,
    n250
  );


  xor
  g896
  (
    n1175,
    n220,
    n173
  );


  xor
  g897
  (
    n805,
    n168,
    n166
  );


  and
  g898
  (
    n1081,
    n224,
    n230
  );


  nor
  g899
  (
    n988,
    n379,
    n244
  );


  or
  g900
  (
    n709,
    n152,
    n173
  );


  nor
  g901
  (
    n689,
    n199,
    n106
  );


  xnor
  g902
  (
    n678,
    n189,
    n340
  );


  xnor
  g903
  (
    n964,
    n278,
    n213
  );


  or
  g904
  (
    n1031,
    n332,
    n381
  );


  xnor
  g905
  (
    n661,
    n366,
    n206
  );


  xnor
  g906
  (
    n1120,
    n319,
    n157
  );


  or
  g907
  (
    n694,
    n338,
    n277
  );


  nor
  g908
  (
    n512,
    n237,
    n352
  );


  nor
  g909
  (
    n459,
    n245,
    n332
  );


  nand
  g910
  (
    n974,
    n139,
    n106
  );


  xnor
  g911
  (
    n878,
    n250,
    n134
  );


  nor
  g912
  (
    n597,
    n116,
    n228
  );


  nor
  g913
  (
    n1105,
    n237,
    n319
  );


  xor
  g914
  (
    n552,
    n324,
    n193
  );


  and
  g915
  (
    n802,
    n253,
    n251
  );


  and
  g916
  (
    n644,
    n234,
    n360
  );


  and
  g917
  (
    n911,
    n197,
    n180
  );


  or
  g918
  (
    n598,
    n219,
    n125
  );


  xnor
  g919
  (
    n1070,
    n122,
    n196
  );


  xnor
  g920
  (
    n497,
    n279,
    n155
  );


  xor
  g921
  (
    n754,
    n244,
    n264
  );


  or
  g922
  (
    n893,
    n223,
    n250
  );


  and
  g923
  (
    n622,
    n144,
    n139
  );


  and
  g924
  (
    n1058,
    n183,
    n172
  );


  nand
  g925
  (
    n844,
    n197,
    n268
  );


  or
  g926
  (
    n553,
    n216,
    n247
  );


  nor
  g927
  (
    n686,
    n118,
    n327
  );


  nor
  g928
  (
    n894,
    n129,
    n185
  );


  nand
  g929
  (
    n1158,
    n215,
    n358
  );


  and
  g930
  (
    n500,
    n217,
    n273
  );


  nor
  g931
  (
    n862,
    n119,
    n385
  );


  xor
  g932
  (
    n696,
    n146,
    n337
  );


  and
  g933
  (
    n962,
    n183,
    n358
  );


  xnor
  g934
  (
    n449,
    n200,
    n316
  );


  and
  g935
  (
    n637,
    n204,
    n269
  );


  or
  g936
  (
    n1047,
    n355,
    n223
  );


  nand
  g937
  (
    n1011,
    n126,
    n109
  );


  xnor
  g938
  (
    n589,
    n145,
    n236
  );


  and
  g939
  (
    KeyWire_0_9,
    n169,
    n292
  );


  or
  g940
  (
    n1080,
    n200,
    n138
  );


  xnor
  g941
  (
    n507,
    n175,
    n179
  );


  not
  g942
  (
    n1039,
    n333
  );


  or
  g943
  (
    n914,
    n106,
    n327
  );


  and
  g944
  (
    n1082,
    n274,
    n242
  );


  xnor
  g945
  (
    n1034,
    n368,
    n181
  );


  xnor
  g946
  (
    n541,
    n380,
    n157
  );


  and
  g947
  (
    n959,
    n274,
    n195
  );


  or
  g948
  (
    n923,
    n365,
    n353
  );


  nor
  g949
  (
    n539,
    n170,
    n145
  );


  xnor
  g950
  (
    n1138,
    n195,
    n369
  );


  and
  g951
  (
    n1077,
    n241,
    n263
  );


  xor
  g952
  (
    n1026,
    n285,
    n372
  );


  xor
  g953
  (
    n463,
    n202,
    n112
  );


  xnor
  g954
  (
    n707,
    n221,
    n180
  );


  nand
  g955
  (
    n1091,
    n281,
    n207
  );


  or
  g956
  (
    n634,
    n378,
    n276
  );


  xor
  g957
  (
    n1036,
    n310,
    n370
  );


  and
  g958
  (
    n999,
    n188,
    n382
  );


  nor
  g959
  (
    n483,
    n293,
    n195
  );


  xor
  g960
  (
    n762,
    n368,
    n162
  );


  nor
  g961
  (
    n445,
    n350,
    n260
  );


  xnor
  g962
  (
    n573,
    n176,
    n348
  );


  nand
  g963
  (
    n1008,
    n248,
    n235
  );


  nor
  g964
  (
    n1139,
    n297,
    n277
  );


  nor
  g965
  (
    n1066,
    n260,
    n274
  );


  nor
  g966
  (
    n1106,
    n331,
    n224
  );


  nor
  g967
  (
    n896,
    n158,
    n361
  );


  nand
  g968
  (
    n976,
    n361,
    n282
  );


  nand
  g969
  (
    n973,
    n122,
    n325
  );


  xor
  g970
  (
    n1045,
    n223,
    n264
  );


  nand
  g971
  (
    n931,
    n317,
    n301
  );


  xnor
  g972
  (
    n443,
    n307,
    n322
  );


  xnor
  g973
  (
    n933,
    n142,
    n267
  );


  xor
  g974
  (
    n1159,
    n322,
    n168
  );


  nor
  g975
  (
    n687,
    n154,
    n344
  );


  nand
  g976
  (
    n841,
    n226,
    n312
  );


  and
  g977
  (
    n744,
    n111,
    n321
  );


  and
  g978
  (
    n511,
    n359,
    n272
  );


  nor
  g979
  (
    KeyWire_0_16,
    n313,
    n126
  );


  xor
  g980
  (
    n671,
    n169,
    n381
  );


  or
  g981
  (
    n708,
    n367,
    n348
  );


  nor
  g982
  (
    n1013,
    n232,
    n165
  );


  xor
  g983
  (
    n1156,
    n179,
    n280
  );


  xor
  g984
  (
    n1023,
    n235,
    n297
  );


  nand
  g985
  (
    n1124,
    n154,
    n120
  );


  xnor
  g986
  (
    n675,
    n354,
    n299
  );


  and
  g987
  (
    n1112,
    n338,
    n185
  );


  xor
  g988
  (
    n522,
    n349,
    n142
  );


  xnor
  g989
  (
    n680,
    n233,
    n180
  );


  nand
  g990
  (
    n714,
    n110,
    n162
  );


  and
  g991
  (
    n470,
    n280,
    n301
  );


  nand
  g992
  (
    n665,
    n259,
    n137
  );


  nor
  g993
  (
    n713,
    n343,
    n279
  );


  xor
  g994
  (
    n748,
    n241,
    n262
  );


  or
  g995
  (
    n615,
    n297,
    n196
  );


  xor
  g996
  (
    n887,
    n246,
    n276
  );


  nor
  g997
  (
    n828,
    n242,
    n171
  );


  and
  g998
  (
    n595,
    n372,
    n201
  );


  or
  g999
  (
    n863,
    n219,
    n362
  );


  xnor
  g1000
  (
    n1090,
    n386,
    n237
  );


  or
  g1001
  (
    n912,
    n138,
    n362
  );


  xnor
  g1002
  (
    n733,
    n286,
    n194
  );


  and
  g1003
  (
    n848,
    n367,
    n336
  );


  nand
  g1004
  (
    n1027,
    n144,
    n209
  );


  and
  g1005
  (
    n825,
    n140,
    n124
  );


  nand
  g1006
  (
    n657,
    n310,
    n210
  );


  xor
  g1007
  (
    n835,
    n298,
    n366
  );


  xor
  g1008
  (
    n850,
    n291,
    n278
  );


  nand
  g1009
  (
    n588,
    n131,
    n239
  );


  or
  g1010
  (
    n603,
    n373,
    n356
  );


  xor
  g1011
  (
    n1123,
    n266,
    n164
  );


  nand
  g1012
  (
    n751,
    n303,
    n376
  );


  nor
  g1013
  (
    n1004,
    n191,
    n221
  );


  and
  g1014
  (
    n910,
    n132,
    n267
  );


  nor
  g1015
  (
    n494,
    n382,
    n383
  );


  nand
  g1016
  (
    n1176,
    n283,
    n148
  );


  xnor
  g1017
  (
    n926,
    n117,
    n258
  );


  xnor
  g1018
  (
    n584,
    n293,
    n347
  );


  xor
  g1019
  (
    n869,
    n269,
    n133
  );


  nand
  g1020
  (
    n670,
    n205,
    n365
  );


  nand
  g1021
  (
    n937,
    n375,
    n363
  );


  nand
  g1022
  (
    n978,
    n354,
    n255
  );


  or
  g1023
  (
    n949,
    n136,
    n135
  );


  nand
  g1024
  (
    n859,
    n109,
    n144
  );


  xnor
  g1025
  (
    n790,
    n309,
    n124
  );


  and
  g1026
  (
    n1078,
    n263,
    n243
  );


  xnor
  g1027
  (
    n1014,
    n339,
    n251
  );


  and
  g1028
  (
    n524,
    n315,
    n254
  );


  or
  g1029
  (
    n1115,
    n345,
    n342
  );


  xnor
  g1030
  (
    n558,
    n368,
    n265
  );


  nor
  g1031
  (
    KeyWire_0_5,
    n220,
    n255
  );


  xor
  g1032
  (
    n884,
    n252,
    n175
  );


  xor
  g1033
  (
    n897,
    n252,
    n224
  );


  xnor
  g1034
  (
    n1182,
    n386,
    n114
  );


  nor
  g1035
  (
    n442,
    n305,
    n201
  );


  nor
  g1036
  (
    n906,
    n286,
    n179
  );


  nand
  g1037
  (
    n837,
    n110,
    n212
  );


  nor
  g1038
  (
    n1130,
    n166,
    n242
  );


  or
  g1039
  (
    n568,
    n208,
    n287
  );


  xor
  g1040
  (
    n525,
    n328,
    n271
  );


  and
  g1041
  (
    n1183,
    n371,
    n304
  );


  or
  g1042
  (
    n1092,
    n171,
    n220
  );


  and
  g1043
  (
    n836,
    n136,
    n351
  );


  and
  g1044
  (
    n951,
    n129,
    n298
  );


  or
  g1045
  (
    n448,
    n350,
    n169
  );


  xor
  g1046
  (
    n1062,
    n345,
    n321
  );


  and
  g1047
  (
    n467,
    n217,
    n329
  );


  nor
  g1048
  (
    n1029,
    n281,
    n381
  );


  xor
  g1049
  (
    n864,
    n187,
    n342
  );


  and
  g1050
  (
    n967,
    n219,
    n294
  );


  xnor
  g1051
  (
    n917,
    n281,
    n305
  );


  xor
  g1052
  (
    n1099,
    n202,
    n135
  );


  xor
  g1053
  (
    n861,
    n131,
    n351
  );


  nand
  g1054
  (
    n764,
    n323,
    n164
  );


  xnor
  g1055
  (
    n1068,
    n135,
    n160
  );


  or
  g1056
  (
    n940,
    n188,
    n205
  );


  nor
  g1057
  (
    n504,
    n155,
    n234
  );


  nand
  g1058
  (
    n685,
    n259,
    n339
  );


  nor
  g1059
  (
    n1143,
    n125,
    n260
  );


  xnor
  g1060
  (
    n866,
    n298,
    n121
  );


  xor
  g1061
  (
    n1018,
    n212,
    n380
  );


  xnor
  g1062
  (
    n692,
    n114,
    n266
  );


  xor
  g1063
  (
    n681,
    n330,
    n198
  );


  and
  g1064
  (
    n632,
    n173,
    n345
  );


  nor
  g1065
  (
    n567,
    n258,
    n214
  );


  nor
  g1066
  (
    n1166,
    n196,
    n231
  );


  or
  g1067
  (
    n875,
    n159,
    n181
  );


  nand
  g1068
  (
    n972,
    n133,
    n230
  );


  and
  g1069
  (
    n902,
    n337,
    n170
  );


  nor
  g1070
  (
    n477,
    n358,
    n197
  );


  or
  g1071
  (
    n945,
    n295,
    n374
  );


  nor
  g1072
  (
    n651,
    n215,
    n228
  );


  or
  g1073
  (
    n1136,
    n173,
    n253
  );


  nor
  g1074
  (
    n551,
    n137,
    n364
  );


  or
  g1075
  (
    n1019,
    n328,
    n357
  );


  and
  g1076
  (
    n581,
    n228,
    n209
  );


  xnor
  g1077
  (
    n882,
    n385,
    n376
  );


  nor
  g1078
  (
    n806,
    n221,
    n175
  );


  or
  g1079
  (
    n1006,
    n170,
    n199
  );


  nand
  g1080
  (
    n907,
    n187,
    n301
  );


  nand
  g1081
  (
    n446,
    n222,
    n149
  );


  nand
  g1082
  (
    n610,
    n333,
    n315
  );


  xnor
  g1083
  (
    n555,
    n218,
    n156
  );


  nand
  g1084
  (
    n1153,
    n316,
    n283
  );


  xnor
  g1085
  (
    n858,
    n284,
    n216
  );


  nor
  g1086
  (
    n779,
    n193,
    n159
  );


  nor
  g1087
  (
    n857,
    n338,
    n357
  );


  or
  g1088
  (
    n784,
    n286,
    n379
  );


  xor
  g1089
  (
    n1101,
    n383,
    n118
  );


  nand
  g1090
  (
    n600,
    n255,
    n361
  );


  xnor
  g1091
  (
    n865,
    n332,
    n117
  );


  or
  g1092
  (
    n688,
    n353,
    n367
  );


  nand
  g1093
  (
    n942,
    n141,
    n114
  );


  xnor
  g1094
  (
    n697,
    n222,
    n315
  );


  xnor
  g1095
  (
    n488,
    n379,
    n119
  );


  nand
  g1096
  (
    n870,
    n343,
    n176
  );


  nor
  g1097
  (
    n482,
    n214,
    n165
  );


  xor
  g1098
  (
    n586,
    n280,
    n255
  );


  nand
  g1099
  (
    n441,
    n326,
    n124
  );


  xor
  g1100
  (
    n1073,
    n362,
    n382
  );


  nand
  g1101
  (
    n1184,
    n183,
    n290
  );


  nor
  g1102
  (
    n660,
    n127,
    n275
  );


  and
  g1103
  (
    n830,
    n377,
    n273
  );


  or
  g1104
  (
    n853,
    n111,
    n370
  );


  xor
  g1105
  (
    n838,
    n366,
    n236
  );


  and
  g1106
  (
    n981,
    n382,
    n367
  );


  xnor
  g1107
  (
    n1134,
    n280,
    n347
  );


  nand
  g1108
  (
    n814,
    n158,
    n235
  );


  and
  g1109
  (
    n529,
    n271,
    n378
  );


  and
  g1110
  (
    n1086,
    n204,
    n184
  );


  xor
  g1111
  (
    n938,
    n265,
    n240
  );


  nand
  g1112
  (
    n1185,
    n172,
    n333
  );


  and
  g1113
  (
    n810,
    n384,
    n247
  );


  nand
  g1114
  (
    n888,
    n132,
    n273
  );


  or
  g1115
  (
    n654,
    n275,
    n126
  );


  nand
  g1116
  (
    n1079,
    n339,
    n208
  );


  xnor
  g1117
  (
    n1037,
    n199,
    n311
  );


  xnor
  g1118
  (
    n943,
    n244,
    n119
  );


  nor
  g1119
  (
    n1152,
    n293,
    n141
  );


  nor
  g1120
  (
    n537,
    n275,
    n256
  );


  or
  g1121
  (
    n980,
    n322,
    n179
  );


  xnor
  g1122
  (
    n668,
    n108,
    n282
  );


  or
  g1123
  (
    n1061,
    n150,
    n314
  );


  xnor
  g1124
  (
    n860,
    n329,
    n287
  );


  and
  g1125
  (
    n774,
    n316,
    n169
  );


  nand
  g1126
  (
    n1126,
    n291,
    n111
  );


  xnor
  g1127
  (
    n735,
    n238,
    n278
  );


  nor
  g1128
  (
    n1125,
    n184,
    n268
  );


  nand
  g1129
  (
    n950,
    n334,
    n112
  );


  nor
  g1130
  (
    n534,
    n308,
    n189
  );


  xnor
  g1131
  (
    n1129,
    n270,
    n156
  );


  xnor
  g1132
  (
    n577,
    n200,
    n125
  );


  or
  g1133
  (
    n1089,
    n321,
    n130
  );


  nand
  g1134
  (
    n1005,
    n308,
    n326
  );


  and
  g1135
  (
    n514,
    n238,
    n293
  );


  nor
  g1136
  (
    n948,
    n238,
    n141
  );


  and
  g1137
  (
    n490,
    n215,
    n139
  );


  nand
  g1138
  (
    n623,
    n298,
    n150
  );


  xnor
  g1139
  (
    n921,
    n213,
    n191
  );


  xnor
  g1140
  (
    n1180,
    n290,
    n373
  );


  and
  g1141
  (
    n956,
    n380,
    n309
  );


  or
  g1142
  (
    n648,
    n343,
    n227
  );


  and
  g1143
  (
    n1064,
    n253,
    n267
  );


  nand
  g1144
  (
    n766,
    n306,
    n236
  );


  or
  g1145
  (
    n617,
    n325,
    n245
  );


  nor
  g1146
  (
    n450,
    n192,
    n360
  );


  xnor
  g1147
  (
    n1177,
    n194,
    n302
  );


  nor
  g1148
  (
    n572,
    n286,
    n113
  );


  nor
  g1149
  (
    n908,
    n303,
    n250
  );


  nor
  g1150
  (
    n1063,
    n252,
    n221
  );


  or
  g1151
  (
    n585,
    n175,
    n225
  );


  or
  g1152
  (
    n1135,
    n202,
    n168
  );


  or
  g1153
  (
    n1033,
    n121,
    n156
  );


  or
  g1154
  (
    n1000,
    n203,
    n337
  );


  and
  g1155
  (
    n781,
    n265,
    n344
  );


  or
  g1156
  (
    n487,
    n155,
    n337
  );


  xor
  g1157
  (
    n1141,
    n239,
    n386
  );


  nor
  g1158
  (
    n968,
    n282,
    n356
  );


  xnor
  g1159
  (
    n1107,
    n202,
    n117
  );


  or
  g1160
  (
    n523,
    n218,
    n323
  );


  or
  g1161
  (
    n1146,
    n205,
    n159
  );


  or
  g1162
  (
    n1028,
    n318,
    n164
  );


  xnor
  g1163
  (
    n559,
    n232,
    n146
  );


  and
  g1164
  (
    n1244,
    n815,
    n397,
    n825,
    n394
  );


  nor
  g1165
  (
    n1380,
    n1045,
    n427,
    n1052,
    n530
  );


  xor
  g1166
  (
    n1301,
    n424,
    n616,
    n774,
    n974
  );


  and
  g1167
  (
    n1368,
    n1009,
    n849,
    n891,
    n719
  );


  xnor
  g1168
  (
    n1330,
    n914,
    n580,
    n499,
    n734
  );


  or
  g1169
  (
    n1313,
    n589,
    n567,
    n994,
    n723
  );


  nor
  g1170
  (
    n1210,
    n421,
    n727,
    n869,
    n647
  );


  or
  g1171
  (
    n1409,
    n928,
    n753,
    n1006,
    n1055
  );


  nor
  g1172
  (
    n1192,
    n395,
    n583,
    n854,
    n962
  );


  and
  g1173
  (
    n1211,
    n870,
    n389,
    n417,
    n388
  );


  xnor
  g1174
  (
    n1319,
    n901,
    n460,
    n1096,
    n427
  );


  or
  g1175
  (
    n1363,
    n400,
    n771,
    n1012,
    n668
  );


  xnor
  g1176
  (
    n1290,
    n561,
    n1021,
    n418,
    n729
  );


  and
  g1177
  (
    n1196,
    n761,
    n415,
    n552,
    n420
  );


  xnor
  g1178
  (
    n1220,
    n767,
    n439,
    n396,
    n388
  );


  nand
  g1179
  (
    n1255,
    n408,
    n1069,
    n593,
    n496
  );


  xor
  g1180
  (
    n1316,
    n844,
    n853,
    n475,
    n483
  );


  xnor
  g1181
  (
    n1304,
    n390,
    n1042,
    n387,
    n1048
  );


  nand
  g1182
  (
    n1324,
    n412,
    n565,
    n795,
    n575
  );


  and
  g1183
  (
    n1295,
    n706,
    n908,
    n425,
    n401
  );


  or
  g1184
  (
    n1187,
    n625,
    n536,
    n760,
    n741
  );


  or
  g1185
  (
    n1205,
    n603,
    n680,
    n398,
    n652
  );


  and
  g1186
  (
    n1361,
    n1098,
    n969,
    n1094,
    n952
  );


  nand
  g1187
  (
    n1217,
    n714,
    n477,
    n971,
    n983
  );


  nor
  g1188
  (
    n1303,
    n820,
    n566,
    n700,
    n1095
  );


  and
  g1189
  (
    n1279,
    n467,
    n389,
    n703,
    n390
  );


  nor
  g1190
  (
    n1404,
    n557,
    n960,
    n717,
    n1000
  );


  xor
  g1191
  (
    n1232,
    n834,
    n1076,
    n429,
    n544
  );


  and
  g1192
  (
    n1200,
    n412,
    n682,
    n421,
    n389
  );


  and
  g1193
  (
    n1401,
    n523,
    n394,
    n412,
    n817
  );


  and
  g1194
  (
    n1348,
    n831,
    n419,
    n521,
    n395
  );


  nand
  g1195
  (
    n1386,
    n400,
    n1044,
    n769,
    n425
  );


  nand
  g1196
  (
    n1389,
    n411,
    n438,
    n440,
    n1083
  );


  or
  g1197
  (
    n1248,
    n404,
    n990,
    n509,
    n396
  );


  nand
  g1198
  (
    n1340,
    n898,
    n1094,
    n980,
    n739
  );


  nand
  g1199
  (
    n1207,
    n1019,
    n392,
    n689,
    n679
  );


  nand
  g1200
  (
    n1325,
    n539,
    n425,
    n393,
    n654
  );


  and
  g1201
  (
    n1281,
    n791,
    n1090,
    n436,
    n942
  );


  and
  g1202
  (
    n1312,
    n744,
    n673,
    n740,
    n1037
  );


  nor
  g1203
  (
    n1241,
    n775,
    n661,
    n592,
    n413
  );


  xnor
  g1204
  (
    n1209,
    n709,
    n404,
    n559,
    n401
  );


  nor
  g1205
  (
    n1294,
    n459,
    n888,
    n401,
    n810
  );


  or
  g1206
  (
    n1407,
    n588,
    n1066,
    n855,
    n443
  );


  xor
  g1207
  (
    n1346,
    n1057,
    n998,
    n1082,
    n683
  );


  nand
  g1208
  (
    n1359,
    n407,
    n428,
    n510,
    n833
  );


  nand
  g1209
  (
    n1345,
    n471,
    n642,
    n394,
    n678
  );


  nor
  g1210
  (
    n1194,
    n594,
    n554,
    n697,
    n1098
  );


  nand
  g1211
  (
    n1395,
    n419,
    n406,
    n798,
    n759
  );


  nor
  g1212
  (
    n1379,
    n395,
    n1016,
    n454,
    n708
  );


  nor
  g1213
  (
    n1240,
    n865,
    n601,
    n958,
    n515
  );


  or
  g1214
  (
    n1267,
    n564,
    n950,
    n821,
    n733
  );


  xor
  g1215
  (
    n1298,
    n413,
    n1051,
    n422,
    n659
  );


  nand
  g1216
  (
    n1362,
    n786,
    n742,
    n961,
    n428
  );


  and
  g1217
  (
    n1375,
    n486,
    n780,
    n414,
    n883
  );


  and
  g1218
  (
    n1253,
    n406,
    n915,
    n646,
    n1094
  );


  xnor
  g1219
  (
    n1302,
    n446,
    n502,
    n437,
    n726
  );


  xor
  g1220
  (
    n1191,
    n822,
    n465,
    n955,
    n713
  );


  nor
  g1221
  (
    n1382,
    n438,
    n781,
    n556,
    n1008
  );


  xnor
  g1222
  (
    n1349,
    n826,
    n438,
    n887,
    n605
  );


  xnor
  g1223
  (
    n1405,
    n524,
    n462,
    n417,
    n976
  );


  xor
  g1224
  (
    n1293,
    n857,
    n1004,
    n492,
    n766
  );


  and
  g1225
  (
    n1305,
    n450,
    n995,
    n435,
    n1068
  );


  xnor
  g1226
  (
    n1383,
    n951,
    n1064,
    n1097,
    n787
  );


  or
  g1227
  (
    n1299,
    n856,
    n830,
    n1059,
    n590
  );


  nand
  g1228
  (
    n1343,
    n639,
    n676,
    n964,
    n868
  );


  xnor
  g1229
  (
    n1402,
    n966,
    n1086,
    n392,
    n527
  );


  xor
  g1230
  (
    n1249,
    n1036,
    n823,
    n688,
    n685
  );


  nor
  g1231
  (
    n1287,
    n432,
    n547,
    n692,
    n681
  );


  nand
  g1232
  (
    n1332,
    n391,
    n428,
    n433,
    n796
  );


  nor
  g1233
  (
    n1351,
    n956,
    n463,
    n610,
    n1063
  );


  xnor
  g1234
  (
    n1310,
    n387,
    n794,
    n402,
    n757
  );


  nor
  g1235
  (
    n1226,
    n1003,
    n526,
    n432,
    n439
  );


  xor
  g1236
  (
    n1308,
    n872,
    n481,
    n430,
    n1038
  );


  and
  g1237
  (
    n1260,
    n1077,
    n484,
    n1096,
    n613
  );


  xor
  g1238
  (
    n1236,
    n408,
    n999,
    n435,
    n416
  );


  or
  g1239
  (
    n1373,
    n779,
    n404,
    n698,
    n967
  );


  xor
  g1240
  (
    n1397,
    n422,
    n568,
    n449,
    n599
  );


  nor
  g1241
  (
    n1213,
    n806,
    n752,
    n412,
    n1020
  );


  xor
  g1242
  (
    n1271,
    n935,
    n453,
    n669,
    n549
  );


  nand
  g1243
  (
    n1352,
    n882,
    n1050,
    n1088,
    n925
  );


  nand
  g1244
  (
    n1289,
    n801,
    n430,
    n848,
    n562
  );


  or
  g1245
  (
    n1268,
    n772,
    n871,
    n1075,
    n890
  );


  xnor
  g1246
  (
    n1365,
    n1098,
    n578,
    n777,
    n945
  );


  xor
  g1247
  (
    n1323,
    n480,
    n847,
    n391,
    n829
  );


  nor
  g1248
  (
    n1403,
    n558,
    n650,
    n436,
    n618
  );


  nor
  g1249
  (
    n1193,
    n420,
    n736,
    n735,
    n691
  );


  xnor
  g1250
  (
    n1276,
    n1025,
    n873,
    n604,
    n858
  );


  and
  g1251
  (
    n1206,
    n665,
    n929,
    n725,
    n405
  );


  or
  g1252
  (
    n1378,
    n756,
    n1097,
    n785,
    n1035
  );


  nand
  g1253
  (
    n1355,
    n429,
    n576,
    n1065,
    n538
  );


  and
  g1254
  (
    n1195,
    n987,
    n694,
    n677,
    n474
  );


  nor
  g1255
  (
    n1297,
    n410,
    n1074,
    n842,
    n528
  );


  and
  g1256
  (
    n1318,
    n867,
    n560,
    n946,
    n904
  );


  nor
  g1257
  (
    n1317,
    n933,
    n516,
    n648,
    n514
  );


  and
  g1258
  (
    n1280,
    n404,
    n411,
    n653,
    n828
  );


  xor
  g1259
  (
    n1254,
    n732,
    n612,
    n434,
    n1072
  );


  or
  g1260
  (
    n1273,
    n396,
    n619,
    n860,
    n405
  );


  or
  g1261
  (
    n1284,
    n436,
    n577,
    n470,
    n1084
  );


  xor
  g1262
  (
    n1203,
    n721,
    n878,
    n921,
    n624
  );


  and
  g1263
  (
    n1272,
    n1085,
    n512,
    n423,
    n455
  );


  xnor
  g1264
  (
    n1322,
    n399,
    n418,
    n451,
    n415
  );


  and
  g1265
  (
    n1367,
    n540,
    n485,
    n953,
    n768
  );


  or
  g1266
  (
    n1222,
    n464,
    n418,
    n424,
    n670
  );


  and
  g1267
  (
    n1366,
    n838,
    n570,
    n1096,
    n818
  );


  xnor
  g1268
  (
    n1335,
    n435,
    n426,
    n490,
    n606
  );


  nor
  g1269
  (
    n1266,
    n393,
    n900,
    n409,
    n968
  );


  or
  g1270
  (
    n1329,
    n816,
    n1091,
    n408,
    n563
  );


  and
  g1271
  (
    n1262,
    n912,
    n926,
    n893,
    n710
  );


  nor
  g1272
  (
    n1228,
    n902,
    n614,
    n1015,
    n846
  );


  xor
  g1273
  (
    n1334,
    n1078,
    n948,
    n1039,
    n494
  );


  xor
  g1274
  (
    n1231,
    n472,
    n413,
    n1089,
    n1060
  );


  and
  g1275
  (
    n1197,
    n1094,
    n529,
    n439,
    n984
  );


  or
  g1276
  (
    n1369,
    n837,
    n448,
    n649,
    n439
  );


  or
  g1277
  (
    n1390,
    n657,
    n415,
    n518,
    n730
  );


  xor
  g1278
  (
    n1229,
    n495,
    n466,
    n411,
    n645
  );


  xor
  g1279
  (
    KeyWire_0_22,
    n1054,
    n1058,
    n972,
    n500
  );


  nand
  g1280
  (
    n1370,
    n758,
    n511,
    n667,
    n398
  );


  and
  g1281
  (
    n1201,
    n635,
    n941,
    n1080,
    n482
  );


  or
  g1282
  (
    KeyWire_0_17,
    n406,
    n546,
    n809,
    n394
  );


  xor
  g1283
  (
    n1326,
    n1007,
    n438,
    n426,
    n399
  );


  and
  g1284
  (
    n1331,
    n731,
    n422,
    n431,
    n437
  );


  xnor
  g1285
  (
    n1384,
    n939,
    n919,
    n585,
    n718
  );


  xor
  g1286
  (
    n1247,
    n416,
    n840,
    n789,
    n1033
  );


  or
  g1287
  (
    n1339,
    n686,
    n423,
    n636,
    n1092
  );


  nand
  g1288
  (
    n1314,
    n551,
    n418,
    n803,
    n487
  );


  and
  g1289
  (
    n1291,
    n991,
    n437,
    n862,
    n609
  );


  xnor
  g1290
  (
    n1278,
    n574,
    n1017,
    n620,
    n419
  );


  xnor
  g1291
  (
    n1342,
    n519,
    n1070,
    n747,
    n937
  );


  or
  g1292
  (
    n1360,
    n392,
    n545,
    n881,
    n550
  );


  nor
  g1293
  (
    n1328,
    n637,
    n1091,
    n947,
    n421
  );


  xnor
  g1294
  (
    n1245,
    n674,
    n808,
    n800,
    n397
  );


  or
  g1295
  (
    n1230,
    n746,
    n410,
    n408,
    n628
  );


  or
  g1296
  (
    n1215,
    n403,
    n695,
    n399,
    n684
  );


  or
  g1297
  (
    n1264,
    n409,
    n936,
    n440,
    n836
  );


  xnor
  g1298
  (
    n1356,
    n861,
    n395,
    n595,
    n985
  );


  xor
  g1299
  (
    n1277,
    n864,
    n387,
    n644,
    n930
  );


  xor
  g1300
  (
    n1337,
    n553,
    n903,
    n1067,
    n824
  );


  and
  g1301
  (
    n1234,
    n993,
    n416,
    n621,
    n1062
  );


  xnor
  g1302
  (
    n1261,
    n720,
    n1095,
    n655,
    n911
  );


  nand
  g1303
  (
    n1258,
    n457,
    n750,
    n434,
    n1093
  );


  and
  g1304
  (
    KeyWire_0_1,
    n444,
    n417,
    n799,
    n1028
  );


  nor
  g1305
  (
    n1186,
    n1013,
    n468,
    n778,
    n392
  );


  nand
  g1306
  (
    n1406,
    n426,
    n701,
    n917,
    n1024
  );


  and
  g1307
  (
    n1243,
    n1031,
    n986,
    n555,
    n894
  );


  xor
  g1308
  (
    n1216,
    n874,
    n715,
    n879,
    n1002
  );


  nor
  g1309
  (
    n1257,
    n745,
    n1026,
    n784,
    n897
  );


  or
  g1310
  (
    n1270,
    n431,
    n743,
    n406,
    n886
  );


  xor
  g1311
  (
    KeyWire_0_8,
    n931,
    n569,
    n520,
    n579
  );


  nor
  g1312
  (
    n1309,
    n841,
    n407,
    n489,
    n397
  );


  nor
  g1313
  (
    n1300,
    n433,
    n790,
    n663,
    n591
  );


  xor
  g1314
  (
    n1259,
    n957,
    n640,
    n602,
    n1046
  );


  xnor
  g1315
  (
    n1198,
    n996,
    n1092,
    n420,
    n923
  );


  nand
  g1316
  (
    n1385,
    n788,
    n419,
    n388,
    n525
  );


  or
  g1317
  (
    n1292,
    n707,
    n420,
    n1093,
    n534
  );


  xnor
  g1318
  (
    n1227,
    n711,
    n1047,
    n814,
    n690
  );


  nand
  g1319
  (
    n1275,
    n633,
    n632,
    n1073,
    n1097
  );


  nor
  g1320
  (
    n1256,
    n413,
    n664,
    n909,
    n476
  );


  nand
  g1321
  (
    n1350,
    n396,
    n429,
    n433,
    n532
  );


  nand
  g1322
  (
    n1283,
    n497,
    n805,
    n573,
    n1061
  );


  nand
  g1323
  (
    n1223,
    n441,
    n922,
    n835,
    n403
  );


  nor
  g1324
  (
    n1321,
    n811,
    n425,
    n533,
    n391
  );


  xor
  g1325
  (
    n1398,
    n498,
    n819,
    n918,
    n437
  );


  or
  g1326
  (
    n1358,
    n617,
    n859,
    n431,
    n399
  );


  xor
  g1327
  (
    n1376,
    n479,
    n1093,
    n458,
    n513
  );


  and
  g1328
  (
    n1237,
    n638,
    n631,
    n1014,
    n1056
  );


  xor
  g1329
  (
    n1371,
    n607,
    n920,
    n1030,
    n863
  );


  or
  g1330
  (
    n1338,
    n1001,
    n748,
    n773,
    n426
  );


  or
  g1331
  (
    n1381,
    n906,
    n1098,
    n813,
    n899
  );


  nor
  g1332
  (
    n1377,
    n792,
    n850,
    n989,
    n749
  );


  and
  g1333
  (
    n1214,
    n400,
    n571,
    n876,
    n505
  );


  nor
  g1334
  (
    n1288,
    n447,
    n409,
    n587,
    n1011
  );


  xor
  g1335
  (
    n1219,
    n866,
    n572,
    n469,
    n401
  );


  xnor
  g1336
  (
    n1218,
    n541,
    n782,
    n1005,
    n584
  );


  or
  g1337
  (
    n1274,
    n409,
    n430,
    n755,
    n827
  );


  nand
  g1338
  (
    n1399,
    n531,
    n988,
    n884,
    n770
  );


  and
  g1339
  (
    n1188,
    n581,
    n390,
    n1040,
    n391
  );


  xor
  g1340
  (
    n1311,
    n506,
    n630,
    n932,
    n1092
  );


  nand
  g1341
  (
    n1372,
    n1091,
    n623,
    n880,
    n537
  );


  xor
  g1342
  (
    n1408,
    n517,
    n738,
    n393,
    n949
  );


  and
  g1343
  (
    n1190,
    n938,
    n429,
    n626,
    n428
  );


  nand
  g1344
  (
    n1251,
    n783,
    n737,
    n493,
    n431
  );


  xor
  g1345
  (
    n1233,
    n776,
    n390,
    n405,
    n597
  );


  nand
  g1346
  (
    n1221,
    n804,
    n975,
    n764,
    n1022
  );


  nor
  g1347
  (
    KeyWire_0_19,
    n456,
    n1010,
    n889,
    n671
  );


  xnor
  g1348
  (
    n1396,
    n845,
    n1071,
    n423,
    n895
  );


  and
  g1349
  (
    n1393,
    n407,
    n944,
    n979,
    n762
  );


  xnor
  g1350
  (
    n1400,
    n716,
    n548,
    n1041,
    n959
  );


  or
  g1351
  (
    n1285,
    n433,
    n797,
    n658,
    n977
  );


  nor
  g1352
  (
    n1327,
    n997,
    n608,
    n852,
    n397
  );


  xnor
  g1353
  (
    n1263,
    n508,
    n542,
    n598,
    n1034
  );


  nand
  g1354
  (
    n1246,
    n666,
    n910,
    n424,
    n622
  );


  nor
  g1355
  (
    n1347,
    n675,
    n600,
    n754,
    n1043
  );


  xnor
  g1356
  (
    n1320,
    n687,
    n491,
    n522,
    n905
  );


  nand
  g1357
  (
    n1315,
    n445,
    n503,
    n927,
    n1023
  );


  and
  g1358
  (
    n1286,
    n722,
    n1095,
    n934,
    n452
  );


  nor
  g1359
  (
    n1204,
    n940,
    n970,
    n807,
    n427
  );


  xor
  g1360
  (
    n1235,
    n1018,
    n403,
    n812,
    n434
  );


  and
  g1361
  (
    n1374,
    n1081,
    n434,
    n414,
    n586
  );


  or
  g1362
  (
    n1252,
    n415,
    n1027,
    n693,
    n965
  );


  nand
  g1363
  (
    n1387,
    n973,
    n704,
    n978,
    n705
  );


  nand
  g1364
  (
    n1336,
    n892,
    n765,
    n436,
    n763
  );


  nor
  g1365
  (
    n1391,
    n913,
    n398,
    n634,
    n660
  );


  or
  g1366
  (
    n1269,
    n924,
    n802,
    n398,
    n582
  );


  xnor
  g1367
  (
    n1242,
    n1096,
    n699,
    n907,
    n410
  );


  and
  g1368
  (
    n1202,
    n627,
    n417,
    n393,
    n435
  );


  xor
  g1369
  (
    n1296,
    n414,
    n832,
    n430,
    n1049
  );


  nor
  g1370
  (
    n1392,
    n402,
    n728,
    n656,
    n1032
  );


  and
  g1371
  (
    n1224,
    n992,
    n672,
    n423,
    n751
  );


  xnor
  g1372
  (
    n1341,
    n1087,
    n388,
    n422,
    n641
  );


  xnor
  g1373
  (
    n1388,
    n982,
    n629,
    n724,
    n461
  );


  nor
  g1374
  (
    n1225,
    n1091,
    n643,
    n543,
    n981
  );


  xor
  g1375
  (
    n1357,
    n389,
    n875,
    n432,
    n403
  );


  xnor
  g1376
  (
    n1306,
    n478,
    n662,
    n1029,
    n488
  );


  nand
  g1377
  (
    n1199,
    n696,
    n851,
    n407,
    n402
  );


  or
  g1378
  (
    n1238,
    n442,
    n424,
    n615,
    n421
  );


  xnor
  g1379
  (
    n1353,
    n402,
    n1095,
    n839,
    n793
  );


  or
  g1380
  (
    n1344,
    n896,
    n414,
    n1053,
    n916
  );


  and
  g1381
  (
    n1239,
    n1092,
    n943,
    n400,
    n427
  );


  or
  g1382
  (
    n1333,
    n535,
    n501,
    n416,
    n387
  );


  and
  g1383
  (
    KeyWire_0_15,
    n611,
    n1093,
    n473,
    n877
  );


  xor
  g1384
  (
    n1282,
    n963,
    n410,
    n596,
    n651
  );


  xor
  g1385
  (
    n1307,
    n954,
    n1079,
    n1097,
    n702
  );


  nor
  g1386
  (
    n1250,
    n885,
    n432,
    n504,
    n405
  );


  and
  g1387
  (
    n1394,
    n712,
    n843,
    n411,
    n507
  );


  buf
  g1388
  (
    n1424,
    n1191
  );


  buf
  g1389
  (
    n1414,
    n1195
  );


  not
  g1390
  (
    n1419,
    n1204
  );


  not
  g1391
  (
    n1413,
    n1198
  );


  buf
  g1392
  (
    n1423,
    n1187
  );


  buf
  g1393
  (
    n1418,
    n1205
  );


  not
  g1394
  (
    n1412,
    n1192
  );


  buf
  g1395
  (
    n1411,
    n1193
  );


  buf
  g1396
  (
    n1422,
    n1189
  );


  not
  g1397
  (
    n1420,
    n1202
  );


  not
  g1398
  (
    n1416,
    n1200
  );


  not
  g1399
  (
    n1421,
    n1194
  );


  buf
  g1400
  (
    n1415,
    n1203
  );


  or
  g1401
  (
    n1410,
    n1190,
    n1196,
    n1186
  );


  xor
  g1402
  (
    n1417,
    n1197,
    n1201,
    n1199,
    n1188
  );


  not
  g1403
  (
    n1432,
    n1218
  );


  buf
  g1404
  (
    n1431,
    n1214
  );


  buf
  g1405
  (
    n1429,
    n1415
  );


  not
  g1406
  (
    n1433,
    n1212
  );


  and
  g1407
  (
    n1428,
    n1414,
    n1207
  );


  or
  g1408
  (
    n1425,
    n1411,
    n1206,
    n1213,
    n1410
  );


  xnor
  g1409
  (
    n1430,
    n1217,
    n1211,
    n1216,
    n1417
  );


  or
  g1410
  (
    n1426,
    n1210,
    n1215,
    n1412,
    n1208
  );


  nand
  g1411
  (
    n1427,
    n1417,
    n1209,
    n1413,
    n1416
  );


  or
  g1412
  (
    n1443,
    n1099,
    n1101,
    n1104,
    n1102
  );


  nor
  g1413
  (
    n1439,
    n1106,
    n1103,
    n1425,
    n1102
  );


  or
  g1414
  (
    n1441,
    n1100,
    n1103,
    n1433
  );


  nor
  g1415
  (
    n1440,
    n1099,
    n1433,
    n1101,
    n1105
  );


  nor
  g1416
  (
    n1434,
    n1429,
    n1104,
    n1431,
    n1428
  );


  or
  g1417
  (
    n1437,
    n1105,
    n1099,
    n1100
  );


  xnor
  g1418
  (
    n1442,
    n1100,
    n1102,
    n1101
  );


  and
  g1419
  (
    n1438,
    n1105,
    n1104,
    n1432,
    n1106
  );


  nor
  g1420
  (
    n1436,
    n1430,
    n1426,
    n1101,
    n1427
  );


  xnor
  g1421
  (
    n1435,
    n1104,
    n1105,
    n1099,
    n1103
  );


  nand
  g1422
  (
    n1472,
    n1320,
    n1306,
    n1442,
    n1228
  );


  or
  g1423
  (
    n1483,
    n1443,
    n1332,
    n1326,
    n1248
  );


  nand
  g1424
  (
    n1457,
    n1303,
    n1438,
    n1254,
    n1436
  );


  xor
  g1425
  (
    n1448,
    n1220,
    n1440,
    n1315,
    n1236
  );


  and
  g1426
  (
    n1458,
    n1286,
    n1258,
    n1443,
    n1271
  );


  nand
  g1427
  (
    n1445,
    n1233,
    n1261,
    n1440,
    n1443
  );


  and
  g1428
  (
    n1453,
    n1439,
    n1243,
    n1279,
    n1316
  );


  or
  g1429
  (
    KeyWire_0_20,
    n1307,
    n1330,
    n1298,
    n1440
  );


  xor
  g1430
  (
    n1452,
    n1317,
    n1305,
    n1308,
    n1256
  );


  or
  g1431
  (
    n1460,
    n1269,
    n1321,
    n1250,
    n1314
  );


  xor
  g1432
  (
    n1450,
    n1294,
    n1439,
    n1438,
    n1435
  );


  nand
  g1433
  (
    n1454,
    n1436,
    n1238,
    n1325,
    n1295
  );


  xnor
  g1434
  (
    n1446,
    n1259,
    n1255,
    n1270,
    n1252
  );


  and
  g1435
  (
    n1463,
    n1290,
    n1323,
    n1226,
    n1328
  );


  xnor
  g1436
  (
    n1469,
    n1297,
    n1435,
    n1240,
    n1231
  );


  nor
  g1437
  (
    n1476,
    n1440,
    n1434,
    n1437,
    n1329
  );


  or
  g1438
  (
    n1464,
    n1230,
    n1227,
    n1237,
    n1241
  );


  xor
  g1439
  (
    n1456,
    n1439,
    n1235,
    n1224,
    n1246
  );


  or
  g1440
  (
    n1468,
    n1229,
    n1437,
    n1434,
    n1242
  );


  xor
  g1441
  (
    n1467,
    n1437,
    n1322,
    n1222,
    n1338
  );


  or
  g1442
  (
    n1462,
    n1337,
    n1301,
    n1435,
    n1223
  );


  xor
  g1443
  (
    n1449,
    n1312,
    n1327,
    n1249,
    n1266
  );


  or
  g1444
  (
    n1461,
    n1436,
    n1309,
    n1442,
    n1273
  );


  and
  g1445
  (
    n1465,
    n1302,
    n1253,
    n1280,
    n1439
  );


  and
  g1446
  (
    n1455,
    n1287,
    n1313,
    n1277,
    n1257
  );


  and
  g1447
  (
    n1481,
    n1438,
    n1251,
    n1324,
    n1267
  );


  or
  g1448
  (
    n1444,
    n1239,
    n1288,
    n1234,
    n1289
  );


  nand
  g1449
  (
    n1447,
    n1225,
    n1434,
    n1300,
    n1438
  );


  nor
  g1450
  (
    n1459,
    n1293,
    n1291,
    n1310,
    n1221
  );


  nor
  g1451
  (
    n1471,
    n1442,
    n1304,
    n1443,
    n1334
  );


  or
  g1452
  (
    n1478,
    n1282,
    n1441,
    n1331
  );


  or
  g1453
  (
    n1470,
    n1296,
    n1247,
    n1319,
    n1299
  );


  and
  g1454
  (
    n1451,
    n1292,
    n1285,
    n1437,
    n1272
  );


  nor
  g1455
  (
    n1479,
    n1268,
    n1219,
    n1275,
    n1274
  );


  nand
  g1456
  (
    n1474,
    n1336,
    n1441,
    n1283,
    n1278
  );


  nor
  g1457
  (
    n1482,
    n1264,
    n1434,
    n1281,
    n1265
  );


  nor
  g1458
  (
    n1475,
    n1436,
    n1442,
    n1244,
    n1245
  );


  xnor
  g1459
  (
    n1480,
    n1311,
    n1262,
    n1263,
    n1232
  );


  or
  g1460
  (
    n1477,
    n1441,
    n1260,
    n1284,
    n1333
  );


  or
  g1461
  (
    n1473,
    n1318,
    n1435,
    n1276,
    n1335
  );


  buf
  g1462
  (
    n1495,
    n1450
  );


  buf
  g1463
  (
    n1505,
    n1347
  );


  not
  g1464
  (
    n1497,
    n1350
  );


  buf
  g1465
  (
    n1494,
    n1450
  );


  buf
  g1466
  (
    n1492,
    n1419
  );


  not
  g1467
  (
    n1496,
    n1452
  );


  buf
  g1468
  (
    n1484,
    n1351
  );


  buf
  g1469
  (
    n1488,
    n1419
  );


  and
  g1470
  (
    n1502,
    n1445,
    n1446
  );


  or
  g1471
  (
    n1487,
    n1358,
    n1339
  );


  nand
  g1472
  (
    n1489,
    n1454,
    n1355,
    n1359,
    n1450
  );


  and
  g1473
  (
    n1498,
    n1364,
    n1453,
    n1361,
    n1365
  );


  nor
  g1474
  (
    n1499,
    n1453,
    n1352,
    n1419,
    n1340
  );


  and
  g1475
  (
    n1506,
    n1421,
    n1422,
    n1454,
    n1341
  );


  or
  g1476
  (
    n1491,
    n1348,
    n1454,
    n1357,
    n1353
  );


  xnor
  g1477
  (
    n1490,
    n1356,
    n1363,
    n1421,
    n1452
  );


  xnor
  g1478
  (
    n1503,
    n1447,
    n1342,
    n1422,
    n1453
  );


  or
  g1479
  (
    n1501,
    n1420,
    n1453,
    n1421,
    n1419
  );


  xnor
  g1480
  (
    n1500,
    n1420,
    n1360,
    n1354,
    n1366
  );


  or
  g1481
  (
    n1508,
    n1418,
    n1368,
    n1451,
    n1444
  );


  nor
  g1482
  (
    n1493,
    n1449,
    n1362,
    n1420,
    n1367
  );


  nand
  g1483
  (
    n1504,
    n1343,
    n1346,
    n1452,
    n1450
  );


  nand
  g1484
  (
    n1507,
    n1349,
    n1451,
    n1345
  );


  nand
  g1485
  (
    n1486,
    n1448,
    n1452,
    n1344,
    n1451
  );


  nor
  g1486
  (
    n1485,
    n1420,
    n1418,
    n1369,
    n1421
  );


  nor
  g1487
  (
    n1535,
    n1474,
    n1467,
    n1473,
    n1462
  );


  nand
  g1488
  (
    n1534,
    n1472,
    n1474,
    n1459,
    n1456
  );


  xnor
  g1489
  (
    n1526,
    n1489,
    n1476,
    n1461,
    n1484
  );


  nor
  g1490
  (
    n1515,
    n1484,
    n1465,
    n1487,
    n1471
  );


  and
  g1491
  (
    n1539,
    n1490,
    n1479,
    n1489,
    n1486
  );


  xor
  g1492
  (
    n1521,
    n1456,
    n1459,
    n1469,
    n1473
  );


  nor
  g1493
  (
    n1538,
    n1485,
    n1486,
    n1466,
    n1464
  );


  and
  g1494
  (
    n1510,
    n1490,
    n1478,
    n1463,
    n1477
  );


  and
  g1495
  (
    n1511,
    n1486,
    n1459,
    n1475,
    n1458
  );


  xnor
  g1496
  (
    n1516,
    n1468,
    n1462,
    n1472,
    n1487
  );


  nand
  g1497
  (
    n1517,
    n1463,
    n1464,
    n1491
  );


  xor
  g1498
  (
    n1528,
    n1458,
    n1463,
    n1460,
    n1461
  );


  or
  g1499
  (
    n1520,
    n1488,
    n1464,
    n1455,
    n1475
  );


  or
  g1500
  (
    n1530,
    n1477,
    n1485,
    n1488,
    n1478
  );


  nand
  g1501
  (
    n1514,
    n1469,
    n1468,
    n1458,
    n1477
  );


  nor
  g1502
  (
    n1532,
    n1456,
    n1461,
    n1472
  );


  nand
  g1503
  (
    n1529,
    n1460,
    n1455,
    n1471,
    n1474
  );


  xor
  g1504
  (
    n1512,
    n1468,
    n1479,
    n1490,
    n1484
  );


  nor
  g1505
  (
    n1524,
    n1478,
    n1492,
    n1464,
    n1488
  );


  xnor
  g1506
  (
    n1527,
    n1462,
    n1475,
    n1489
  );


  nor
  g1507
  (
    n1509,
    n1460,
    n1487,
    n1469,
    n1465
  );


  nor
  g1508
  (
    n1541,
    n1491,
    n1455,
    n1467,
    n1457
  );


  nand
  g1509
  (
    n1525,
    n1457,
    n1471,
    n1478
  );


  nand
  g1510
  (
    n1513,
    n1467,
    n1454,
    n1485,
    n1487
  );


  nor
  g1511
  (
    n1536,
    n1484,
    n1458,
    n1476,
    n1470
  );


  nor
  g1512
  (
    n1523,
    n1474,
    n1457,
    n1473,
    n1469
  );


  nand
  g1513
  (
    n1522,
    n1465,
    n1463,
    n1462,
    n1461
  );


  nor
  g1514
  (
    n1518,
    n1473,
    n1486,
    n1465,
    n1466
  );


  xnor
  g1515
  (
    n1540,
    n1457,
    n1466,
    n1485,
    n1455
  );


  nor
  g1516
  (
    n1519,
    n1476,
    n1470,
    n1477,
    n1488
  );


  nor
  g1517
  (
    n1531,
    n1470,
    n1475,
    n1491,
    n1490
  );


  and
  g1518
  (
    n1533,
    n1476,
    n1459,
    n1460,
    n1470
  );


  nand
  g1519
  (
    n1537,
    n1456,
    n1467,
    n1468,
    n1466
  );


  buf
  g1520
  (
    n1543,
    n1107
  );


  buf
  g1521
  (
    n1542,
    n1108
  );


  not
  g1522
  (
    n1562,
    n1482
  );


  not
  g1523
  (
    n1549,
    n1494
  );


  not
  g1524
  (
    n1557,
    n1494
  );


  buf
  g1525
  (
    n1550,
    n1520
  );


  xnor
  g1526
  (
    n1544,
    n1378,
    n1495,
    n1110,
    n1107
  );


  nand
  g1527
  (
    n1564,
    n1531,
    n1522,
    n1480,
    n1521
  );


  xor
  g1528
  (
    n1554,
    n1377,
    n1109,
    n1513,
    n1482
  );


  nand
  g1529
  (
    n1545,
    n1480,
    n1374,
    n1106,
    n1108
  );


  xnor
  g1530
  (
    n1558,
    n1375,
    n1524,
    n1494,
    n1109
  );


  nand
  g1531
  (
    n1555,
    n1514,
    n1493,
    n1371,
    n1523
  );


  nor
  g1532
  (
    n1561,
    n1370,
    n1516,
    n1532,
    n1108
  );


  and
  g1533
  (
    n1548,
    n1495,
    n1492,
    n1511,
    n1479
  );


  xor
  g1534
  (
    n1559,
    n1493,
    n1519,
    n1108,
    n1481
  );


  xor
  g1535
  (
    n1553,
    n1376,
    n1493,
    n1527,
    n1492
  );


  xnor
  g1536
  (
    n1556,
    n1494,
    n1109,
    n1517,
    n1480
  );


  nor
  g1537
  (
    n1547,
    n1515,
    n1530,
    n1510,
    n1481
  );


  and
  g1538
  (
    n1551,
    n1110,
    n1107,
    n1526
  );


  and
  g1539
  (
    n1563,
    n1481,
    n1373,
    n1512,
    n1493
  );


  or
  g1540
  (
    n1546,
    n1372,
    n1492,
    n1529,
    n1528
  );


  and
  g1541
  (
    n1552,
    n1518,
    n1481,
    n1525,
    n1479
  );


  nor
  g1542
  (
    n1560,
    n1106,
    n1109,
    n1480,
    n1482
  );


  not
  g1543
  (
    n1571,
    n1556
  );


  not
  g1544
  (
    n1569,
    n1560
  );


  not
  g1545
  (
    n1566,
    n1483
  );


  buf
  g1546
  (
    n1570,
    n1482
  );


  buf
  g1547
  (
    n1568,
    n1483
  );


  or
  g1548
  (
    n1567,
    n1557,
    n1483,
    n1554
  );


  and
  g1549
  (
    n1565,
    n1483,
    n1559,
    n1555,
    n1558
  );


  xnor
  g1550
  (
    n1573,
    n1567,
    n1571,
    n1570,
    n1569
  );


  xnor
  g1551
  (
    n1572,
    n1508,
    n1496,
    n1502,
    n1506
  );


  xnor
  g1552
  (
    n1595,
    n1567,
    n1499,
    n1386,
    n1569
  );


  nor
  g1553
  (
    n1574,
    n1500,
    n1498,
    n1504,
    n1570
  );


  and
  g1554
  (
    n1589,
    n1502,
    n1500,
    n1566,
    n1506
  );


  nor
  g1555
  (
    n1587,
    n1498,
    n1499,
    n1561,
    n1568
  );


  xor
  g1556
  (
    n1594,
    n1381,
    n1396,
    n1504,
    n1507
  );


  and
  g1557
  (
    n1576,
    n1394,
    n1571,
    n1495,
    n1563
  );


  and
  g1558
  (
    n1591,
    n1505,
    n1569,
    n1570,
    n1568
  );


  nor
  g1559
  (
    n1585,
    n1395,
    n1497,
    n1496,
    n1502
  );


  nor
  g1560
  (
    n1582,
    n1507,
    n1380,
    n1500,
    n1499
  );


  xor
  g1561
  (
    n1580,
    n1389,
    n1503,
    n1567,
    n1566
  );


  xor
  g1562
  (
    n1590,
    n1390,
    n1570,
    n1571,
    n1505
  );


  and
  g1563
  (
    n1588,
    n1564,
    n1497,
    n1498,
    n1495
  );


  nand
  g1564
  (
    n1583,
    n1562,
    n1566,
    n1379,
    n1503
  );


  and
  g1565
  (
    n1596,
    n1397,
    n1569,
    n1571,
    n1392
  );


  nor
  g1566
  (
    n1578,
    n1501,
    n1508,
    n1393
  );


  nand
  g1567
  (
    n1592,
    n1506,
    n1505,
    n1565,
    n1503
  );


  xor
  g1568
  (
    n1581,
    n1383,
    n1387,
    n1507,
    n1502
  );


  xnor
  g1569
  (
    n1593,
    n1504,
    n1499,
    n1565,
    n1382
  );


  xor
  g1570
  (
    n1597,
    n1385,
    n1388,
    n1501,
    n1505
  );


  or
  g1571
  (
    n1577,
    n1503,
    n1568,
    n1508,
    n1501
  );


  xnor
  g1572
  (
    n1575,
    n1507,
    n1497,
    n1384
  );


  or
  g1573
  (
    n1584,
    n1566,
    n1501,
    n1391,
    n1506
  );


  nor
  g1574
  (
    n1586,
    n1568,
    n1398,
    n1504,
    n1496
  );


  xor
  g1575
  (
    n1579,
    n1567,
    n1496,
    n1498,
    n1500
  );


  nand
  g1576
  (
    n1647,
    n1176,
    n1121,
    n1170,
    n1135
  );


  nor
  g1577
  (
    n1652,
    n1119,
    n1541,
    n1597,
    n1591
  );


  or
  g1578
  (
    n1624,
    n1133,
    n1593,
    n1580,
    n1594
  );


  and
  g1579
  (
    n1608,
    n1167,
    n1161,
    n1574,
    n1165
  );


  and
  g1580
  (
    n1694,
    n1585,
    n1118,
    n1588,
    n1576
  );


  nand
  g1581
  (
    n1629,
    n1586,
    n1592,
    n1176,
    n1164
  );


  and
  g1582
  (
    n1659,
    n1150,
    n1588,
    n1117,
    n1169
  );


  and
  g1583
  (
    n1661,
    n1580,
    n1184,
    n1579,
    n1593
  );


  xor
  g1584
  (
    n1695,
    n1153,
    n1145,
    n1594,
    n1154
  );


  and
  g1585
  (
    n1670,
    n1581,
    n1169,
    n1138,
    n1177
  );


  xnor
  g1586
  (
    n1658,
    n1589,
    n1183,
    n1157,
    n1572
  );


  nor
  g1587
  (
    n1649,
    n1156,
    n1152,
    n1179,
    n1537
  );


  xnor
  g1588
  (
    n1654,
    n1538,
    n1168,
    n1172,
    n1121
  );


  nand
  g1589
  (
    n1602,
    n1167,
    n1577,
    n1182,
    n1179
  );


  nand
  g1590
  (
    n1611,
    n1120,
    n1112,
    n1184
  );


  and
  g1591
  (
    n1692,
    n1127,
    n1535,
    n1130,
    n1128
  );


  and
  g1592
  (
    n1603,
    n1140,
    n1139,
    n1144,
    n1154
  );


  xor
  g1593
  (
    n1599,
    n1130,
    n1150,
    n1125,
    n1591
  );


  and
  g1594
  (
    n1648,
    n1180,
    n1124,
    n1174,
    n1132
  );


  nor
  g1595
  (
    n1623,
    n1116,
    n1165,
    n1173,
    n1140
  );


  xnor
  g1596
  (
    n1617,
    n1588,
    n1172,
    n1585,
    n1160
  );


  nor
  g1597
  (
    n1598,
    n1156,
    n1144,
    n1178,
    n1576
  );


  nor
  g1598
  (
    n1625,
    n1575,
    n1127,
    n1175,
    n1170
  );


  xor
  g1599
  (
    n1668,
    n1584,
    n1169,
    n1574,
    n1161
  );


  or
  g1600
  (
    n1635,
    n1140,
    n1112,
    n1180,
    n1157
  );


  xnor
  g1601
  (
    n1605,
    n1580,
    n1584,
    n1124,
    n1123
  );


  or
  g1602
  (
    n1637,
    n1144,
    n1593,
    n1132,
    n1182
  );


  nor
  g1603
  (
    n1679,
    n1117,
    n440,
    n1153,
    n1110
  );


  xnor
  g1604
  (
    n1685,
    n1158,
    n1155,
    n1597,
    n1582
  );


  nand
  g1605
  (
    n1696,
    n1573,
    n1167,
    n1158,
    n1168
  );


  nor
  g1606
  (
    n1687,
    n1143,
    n1119,
    n1579,
    n1175
  );


  nand
  g1607
  (
    n1631,
    n1539,
    n1126,
    n1592,
    n1164
  );


  and
  g1608
  (
    n1664,
    n1181,
    n1593,
    n1131,
    n1148
  );


  xor
  g1609
  (
    n1639,
    n1540,
    n1576,
    n1121,
    n1594
  );


  xnor
  g1610
  (
    n1622,
    n1174,
    n1148,
    n1164,
    n1151
  );


  nand
  g1611
  (
    n1657,
    n1146,
    n1162,
    n1118,
    n1172
  );


  or
  g1612
  (
    n1690,
    n1583,
    n1159,
    n1183,
    n1141
  );


  xnor
  g1613
  (
    n1650,
    n1166,
    n1163,
    n1581,
    n1135
  );


  nor
  g1614
  (
    n1600,
    n1125,
    n1156,
    n1577,
    n1138
  );


  nand
  g1615
  (
    n1691,
    n1179,
    n1166,
    n1162,
    n1168
  );


  nand
  g1616
  (
    n1613,
    n1119,
    n1124,
    n1578,
    n1577
  );


  nor
  g1617
  (
    n1698,
    n1150,
    n1122,
    n1151,
    n1153
  );


  nor
  g1618
  (
    n1627,
    n1117,
    n1163,
    n1148,
    n1173
  );


  xnor
  g1619
  (
    n1686,
    n1157,
    n1131,
    n1143,
    n1129
  );


  nor
  g1620
  (
    n1630,
    n1148,
    n1137,
    n1136,
    n1163
  );


  nand
  g1621
  (
    n1675,
    n1580,
    n1133,
    n1163,
    n1126
  );


  nor
  g1622
  (
    n1628,
    n1581,
    n1577,
    n1126,
    n1113
  );


  and
  g1623
  (
    n1666,
    n1118,
    n1178,
    n1127,
    n1154
  );


  and
  g1624
  (
    n1607,
    n1578,
    n440,
    n1132,
    n1176
  );


  xnor
  g1625
  (
    n1669,
    n1144,
    n1152,
    n1587,
    n1575
  );


  xnor
  g1626
  (
    n1663,
    n1136,
    n1167,
    n1578,
    n1114
  );


  nand
  g1627
  (
    n1681,
    n1171,
    n1142,
    n1124,
    n1152
  );


  and
  g1628
  (
    n1674,
    n1117,
    n1177,
    n1584,
    n1119
  );


  nor
  g1629
  (
    n1609,
    n1156,
    n1175,
    n1130,
    n1111
  );


  xor
  g1630
  (
    n1653,
    n1114,
    n1154,
    n1592,
    n1152
  );


  or
  g1631
  (
    n1644,
    n1185,
    n1181,
    n1590,
    n1139
  );


  xor
  g1632
  (
    n1688,
    n1184,
    n1149,
    n1123,
    n1583
  );


  and
  g1633
  (
    n1615,
    n1122,
    n1181,
    n1146,
    n1134
  );


  nand
  g1634
  (
    n1667,
    n1121,
    n1138,
    n1184,
    n1155
  );


  xnor
  g1635
  (
    n1683,
    n1161,
    n1115,
    n1575,
    n1590
  );


  or
  g1636
  (
    n1636,
    n1595,
    n1125,
    n1142,
    n1164
  );


  xnor
  g1637
  (
    n1651,
    n1120,
    n1134,
    n1182,
    n1172
  );


  or
  g1638
  (
    n1643,
    n1536,
    n1111,
    n1178,
    n1143
  );


  or
  g1639
  (
    n1665,
    n1183,
    n1113,
    n1125,
    n1595
  );


  xor
  g1640
  (
    n1660,
    n1572,
    n1585,
    n1159,
    n1128
  );


  nand
  g1641
  (
    n1677,
    n1146,
    n1134,
    n1149,
    n1123
  );


  or
  g1642
  (
    n1678,
    n1131,
    n1171,
    n1582,
    n1138
  );


  xnor
  g1643
  (
    n1640,
    n1145,
    n1116,
    n1136
  );


  xnor
  g1644
  (
    n1645,
    n1183,
    n1147,
    n1173,
    n1111
  );


  or
  g1645
  (
    n1693,
    n1140,
    n1129,
    n1590,
    n1596
  );


  nand
  g1646
  (
    n1699,
    n1151,
    n1139,
    n1594,
    n1135
  );


  and
  g1647
  (
    n1618,
    n1122,
    n1177,
    n1171,
    n1113
  );


  nor
  g1648
  (
    n1633,
    n1137,
    n1141,
    n1133,
    n1166
  );


  and
  g1649
  (
    n1610,
    n1166,
    n1578,
    n1584,
    n1173
  );


  and
  g1650
  (
    n1616,
    n1574,
    n1586,
    n1589
  );


  nor
  g1651
  (
    n1689,
    n1115,
    n1134,
    n1534,
    n1177
  );


  xnor
  g1652
  (
    n1626,
    n1159,
    n1591,
    n1137,
    n1573
  );


  nand
  g1653
  (
    n1621,
    n1162,
    n1123,
    n1115,
    n1174
  );


  nand
  g1654
  (
    n1684,
    n1158,
    n1158,
    n1159,
    n1114
  );


  nand
  g1655
  (
    n1606,
    n1129,
    n1160,
    n1533,
    n1592
  );


  or
  g1656
  (
    n1614,
    n1155,
    n1174,
    n1131,
    n1596
  );


  or
  g1657
  (
    n1672,
    n1590,
    n1168,
    n1595,
    n1576
  );


  xnor
  g1658
  (
    n1673,
    n1582,
    n1160,
    n1596,
    n1170
  );


  or
  g1659
  (
    n1612,
    n1575,
    n1157,
    n1585,
    n1147
  );


  and
  g1660
  (
    n1619,
    n1128,
    n1583,
    n1579,
    n1147
  );


  nand
  g1661
  (
    n1656,
    n1149,
    n1135,
    n1120,
    n1155
  );


  and
  g1662
  (
    n1701,
    n1120,
    n1149,
    n1153,
    n1113
  );


  or
  g1663
  (
    n1620,
    n1129,
    n1182,
    n1581,
    n1130
  );


  nor
  g1664
  (
    n1634,
    n1141,
    n1180,
    n1165,
    n1145
  );


  xor
  g1665
  (
    n1662,
    n1147,
    n1118,
    n1591,
    n1572
  );


  nor
  g1666
  (
    n1646,
    n1573,
    n1597,
    n1574,
    n1146
  );


  or
  g1667
  (
    n1682,
    n1185,
    n1110,
    n1111,
    n1171
  );


  xor
  g1668
  (
    n1632,
    n1126,
    n1181,
    n1136,
    n1133
  );


  and
  g1669
  (
    n1700,
    n1115,
    n1587,
    n1589,
    n1114
  );


  or
  g1670
  (
    n1601,
    n1165,
    n1145,
    n1142,
    n1143
  );


  xnor
  g1671
  (
    n1655,
    n1179,
    n1572,
    n1150,
    n1586
  );


  nand
  g1672
  (
    n1604,
    n1582,
    n1587,
    n1178,
    n1596
  );


  nor
  g1673
  (
    n1642,
    n1127,
    n1597,
    n1587,
    n1162
  );


  and
  g1674
  (
    n1676,
    n1586,
    n1139,
    n1176,
    n1141
  );


  xor
  g1675
  (
    n1680,
    n1579,
    n1583,
    n1122,
    n1161
  );


  nor
  g1676
  (
    n1671,
    n1595,
    n1128,
    n1132,
    n1160
  );


  or
  g1677
  (
    n1638,
    n1588,
    n1185,
    n1116,
    n1112
  );


  or
  g1678
  (
    n1641,
    n1573,
    n1175,
    n1170,
    n1137
  );


  xnor
  g1679
  (
    n1697,
    n1142,
    n1169,
    n1151,
    n1180
  );


  not
  g1680
  (
    n1706,
    n1611
  );


  buf
  g1681
  (
    n1702,
    n1600
  );


  buf
  g1682
  (
    n1719,
    n1604
  );


  not
  g1683
  (
    n1705,
    n1608
  );


  buf
  g1684
  (
    n1707,
    n1612
  );


  buf
  g1685
  (
    n1703,
    n1606
  );


  not
  g1686
  (
    n1717,
    n1609
  );


  not
  g1687
  (
    n1713,
    n1598
  );


  not
  g1688
  (
    n1716,
    n1603
  );


  not
  g1689
  (
    n1704,
    n1615
  );


  buf
  g1690
  (
    n1712,
    n1602
  );


  buf
  g1691
  (
    n1714,
    n1607
  );


  not
  g1692
  (
    n1718,
    n1601
  );


  not
  g1693
  (
    n1708,
    n1614
  );


  buf
  g1694
  (
    n1709,
    n1613
  );


  buf
  g1695
  (
    n1710,
    n1599
  );


  buf
  g1696
  (
    n1711,
    n1610
  );


  buf
  g1697
  (
    n1715,
    n1605
  );


  xor
  g1698
  (
    n1738,
    n1642,
    n1653,
    n1713,
    n1647
  );


  xnor
  g1699
  (
    n1749,
    n1621,
    n1710,
    n1652,
    n1631
  );


  nand
  g1700
  (
    n1785,
    n1626,
    n1656,
    n1644,
    n1719
  );


  nand
  g1701
  (
    n1776,
    n1711,
    n1669,
    n1653,
    n1646
  );


  xnor
  g1702
  (
    n1744,
    n1671,
    n1649,
    n1639,
    n1642
  );


  nor
  g1703
  (
    n1758,
    n1670,
    n1645,
    n1637,
    n1659
  );


  nor
  g1704
  (
    n1737,
    n1638,
    n1660,
    n1636,
    n1710
  );


  nor
  g1705
  (
    n1781,
    n1668,
    n1623,
    n1713,
    n1656
  );


  and
  g1706
  (
    n1740,
    n1643,
    n1656,
    n1621,
    n1666
  );


  xor
  g1707
  (
    n1787,
    n1633,
    n1640,
    n1661
  );


  or
  g1708
  (
    n1771,
    n1629,
    n1651,
    n1616,
    n1638
  );


  xor
  g1709
  (
    n1750,
    n1644,
    n1647,
    n1667,
    n1653
  );


  and
  g1710
  (
    n1767,
    n1657,
    n1643,
    n1654,
    n1710
  );


  or
  g1711
  (
    n1784,
    n1718,
    n1637,
    n1632,
    n1716
  );


  nor
  g1712
  (
    n1726,
    n1652,
    n1662,
    n1650,
    n1717
  );


  nand
  g1713
  (
    n1772,
    n1715,
    n1642,
    n1664,
    n1703
  );


  xnor
  g1714
  (
    KeyWire_0_24,
    n1718,
    n1672,
    n1709,
    n1651
  );


  and
  g1715
  (
    n1735,
    n1707,
    n1657,
    n1624,
    n1643
  );


  nand
  g1716
  (
    n1762,
    n1704,
    n1673,
    n1666,
    n1703
  );


  nand
  g1717
  (
    n1760,
    n1632,
    n1627,
    n1626,
    n1652
  );


  and
  g1718
  (
    n1761,
    n1648,
    n1712,
    n1635
  );


  xnor
  g1719
  (
    n1745,
    n1626,
    n1623,
    n1705,
    n1631
  );


  or
  g1720
  (
    n1747,
    n1649,
    n1672,
    n1652,
    n1634
  );


  nor
  g1721
  (
    n1770,
    n1655,
    n1635,
    n1639,
    n1629
  );


  nor
  g1722
  (
    n1754,
    n1648,
    n1640,
    n1620,
    n1717
  );


  or
  g1723
  (
    n1777,
    n1665,
    n1648,
    n1627,
    n1622
  );


  or
  g1724
  (
    n1786,
    n1708,
    n1708,
    n1634,
    n1705
  );


  xnor
  g1725
  (
    n1734,
    n1657,
    n1717,
    n1715,
    n1671
  );


  or
  g1726
  (
    n1743,
    n1632,
    n1658,
    n1648,
    n1636
  );


  nand
  g1727
  (
    n1728,
    n1642,
    n1662,
    n1635,
    n1668
  );


  nand
  g1728
  (
    n1779,
    n1630,
    n1624,
    n1670,
    n1638
  );


  nand
  g1729
  (
    n1736,
    n1634,
    n1707,
    n1626,
    n1668
  );


  xnor
  g1730
  (
    n1722,
    n1655,
    n1655,
    n1625,
    n1649
  );


  nor
  g1731
  (
    n1766,
    n1702,
    n1620,
    n1628,
    n1719
  );


  xnor
  g1732
  (
    n1765,
    n1650,
    n1708,
    n1631,
    n1663
  );


  and
  g1733
  (
    n1723,
    n1711,
    n1645,
    n1660,
    n1709
  );


  nand
  g1734
  (
    n1759,
    n1667,
    n1639,
    n1660,
    n1705
  );


  nand
  g1735
  (
    n1783,
    n1627,
    n1659,
    n1651,
    n1641
  );


  xnor
  g1736
  (
    n1763,
    n1714,
    n1672,
    n1665,
    n1647
  );


  nand
  g1737
  (
    n1741,
    n1673,
    n1624,
    n1704
  );


  or
  g1738
  (
    n1746,
    n1633,
    n1719,
    n1711,
    n1630
  );


  nand
  g1739
  (
    n1757,
    n1702,
    n1715,
    n1651,
    n1646
  );


  or
  g1740
  (
    n1788,
    n1637,
    n1713,
    n1716,
    n1668
  );


  nor
  g1741
  (
    n1721,
    n1630,
    n1716,
    n1646,
    n1623
  );


  nor
  g1742
  (
    n1751,
    n1624,
    n1656,
    n1646,
    n1622
  );


  nand
  g1743
  (
    n1768,
    n1640,
    n1670,
    n1713,
    n1665
  );


  nor
  g1744
  (
    n1756,
    n1629,
    n1663,
    n1669,
    n1622
  );


  nor
  g1745
  (
    n1720,
    n1709,
    n1706,
    n1660,
    n1659
  );


  nor
  g1746
  (
    n1778,
    n1719,
    n1641,
    n1630,
    n1658
  );


  or
  g1747
  (
    KeyWire_0_31,
    n1634,
    n1706,
    n1710,
    n1654
  );


  or
  g1748
  (
    n1742,
    n1640,
    n1669,
    n1703,
    n1661
  );


  nand
  g1749
  (
    n1780,
    n1659,
    n1662,
    n1666,
    n1703
  );


  and
  g1750
  (
    n1790,
    n1669,
    n1705,
    n1670,
    n1625
  );


  xor
  g1751
  (
    n1773,
    n1633,
    n1628,
    n1623,
    n1711
  );


  xnor
  g1752
  (
    n1748,
    n1714,
    n1658,
    n1715,
    n1621
  );


  or
  g1753
  (
    n1739,
    n1636,
    n1717,
    n1625,
    n1657
  );


  xnor
  g1754
  (
    n1755,
    n1672,
    n1637,
    n1664,
    n1632
  );


  xnor
  g1755
  (
    n1782,
    n1628,
    n1639,
    n1661,
    n1654
  );


  nor
  g1756
  (
    n1775,
    n1628,
    n1625,
    n1641,
    n1636
  );


  or
  g1757
  (
    n1753,
    n1631,
    n1635,
    n1618,
    n1702
  );


  or
  g1758
  (
    n1724,
    n1718,
    n1650,
    n1714,
    n1638
  );


  or
  g1759
  (
    KeyWire_0_27,
    n1650,
    n1663,
    n1716,
    n1621
  );


  and
  g1760
  (
    n1733,
    n1707,
    n1712,
    n1718,
    n1644
  );


  and
  g1761
  (
    n1789,
    n1629,
    n1617,
    n1666,
    n1671
  );


  and
  g1762
  (
    n1752,
    n1627,
    n1645,
    n1662,
    n1653
  );


  xnor
  g1763
  (
    n1769,
    n1665,
    n1647,
    n1619,
    n1714
  );


  or
  g1764
  (
    n1730,
    n1654,
    n1649,
    n1633,
    n1658
  );


  nor
  g1765
  (
    n1774,
    n1667,
    n1712,
    n1664,
    n1622
  );


  or
  g1766
  (
    n1764,
    n1704,
    n1643,
    n1644,
    n1671
  );


  nor
  g1767
  (
    n1729,
    n1708,
    n1709,
    n1645,
    n1655
  );


  xnor
  g1768
  (
    n1727,
    n1664,
    n1667,
    n1663,
    n1641
  );


  nand
  g1769
  (
    n1791,
    n1707,
    n1706,
    n1702
  );


  not
  g1770
  (
    n1792,
    n1724
  );


  not
  g1771
  (
    n1793,
    n1404
  );


  xnor
  g1772
  (
    n1796,
    n1722,
    n1402,
    n1400,
    n1405
  );


  xor
  g1773
  (
    n1794,
    n1407,
    n1723,
    n1399,
    n1403
  );


  or
  g1774
  (
    n1795,
    n1720,
    n1401,
    n1406,
    n1721
  );


  not
  g1775
  (
    n1806,
    n1794
  );


  buf
  g1776
  (
    n1799,
    n1793
  );


  buf
  g1777
  (
    n1801,
    n1793
  );


  buf
  g1778
  (
    n1800,
    n1792
  );


  not
  g1779
  (
    n1804,
    n1793
  );


  not
  g1780
  (
    n1797,
    n1792
  );


  not
  g1781
  (
    n1802,
    n1792
  );


  not
  g1782
  (
    n1803,
    n1792
  );


  not
  g1783
  (
    n1805,
    n1793
  );


  not
  g1784
  (
    n1798,
    n1794
  );


  xnor
  g1785
  (
    n1816,
    n1679,
    n1687,
    n1798
  );


  xor
  g1786
  (
    n1822,
    n1680,
    n1693,
    n1692,
    n1681
  );


  or
  g1787
  (
    n1821,
    n1678,
    n1423,
    n1677,
    n1797
  );


  nor
  g1788
  (
    n1818,
    n1695,
    n1676,
    n1804,
    n1690
  );


  xor
  g1789
  (
    n1809,
    n1695,
    n1680,
    n1806,
    n1690
  );


  and
  g1790
  (
    n1844,
    n1802,
    n1698,
    n1674,
    n1690
  );


  nor
  g1791
  (
    n1845,
    n1801,
    n1800,
    n1678,
    n1796
  );


  nand
  g1792
  (
    n1831,
    n1422,
    n1806,
    n1688,
    n1796
  );


  or
  g1793
  (
    n1819,
    n1795,
    n1802,
    n1682,
    n1799
  );


  and
  g1794
  (
    n1827,
    n1684,
    n1697,
    n1683,
    n1694
  );


  or
  g1795
  (
    n1838,
    n1686,
    n1687,
    n1684,
    n1802
  );


  and
  g1796
  (
    n1836,
    n1805,
    n1806,
    n1800,
    n1675
  );


  nor
  g1797
  (
    n1835,
    n1677,
    n1681,
    n1423,
    n1679
  );


  xor
  g1798
  (
    n1823,
    n1798,
    n1675,
    n1803,
    n1805
  );


  xnor
  g1799
  (
    n1832,
    n1684,
    n1696,
    n1693,
    n1690
  );


  nor
  g1800
  (
    n1810,
    n1796,
    n1685,
    n1802,
    n1699
  );


  xor
  g1801
  (
    n1807,
    n1683,
    n1698,
    n1689
  );


  and
  g1802
  (
    n1841,
    n1693,
    n1689,
    n1684,
    n1678
  );


  nand
  g1803
  (
    n1817,
    n1683,
    n1799,
    n1685,
    n1699
  );


  and
  g1804
  (
    n1839,
    n1797,
    n1692,
    n1680,
    n1685
  );


  xor
  g1805
  (
    n1837,
    n1801,
    n1798,
    n1696,
    n1800
  );


  xnor
  g1806
  (
    n1829,
    n1677,
    n1676,
    n1683,
    n1682
  );


  or
  g1807
  (
    n1846,
    n1685,
    n1694,
    n1797,
    n1795
  );


  and
  g1808
  (
    n1840,
    n1797,
    n1673,
    n1675,
    n1409
  );


  xnor
  g1809
  (
    n1833,
    n1694,
    n1682,
    n1798,
    n1686
  );


  and
  g1810
  (
    n1815,
    n1686,
    n1682,
    n1674,
    n1676
  );


  or
  g1811
  (
    n1820,
    n1681,
    n1805,
    n1696,
    n1794
  );


  nand
  g1812
  (
    n1808,
    n1803,
    n1794,
    n1689,
    n1799
  );


  xor
  g1813
  (
    n1825,
    n1677,
    n1692,
    n1799,
    n1695
  );


  nand
  g1814
  (
    n1842,
    n1679,
    n1804,
    n1675,
    n1796
  );


  xnor
  g1815
  (
    n1834,
    n1697,
    n1697,
    n1804,
    n1678
  );


  and
  g1816
  (
    n1824,
    n1680,
    n1691,
    n1803,
    n1686
  );


  and
  g1817
  (
    n1843,
    n1691,
    n1795,
    n1674,
    n1803
  );


  nand
  g1818
  (
    n1812,
    n1795,
    n1691,
    n1805,
    n1800
  );


  nor
  g1819
  (
    n1826,
    n1696,
    n1801,
    n1674
  );


  nor
  g1820
  (
    n1828,
    n1408,
    n1422,
    n1688,
    n1697
  );


  or
  g1821
  (
    n1813,
    n1691,
    n1681,
    n1679,
    n1692
  );


  nand
  g1822
  (
    n1811,
    n1676,
    n1806,
    n1695,
    n1694
  );


  nand
  g1823
  (
    n1814,
    n1687,
    n1688,
    n1673
  );


  and
  g1824
  (
    n1830,
    n1693,
    n1698,
    n1804
  );


  or
  g1825
  (
    n1850,
    n1789,
    n1423,
    n1726,
    n1736
  );


  xnor
  g1826
  (
    n1901,
    n1843,
    n1776,
    n1767,
    n1765
  );


  and
  g1827
  (
    n1879,
    n1824,
    n1771,
    n1839,
    n1744
  );


  nor
  g1828
  (
    n1858,
    n1770,
    n1839,
    n1844,
    n1774
  );


  xnor
  g1829
  (
    n1903,
    n1757,
    n1812,
    n1766,
    n1782
  );


  nand
  g1830
  (
    n1854,
    n1843,
    n1700,
    n1790,
    n1759
  );


  nand
  g1831
  (
    n1853,
    n1774,
    n1839,
    n1791,
    n1752
  );


  xor
  g1832
  (
    n1863,
    n1770,
    n1807,
    n1781,
    n1766
  );


  and
  g1833
  (
    n1870,
    n1832,
    n1840,
    n1787,
    n1829
  );


  and
  g1834
  (
    n1877,
    n1780,
    n1783,
    n1846,
    n1756
  );


  nor
  g1835
  (
    n1880,
    n1783,
    n1776,
    n1775,
    n1761
  );


  nor
  g1836
  (
    n1871,
    n1768,
    n1816,
    n1759,
    n1748
  );


  xor
  g1837
  (
    n1866,
    n1846,
    n1762,
    n1827,
    n1787
  );


  nand
  g1838
  (
    n1896,
    n1734,
    n1783,
    n1745,
    n1791
  );


  or
  g1839
  (
    n1876,
    n1700,
    n1766,
    n1842,
    n1746
  );


  or
  g1840
  (
    n1900,
    n1701,
    n1780,
    n1844,
    n1699
  );


  nand
  g1841
  (
    n1886,
    n1843,
    n1770,
    n1185,
    n1783
  );


  or
  g1842
  (
    n1860,
    n1815,
    n1820,
    n1830,
    n1784
  );


  nor
  g1843
  (
    n1847,
    n1786,
    n1842,
    n1701,
    n1845
  );


  xor
  g1844
  (
    n1907,
    n1424,
    n1777,
    n1728,
    n1775
  );


  and
  g1845
  (
    n1872,
    n1841,
    n1767,
    n1821,
    n1752
  );


  xor
  g1846
  (
    n1867,
    n1765,
    n1729,
    n1779,
    n1778
  );


  nor
  g1847
  (
    n1851,
    n1788,
    n1743,
    n1838,
    n1828
  );


  xor
  g1848
  (
    n1874,
    n1767,
    n1762,
    n1763,
    n1751
  );


  nor
  g1849
  (
    n1887,
    n1841,
    n1760,
    n1772
  );


  and
  g1850
  (
    n1906,
    n1727,
    n1751,
    n1761,
    n1760
  );


  and
  g1851
  (
    n1904,
    n1845,
    n1740,
    n1782
  );


  nor
  g1852
  (
    n1885,
    n1755,
    n1790,
    n1846,
    n1754
  );


  xor
  g1853
  (
    n1892,
    n1785,
    n1788,
    n1843,
    n1758
  );


  nand
  g1854
  (
    n1852,
    n1774,
    n1765,
    n1823,
    n1759
  );


  and
  g1855
  (
    n1910,
    n1773,
    n1810,
    n1771,
    n1808
  );


  and
  g1856
  (
    n1848,
    n1777,
    n1771,
    n1749,
    n1731
  );


  nor
  g1857
  (
    n1897,
    n1834,
    n1764,
    n1833,
    n1760
  );


  or
  g1858
  (
    n1856,
    n1779,
    n1742,
    n1701,
    n105
  );


  xor
  g1859
  (
    n1883,
    n1840,
    n1791,
    n1789,
    n1738
  );


  xor
  g1860
  (
    n1884,
    n1768,
    n1753,
    n1779,
    n1781
  );


  nor
  g1861
  (
    n1909,
    n1700,
    n1763,
    n1769,
    n1699
  );


  xnor
  g1862
  (
    n1902,
    n1763,
    n1769,
    n1735,
    n1701
  );


  and
  g1863
  (
    n1862,
    n1778,
    n1840,
    n1756,
    n1733
  );


  xor
  g1864
  (
    n1881,
    n1781,
    n1775,
    n1786,
    n1845
  );


  or
  g1865
  (
    n1895,
    n1725,
    n1784,
    n1773,
    n1776
  );


  nor
  g1866
  (
    n1908,
    n1780,
    n1772,
    n1839,
    n1785
  );


  nand
  g1867
  (
    n1893,
    n1825,
    n1819,
    n1770,
    n1768
  );


  xnor
  g1868
  (
    n1873,
    n1774,
    n1785,
    n1846,
    n1754
  );


  xnor
  g1869
  (
    n1864,
    n1814,
    n1784,
    n1775,
    n1768
  );


  and
  g1870
  (
    n1859,
    n1755,
    n1764,
    n1778,
    n1788
  );


  nor
  g1871
  (
    n1889,
    n1790,
    n1741,
    n1842,
    n1844
  );


  nand
  g1872
  (
    n1857,
    n1730,
    n1777,
    n1787,
    n1764
  );


  nor
  g1873
  (
    n1849,
    n1781,
    n1780,
    n1836,
    n1813
  );


  xor
  g1874
  (
    n1891,
    n1818,
    n1835,
    n1786,
    n1784
  );


  or
  g1875
  (
    KeyWire_0_26,
    n1778,
    n1809,
    n1424,
    n1767
  );


  xor
  g1876
  (
    n1875,
    n1817,
    n1769,
    n1837,
    n1840
  );


  xor
  g1877
  (
    n1894,
    n1772,
    n1773,
    n1789,
    n1841
  );


  nand
  g1878
  (
    n1868,
    n1811,
    n1737,
    n1761,
    n1782
  );


  nor
  g1879
  (
    n1861,
    n1700,
    n1762,
    n1773,
    n1785
  );


  and
  g1880
  (
    n1905,
    n1788,
    n1759,
    n1822,
    n1423
  );


  xnor
  g1881
  (
    n1890,
    n1845,
    n1424,
    n1779,
    n1750
  );


  xnor
  g1882
  (
    n1882,
    n1776,
    n1757,
    n1769,
    n1787
  );


  nand
  g1883
  (
    n1878,
    n1765,
    n1842,
    n1771,
    n1760
  );


  xor
  g1884
  (
    n1898,
    n1791,
    n1753,
    n1747,
    n1764
  );


  nor
  g1885
  (
    n1869,
    n1739,
    n1766,
    n1761,
    n1732
  );


  xnor
  g1886
  (
    n1899,
    n1826,
    n1786,
    n1424,
    n1777
  );


  or
  g1887
  (
    KeyWire_0_30,
    n1762,
    n1841,
    n1831,
    n1763
  );


  and
  g1888
  (
    n1888,
    n1789,
    n1844,
    n1758,
    n1790
  );


  nand
  g1889
  (
    n1913,
    n1888,
    n1871,
    n1877,
    n1848
  );


  nand
  g1890
  (
    n1914,
    n1897,
    n1852,
    n1890,
    n1895
  );


  or
  g1891
  (
    n1912,
    n1853,
    n1859,
    n1867,
    n1874
  );


  xnor
  g1892
  (
    n1926,
    n1858,
    n1862,
    n1850,
    n1902
  );


  nor
  g1893
  (
    n1916,
    n1884,
    n1881,
    n1847,
    n1898
  );


  xnor
  g1894
  (
    n1921,
    n1866,
    n1875,
    n1851,
    n1878
  );


  and
  g1895
  (
    n1925,
    n1856,
    n1880,
    n1908,
    n1901
  );


  or
  g1896
  (
    n1911,
    n1886,
    n1868,
    n1879,
    n1860
  );


  xnor
  g1897
  (
    n1923,
    n1887,
    n1904,
    n1873,
    n1883
  );


  xnor
  g1898
  (
    n1917,
    n1861,
    n1907,
    n1900,
    n1865
  );


  xor
  g1899
  (
    n1918,
    n1903,
    n1882,
    n1910,
    n1864
  );


  and
  g1900
  (
    n1915,
    n1893,
    n1892,
    n1863,
    n1855
  );


  nor
  g1901
  (
    n1919,
    n1894,
    n1899,
    n1896,
    n1857
  );


  nor
  g1902
  (
    n1922,
    n1854,
    n1870,
    n1906,
    n1891
  );


  or
  g1903
  (
    n1924,
    n1869,
    n1905,
    n1889,
    n1876
  );


  xnor
  g1904
  (
    n1920,
    n1909,
    n1885,
    n1849,
    n1872
  );


  xor
  KeyGate_0_0
  (
    n92,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1208,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n173,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n420,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n27,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n650,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n31,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1067,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1189,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1142,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n969,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n502,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n601,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n562,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n263,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1364,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n772,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1212,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n557,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n1354,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1466,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n279,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n1265,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n820,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1732,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n518,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1865,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1731,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n737,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n216,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1855,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1725,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

