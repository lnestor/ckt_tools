// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_44 written by SynthGen on 2021/04/05 11:08:37
module Stat_100_44( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n112, n113, n114, n123, n105, n101, n122, n111,
 n115, n119, n110, n131, n103, n107, n109, n129,
 n116, n106, n128, n132, n130, n125, n120, n117,
 n118, n126, n127, n104, n121, n108, n102, n124);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n112, n113, n114, n123, n105, n101, n122, n111,
 n115, n119, n110, n131, n103, n107, n109, n129,
 n116, n106, n128, n132, n130, n125, n120, n117,
 n118, n126, n127, n104, n121, n108, n102, n124;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100;

not  g0 (n45, n19);
buf  g1 (n88, n21);
not  g2 (n39, n22);
not  g3 (n74, n18);
buf  g4 (n77, n31);
buf  g5 (n65, n6);
not  g6 (n71, n1);
not  g7 (n72, n25);
not  g8 (n75, n8);
buf  g9 (n70, n28);
buf  g10 (n82, n26);
not  g11 (n78, n32);
buf  g12 (n37, n20);
not  g13 (n46, n27);
buf  g14 (n84, n23);
not  g15 (n63, n15);
not  g16 (n50, n13);
not  g17 (n49, n27);
buf  g18 (n48, n3);
not  g19 (n60, n29);
buf  g20 (n33, n11);
not  g21 (n34, n29);
buf  g22 (n51, n14);
not  g23 (n52, n4);
not  g24 (n38, n27);
buf  g25 (n68, n23);
not  g26 (n85, n30);
not  g27 (n73, n25);
buf  g28 (n36, n24);
not  g29 (n55, n5);
buf  g30 (n43, n16);
not  g31 (n80, n28);
not  g32 (n86, n21);
buf  g33 (n66, n9);
buf  g34 (n76, n17);
not  g35 (n56, n29);
buf  g36 (n61, n21);
buf  g37 (n35, n32);
not  g38 (n79, n31);
buf  g39 (n83, n26);
buf  g40 (n58, n7);
not  g41 (n57, n24);
not  g42 (n41, n10);
buf  g43 (n40, n30);
buf  g44 (n69, n26);
buf  g45 (n54, n31);
buf  g46 (n47, n12);
buf  g47 (n64, n23);
buf  g48 (n62, n30);
buf  g49 (n81, n25);
buf  g50 (n44, n22);
buf  g51 (n87, n24);
buf  g52 (n53, n22);
buf  g53 (n42, n28);
buf  g54 (n59, n32);
buf  g55 (n67, n2);
buf  g56 (n91, n38);
not  g57 (n92, n36);
buf  g58 (n89, n34);
and  g59 (n90, n33, n35, n37);
not  g60 (n95, n91);
buf  g61 (n93, n90);
buf  g62 (n98, n92);
buf  g63 (n100, n92);
not  g64 (n97, n92);
not  g65 (n96, n91);
not  g66 (n94, n91);
buf  g67 (n99, n89);
xnor g68 (n127, n98, n75, n97, n54);
xor  g69 (n103, n69, n56, n62, n85);
or   g70 (n126, n88, n76, n63, n68);
and  g71 (n128, n100, n96, n45, n93);
xnor g72 (n113, n74, n51, n52, n76);
and  g73 (n129, n84, n99, n66);
xnor g74 (n118, n82, n44, n86, n88);
and  g75 (n114, n96, n98, n75, n70);
xor  g76 (n125, n81, n53, n66, n97);
nand g77 (n117, n71, n73, n79);
and  g78 (n123, n79, n72, n88);
nand g79 (n124, n43, n71, n95, n85);
xnor g80 (n119, n100, n81, n60, n94);
and  g81 (n104, n87, n66, n42, n86);
nand g82 (n132, n93, n69, n94, n77);
xnor g83 (n111, n76, n67, n70, n80);
xnor g84 (n107, n83, n82, n95, n77);
xnor g85 (n109, n99, n94, n82, n65);
or   g86 (n115, n98, n79, n49, n68);
xnor g87 (n121, n80, n50, n93, n68);
nand g88 (n101, n78, n99, n95, n41);
or   g89 (n110, n98, n78, n61, n100);
nand g90 (n131, n80, n40, n94, n78);
or   g91 (n112, n59, n48, n97, n58);
nand g92 (n105, n86, n46, n84, n81);
xnor g93 (n122, n97, n67, n39, n64);
xor  g94 (n108, n95, n75, n47, n70);
and  g95 (n120, n57, n87, n73, n96);
or   g96 (n130, n55, n69, n87, n100);
nand g97 (n116, n74, n85, n84, n96);
nand g98 (n106, n93, n67, n77, n74);
or   g99 (n102, n71, n83, n72);
endmodule
