// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_2799_38_8 written by SynthGen on 2021/06/15 15:06:09
module Stat_2799_38_8( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34,
 n1096, n1093, n1094, n1081, n1101, n1083, n1099, n1092,
 n1097, n1098, n1079, n1082, n1078, n1088, n1103, n1091,
 n2636, n2813, n2809, n2806, n2803, n2814, n2811, n2800,
 n2805, n2804, n2799, n2796, n2810, n2812, n2808, n2801,
 n2815, n2833);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34;

output n1096, n1093, n1094, n1081, n1101, n1083, n1099, n1092,
 n1097, n1098, n1079, n1082, n1078, n1088, n1103, n1091,
 n2636, n2813, n2809, n2806, n2803, n2814, n2811, n2800,
 n2805, n2804, n2799, n2796, n2810, n2812, n2808, n2801,
 n2815, n2833;

wire n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n487, n488, n489, n490,
 n491, n492, n493, n494, n495, n496, n497, n498,
 n499, n500, n501, n502, n503, n504, n505, n506,
 n507, n508, n509, n510, n511, n512, n513, n514,
 n515, n516, n517, n518, n519, n520, n521, n522,
 n523, n524, n525, n526, n527, n528, n529, n530,
 n531, n532, n533, n534, n535, n536, n537, n538,
 n539, n540, n541, n542, n543, n544, n545, n546,
 n547, n548, n549, n550, n551, n552, n553, n554,
 n555, n556, n557, n558, n559, n560, n561, n562,
 n563, n564, n565, n566, n567, n568, n569, n570,
 n571, n572, n573, n574, n575, n576, n577, n578,
 n579, n580, n581, n582, n583, n584, n585, n586,
 n587, n588, n589, n590, n591, n592, n593, n594,
 n595, n596, n597, n598, n599, n600, n601, n602,
 n603, n604, n605, n606, n607, n608, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n660, n661, n662, n663, n664, n665, n666,
 n667, n668, n669, n670, n671, n672, n673, n674,
 n675, n676, n677, n678, n679, n680, n681, n682,
 n683, n684, n685, n686, n687, n688, n689, n690,
 n691, n692, n693, n694, n695, n696, n697, n698,
 n699, n700, n701, n702, n703, n704, n705, n706,
 n707, n708, n709, n710, n711, n712, n713, n714,
 n715, n716, n717, n718, n719, n720, n721, n722,
 n723, n724, n725, n726, n727, n728, n729, n730,
 n731, n732, n733, n734, n735, n736, n737, n738,
 n739, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1080, n1084, n1085, n1086, n1087,
 n1089, n1090, n1095, n1100, n1102, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
 n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026,
 n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
 n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
 n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
 n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
 n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066,
 n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
 n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
 n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
 n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
 n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106,
 n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
 n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
 n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
 n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
 n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146,
 n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
 n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
 n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
 n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
 n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186,
 n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
 n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
 n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
 n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
 n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226,
 n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
 n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
 n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
 n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
 n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266,
 n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
 n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
 n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
 n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
 n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306,
 n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
 n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
 n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
 n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
 n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346,
 n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
 n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
 n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
 n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
 n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386,
 n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
 n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
 n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
 n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
 n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426,
 n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
 n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
 n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
 n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
 n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466,
 n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
 n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
 n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
 n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
 n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506,
 n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
 n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
 n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
 n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
 n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546,
 n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
 n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
 n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
 n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
 n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586,
 n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
 n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
 n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
 n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
 n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626,
 n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
 n2635, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
 n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
 n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
 n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
 n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675,
 n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
 n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
 n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
 n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
 n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715,
 n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
 n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
 n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
 n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
 n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
 n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
 n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
 n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
 n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
 n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795,
 n2797, n2798, n2802, n2807, n2816, n2817, n2818, n2819,
 n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
 n2828, n2829, n2830, n2831, n2832;

buf  g0 (n65, n16);
buf  g1 (n92, n11);
buf  g2 (n42, n26);
buf  g3 (n58, n12);
buf  g4 (n86, n26);
not  g5 (n41, n21);
buf  g6 (n85, n24);
not  g7 (n110, n12);
buf  g8 (n109, n19);
not  g9 (n38, n15);
buf  g10 (n75, n19);
buf  g11 (n68, n19);
buf  g12 (n117, n6);
buf  g13 (n91, n10);
buf  g14 (n48, n9);
buf  g15 (n81, n20);
not  g16 (n49, n10);
not  g17 (n35, n21);
not  g18 (n73, n16);
buf  g19 (n37, n13);
buf  g20 (n113, n20);
buf  g21 (n96, n12);
not  g22 (n83, n22);
not  g23 (n59, n20);
buf  g24 (n43, n12);
buf  g25 (n57, n4);
buf  g26 (n112, n18);
not  g27 (n54, n19);
buf  g28 (n114, n17);
not  g29 (n51, n25);
buf  g30 (n105, n22);
not  g31 (n111, n11);
not  g32 (n93, n20);
not  g33 (n63, n18);
buf  g34 (n104, n24);
not  g35 (n107, n17);
not  g36 (n56, n9);
buf  g37 (n95, n17);
not  g38 (n108, n11);
buf  g39 (n106, n18);
buf  g40 (n101, n2);
buf  g41 (n62, n26);
not  g42 (n78, n14);
buf  g43 (n71, n25);
not  g44 (n66, n23);
buf  g45 (n72, n18);
buf  g46 (n46, n13);
buf  g47 (n40, n15);
not  g48 (n80, n23);
buf  g49 (n94, n24);
not  g50 (n53, n10);
not  g51 (n89, n27);
buf  g52 (n87, n25);
not  g53 (n44, n5);
not  g54 (n70, n3);
buf  g55 (n55, n15);
buf  g56 (n47, n9);
buf  g57 (n67, n15);
buf  g58 (n84, n16);
not  g59 (n45, n8);
buf  g60 (n52, n27);
not  g61 (n39, n14);
buf  g62 (n88, n22);
buf  g63 (n74, n25);
buf  g64 (n60, n21);
not  g65 (n102, n23);
buf  g66 (n79, n23);
not  g67 (n100, n10);
buf  g68 (n103, n22);
not  g69 (n77, n26);
buf  g70 (n64, n14);
buf  g71 (n90, n1);
not  g72 (n115, n14);
buf  g73 (n118, n27);
buf  g74 (n116, n13);
buf  g75 (n36, n27);
not  g76 (n98, n21);
not  g77 (n76, n13);
not  g78 (n50, n7);
not  g79 (n97, n11);
buf  g80 (n82, n16);
not  g81 (n61, n24);
buf  g82 (n69, n17);
not  g83 (n99, n9);
buf  g84 (n398, n36);
not  g85 (n148, n102);
buf  g86 (n166, n109);
not  g87 (n188, n99);
buf  g88 (n344, n107);
buf  g89 (n200, n47);
not  g90 (n330, n89);
buf  g91 (n365, n47);
not  g92 (n401, n89);
not  g93 (n159, n76);
not  g94 (n302, n96);
buf  g95 (n278, n82);
buf  g96 (n342, n114);
buf  g97 (n238, n92);
buf  g98 (n300, n113);
not  g99 (n217, n37);
buf  g100 (n297, n90);
buf  g101 (n237, n105);
buf  g102 (n262, n40);
not  g103 (n431, n90);
buf  g104 (n241, n59);
buf  g105 (n204, n77);
not  g106 (n150, n106);
not  g107 (n301, n92);
not  g108 (n266, n82);
not  g109 (n199, n98);
not  g110 (n126, n106);
buf  g111 (n231, n84);
not  g112 (n163, n48);
not  g113 (n119, n97);
buf  g114 (n140, n74);
buf  g115 (n404, n78);
buf  g116 (n289, n64);
not  g117 (n244, n95);
not  g118 (n201, n89);
not  g119 (n338, n55);
buf  g120 (n160, n44);
buf  g121 (n189, n40);
buf  g122 (n240, n110);
not  g123 (n390, n69);
not  g124 (n259, n81);
buf  g125 (n320, n36);
buf  g126 (n382, n68);
not  g127 (n333, n88);
not  g128 (n247, n78);
buf  g129 (n412, n85);
buf  g130 (n303, n104);
buf  g131 (n352, n53);
buf  g132 (n357, n56);
not  g133 (n285, n41);
not  g134 (n232, n43);
not  g135 (n314, n73);
buf  g136 (n161, n98);
not  g137 (n206, n54);
buf  g138 (n326, n88);
not  g139 (n324, n68);
buf  g140 (n318, n49);
buf  g141 (n393, n43);
not  g142 (n235, n67);
not  g143 (n197, n56);
buf  g144 (n293, n49);
buf  g145 (n178, n113);
buf  g146 (n413, n92);
not  g147 (n378, n66);
not  g148 (n146, n76);
not  g149 (n355, n39);
buf  g150 (n423, n79);
not  g151 (n251, n102);
buf  g152 (n164, n114);
buf  g153 (n187, n83);
buf  g154 (n429, n97);
buf  g155 (n306, n63);
not  g156 (n373, n61);
not  g157 (n286, n108);
not  g158 (n220, n45);
buf  g159 (n135, n77);
buf  g160 (n349, n98);
buf  g161 (n127, n44);
not  g162 (n131, n53);
buf  g163 (n133, n54);
not  g164 (n215, n90);
buf  g165 (n253, n84);
buf  g166 (n249, n57);
buf  g167 (n172, n61);
buf  g168 (n417, n68);
buf  g169 (n151, n65);
buf  g170 (n122, n58);
not  g171 (n292, n55);
not  g172 (n261, n75);
not  g173 (n363, n104);
buf  g174 (n385, n58);
not  g175 (n192, n87);
not  g176 (n228, n85);
buf  g177 (n359, n80);
not  g178 (n136, n100);
buf  g179 (n339, n111);
buf  g180 (n134, n77);
not  g181 (n351, n41);
not  g182 (n145, n83);
buf  g183 (n291, n87);
buf  g184 (n422, n40);
buf  g185 (n380, n80);
buf  g186 (n399, n82);
not  g187 (n364, n51);
not  g188 (n316, n46);
not  g189 (n190, n46);
not  g190 (n130, n76);
buf  g191 (n275, n66);
buf  g192 (n198, n95);
buf  g193 (n202, n52);
buf  g194 (n386, n75);
not  g195 (n222, n69);
not  g196 (n230, n72);
not  g197 (n208, n36);
not  g198 (n180, n94);
buf  g199 (n205, n42);
buf  g200 (n141, n66);
not  g201 (n157, n79);
buf  g202 (n265, n93);
buf  g203 (n371, n39);
not  g204 (n125, n47);
buf  g205 (n287, n86);
not  g206 (n258, n90);
buf  g207 (n418, n38);
buf  g208 (n337, n94);
buf  g209 (n298, n93);
not  g210 (n277, n73);
not  g211 (n193, n100);
buf  g212 (n271, n71);
not  g213 (n165, n61);
not  g214 (n402, n80);
buf  g215 (n432, n74);
buf  g216 (n227, n103);
not  g217 (n169, n101);
not  g218 (n281, n36);
not  g219 (n213, n78);
not  g220 (n274, n40);
not  g221 (n149, n86);
buf  g222 (n394, n69);
not  g223 (n327, n64);
not  g224 (n255, n46);
buf  g225 (n374, n114);
not  g226 (n174, n65);
buf  g227 (n354, n68);
buf  g228 (n389, n109);
buf  g229 (n435, n59);
buf  g230 (n311, n72);
not  g231 (n284, n101);
buf  g232 (n283, n105);
buf  g233 (n321, n106);
buf  g234 (n310, n67);
buf  g235 (n309, n108);
buf  g236 (n436, n84);
buf  g237 (n438, n35);
not  g238 (n264, n85);
buf  g239 (n167, n86);
buf  g240 (n124, n70);
buf  g241 (n425, n35);
buf  g242 (n356, n113);
buf  g243 (n183, n58);
not  g244 (n223, n41);
buf  g245 (n366, n112);
not  g246 (n279, n52);
buf  g247 (n225, n91);
buf  g248 (n129, n37);
buf  g249 (n384, n88);
not  g250 (n252, n53);
not  g251 (n335, n99);
not  g252 (n362, n101);
buf  g253 (n211, n107);
not  g254 (n368, n79);
buf  g255 (n391, n99);
buf  g256 (n319, n42);
not  g257 (n154, n95);
not  g258 (n430, n52);
buf  g259 (n137, n63);
not  g260 (n269, n62);
not  g261 (n409, n104);
not  g262 (n143, n46);
buf  g263 (n236, n60);
buf  g264 (n392, n47);
buf  g265 (n170, n64);
not  g266 (n305, n63);
buf  g267 (n132, n78);
buf  g268 (n280, n35);
not  g269 (n340, n54);
buf  g270 (n139, n56);
buf  g271 (n176, n57);
buf  g272 (n214, n95);
not  g273 (n332, n65);
buf  g274 (n290, n45);
buf  g275 (n334, n86);
buf  g276 (n216, n103);
buf  g277 (n144, n72);
not  g278 (n294, n110);
not  g279 (n379, n110);
buf  g280 (n186, n60);
buf  g281 (n406, n111);
not  g282 (n307, n49);
not  g283 (n348, n103);
buf  g284 (n181, n50);
not  g285 (n155, n110);
buf  g286 (n194, n109);
buf  g287 (n218, n37);
buf  g288 (n196, n113);
buf  g289 (n168, n83);
not  g290 (n171, n74);
not  g291 (n428, n104);
buf  g292 (n203, n57);
buf  g293 (n325, n48);
not  g294 (n239, n77);
not  g295 (n424, n38);
buf  g296 (n345, n63);
buf  g297 (n153, n83);
buf  g298 (n234, n103);
not  g299 (n317, n72);
not  g300 (n185, n114);
not  g301 (n437, n98);
not  g302 (n120, n81);
buf  g303 (n147, n94);
buf  g304 (n175, n56);
not  g305 (n347, n105);
buf  g306 (n245, n69);
not  g307 (n123, n62);
not  g308 (n191, n76);
not  g309 (n254, n45);
not  g310 (n250, n70);
not  g311 (n427, n88);
buf  g312 (n350, n81);
buf  g313 (n387, n108);
not  g314 (n376, n96);
not  g315 (n407, n80);
buf  g316 (n256, n65);
not  g317 (n397, n37);
not  g318 (n403, n99);
buf  g319 (n388, n107);
buf  g320 (n336, n102);
buf  g321 (n182, n112);
buf  g322 (n346, n44);
buf  g323 (n260, n59);
buf  g324 (n246, n48);
not  g325 (n268, n50);
not  g326 (n273, n59);
not  g327 (n304, n39);
buf  g328 (n400, n38);
buf  g329 (n361, n91);
buf  g330 (n395, n89);
not  g331 (n242, n44);
not  g332 (n410, n74);
not  g333 (n226, n61);
not  g334 (n343, n87);
buf  g335 (n426, n52);
buf  g336 (n312, n92);
not  g337 (n179, n67);
buf  g338 (n315, n85);
not  g339 (n381, n42);
not  g340 (n370, n55);
not  g341 (n162, n93);
buf  g342 (n323, n87);
buf  g343 (n184, n48);
buf  g344 (n331, n73);
buf  g345 (n377, n60);
buf  g346 (n243, n79);
not  g347 (n341, n107);
buf  g348 (n408, n42);
buf  g349 (n248, n102);
buf  g350 (n414, n82);
buf  g351 (n322, n51);
not  g352 (n420, n96);
not  g353 (n128, n111);
not  g354 (n229, n43);
buf  g355 (n353, n73);
buf  g356 (n207, n49);
not  g357 (n360, n100);
buf  g358 (n416, n70);
not  g359 (n329, n50);
not  g360 (n419, n62);
buf  g361 (n267, n97);
not  g362 (n173, n94);
buf  g363 (n257, n91);
not  g364 (n375, n84);
buf  g365 (n142, n106);
not  g366 (n383, n35);
not  g367 (n313, n62);
not  g368 (n308, n111);
buf  g369 (n396, n51);
not  g370 (n296, n55);
not  g371 (n405, n112);
not  g372 (n212, n50);
not  g373 (n299, n71);
not  g374 (n282, n71);
buf  g375 (n272, n60);
not  g376 (n138, n66);
buf  g377 (n121, n108);
buf  g378 (n433, n70);
not  g379 (n270, n64);
buf  g380 (n263, n105);
buf  g381 (n233, n81);
buf  g382 (n156, n67);
buf  g383 (n369, n71);
buf  g384 (n358, n93);
not  g385 (n224, n58);
not  g386 (n276, n112);
buf  g387 (n210, n97);
buf  g388 (n221, n101);
not  g389 (n411, n96);
not  g390 (n372, n51);
buf  g391 (n415, n43);
buf  g392 (n328, n38);
not  g393 (n434, n41);
buf  g394 (n367, n75);
buf  g395 (n152, n54);
not  g396 (n219, n91);
buf  g397 (n158, n45);
buf  g398 (n295, n57);
not  g399 (n195, n53);
not  g400 (n421, n75);
buf  g401 (n209, n100);
not  g402 (n177, n109);
buf  g403 (n288, n39);
not  g404 (n618, n163);
not  g405 (n517, n152);
buf  g406 (n647, n156);
buf  g407 (n502, n139);
buf  g408 (n644, n124);
not  g409 (n514, n132);
buf  g410 (n612, n155);
buf  g411 (n613, n153);
not  g412 (n633, n166);
buf  g413 (n628, n145);
buf  g414 (n486, n151);
buf  g415 (n506, n121);
buf  g416 (n464, n146);
buf  g417 (n571, n170);
not  g418 (n573, n140);
not  g419 (n465, n120);
not  g420 (n619, n169);
buf  g421 (n593, n151);
buf  g422 (n615, n128);
buf  g423 (n459, n132);
buf  g424 (n575, n161);
not  g425 (n663, n138);
not  g426 (n559, n136);
buf  g427 (n590, n139);
not  g428 (n574, n125);
not  g429 (n544, n144);
buf  g430 (n478, n169);
buf  g431 (n538, n131);
not  g432 (n599, n148);
not  g433 (n651, n180);
buf  g434 (n582, n128);
buf  g435 (n454, n158);
buf  g436 (n462, n156);
buf  g437 (n659, n153);
buf  g438 (n626, n164);
buf  g439 (n585, n142);
buf  g440 (n529, n134);
not  g441 (n568, n167);
not  g442 (n449, n154);
buf  g443 (n584, n142);
buf  g444 (n600, n171);
not  g445 (n481, n122);
not  g446 (n472, n131);
buf  g447 (n662, n157);
not  g448 (n521, n124);
buf  g449 (n439, n124);
buf  g450 (n564, n126);
buf  g451 (n455, n166);
not  g452 (n623, n172);
buf  g453 (n587, n178);
not  g454 (n475, n177);
not  g455 (n492, n176);
buf  g456 (n441, n180);
not  g457 (n460, n136);
buf  g458 (n639, n180);
not  g459 (n646, n140);
buf  g460 (n669, n130);
not  g461 (n589, n132);
not  g462 (n624, n163);
not  g463 (n607, n179);
not  g464 (n643, n161);
not  g465 (n658, n140);
not  g466 (n550, n171);
buf  g467 (n660, n160);
buf  g468 (n510, n142);
buf  g469 (n503, n126);
not  g470 (n520, n125);
not  g471 (n572, n157);
not  g472 (n534, n164);
buf  g473 (n665, n165);
not  g474 (n526, n171);
buf  g475 (n484, n150);
buf  g476 (n483, n128);
buf  g477 (n451, n143);
not  g478 (n542, n119);
not  g479 (n604, n174);
not  g480 (n489, n174);
buf  g481 (n597, n148);
not  g482 (n594, n145);
not  g483 (n499, n149);
not  g484 (n448, n171);
not  g485 (n562, n145);
not  g486 (n527, n168);
buf  g487 (n567, n160);
buf  g488 (n553, n125);
not  g489 (n504, n140);
not  g490 (n555, n160);
buf  g491 (n598, n154);
buf  g492 (n603, n133);
buf  g493 (n557, n180);
not  g494 (n479, n177);
buf  g495 (n523, n179);
not  g496 (n476, n160);
buf  g497 (n609, n159);
buf  g498 (n463, n131);
not  g499 (n549, n134);
buf  g500 (n657, n147);
buf  g501 (n591, n144);
not  g502 (n588, n169);
not  g503 (n471, n135);
not  g504 (n636, n133);
not  g505 (n530, n144);
not  g506 (n495, n136);
not  g507 (n480, n159);
buf  g508 (n511, n137);
not  g509 (n668, n127);
not  g510 (n494, n162);
buf  g511 (n488, n155);
buf  g512 (n580, n178);
not  g513 (n616, n149);
buf  g514 (n563, n155);
buf  g515 (n501, n139);
not  g516 (n457, n127);
buf  g517 (n522, n129);
not  g518 (n490, n155);
buf  g519 (n664, n166);
buf  g520 (n453, n165);
not  g521 (n440, n177);
not  g522 (n491, n137);
not  g523 (n535, n178);
buf  g524 (n601, n147);
buf  g525 (n508, n172);
buf  g526 (n512, n167);
buf  g527 (n645, n174);
not  g528 (n654, n156);
not  g529 (n583, n135);
buf  g530 (n606, n129);
not  g531 (n469, n168);
buf  g532 (n498, n127);
buf  g533 (n671, n138);
not  g534 (n634, n149);
not  g535 (n631, n173);
not  g536 (n608, n178);
not  g537 (n466, n175);
buf  g538 (n630, n170);
not  g539 (n637, n173);
buf  g540 (n620, n147);
buf  g541 (n565, n170);
not  g542 (n497, n123);
not  g543 (n586, n128);
buf  g544 (n541, n150);
not  g545 (n496, n142);
buf  g546 (n477, n167);
buf  g547 (n470, n153);
not  g548 (n592, n154);
not  g549 (n546, n143);
buf  g550 (n445, n175);
buf  g551 (n461, n145);
buf  g552 (n667, n143);
not  g553 (n536, n125);
buf  g554 (n524, n173);
buf  g555 (n493, n176);
buf  g556 (n458, n135);
not  g557 (n570, n134);
not  g558 (n670, n163);
buf  g559 (n537, n162);
not  g560 (n482, n159);
buf  g561 (n532, n146);
not  g562 (n487, n164);
buf  g563 (n595, n152);
not  g564 (n611, n166);
not  g565 (n622, n149);
buf  g566 (n577, n144);
buf  g567 (n632, n162);
not  g568 (n648, n137);
buf  g569 (n543, n158);
not  g570 (n548, n134);
buf  g571 (n610, n141);
not  g572 (n525, n132);
not  g573 (n578, n165);
buf  g574 (n561, n139);
not  g575 (n468, n159);
buf  g576 (n638, n152);
not  g577 (n450, n176);
not  g578 (n500, n138);
buf  g579 (n452, n126);
buf  g580 (n473, n151);
not  g581 (n539, n146);
not  g582 (n518, n158);
buf  g583 (n528, n143);
buf  g584 (n569, n146);
not  g585 (n516, n169);
buf  g586 (n554, n141);
buf  g587 (n444, n152);
buf  g588 (n655, n133);
buf  g589 (n579, n138);
not  g590 (n629, n167);
not  g591 (n661, n148);
buf  g592 (n649, n165);
not  g593 (n625, n147);
buf  g594 (n545, n175);
not  g595 (n446, n168);
buf  g596 (n653, n157);
buf  g597 (n485, n173);
buf  g598 (n656, n130);
buf  g599 (n641, n148);
buf  g600 (n560, n162);
not  g601 (n605, n179);
buf  g602 (n617, n156);
buf  g603 (n547, n130);
not  g604 (n507, n151);
not  g605 (n552, n130);
not  g606 (n614, n131);
buf  g607 (n531, n158);
buf  g608 (n576, n137);
not  g609 (n558, n127);
buf  g610 (n443, n129);
buf  g611 (n505, n126);
buf  g612 (n566, n168);
not  g613 (n640, n154);
buf  g614 (n519, n150);
not  g615 (n666, n124);
buf  g616 (n515, n157);
not  g617 (n447, n141);
not  g618 (n467, n174);
not  g619 (n602, n141);
not  g620 (n540, n136);
not  g621 (n509, n129);
buf  g622 (n556, n161);
not  g623 (n621, n175);
not  g624 (n581, n170);
not  g625 (n642, n153);
not  g626 (n442, n150);
not  g627 (n551, n164);
not  g628 (n533, n133);
buf  g629 (n635, n135);
not  g630 (n456, n172);
not  g631 (n513, n172);
not  g632 (n627, n161);
buf  g633 (n596, n179);
not  g634 (n474, n163);
not  g635 (n652, n177);
not  g636 (n650, n176);
buf  g637 (n768, n582);
buf  g638 (n852, n619);
not  g639 (n761, n462);
buf  g640 (n774, n606);
buf  g641 (n690, n506);
buf  g642 (n726, n587);
buf  g643 (n707, n498);
not  g644 (n853, n590);
buf  g645 (n706, n538);
buf  g646 (n851, n508);
buf  g647 (n712, n535);
not  g648 (n672, n605);
not  g649 (n734, n567);
not  g650 (n718, n549);
not  g651 (n795, n530);
buf  g652 (n756, n560);
not  g653 (n778, n569);
not  g654 (n826, n621);
buf  g655 (n708, n449);
not  g656 (n765, n474);
buf  g657 (n735, n574);
not  g658 (n855, n183);
not  g659 (n847, n618);
not  g660 (n783, n604);
not  g661 (n822, n575);
not  g662 (n683, n456);
buf  g663 (n837, n531);
buf  g664 (n730, n545);
not  g665 (n695, n473);
not  g666 (n757, n623);
buf  g667 (n773, n602);
buf  g668 (n728, n572);
not  g669 (n723, n558);
not  g670 (n766, n581);
buf  g671 (n791, n517);
buf  g672 (n850, n520);
not  g673 (n770, n551);
buf  g674 (n680, n584);
buf  g675 (n842, n442);
buf  g676 (n737, n599);
buf  g677 (n789, n591);
not  g678 (n781, n555);
buf  g679 (n772, n493);
buf  g680 (n785, n532);
not  g681 (n694, n501);
not  g682 (n720, n479);
buf  g683 (n691, n464);
buf  g684 (n818, n475);
buf  g685 (n716, n613);
buf  g686 (n703, n446);
not  g687 (n701, n497);
not  g688 (n752, n597);
buf  g689 (n696, n593);
buf  g690 (n814, n554);
buf  g691 (n678, n482);
not  g692 (n674, n559);
buf  g693 (n760, n477);
buf  g694 (n697, n612);
not  g695 (n699, n458);
not  g696 (n856, n463);
buf  g697 (n688, n489);
not  g698 (n704, n607);
not  g699 (n709, n546);
not  g700 (n838, n483);
buf  g701 (n831, n588);
buf  g702 (n762, n585);
buf  g703 (n724, n445);
not  g704 (n857, n443);
buf  g705 (n802, n514);
buf  g706 (n820, n440);
not  g707 (n763, n598);
not  g708 (n731, n451);
buf  g709 (n854, n523);
buf  g710 (n817, n529);
buf  g711 (n788, n183);
not  g712 (n733, n571);
buf  g713 (n848, n488);
not  g714 (n815, n541);
not  g715 (n796, n492);
buf  g716 (n813, n595);
buf  g717 (n767, n609);
buf  g718 (n845, n548);
not  g719 (n829, n499);
not  g720 (n754, n533);
not  g721 (n685, n527);
buf  g722 (n780, n544);
not  g723 (n828, n573);
buf  g724 (n790, n181);
not  g725 (n849, n615);
buf  g726 (n782, n600);
not  g727 (n825, n563);
not  g728 (n816, n470);
buf  g729 (n810, n182);
not  g730 (n808, n510);
buf  g731 (n710, n570);
buf  g732 (n753, n448);
not  g733 (n732, n511);
not  g734 (n744, n608);
not  g735 (n715, n586);
not  g736 (n755, n580);
buf  g737 (n841, n518);
not  g738 (n804, n181);
not  g739 (n806, n486);
not  g740 (n677, n491);
not  g741 (n747, n450);
buf  g742 (n809, n500);
not  g743 (n713, n515);
buf  g744 (n681, n471);
not  g745 (n799, n543);
buf  g746 (n751, n534);
buf  g747 (n798, n496);
not  g748 (n811, n610);
buf  g749 (n693, n579);
buf  g750 (n833, n444);
not  g751 (n832, n526);
buf  g752 (n702, n182);
buf  g753 (n745, n616);
not  g754 (n673, n181);
buf  g755 (n729, n461);
buf  g756 (n839, n550);
not  g757 (n801, n553);
not  g758 (n721, n457);
buf  g759 (n705, n460);
not  g760 (n758, n184);
not  g761 (n794, n596);
not  g762 (n741, n452);
not  g763 (n675, n502);
not  g764 (n846, n577);
not  g765 (n700, n505);
buf  g766 (n819, n441);
buf  g767 (n771, n614);
buf  g768 (n687, n495);
buf  g769 (n684, n611);
not  g770 (n821, n182);
not  g771 (n746, n542);
buf  g772 (n787, n524);
buf  g773 (n830, n184);
not  g774 (n844, n557);
not  g775 (n714, n472);
buf  g776 (n823, n183);
buf  g777 (n692, n447);
not  g778 (n776, n181);
not  g779 (n722, n552);
not  g780 (n800, n576);
buf  g781 (n807, n484);
buf  g782 (n786, n439);
buf  g783 (n779, n453);
not  g784 (n805, n528);
buf  g785 (n764, n556);
not  g786 (n736, n561);
buf  g787 (n717, n583);
not  g788 (n686, n513);
not  g789 (n834, n622);
not  g790 (n749, n455);
buf  g791 (n676, n522);
buf  g792 (n727, n494);
not  g793 (n738, n624);
buf  g794 (n740, n485);
not  g795 (n797, n459);
not  g796 (n750, n519);
not  g797 (n682, n467);
buf  g798 (n743, n465);
buf  g799 (n759, n183);
not  g800 (n843, n568);
not  g801 (n742, n578);
not  g802 (n792, n487);
not  g803 (n725, n620);
buf  g804 (n835, n601);
buf  g805 (n803, n564);
not  g806 (n698, n539);
buf  g807 (n739, n566);
not  g808 (n775, n466);
buf  g809 (n777, n184);
not  g810 (n793, n537);
buf  g811 (n769, n469);
not  g812 (n689, n562);
not  g813 (n719, n476);
not  g814 (n840, n565);
not  g815 (n836, n182);
buf  g816 (n812, n490);
buf  g817 (n748, n509);
xnor g818 (n679, n516, n589, n512, n536);
or   g819 (n784, n547, n454, n540, n478);
nand g820 (n827, n481, n525, n592, n504);
nand g821 (n824, n521, n594, n468, n603);
or   g822 (n711, n503, n480, n507, n617);
not  g823 (n934, n851);
buf  g824 (n972, n778);
buf  g825 (n986, n702);
buf  g826 (n932, n852);
not  g827 (n979, n733);
buf  g828 (n889, n781);
buf  g829 (n897, n847);
not  g830 (n1048, n845);
not  g831 (n874, n796);
buf  g832 (n859, n716);
not  g833 (n890, n815);
not  g834 (n871, n776);
not  g835 (n1014, n843);
not  g836 (n1001, n854);
not  g837 (n1012, n693);
buf  g838 (n914, n808);
not  g839 (n900, n775);
not  g840 (n1076, n784);
not  g841 (n1074, n761);
not  g842 (n1052, n748);
not  g843 (n868, n727);
buf  g844 (n994, n725);
not  g845 (n1059, n821);
not  g846 (n931, n842);
not  g847 (n960, n850);
not  g848 (n1041, n760);
not  g849 (n1055, n786);
not  g850 (n1009, n852);
buf  g851 (n891, n851);
buf  g852 (n1043, n831);
not  g853 (n1040, n814);
buf  g854 (n950, n772);
not  g855 (n995, n756);
not  g856 (n964, n745);
buf  g857 (n1021, n717);
not  g858 (n901, n840);
buf  g859 (n865, n833);
buf  g860 (n872, n854);
not  g861 (n862, n798);
not  g862 (n913, n741);
not  g863 (n881, n836);
buf  g864 (n884, n724);
not  g865 (n1034, n847);
buf  g866 (n1003, n707);
buf  g867 (n992, n758);
buf  g868 (n894, n825);
not  g869 (n879, n828);
buf  g870 (n1030, n835);
buf  g871 (n880, n843);
not  g872 (n1071, n739);
not  g873 (n915, n714);
not  g874 (n1047, n845);
buf  g875 (n1016, n807);
buf  g876 (n858, n783);
not  g877 (n910, n742);
buf  g878 (n998, n804);
not  g879 (n967, n851);
not  g880 (n930, n848);
buf  g881 (n990, n802);
not  g882 (n916, n734);
buf  g883 (n941, n843);
not  g884 (n938, n803);
buf  g885 (n878, n845);
buf  g886 (n999, n846);
not  g887 (n963, n782);
buf  g888 (n1020, n826);
not  g889 (n937, n834);
not  g890 (n952, n847);
not  g891 (n873, n785);
not  g892 (n985, n699);
buf  g893 (n924, n747);
buf  g894 (n1004, n822);
not  g895 (n1028, n752);
not  g896 (n1049, n681);
buf  g897 (n1066, n841);
buf  g898 (n1035, n844);
not  g899 (n954, n736);
not  g900 (n961, n695);
not  g901 (n885, n771);
buf  g902 (n1029, n837);
not  g903 (n1070, n812);
buf  g904 (n898, n843);
buf  g905 (n923, n692);
not  g906 (n1036, n682);
buf  g907 (n942, n749);
not  g908 (n971, n746);
buf  g909 (n975, n751);
buf  g910 (n1019, n845);
not  g911 (n958, n844);
not  g912 (n918, n811);
buf  g913 (n907, n792);
not  g914 (n1015, n672);
buf  g915 (n1044, n677);
not  g916 (n870, n678);
not  g917 (n991, n706);
buf  g918 (n1011, n766);
buf  g919 (n1031, n721);
buf  g920 (n949, n787);
buf  g921 (n1045, n810);
not  g922 (n1072, n852);
buf  g923 (n1053, n732);
not  g924 (n1051, n853);
not  g925 (n981, n842);
not  g926 (n939, n846);
not  g927 (n953, n675);
buf  g928 (n983, n759);
buf  g929 (n1022, n838);
buf  g930 (n887, n743);
not  g931 (n976, n848);
not  g932 (n989, n819);
buf  g933 (n863, n849);
buf  g934 (n929, n780);
buf  g935 (n1018, n813);
not  g936 (n946, n824);
buf  g937 (n987, n685);
not  g938 (n1037, n701);
buf  g939 (n997, n839);
buf  g940 (n1067, n790);
buf  g941 (n921, n823);
not  g942 (n955, n767);
not  g943 (n1000, n729);
not  g944 (n1063, n723);
not  g945 (n1002, n797);
not  g946 (n974, n846);
not  g947 (n917, n686);
buf  g948 (n1017, n673);
buf  g949 (n1024, n849);
buf  g950 (n877, n853);
not  g951 (n1013, n737);
not  g952 (n1023, n849);
not  g953 (n927, n755);
not  g954 (n1027, n712);
buf  g955 (n968, n700);
not  g956 (n1077, n799);
not  g957 (n965, n805);
buf  g958 (n912, n697);
buf  g959 (n1007, n816);
not  g960 (n1039, n710);
not  g961 (n933, n719);
not  g962 (n948, n853);
not  g963 (n1064, n680);
buf  g964 (n977, n684);
not  g965 (n902, n709);
buf  g966 (n899, n750);
buf  g967 (n919, n730);
not  g968 (n1046, n718);
not  g969 (n982, n842);
buf  g970 (n969, n720);
buf  g971 (n1054, n764);
buf  g972 (n945, n689);
buf  g973 (n1008, n705);
not  g974 (n970, n846);
not  g975 (n886, n687);
not  g976 (n882, n852);
not  g977 (n876, n691);
buf  g978 (n943, n830);
buf  g979 (n966, n740);
not  g980 (n1057, n806);
buf  g981 (n909, n817);
buf  g982 (n978, n777);
not  g983 (n1069, n844);
buf  g984 (n888, n731);
buf  g985 (n922, n768);
not  g986 (n936, n850);
buf  g987 (n1075, n793);
buf  g988 (n957, n769);
not  g989 (n1058, n844);
buf  g990 (n996, n690);
buf  g991 (n867, n849);
buf  g992 (n908, n801);
buf  g993 (n993, n791);
buf  g994 (n905, n795);
buf  g995 (n1006, n676);
buf  g996 (n861, n757);
not  g997 (n956, n850);
buf  g998 (n973, n735);
not  g999 (n904, n722);
buf  g1000 (n911, n726);
buf  g1001 (n944, n773);
buf  g1002 (n903, n744);
buf  g1003 (n951, n711);
buf  g1004 (n860, n851);
not  g1005 (n925, n694);
buf  g1006 (n1050, n789);
not  g1007 (n906, n708);
buf  g1008 (n1026, n774);
not  g1009 (n1073, n698);
buf  g1010 (n1065, n738);
buf  g1011 (n896, n762);
buf  g1012 (n1033, n763);
buf  g1013 (n1060, n818);
not  g1014 (n988, n704);
not  g1015 (n980, n674);
buf  g1016 (n1005, n715);
not  g1017 (n1010, n703);
not  g1018 (n866, n848);
buf  g1019 (n1025, n770);
not  g1020 (n1038, n842);
buf  g1021 (n926, n713);
buf  g1022 (n1056, n794);
not  g1023 (n1061, n820);
not  g1024 (n935, n779);
buf  g1025 (n892, n679);
not  g1026 (n864, n829);
not  g1027 (n928, n850);
not  g1028 (n962, n788);
buf  g1029 (n984, n827);
not  g1030 (n1032, n688);
buf  g1031 (n875, n848);
buf  g1032 (n1062, n809);
buf  g1033 (n1042, n728);
not  g1034 (n895, n754);
buf  g1035 (n920, n765);
not  g1036 (n947, n832);
buf  g1037 (n893, n683);
buf  g1038 (n869, n800);
not  g1039 (n959, n696);
not  g1040 (n883, n753);
buf  g1041 (n940, n853);
not  g1042 (n1068, n847);
nand g1043 (n1098, n890, n916);
xor  g1044 (n1102, n912, n879, n917, n915);
nand g1045 (n1090, n920, n896, n860, n918);
xnor g1046 (n1081, n917, n863, n886, n915);
nand g1047 (n1079, n913, n914, n903, n910);
xnor g1048 (n1087, n913, n911, n876, n916);
or   g1049 (n1095, n906, n872, n870, n894);
and  g1050 (n1086, n920, n887, n902, n911);
xnor g1051 (n1093, n888, n910, n854, n884);
nand g1052 (n1100, n918, n919, n920, n877);
and  g1053 (n1084, n892, n905, n909);
or   g1054 (n1101, n880, n914, n910);
xor  g1055 (n1091, n891, n878, n900, n893);
xnor g1056 (n1085, n918, n881, n921, n901);
xnor g1057 (n1094, n913, n912, n911, n919);
xor  g1058 (n1097, n874, n869, n859, n919);
nand g1059 (n1080, n913, n883, n904, n889);
xor  g1060 (n1099, n858, n868, n916, n895);
xor  g1061 (n1078, n898, n871, n899, n915);
nand g1062 (n1089, n907, n864, n909, n920);
and  g1063 (n1092, n914, n912, n865);
xor  g1064 (n1082, n910, n916, n866, n854);
and  g1065 (n1088, n911, n915, n861, n918);
xor  g1066 (n1083, n873, n875, n908, n862);
nor  g1067 (n1103, n885, n867, n882, n897);
xnor g1068 (n1096, n909, n919, n917);
nand g1069 (n1104, n923, n1101);
xnor g1070 (n1106, n922, n1094);
and  g1071 (n1107, n922, n1102);
nor  g1072 (n1112, n922, n921);
xor  g1073 (n1105, n921, n922);
and  g1074 (n1111, n923, n1097);
nand g1075 (n1113, n1100, n1095);
and  g1076 (n1109, n1103, n923);
or   g1077 (n1110, n1096, n921);
or   g1078 (n1108, n1098, n1099);
not  g1079 (n1124, n1107);
not  g1080 (n1122, n1105);
buf  g1081 (n1119, n1106);
not  g1082 (n1120, n1105);
not  g1083 (n1115, n1107);
not  g1084 (n1114, n1104);
not  g1085 (n1118, n1106);
buf  g1086 (n1123, n1106);
buf  g1087 (n1117, n1105);
buf  g1088 (n1126, n1104);
not  g1089 (n1125, n1104);
not  g1090 (n1116, n1105);
buf  g1091 (n1127, n1104);
buf  g1092 (n1121, n1106);
not  g1093 (n1169, n1126);
not  g1094 (n1183, n1116);
buf  g1095 (n1178, n1122);
buf  g1096 (n1176, n1115);
buf  g1097 (n1168, n1121);
not  g1098 (n1161, n1123);
not  g1099 (n1150, n1121);
not  g1100 (n1140, n1117);
not  g1101 (n1137, n1120);
buf  g1102 (n1133, n1118);
not  g1103 (n1136, n1121);
buf  g1104 (n1154, n1127);
buf  g1105 (n1152, n1122);
not  g1106 (n1160, n1119);
buf  g1107 (n1173, n1126);
buf  g1108 (n1132, n1127);
buf  g1109 (n1165, n1120);
buf  g1110 (n1148, n1126);
not  g1111 (n1179, n1123);
not  g1112 (n1134, n1116);
not  g1113 (n1159, n1114);
buf  g1114 (n1139, n1127);
not  g1115 (n1143, n1124);
not  g1116 (n1141, n1119);
not  g1117 (n1162, n1123);
buf  g1118 (n1142, n1120);
not  g1119 (n1138, n1114);
not  g1120 (n1131, n1119);
buf  g1121 (n1129, n1115);
buf  g1122 (n1182, n1122);
buf  g1123 (n1157, n1114);
buf  g1124 (n1128, n1127);
buf  g1125 (n1156, n1114);
buf  g1126 (n1158, n1118);
not  g1127 (n1151, n1116);
not  g1128 (n1153, n1124);
not  g1129 (n1164, n1125);
not  g1130 (n1174, n1118);
not  g1131 (n1171, n1125);
buf  g1132 (n1180, n1125);
buf  g1133 (n1149, n1115);
not  g1134 (n1163, n1124);
not  g1135 (n1135, n1124);
buf  g1136 (n1170, n1118);
buf  g1137 (n1177, n1121);
not  g1138 (n1167, n1117);
not  g1139 (n1175, n1123);
buf  g1140 (n1144, n1122);
buf  g1141 (n1130, n1115);
buf  g1142 (n1172, n1117);
buf  g1143 (n1146, n1120);
buf  g1144 (n1155, n1126);
not  g1145 (n1166, n1117);
buf  g1146 (n1181, n1125);
not  g1147 (n1147, n1119);
buf  g1148 (n1145, n1116);
not  g1149 (n1185, n1135);
not  g1150 (n1256, n1136);
buf  g1151 (n1263, n1128);
buf  g1152 (n1260, n1140);
not  g1153 (n1190, n1143);
buf  g1154 (n1230, n1138);
buf  g1155 (n1234, n1128);
buf  g1156 (n1239, n1134);
buf  g1157 (n1224, n1146);
buf  g1158 (n1205, n1129);
not  g1159 (n1248, n1132);
buf  g1160 (n1213, n1140);
buf  g1161 (n1210, n1139);
buf  g1162 (n1227, n1129);
buf  g1163 (n1225, n1136);
not  g1164 (n1219, n1141);
not  g1165 (n1212, n1129);
not  g1166 (n1232, n1133);
not  g1167 (n1257, n1147);
not  g1168 (n1197, n1130);
not  g1169 (n1246, n1131);
not  g1170 (n1218, n1140);
not  g1171 (n1199, n1135);
buf  g1172 (n1245, n1131);
not  g1173 (n1184, n1142);
not  g1174 (n1223, n1133);
not  g1175 (n1233, n1130);
not  g1176 (n1189, n1146);
buf  g1177 (n1258, n1141);
buf  g1178 (n1240, n1142);
not  g1179 (n1220, n1147);
not  g1180 (n1250, n1138);
not  g1181 (n1254, n1147);
buf  g1182 (n1215, n1130);
buf  g1183 (n1195, n1146);
not  g1184 (n1186, n1144);
not  g1185 (n1259, n1144);
not  g1186 (n1192, n1133);
buf  g1187 (n1255, n1142);
not  g1188 (n1236, n1139);
buf  g1189 (n1251, n1129);
buf  g1190 (n1262, n1142);
buf  g1191 (n1222, n1139);
not  g1192 (n1243, n1145);
not  g1193 (n1217, n1141);
not  g1194 (n1206, n1138);
buf  g1195 (n1191, n1144);
not  g1196 (n1207, n1144);
buf  g1197 (n1211, n1137);
buf  g1198 (n1209, n1134);
not  g1199 (n1238, n1135);
not  g1200 (n1196, n1145);
not  g1201 (n1249, n1136);
not  g1202 (n1198, n1128);
not  g1203 (n1193, n1146);
buf  g1204 (n1242, n1135);
not  g1205 (n1194, n1140);
buf  g1206 (n1202, n1143);
buf  g1207 (n1235, n1131);
buf  g1208 (n1247, n1130);
not  g1209 (n1187, n1132);
buf  g1210 (n1241, n1132);
not  g1211 (n1221, n1137);
not  g1212 (n1226, n1134);
buf  g1213 (n1253, n1145);
not  g1214 (n1188, n1138);
buf  g1215 (n1237, n1143);
not  g1216 (n1252, n1139);
not  g1217 (n1204, n1128);
buf  g1218 (n1229, n1131);
not  g1219 (n1216, n1147);
buf  g1220 (n1231, n1134);
buf  g1221 (n1200, n1137);
buf  g1222 (n1201, n1143);
not  g1223 (n1261, n1136);
not  g1224 (n1244, n1137);
buf  g1225 (n1214, n1133);
buf  g1226 (n1208, n1145);
not  g1227 (n1228, n1132);
not  g1228 (n1203, n1141);
buf  g1229 (n1551, n29);
buf  g1230 (n1404, n1160);
buf  g1231 (n1350, n1255);
not  g1232 (n1382, n1200);
buf  g1233 (n1453, n924);
not  g1234 (n1267, n186);
not  g1235 (n1405, n1263);
not  g1236 (n1386, n1154);
not  g1237 (n1412, n1222);
not  g1238 (n1302, n1242);
buf  g1239 (n1339, n1174);
not  g1240 (n1318, n1169);
not  g1241 (n1288, n1225);
not  g1242 (n1450, n1248);
buf  g1243 (n1526, n185);
not  g1244 (n1313, n1211);
buf  g1245 (n1373, n29);
buf  g1246 (n1452, n1206);
not  g1247 (n1272, n1178);
not  g1248 (n1304, n1203);
not  g1249 (n1299, n1165);
buf  g1250 (n1518, n1160);
not  g1251 (n1457, n1218);
not  g1252 (n1578, n1185);
not  g1253 (n1490, n926);
buf  g1254 (n1265, n857);
buf  g1255 (n1466, n1206);
buf  g1256 (n1371, n1204);
not  g1257 (n1414, n1184);
buf  g1258 (n1550, n925);
buf  g1259 (n1446, n1223);
not  g1260 (n1555, n857);
buf  g1261 (n1530, n1234);
buf  g1262 (n1368, n1159);
not  g1263 (n1338, n1246);
buf  g1264 (n1417, n30);
buf  g1265 (n1568, n1192);
buf  g1266 (n1311, n1168);
buf  g1267 (n1362, n1260);
not  g1268 (n1547, n1253);
not  g1269 (n1432, n28);
buf  g1270 (n1374, n1168);
not  g1271 (n1381, n1251);
not  g1272 (n1308, n1241);
buf  g1273 (n1325, n1183);
not  g1274 (n1482, n31);
buf  g1275 (n1331, n1160);
buf  g1276 (n1460, n855);
buf  g1277 (n1438, n1151);
not  g1278 (n1495, n1171);
buf  g1279 (n1275, n1195);
buf  g1280 (n1473, n1209);
buf  g1281 (n1561, n1216);
not  g1282 (n1570, n1186);
not  g1283 (n1581, n1220);
buf  g1284 (n1556, n1153);
buf  g1285 (n1546, n1242);
buf  g1286 (n1310, n1226);
not  g1287 (n1497, n855);
not  g1288 (n1408, n29);
buf  g1289 (n1538, n1227);
not  g1290 (n1341, n1232);
not  g1291 (n1485, n1260);
not  g1292 (n1360, n1162);
not  g1293 (n1477, n1200);
buf  g1294 (n1471, n626);
not  g1295 (n1300, n1181);
not  g1296 (n1503, n1233);
buf  g1297 (n1519, n1194);
not  g1298 (n1549, n1232);
buf  g1299 (n1456, n1214);
buf  g1300 (n1296, n1261);
not  g1301 (n1527, n1163);
buf  g1302 (n1552, n630);
not  g1303 (n1539, n1244);
not  g1304 (n1291, n1228);
buf  g1305 (n1448, n1193);
buf  g1306 (n1491, n1213);
buf  g1307 (n1565, n1168);
not  g1308 (n1294, n1252);
buf  g1309 (n1274, n1173);
buf  g1310 (n1461, n31);
buf  g1311 (n1326, n1204);
not  g1312 (n1402, n1178);
buf  g1313 (n1483, n1191);
buf  g1314 (n1455, n1242);
buf  g1315 (n1467, n1150);
buf  g1316 (n1280, n1213);
not  g1317 (n1337, n1153);
buf  g1318 (n1501, n1174);
buf  g1319 (n1564, n1233);
buf  g1320 (n1306, n1167);
not  g1321 (n1352, n1204);
not  g1322 (n1582, n1180);
not  g1323 (n1447, n1161);
buf  g1324 (n1433, n1198);
buf  g1325 (n1378, n1250);
not  g1326 (n1445, n1225);
not  g1327 (n1364, n1165);
not  g1328 (n1407, n1233);
not  g1329 (n1524, n1258);
not  g1330 (n1506, n186);
not  g1331 (n1298, n1182);
not  g1332 (n1428, n1240);
buf  g1333 (n1369, n1185);
buf  g1334 (n1573, n1167);
not  g1335 (n1282, n1177);
buf  g1336 (n1545, n1241);
buf  g1337 (n1492, n1212);
not  g1338 (n1421, n1244);
not  g1339 (n1301, n1228);
buf  g1340 (n1354, n1152);
buf  g1341 (n1328, n1175);
not  g1342 (n1356, n1221);
buf  g1343 (n1419, n1187);
not  g1344 (n1383, n1195);
buf  g1345 (n1489, n1186);
buf  g1346 (n1554, n1263);
not  g1347 (n1580, n1252);
not  g1348 (n1520, n1199);
buf  g1349 (n1523, n1238);
not  g1350 (n1416, n1166);
buf  g1351 (n1397, n1261);
not  g1352 (n1476, n1233);
not  g1353 (n1384, n1208);
not  g1354 (n1387, n1153);
not  g1355 (n1474, n1194);
not  g1356 (n1403, n1185);
buf  g1357 (n1572, n1182);
buf  g1358 (n1349, n1194);
buf  g1359 (n1444, n1174);
not  g1360 (n1425, n1200);
not  g1361 (n1345, n1251);
not  g1362 (n1398, n1230);
not  g1363 (n1516, n856);
not  g1364 (n1499, n1221);
not  g1365 (n1393, n1198);
not  g1366 (n1353, n1208);
buf  g1367 (n1576, n1212);
not  g1368 (n1422, n1185);
not  g1369 (n1470, n1191);
buf  g1370 (n1424, n1231);
buf  g1371 (n1420, n631);
buf  g1372 (n1312, n1244);
buf  g1373 (n1577, n1163);
not  g1374 (n1537, n28);
not  g1375 (n1363, n1202);
buf  g1376 (n1329, n1170);
not  g1377 (n1367, n1188);
not  g1378 (n1320, n1189);
buf  g1379 (n1479, n1186);
buf  g1380 (n1449, n1263);
not  g1381 (n1463, n1163);
not  g1382 (n1451, n1205);
not  g1383 (n1400, n1209);
buf  g1384 (n1468, n1157);
not  g1385 (n1287, n1173);
buf  g1386 (n1548, n1201);
not  g1387 (n1500, n1191);
buf  g1388 (n1544, n1180);
not  g1389 (n1284, n1158);
buf  g1390 (n1285, n1171);
not  g1391 (n1567, n1219);
buf  g1392 (n1351, n1173);
buf  g1393 (n1563, n1190);
buf  g1394 (n1542, n1239);
not  g1395 (n1507, n1178);
buf  g1396 (n1279, n1158);
buf  g1397 (n1528, n856);
buf  g1398 (n1543, n1258);
buf  g1399 (n1406, n1215);
buf  g1400 (n1372, n1262);
not  g1401 (n1493, n1254);
buf  g1402 (n1512, n1162);
not  g1403 (n1270, n1156);
not  g1404 (n1347, n1244);
buf  g1405 (n1439, n856);
not  g1406 (n1511, n1193);
buf  g1407 (n1380, n925);
not  g1408 (n1395, n1180);
buf  g1409 (n1464, n1246);
not  g1410 (n1323, n1235);
not  g1411 (n1437, n1258);
not  g1412 (n1531, n1239);
not  g1413 (n1436, n1256);
buf  g1414 (n1293, n1151);
not  g1415 (n1553, n1245);
not  g1416 (n1342, n1189);
buf  g1417 (n1264, n1197);
buf  g1418 (n1566, n924);
not  g1419 (n1303, n185);
buf  g1420 (n1391, n1256);
not  g1421 (n1388, n1255);
buf  g1422 (n1361, n1254);
not  g1423 (n1305, n1259);
buf  g1424 (n1319, n1217);
not  g1425 (n1469, n1259);
buf  g1426 (n1557, n28);
buf  g1427 (n1376, n1171);
buf  g1428 (n1533, n1151);
not  g1429 (n1558, n1184);
not  g1430 (n1583, n1212);
buf  g1431 (n1454, n1254);
not  g1432 (n1509, n1219);
not  g1433 (n1399, n1157);
buf  g1434 (n1266, n1236);
buf  g1435 (n1486, n1182);
not  g1436 (n1307, n1194);
not  g1437 (n1559, n1225);
not  g1438 (n1346, n1228);
buf  g1439 (n1348, n925);
not  g1440 (n1314, n1192);
buf  g1441 (n1475, n1159);
not  g1442 (n1434, n1231);
buf  g1443 (n1276, n1159);
buf  g1444 (n1327, n1175);
not  g1445 (n1309, n1184);
not  g1446 (n1579, n30);
buf  g1447 (n1357, n1225);
buf  g1448 (n1278, n1238);
not  g1449 (n1286, n1251);
not  g1450 (n1535, n1197);
not  g1451 (n1340, n1170);
not  g1452 (n1478, n30);
buf  g1453 (n1401, n1157);
buf  g1454 (n1459, n1150);
buf  g1455 (n1332, n1222);
not  g1456 (n1514, n1237);
buf  g1457 (n1295, n1211);
not  g1458 (n1440, n1238);
not  g1459 (n1508, n1229);
not  g1460 (n1441, n1170);
buf  g1461 (n1560, n1224);
not  g1462 (n1515, n1196);
not  g1463 (n1529, n185);
buf  g1464 (n1370, n1263);
buf  g1465 (n1442, n1196);
not  g1466 (n1430, n1236);
not  g1467 (n1375, n1176);
buf  g1468 (n1496, n1201);
buf  g1469 (n1336, n1235);
buf  g1470 (n1394, n1235);
buf  g1471 (n1510, n1189);
buf  g1472 (n1431, n1156);
buf  g1473 (n1290, n1215);
buf  g1474 (n1494, n1261);
not  g1475 (n1481, n1205);
not  g1476 (n1324, n1210);
not  g1477 (n1410, n1220);
not  g1478 (n1385, n1191);
buf  g1479 (n1484, n1155);
buf  g1480 (n1504, n1230);
buf  g1481 (n1502, n1214);
not  g1482 (n1289, n1213);
not  g1483 (n1498, n1154);
not  g1484 (n1426, n1235);
xnor g1485 (n1571, n1260, n924, n1226, n855);
xor  g1486 (n1521, n1152, n1154, n1221, n1215);
nor  g1487 (n1458, n1228, n1149, n1217, n1148);
or   g1488 (n1513, n1216, n30, n1259, n1155);
or   g1489 (n1443, n1172, n1253, n1149, n923);
xor  g1490 (n1321, n1261, n1226, n1166, n1239);
or   g1491 (n1562, n1216, n1210, n1187, n1207);
and  g1492 (n1396, n1248, n1167, n1252, n1148);
nor  g1493 (n1377, n1203, n1248, n1162, n1166);
and  g1494 (n1472, n1210, n1195, n1246, n1192);
xor  g1495 (n1355, n1179, n1168, n1176, n1206);
and  g1496 (n1423, n1196, n1205, n1207, n1223);
xnor g1497 (n1392, n1201, n29, n1209, n625);
nand g1498 (n1317, n1257, n628, n1203, n1240);
xnor g1499 (n1522, n1262, n1213, n1222, n1181);
or   g1500 (n1273, n1219, n1227, n1164, n1257);
xnor g1501 (n1358, n1153, n1249, n1250, n1247);
and  g1502 (n1365, n1158, n1190, n1188);
and  g1503 (n1322, n1258, n1155, n1246, n856);
and  g1504 (n1517, n1170, n1157, n1253, n1175);
xor  g1505 (n1315, n1251, n1197, n1252, n1227);
xor  g1506 (n1536, n1234, n1155, n1177, n1220);
xor  g1507 (n1379, n28, n1219, n1193, n1241);
or   g1508 (n1409, n1243, n1202, n31, n1212);
and  g1509 (n1541, n1257, n627, n1149, n1224);
nor  g1510 (n1344, n1172, n1159, n1204, n1163);
xnor g1511 (n1283, n1179, n1209, n1237, n1169);
and  g1512 (n1525, n855, n1243, n1217, n1208);
xor  g1513 (n1271, n1180, n1247, n1211, n31);
or   g1514 (n1534, n1152, n1249, n1224, n1150);
xor  g1515 (n1487, n1177, n1220, n1237, n1187);
and  g1516 (n1390, n1256, n1238, n1150, n1229);
or   g1517 (n1575, n1214, n1193, n186, n1232);
or   g1518 (n1488, n1190, n1240, n1262, n1216);
and  g1519 (n1418, n1164, n1161, n1156, n629);
and  g1520 (n1532, n1202, n1254, n1223, n1259);
and  g1521 (n1411, n1210, n1224, n1158, n1236);
or   g1522 (n1569, n1223, n1232, n1255, n1160);
nand g1523 (n1462, n1255, n1152, n1182, n1250);
xnor g1524 (n1427, n1218, n1196, n1215, n1195);
or   g1525 (n1297, n1211, n1234, n1226, n1179);
nand g1526 (n1366, n1148, n924, n1243, n1186);
nand g1527 (n1292, n1239, n1218, n1189, n1175);
xnor g1528 (n1505, n1248, n1164, n1262, n1245);
nand g1529 (n1540, n1166, n1236, n1245, n1176);
or   g1530 (n1389, n1154, n1231, n1169, n1222);
xnor g1531 (n1330, n1198, n1199, n1165);
xnor g1532 (n1343, n1230, n1203, n1253, n1242);
nand g1533 (n1429, n1199, n1162, n1240, n1188);
nand g1534 (n1480, n1176, n1217, n1249, n1243);
nand g1535 (n1465, n1178, n1245, n1207, n1260);
or   g1536 (n1333, n1214, n1257, n1172, n1206);
nor  g1537 (n1413, n1181, n184, n1177, n1174);
xnor g1538 (n1415, n1200, n925, n1202, n1172);
nand g1539 (n1281, n1149, n1221, n1218, n1247);
or   g1540 (n1574, n1227, n1198, n1231, n1234);
xor  g1541 (n1334, n1247, n1197, n1192, n1229);
and  g1542 (n1359, n1171, n1250, n1179, n1164);
xor  g1543 (n1277, n1201, n1161, n1237, n1156);
or   g1544 (n1268, n1161, n1184, n1188, n1151);
xnor g1545 (n1435, n1173, n185, n1249, n1148);
and  g1546 (n1269, n1207, n1169, n1241, n1229);
and  g1547 (n1316, n1230, n1256, n1187, n1165);
xor  g1548 (n1335, n1181, n1208, n1205, n1167);
buf  g1549 (n1647, n1527);
buf  g1550 (n1609, n1390);
not  g1551 (n1606, n1400);
buf  g1552 (n1598, n1439);
xor  g1553 (n1601, n1312, n1298, n1415, n1412);
nand g1554 (n1644, n1276, n1268, n1267, n1525);
xnor g1555 (n1615, n1550, n1338, n1314, n1562);
nand g1556 (n1627, n1552, n1531, n1519, n1311);
nor  g1557 (n1585, n1304, n1451, n1349, n1430);
nand g1558 (n1653, n1378, n1423, n1453, n1508);
nor  g1559 (n1628, n1334, n1345, n1364, n1470);
xnor g1560 (n1587, n1461, n1385, n1353, n1476);
and  g1561 (n1654, n1506, n1362, n1530, n1421);
xnor g1562 (n1618, n1460, n1330, n1542, n1436);
or   g1563 (n1607, n1283, n1486, n1343, n1501);
xnor g1564 (n1588, n1479, n1422, n1522, n1472);
and  g1565 (n1634, n1328, n1544, n1492, n1310);
nand g1566 (n1643, n1265, n1469, n1517, n1288);
xnor g1567 (n1636, n1358, n1316, n1271, n1555);
nor  g1568 (n1617, n1455, n1402, n1429, n1511);
xnor g1569 (n1646, n1295, n1566, n1322, n1351);
and  g1570 (n1599, n1357, n1290, n1496, n1464);
xor  g1571 (n1640, n1266, n1388, n1306, n1431);
xnor g1572 (n1611, n1485, n1286, n1404, n1493);
xnor g1573 (n1593, n1292, n1512, n1277, n1375);
nor  g1574 (n1650, n1494, n1384, n1433, n1284);
xor  g1575 (n1602, n1434, n1545, n1293, n1547);
nor  g1576 (n1660, n1406, n1294, n1326, n1373);
nor  g1577 (n1608, n1559, n1363, n1541, n1321);
xnor g1578 (n1603, n1513, n1305, n1318, n1368);
nand g1579 (n1641, n1346, n1341, n1564, n1468);
xor  g1580 (n1614, n1432, n1337, n1323, n1274);
xor  g1581 (n1651, n1269, n1481, n1457, n1380);
xor  g1582 (n1597, n1425, n1370, n1300, n1336);
xor  g1583 (n1635, n1355, n1567, n1440, n1401);
xor  g1584 (n1633, n1532, n1424, n1394, n1372);
xor  g1585 (n1655, n1483, n1543, n1369, n1320);
xnor g1586 (n1658, n1399, n1379, n1340, n1443);
nand g1587 (n1652, n1319, n1374, n1315, n1278);
xor  g1588 (n1592, n1462, n1488, n1471, n1264);
or   g1589 (n1590, n1503, n1350, n1551, n1409);
or   g1590 (n1604, n1445, n1565, n1285, n1504);
nand g1591 (n1624, n1395, n1407, n1447, n1308);
xor  g1592 (n1629, n1392, n1299, n1487, n1301);
nor  g1593 (n1616, n1507, n1520, n1495, n1497);
nand g1594 (n1659, n1414, n1490, n1556, n1523);
nand g1595 (n1594, n1441, n1307, n1427, n1417);
and  g1596 (n1625, n1563, n1475, n1448, n1291);
and  g1597 (n1648, n1324, n1333, n1500, n1325);
or   g1598 (n1642, n1477, n1482, n1289, n1459);
or   g1599 (n1600, n1529, n1515, n1389, n1317);
nand g1600 (n1630, n1474, n1332, n1365, n1270);
nor  g1601 (n1638, n1393, n1539, n1366, n1377);
nor  g1602 (n1639, n1383, n1456, n1327, n1275);
nand g1603 (n1626, n1272, n1449, n1331, n1282);
xnor g1604 (n1622, n1463, n1518, n1418, n1533);
and  g1605 (n1605, n1302, n1398, n1498, n1538);
and  g1606 (n1657, n1381, n1521, n1410, n1524);
nand g1607 (n1591, n1281, n1465, n1348, n1403);
and  g1608 (n1612, n1347, n1480, n1280, n1554);
and  g1609 (n1661, n1419, n1534, n1473, n1558);
nor  g1610 (n1584, n1557, n1467, n1450, n1526);
nand g1611 (n1619, n1478, n1397, n1489, n1367);
and  g1612 (n1649, n1413, n1499, n1386, n1505);
and  g1613 (n1645, n1510, n1303, n1502, n1491);
and  g1614 (n1621, n1454, n1458, n1335, n1438);
nand g1615 (n1631, n1428, n1391, n1411, n1553);
xor  g1616 (n1620, n1420, n1273, n1396, n1446);
xnor g1617 (n1589, n1387, n1329, n1540, n1452);
xor  g1618 (n1623, n1354, n1426, n1466, n1287);
and  g1619 (n1662, n1309, n1514, n1376, n1342);
nand g1620 (n1595, n1382, n1560, n1437, n1535);
nor  g1621 (n1610, n1405, n1561, n1537, n1548);
or   g1622 (n1632, n1361, n1371, n1536, n1296);
or   g1623 (n1586, n1344, n1444, n1360, n1484);
xnor g1624 (n1613, n1442, n1435, n1408, n1549);
nand g1625 (n1637, n1313, n1509, n1352, n1416);
and  g1626 (n1596, n1359, n1339, n1297, n1546);
xnor g1627 (n1656, n1516, n1528, n1356, n1279);
nor  g1628 (n1669, n1590, n1615, n1639, n1630);
nand g1629 (n1679, n1605, n1635, n1584, n1633);
xor  g1630 (n1663, n1622, n1625, n1610, n1599);
and  g1631 (n1671, n1614, n1598, n1640, n1629);
nand g1632 (n1673, n1604, n1612, n1613, n1592);
or   g1633 (n1676, n1650, n1607, n1593, n1602);
xnor g1634 (n1677, n1619, n1617, n1611, n1618);
xor  g1635 (n1665, n1636, n1642, n1588, n1647);
nor  g1636 (n1672, n1587, n1623, n1603, n1594);
or   g1637 (n1667, n1632, n1627, n1651, n1591);
nor  g1638 (n1668, n1626, n1638, n1637, n1597);
nor  g1639 (n1664, n1645, n1585, n1589, n1631);
and  g1640 (n1675, n1600, n1620, n1595, n1644);
xor  g1641 (n1666, n1621, n1634, n1601, n1641);
and  g1642 (n1678, n1586, n1609, n1596, n1606);
xnor g1643 (n1670, n1649, n1608, n1628, n1624);
or   g1644 (n1674, n1616, n1643, n1646, n1648);
buf  g1645 (n1684, n1665);
not  g1646 (n1680, n1664);
buf  g1647 (n1685, n1667);
not  g1648 (n1687, n1663);
not  g1649 (n1686, n1672);
buf  g1650 (n1683, n1670);
buf  g1651 (n1681, n1669);
not  g1652 (n1689, n1671);
not  g1653 (n1688, n1666);
buf  g1654 (n1682, n1668);
buf  g1655 (n1703, n633);
not  g1656 (n1717, n1688);
buf  g1657 (n1698, n645);
buf  g1658 (n1690, n634);
buf  g1659 (n1710, n1686);
buf  g1660 (n1724, n1680);
not  g1661 (n1723, n1684);
not  g1662 (n1693, n654);
buf  g1663 (n1694, n639);
not  g1664 (n1727, n667);
buf  g1665 (n1704, n1687);
not  g1666 (n1713, n635);
not  g1667 (n1695, n1683);
not  g1668 (n1696, n666);
not  g1669 (n1708, n1685);
not  g1670 (n1701, n1685);
buf  g1671 (n1721, n1684);
buf  g1672 (n1720, n657);
buf  g1673 (n1697, n1684);
buf  g1674 (n1702, n1686);
not  g1675 (n1719, n638);
not  g1676 (n1715, n1684);
not  g1677 (n1699, n1653);
not  g1678 (n1725, n1688);
xnor g1679 (n1706, n1687, n653);
and  g1680 (n1729, n662, n659);
nor  g1681 (n1712, n1678, n641, n1688, n649);
or   g1682 (n1705, n1682, n1680, n642, n1689);
or   g1683 (n1716, n644, n640, n651, n647);
xnor g1684 (n1726, n1676, n1675, n1682, n663);
xor  g1685 (n1722, n1689, n1681, n1686, n1683);
and  g1686 (n1691, n1673, n1674, n1677, n643);
xnor g1687 (n1707, n646, n1683, n1681, n660);
nand g1688 (n1728, n655, n1682, n1687);
or   g1689 (n1714, n1681, n1680, n648, n632);
nor  g1690 (n1692, n1685, n1689, n1687, n658);
or   g1691 (n1700, n1686, n1685, n650, n661);
nand g1692 (n1709, n1680, n656, n652, n1681);
xor  g1693 (n1711, n1652, n1689, n1688, n664);
xor  g1694 (n1718, n1683, n665, n637, n636);
buf  g1695 (n1740, n1722);
not  g1696 (n1755, n1699);
not  g1697 (n1831, n1704);
buf  g1698 (n1803, n1695);
buf  g1699 (n1823, n1695);
buf  g1700 (n1838, n1700);
not  g1701 (n1839, n1727);
buf  g1702 (n1786, n1715);
not  g1703 (n1781, n1712);
buf  g1704 (n1738, n1695);
buf  g1705 (n1826, n1704);
buf  g1706 (n1788, n1695);
buf  g1707 (n1867, n1706);
buf  g1708 (n1856, n1712);
not  g1709 (n1881, n1703);
not  g1710 (n1864, n1697);
not  g1711 (n1758, n1709);
not  g1712 (n1878, n1719);
buf  g1713 (n1853, n1696);
buf  g1714 (n1808, n1722);
buf  g1715 (n1733, n1690);
buf  g1716 (n1884, n1709);
not  g1717 (n1837, n1706);
buf  g1718 (n1807, n1705);
buf  g1719 (n1742, n1712);
buf  g1720 (n1730, n1718);
buf  g1721 (n1885, n1725);
buf  g1722 (n1832, n1708);
not  g1723 (n1815, n1703);
buf  g1724 (n1783, n1723);
buf  g1725 (n1756, n1706);
buf  g1726 (n1799, n1729);
buf  g1727 (n1746, n1723);
not  g1728 (n1888, n1718);
buf  g1729 (n1850, n1702);
buf  g1730 (n1735, n1728);
not  g1731 (n1879, n1694);
not  g1732 (n1858, n1699);
not  g1733 (n1772, n1702);
not  g1734 (n1882, n1710);
not  g1735 (n1745, n1713);
not  g1736 (n1886, n1707);
not  g1737 (n1834, n1691);
not  g1738 (n1845, n1708);
buf  g1739 (n1842, n1702);
not  g1740 (n1859, n1703);
buf  g1741 (n1748, n1696);
buf  g1742 (n1741, n1698);
not  g1743 (n1801, n1701);
not  g1744 (n1804, n1694);
not  g1745 (n1794, n1691);
buf  g1746 (n1795, n1707);
not  g1747 (n1734, n1716);
buf  g1748 (n1743, n1690);
not  g1749 (n1852, n1720);
buf  g1750 (n1861, n1712);
not  g1751 (n1863, n1728);
not  g1752 (n1784, n1699);
not  g1753 (n1793, n1727);
buf  g1754 (n1851, n1729);
not  g1755 (n1777, n1701);
not  g1756 (n1820, n1692);
not  g1757 (n1887, n1727);
not  g1758 (n1849, n1710);
buf  g1759 (n1822, n1692);
buf  g1760 (n1775, n1692);
not  g1761 (n1785, n1691);
not  g1762 (n1806, n1711);
not  g1763 (n1821, n1729);
not  g1764 (n1813, n1697);
not  g1765 (n1875, n1717);
not  g1766 (n1780, n1698);
not  g1767 (n1857, n1726);
buf  g1768 (n1761, n1699);
not  g1769 (n1865, n1694);
not  g1770 (n1855, n1723);
buf  g1771 (n1868, n1720);
buf  g1772 (n1848, n1698);
buf  g1773 (n1765, n1714);
buf  g1774 (n1872, n1705);
buf  g1775 (n1790, n1713);
buf  g1776 (n1869, n1718);
not  g1777 (n1854, n1711);
buf  g1778 (n1843, n1719);
not  g1779 (n1802, n1724);
not  g1780 (n1873, n1722);
buf  g1781 (n1862, n1715);
not  g1782 (n1762, n1696);
not  g1783 (n1824, n1715);
buf  g1784 (n1825, n1710);
buf  g1785 (n1744, n1726);
buf  g1786 (n1754, n1697);
not  g1787 (n1880, n1701);
buf  g1788 (n1766, n1702);
buf  g1789 (n1866, n1714);
buf  g1790 (n1796, n857);
not  g1791 (n1827, n1713);
not  g1792 (n1764, n1694);
buf  g1793 (n1809, n1728);
not  g1794 (n1776, n1724);
buf  g1795 (n1874, n1705);
not  g1796 (n1844, n1721);
buf  g1797 (n1847, n1693);
not  g1798 (n1750, n1701);
buf  g1799 (n1751, n1726);
buf  g1800 (n1816, n1700);
not  g1801 (n1774, n1691);
buf  g1802 (n1778, n1700);
not  g1803 (n1763, n1721);
not  g1804 (n1768, n1703);
buf  g1805 (n1773, n1708);
buf  g1806 (n1828, n1718);
buf  g1807 (n1759, n1693);
buf  g1808 (n1791, n1717);
not  g1809 (n1883, n1720);
not  g1810 (n1732, n1715);
buf  g1811 (n1889, n1721);
not  g1812 (n1836, n1714);
not  g1813 (n1810, n1716);
buf  g1814 (n1818, n1725);
not  g1815 (n1737, n1704);
buf  g1816 (n1792, n1711);
buf  g1817 (n1760, n1706);
not  g1818 (n1870, n1707);
not  g1819 (n1846, n1692);
not  g1820 (n1747, n1693);
not  g1821 (n1779, n1716);
not  g1822 (n1767, n1721);
buf  g1823 (n1811, n1698);
buf  g1824 (n1840, n1717);
not  g1825 (n1877, n1710);
not  g1826 (n1770, n1717);
not  g1827 (n1805, n1709);
not  g1828 (n1797, n1704);
buf  g1829 (n1833, n1700);
buf  g1830 (n1739, n1697);
not  g1831 (n1860, n1720);
not  g1832 (n1736, n1708);
not  g1833 (n1782, n1719);
not  g1834 (n1817, n1724);
not  g1835 (n1814, n1729);
not  g1836 (n1731, n1716);
not  g1837 (n1787, n1714);
not  g1838 (n1749, n1693);
not  g1839 (n1876, n1719);
buf  g1840 (n1753, n1705);
not  g1841 (n1771, n1725);
buf  g1842 (n1841, n1707);
not  g1843 (n1835, n1713);
not  g1844 (n1789, n1728);
not  g1845 (n1830, n1696);
buf  g1846 (n1769, n1725);
buf  g1847 (n1812, n1690);
not  g1848 (n1819, n1711);
not  g1849 (n1752, n1726);
buf  g1850 (n1829, n1722);
buf  g1851 (n1800, n1724);
not  g1852 (n1757, n1723);
not  g1853 (n1871, n1727);
or   g1854 (n1798, n1709, n1690);
xor  g1855 (n1977, n420, n1068);
xor  g1856 (n2004, n1041, n974);
nor  g1857 (n2389, n1785, n1777);
xnor g1858 (n2068, n1821, n348);
xnor g1859 (n2166, n1075, n1802);
nor  g1860 (n2069, n1021, n285);
nor  g1861 (n2343, n960, n935);
nor  g1862 (n1917, n1005, n1794);
xnor g1863 (n1983, n1874, n1015);
or   g1864 (n2034, n1812, n1794);
or   g1865 (n1971, n1056, n1065);
xor  g1866 (n2273, n235, n356);
nor  g1867 (n2285, n363, n1756);
xor  g1868 (n2199, n253, n952);
nor  g1869 (n2469, n1016, n312);
nor  g1870 (n2356, n1804, n1877);
nand g1871 (n2184, n1011, n1818);
nor  g1872 (n2264, n278, n1885);
xor  g1873 (n2042, n248, n1889);
xnor g1874 (n2169, n425, n1004);
xnor g1875 (n2116, n1886, n1754);
nor  g1876 (n2336, n1740, n1804);
nand g1877 (n1899, n363, n1840);
nor  g1878 (n2431, n392, n979);
or   g1879 (n2505, n432, n1817);
or   g1880 (n2339, n287, n928);
and  g1881 (n2181, n999, n382);
nor  g1882 (n1957, n432, n1058);
nor  g1883 (n2050, n949, n1010);
nor  g1884 (n2293, n211, n1737);
nand g1885 (n2299, n215, n359);
xor  g1886 (n2115, n265, n1837);
and  g1887 (n2269, n1052, n343);
or   g1888 (n1914, n1802, n256);
or   g1889 (n2525, n1831, n1810);
nand g1890 (n2032, n1869, n1842);
and  g1891 (n2151, n1850, n296);
and  g1892 (n2500, n1072, n248);
or   g1893 (n2270, n1776, n1743);
xor  g1894 (n1979, n958, n1854);
nand g1895 (n2320, n1806, n411);
xnor g1896 (n2003, n363, n1886);
and  g1897 (n2248, n219, n931);
xor  g1898 (n2242, n198, n1858);
and  g1899 (n2489, n1884, n341);
and  g1900 (n2000, n401, n205);
nor  g1901 (n2194, n403, n315);
or   g1902 (n2046, n1072, n1034);
nand g1903 (n2124, n266, n327);
and  g1904 (n2377, n1781, n266);
nand g1905 (n2476, n1829, n1767);
xnor g1906 (n2503, n978, n334);
xor  g1907 (n2102, n1837, n398);
nand g1908 (n2175, n1032, n1065);
or   g1909 (n2197, n1768, n1812);
nand g1910 (n2100, n356, n943);
xnor g1911 (n2423, n398, n194);
buf  g1912 (n1909, n286);
xnor g1913 (n2160, n930, n1038);
xor  g1914 (n2443, n972, n1795);
nor  g1915 (n2008, n249, n1028);
or   g1916 (n2494, n345, n955);
nor  g1917 (n2061, n320, n1016);
xor  g1918 (n2385, n303, n1027);
or   g1919 (n2258, n271, n325);
xor  g1920 (n2457, n1821, n1787);
xnor g1921 (n2452, n929, n1801);
nand g1922 (n2238, n435, n308);
nor  g1923 (n2453, n402, n372);
or   g1924 (n2417, n1885, n413);
nand g1925 (n2018, n313, n332);
or   g1926 (n2023, n1884, n201);
nand g1927 (n1916, n1820, n380);
nor  g1928 (n2394, n333, n1755);
xor  g1929 (n2393, n204, n228);
xnor g1930 (n1951, n299, n433);
nor  g1931 (n1941, n1730, n1881);
nand g1932 (n2435, n1819, n324);
nor  g1933 (n1986, n429, n238);
xnor g1934 (n2308, n1740, n229);
or   g1935 (n2421, n1844, n262);
xor  g1936 (n2335, n1860, n257);
xor  g1937 (n2297, n1879, n1040);
xor  g1938 (n1935, n265, n410);
xnor g1939 (n2054, n1814, n1766);
or   g1940 (n2322, n1810, n1774);
nand g1941 (n2515, n276, n1867);
xor  g1942 (n2284, n230, n394);
or   g1943 (n2463, n1014, n1738);
xor  g1944 (n2526, n942, n1882);
or   g1945 (n2304, n1878, n390);
xnor g1946 (n2055, n248, n193);
xnor g1947 (n1944, n233, n222);
nand g1948 (n2480, n197, n1843);
xor  g1949 (n2048, n1865, n321);
xnor g1950 (n2448, n254, n1853);
and  g1951 (n2117, n1801, n964);
xor  g1952 (n2404, n371, n187);
nand g1953 (n2092, n1065, n1799);
and  g1954 (n2060, n408, n1750);
xnor g1955 (n1991, n1009, n290);
xor  g1956 (n1963, n989, n965);
or   g1957 (n2047, n213, n986);
nor  g1958 (n2462, n359, n955);
xor  g1959 (n2358, n1870, n206);
and  g1960 (n2298, n1075, n405);
and  g1961 (n2075, n215, n1027);
nand g1962 (n2073, n1834, n319);
xnor g1963 (n2195, n1785, n946);
and  g1964 (n1946, n1064, n1841);
nor  g1965 (n2510, n427, n233);
xor  g1966 (n1936, n207, n950);
and  g1967 (n2130, n262, n1751);
xor  g1968 (n1985, n365, n1789);
or   g1969 (n2162, n233, n963);
xnor g1970 (n2450, n269, n1039);
xnor g1971 (n2326, n997, n337);
and  g1972 (n2342, n1856, n225);
nand g1973 (n1938, n936, n999);
and  g1974 (n2159, n367, n345);
nor  g1975 (n1960, n416, n1809);
or   g1976 (n2044, n332, n1800);
or   g1977 (n2466, n1821, n933);
xor  g1978 (n2498, n356, n1741);
nand g1979 (n2148, n370, n295);
and  g1980 (n2267, n1813, n303);
nand g1981 (n1892, n292, n1045);
and  g1982 (n2274, n1016, n289);
xnor g1983 (n2375, n237, n1039);
xor  g1984 (n2093, n329, n339);
and  g1985 (n1891, n1058, n267);
xnor g1986 (n2209, n334, n1794);
or   g1987 (n2218, n196, n1866);
and  g1988 (n1990, n1877, n251);
xnor g1989 (n2152, n326, n1869);
xnor g1990 (n2170, n239, n1021);
nor  g1991 (n2200, n419, n1806);
nor  g1992 (n2187, n231, n366);
nand g1993 (n2106, n257, n1029);
and  g1994 (n2366, n411, n352);
xnor g1995 (n2324, n1797, n322);
nor  g1996 (n2229, n967, n263);
xor  g1997 (n2286, n1888, n1841);
xnor g1998 (n2529, n281, n1059);
xor  g1999 (n2350, n236, n1737);
nand g2000 (n2312, n1836, n932);
nor  g2001 (n2316, n952, n1039);
xor  g2002 (n2268, n374, n244);
nand g2003 (n2058, n962, n1887);
or   g2004 (n2513, n294, n288);
and  g2005 (n2438, n1753, n408);
xor  g2006 (n1981, n282, n339);
xor  g2007 (n2344, n980, n305);
nor  g2008 (n2427, n1774, n1732);
and  g2009 (n2070, n268, n1815);
and  g2010 (n2460, n1812, n948);
nand g2011 (n2329, n199, n316);
xor  g2012 (n1978, n316, n377);
nand g2013 (n2137, n1788, n280);
nor  g2014 (n2294, n986, n1754);
nor  g2015 (n2487, n361, n1803, n1004, n249);
or   g2016 (n2030, n1759, n365, n286, n1843);
xnor g2017 (n2085, n1039, n402, n1015, n1868);
xor  g2018 (n2262, n1885, n970, n415, n423);
or   g2019 (n2119, n425, n1858, n1760, n421);
and  g2020 (n2190, n970, n211, n216, n292);
nor  g2021 (n2244, n276, n943, n1060, n286);
xor  g2022 (n1900, n401, n1035, n1008, n1058);
or   g2023 (n2400, n1028, n1035, n1831, n1886);
xor  g2024 (n2178, n930, n969, n1783, n939);
xor  g2025 (n2519, n236, n1052, n246, n383);
xnor g2026 (n2311, n428, n230, n934, n1782);
or   g2027 (n2120, n1839, n314, n1805, n377);
xor  g2028 (n2246, n1836, n241, n1856, n407);
or   g2029 (n2402, n361, n1054, n387, n347);
nor  g2030 (n2396, n406, n981, n1817, n1022);
or   g2031 (n2517, n1055, n408, n1749, n279);
nor  g2032 (n1923, n967, n382, n287, n321);
nor  g2033 (n2038, n366, n1770, n384, n288);
or   g2034 (n2332, n967, n982, n994, n1873);
xnor g2035 (n2094, n1791, n1756, n1796, n331);
nand g2036 (n2360, n400, n358, n234, n1842);
xor  g2037 (n2378, n1820, n282, n211, n937);
nor  g2038 (n2414, n304, n1888, n1827, n938);
and  g2039 (n2007, n341, n1847, n1785, n1012);
nor  g2040 (n2341, n365, n978, n1074, n1020);
nand g2041 (n2031, n282, n310, n995, n373);
and  g2042 (n2129, n376, n1025, n215, n367);
xnor g2043 (n2074, n988, n400, n336, n998);
or   g2044 (n2216, n323, n927, n1772, n206);
xor  g2045 (n2279, n301, n327, n339, n371);
nor  g2046 (n2521, n1865, n340, n961, n389);
or   g2047 (n2451, n931, n191, n263, n1734);
xor  g2048 (n2318, n1831, n332, n1061, n940);
nand g2049 (n1964, n288, n204, n1011, n1049);
and  g2050 (n2499, n418, n196, n295, n1006);
xor  g2051 (n2348, n993, n977, n359, n422);
nor  g2052 (n2391, n1786, n1772, n274, n1872);
nor  g2053 (n1956, n1069, n1020, n423, n362);
nand g2054 (n1931, n992, n333, n206, n937);
or   g2055 (n2002, n428, n956, n1817, n965);
nand g2056 (n2223, n1057, n1864, n1755, n1034);
nor  g2057 (n2025, n264, n247, n990);
and  g2058 (n2384, n1048, n1763, n1825, n1762);
nor  g2059 (n2006, n371, n403, n240, n311);
nand g2060 (n1933, n427, n1068, n313, n1738);
xor  g2061 (n1897, n412, n1007, n295, n337);
xnor g2062 (n1911, n1066, n338, n380, n1062);
xnor g2063 (n2493, n1021, n194, n1784, n374);
and  g2064 (n2368, n210, n357, n1766, n1848);
and  g2065 (n2024, n930, n203, n976, n1824);
nor  g2066 (n2428, n256, n208, n220, n217);
nand g2067 (n2454, n1055, n188, n1814, n935);
xor  g2068 (n2147, n1808, n1058, n1753, n291);
xnor g2069 (n1943, n966, n329, n1047, n1738);
or   g2070 (n2330, n1764, n1768, n214, n414);
xor  g2071 (n2399, n1003, n253, n319, n1811);
nor  g2072 (n2520, n193, n328, n1036, n1758);
xnor g2073 (n2020, n958, n349, n194, n1049);
or   g2074 (n2126, n335, n372, n225, n962);
nor  g2075 (n1950, n247, n1735, n261, n1042);
or   g2076 (n2084, n1053, n975, n198, n290);
or   g2077 (n1905, n1863, n1775, n418, n352);
or   g2078 (n2280, n1871, n201, n275, n1743);
nor  g2079 (n2091, n230, n1774, n431, n317);
nand g2080 (n2205, n280, n1008, n1055, n366);
or   g2081 (n2259, n386, n1846, n1741, n344);
or   g2082 (n2283, n339, n974, n396, n1811);
xnor g2083 (n2057, n1796, n292, n1068, n434);
or   g2084 (n2108, n1765, n216, n298, n407);
xnor g2085 (n2183, n953, n940, n372, n1061);
nand g2086 (n1893, n324, n949, n1044, n390);
or   g2087 (n1918, n1004, n431, n293, n1052);
xor  g2088 (n2225, n370, n349, n1014, n348);
xnor g2089 (n2219, n351, n427, n410, n1837);
and  g2090 (n2440, n221, n1051, n234, n947);
xor  g2091 (n2104, n375, n220, n358, n1059);
xor  g2092 (n1902, n1735, n323, n370, n972);
xor  g2093 (n2227, n992, n1736, n1030, n276);
nor  g2094 (n1945, n344, n1070, n1829, n429);
nand g2095 (n2412, n225, n208, n1732, n968);
xor  g2096 (n2077, n228, n203, n1027, n189);
nor  g2097 (n2028, n932, n307, n420, n259);
xor  g2098 (n2101, n254, n1833, n336, n1775);
nor  g2099 (n2482, n1806, n393, n229, n219);
or   g2100 (n2522, n324, n1798, n1072, n280);
or   g2101 (n1934, n1001, n298, n211, n1020);
xnor g2102 (n2413, n1003, n1070, n1756, n309);
nand g2103 (n2239, n359, n226, n1861, n980);
nand g2104 (n2064, n939, n267, n210, n235);
xor  g2105 (n2253, n1061, n1790, n1066, n341);
nand g2106 (n2206, n1758, n1748, n995, n299);
xnor g2107 (n2359, n203, n394, n208, n354);
xor  g2108 (n2035, n325, n273, n222, n258);
and  g2109 (n2271, n1744, n353, n966, n404);
xnor g2110 (n2191, n435, n279, n347, n255);
nand g2111 (n2523, n965, n1763, n268, n336);
nand g2112 (n1925, n237, n241, n1771, n1049);
nor  g2113 (n2107, n260, n995, n1769, n333);
nor  g2114 (n2082, n217, n1825, n1027, n196);
nor  g2115 (n1955, n936, n402, n334, n974);
nand g2116 (n2173, n239, n941, n1872, n435);
xor  g2117 (n1948, n269, n1870, n1013, n346);
nand g2118 (n2365, n369, n433, n941, n305);
nor  g2119 (n2468, n373, n310, n432, n255);
xor  g2120 (n2347, n1777, n195, n424, n369);
xor  g2121 (n1896, n926, n1063, n1031, n413);
nor  g2122 (n2153, n926, n949, n1038, n213);
xor  g2123 (n1987, n1834, n1862, n1030, n1769);
nand g2124 (n2235, n1787, n335, n1742, n1883);
nor  g2125 (n2289, n397, n985, n944, n374);
xnor g2126 (n2163, n1067, n944, n1032, n946);
xnor g2127 (n2333, n238, n1855, n1854, n1767);
xnor g2128 (n2449, n948, n957, n1850, n266);
nor  g2129 (n2252, n1816, n285, n969, n1773);
xor  g2130 (n2123, n214, n1745, n935, n1824);
nand g2131 (n1996, n1779, n1069, n1739, n1816);
or   g2132 (n2033, n1840, n213, n188, n196);
and  g2133 (n2490, n381, n212, n235, n260);
xnor g2134 (n2319, n982, n414, n224, n381);
and  g2135 (n2217, n1852, n1018, n1046, n332);
nor  g2136 (n2281, n1075, n295, n408, n218);
nor  g2137 (n2145, n424, n394, n1016, n1764);
xor  g2138 (n2478, n228, n1789, n1019, n959);
nand g2139 (n2243, n277, n1776, n1025, n407);
or   g2140 (n2346, n935, n945, n957, n205);
or   g2141 (n2247, n1855, n397, n1813, n1071);
xnor g2142 (n1907, n401, n409, n376, n256);
nand g2143 (n2370, n1848, n1059, n205, n1751);
xnor g2144 (n2171, n245, n952, n1018, n392);
and  g2145 (n2226, n1768, n207, n1010, n323);
xnor g2146 (n2097, n1760, n403, n954, n926);
or   g2147 (n2131, n1803, n341, n1875, n961);
nand g2148 (n2232, n434, n320, n981, n186);
and  g2149 (n2302, n299, n1830, n1849, n262);
and  g2150 (n2265, n425, n1773, n398, n1029);
or   g2151 (n2439, n387, n237, n1832, n1788);
nand g2152 (n2441, n1853, n1074, n1758, n1007);
or   g2153 (n2250, n1008, n240, n1751, n1047);
and  g2154 (n1966, n268, n947, n214, n291);
nor  g2155 (n2313, n999, n1786, n971, n980);
xor  g2156 (n2207, n1765, n430, n279, n1777);
or   g2157 (n1994, n1069, n975, n346, n348);
xnor g2158 (n2372, n1050, n267, n1019, n1747);
and  g2159 (n2155, n1797, n1837, n220, n360);
xnor g2160 (n2432, n1024, n1829, n197, n1878);
or   g2161 (n2354, n951, n958, n1022, n403);
and  g2162 (n2127, n1780, n310, n251, n285);
nand g2163 (n2256, n331, n1731, n223);
nand g2164 (n1895, n1752, n257, n311, n988);
nand g2165 (n1988, n1005, n1803, n326, n232);
nand g2166 (n2087, n243, n356, n1075, n1878);
xnor g2167 (n2437, n417, n319, n1753, n212);
nor  g2168 (n2338, n1781, n1827, n1013, n412);
and  g2169 (n2276, n396, n379, n936, n351);
nor  g2170 (n2374, n269, n1760, n1733, n1734);
or   g2171 (n2357, n224, n283, n1850, n1849);
xnor g2172 (n2506, n296, n1036, n391, n1043);
nand g2173 (n2049, n1060, n1848, n210, n1852);
nand g2174 (n2041, n1880, n1072, n1815, n225);
or   g2175 (n1928, n1732, n1863, n238, n413);
xor  g2176 (n2459, n424, n321, n928, n977);
and  g2177 (n2485, n1076, n292, n987, n192);
and  g2178 (n2424, n417, n344, n1748, n289);
nand g2179 (n1953, n938, n191, n274, n283);
nand g2180 (n2501, n353, n357, n1792, n987);
or   g2181 (n1904, n351, n216, n1816, n1025);
and  g2182 (n2418, n307, n932, n293, n1831);
and  g2183 (n2349, n395, n342, n1003, n1788);
nand g2184 (n2168, n249, n1057, n1011, n397);
xor  g2185 (n2484, n380, n1881, n1809, n251);
and  g2186 (n2081, n1042, n1040, n975, n979);
xnor g2187 (n2508, n270, n241, n1826, n1025);
nand g2188 (n2158, n276, n928, n323, n1739);
xor  g2189 (n2472, n384, n363, n953, n400);
or   g2190 (n2327, n1870, n288, n387, n1835);
or   g2191 (n2376, n928, n1793, n431, n217);
xnor g2192 (n2416, n202, n191, n355, n209);
xnor g2193 (n2380, n231, n1054, n1755, n1761);
xnor g2194 (n2328, n1037, n1807, n1762, n1752);
and  g2195 (n2052, n1789, n189, n377, n1818);
nor  g2196 (n2185, n1747, n404, n992, n304);
nand g2197 (n1898, n1783, n1868, n1808, n996);
nand g2198 (n2134, n1779, n1074, n972, n373);
nand g2199 (n2481, n384, n936, n1731, n1841);
xor  g2200 (n2056, n1045, n1889, n239, n1875);
xor  g2201 (n2371, n1845, n998, n380, n379);
nor  g2202 (n2213, n1073, n250, n1060, n1787);
nor  g2203 (n2110, n297, n338, n1869, n950);
and  g2204 (n1999, n1776, n970, n259, n284);
xor  g2205 (n2066, n315, n342, n1008, n368);
xor  g2206 (n2507, n1749, n308, n367, n1773);
nand g2207 (n2410, n349, n1067, n1010, n1062);
and  g2208 (n2063, n1005, n1042, n1800, n1820);
xnor g2209 (n2111, n266, n382, n192, n942);
xor  g2210 (n2470, n1048, n1003, n1037, n221);
or   g2211 (n2233, n1748, n1859, n309, n1033);
xnor g2212 (n2121, n429, n1882, n430, n1822);
xnor g2213 (n2383, n1833, n410, n1860, n1853);
nor  g2214 (n2078, n326, n1069, n1009, n192);
xor  g2215 (n1959, n360, n1784, n1877, n1026);
nand g2216 (n2221, n273, n950, n1733, n1846);
and  g2217 (n2364, n1055, n325, n1041, n1015);
and  g2218 (n2495, n216, n1795, n424, n1051);
nand g2219 (n1937, n976, n308, n261, n995);
or   g2220 (n2408, n328, n1029, n1774, n261);
and  g2221 (n2420, n434, n250, n1074, n207);
nand g2222 (n2296, n971, n241, n245, n346);
xnor g2223 (n2231, n1879, n957, n385, n963);
nor  g2224 (n1930, n1819, n991, n197, n1888);
xnor g2225 (n1913, n1784, n1045, n1031, n970);
nand g2226 (n2351, n1754, n265, n1791, n1076);
xor  g2227 (n2133, n430, n1810, n243, n272);
nand g2228 (n2465, n1030, n1866, n1863, n187);
xnor g2229 (n2405, n1786, n381, n1828, n227);
and  g2230 (n2401, n1880, n284, n253, n1868);
xnor g2231 (n2202, n1867, n1000, n1799, n1840);
nor  g2232 (n2369, n1813, n326, n190, n300);
xnor g2233 (n2222, n388, n318, n316, n1743);
nand g2234 (n2300, n376, n396, n975, n242);
xnor g2235 (n2086, n252, n409, n964, n378);
nor  g2236 (n2203, n419, n965, n252, n351);
xnor g2237 (n2340, n1830, n272, n1036, n1771);
xor  g2238 (n2180, n939, n313, n1740, n1879);
xnor g2239 (n2136, n973, n939, n1833, n1014);
or   g2240 (n2367, n1809, n229, n245, n1062);
or   g2241 (n2288, n328, n379, n1778, n240);
or   g2242 (n1921, n364, n978, n203, n938);
and  g2243 (n2198, n189, n309, n962, n1787);
or   g2244 (n2036, n230, n1839, n388, n406);
and  g2245 (n2090, n312, n982, n930, n239);
nor  g2246 (n2255, n338, n404, n961, n980);
or   g2247 (n2483, n1766, n983, n297, n1857);
xnor g2248 (n2511, n934, n270, n1859, n1040);
and  g2249 (n2021, n385, n343, n960, n317);
or   g2250 (n2037, n940, n245, n316, n1758);
xor  g2251 (n2492, n1045, n985, n969, n1741);
or   g2252 (n1998, n317, n345, n375, n1790);
and  g2253 (n2305, n354, n415, n1736, n945);
xor  g2254 (n2390, n234, n430, n261, n391);
and  g2255 (n2310, n1864, n1011, n1867, n300);
xnor g2256 (n2177, n944, n1007, n416, n1800);
and  g2257 (n2188, n1791, n1886, n1746, n336);
xnor g2258 (n2122, n1848, n238, n1744, n1808);
xor  g2259 (n2355, n340, n347, n1828, n1004);
nor  g2260 (n2398, n1836, n1057, n1864, n229);
and  g2261 (n2409, n389, n1878, n1869, n294);
or   g2262 (n2352, n1851, n1760, n1766, n278);
nand g2263 (n2109, n422, n1856, n1073, n357);
nor  g2264 (n2415, n388, n1740, n417, n1013);
nor  g2265 (n2512, n932, n994, n284, n950);
nand g2266 (n2446, n419, n415, n426, n300);
xnor g2267 (n2154, n315, n399, n1826, n215);
nor  g2268 (n2105, n1023, n1822, n1797, n1024);
nor  g2269 (n1912, n1030, n369, n236, n350);
xnor g2270 (n2257, n287, n294, n1019, n1773);
nand g2271 (n2228, n1071, n979, n399, n418);
xnor g2272 (n1989, n1866, n963, n1881, n959);
nor  g2273 (n1942, n318, n382, n1012, n426);
nand g2274 (n2099, n222, n991, n259, n1805);
nor  g2275 (n1940, n262, n264, n416, n951);
or   g2276 (n2471, n1847, n344, n1053, n1761);
xor  g2277 (n1993, n1052, n273, n429, n1739);
nand g2278 (n2240, n997, n1862, n1046, n223);
nand g2279 (n2301, n289, n378, n1806, n277);
nor  g2280 (n1972, n218, n1071, n985, n1026);
nor  g2281 (n1903, n376, n1744, n1044, n1776);
xnor g2282 (n2143, n1051, n1859, n1847, n281);
nand g2283 (n2164, n954, n307, n416, n1037);
nand g2284 (n2208, n1064, n374, n391, n1851);
xnor g2285 (n2071, n973, n249, n360, n320);
or   g2286 (n2045, n435, n1762, n219, n953);
xor  g2287 (n2516, n330, n951, n390, n1813);
xnor g2288 (n2027, n1026, n396, n1844, n1843);
and  g2289 (n2179, n1819, n1733, n957, n361);
xor  g2290 (n2275, n350, n1822, n246, n1750);
nand g2291 (n2473, n256, n335, n224, n1764);
and  g2292 (n2089, n1064, n1876, n1849, n1877);
xnor g2293 (n2434, n1874, n988, n1836, n265);
and  g2294 (n2072, n242, n937, n954, n927);
and  g2295 (n2303, n194, n1873, n1876, n201);
xor  g2296 (n2017, n1889, n1882, n1043, n1796);
nand g2297 (n2112, n1034, n273, n1000, n1875);
nand g2298 (n1920, n934, n303, n221, n1815);
xor  g2299 (n1958, n1017, n306, n1792, n302);
xnor g2300 (n2514, n1012, n1038, n270, n983);
xor  g2301 (n1962, n1054, n417, n938, n1889);
nand g2302 (n2386, n240, n192, n1757, n324);
xnor g2303 (n2059, n948, n294, n189, n258);
and  g2304 (n2426, n318, n973, n322, n381);
xnor g2305 (n1968, n1046, n212, n1876);
or   g2306 (n2149, n204, n946, n253, n956);
xnor g2307 (n2456, n362, n298, n960, n325);
nand g2308 (n2096, n941, n1022, n927, n1803);
nand g2309 (n1929, n343, n428, n1819, n243);
nor  g2310 (n2079, n978, n355, n1747, n327);
or   g2311 (n2156, n972, n302, n1825, n1735);
and  g2312 (n2406, n303, n1054, n1770, n1845);
or   g2313 (n2039, n338, n961, n1804, n1043);
nor  g2314 (n2395, n313, n1786, n976, n187);
nand g2315 (n1915, n969, n394, n1832, n1846);
xnor g2316 (n2323, n1769, n1747, n1845, n1820);
and  g2317 (n2182, n1017, n971, n1736, n277);
xor  g2318 (n2114, n1756, n994, n195, n304);
xnor g2319 (n2509, n422, n984, n1032, n198);
or   g2320 (n2411, n352, n1761, n297, n202);
xnor g2321 (n2295, n1009, n218, n254, n1028);
xnor g2322 (n2014, n1732, n1012, n1823, n966);
nor  g2323 (n2214, n929, n385, n1779, n1031);
or   g2324 (n2140, n1838, n991, n255, n1070);
or   g2325 (n2419, n274, n1887, n1737, n1818);
xnor g2326 (n2118, n1730, n377, n191, n235);
nor  g2327 (n2132, n1790, n1858, n287, n312);
and  g2328 (n2236, n353, n228, n1029, n309);
or   g2329 (n2309, n1033, n953, n405, n348);
xor  g2330 (n2026, n252, n1015, n1812, n1006);
xor  g2331 (n2353, n222, n368, n1017, n233);
nand g2332 (n2455, n283, n384, n433, n219);
xor  g2333 (n1984, n940, n1024, n368, n226);
or   g2334 (n2436, n1739, n322, n277, n1781);
nand g2335 (n1973, n350, n1750, n989, n1057);
or   g2336 (n2249, n1844, n1834, n297, n247);
nor  g2337 (n1975, n1792, n193, n955, n291);
and  g2338 (n2497, n1799, n1838, n1048, n268);
and  g2339 (n2263, n1000, n1020, n1021, n1802);
nand g2340 (n2266, n1041, n1009, n943, n1763);
xor  g2341 (n2425, n1784, n982, n929, n355);
and  g2342 (n2144, n1807, n1801, n1823, n989);
xor  g2343 (n1995, n955, n1797, n1883, n1865);
or   g2344 (n1969, n346, n199, n244, n941);
xnor g2345 (n2290, n200, n1808, n1782, n1041);
and  g2346 (n2461, n990, n398, n1063, n311);
and  g2347 (n2224, n1871, n1031, n1857, n406);
xor  g2348 (n2019, n1826, n1853, n411, n281);
xnor g2349 (n1927, n984, n1750, n1793, n1849);
or   g2350 (n2076, n985, n399, n964, n275);
nand g2351 (n2321, n959, n1842, n956, n393);
nand g2352 (n2382, n1802, n996, n232, n259);
xnor g2353 (n2488, n232, n1778, n1798, n379);
and  g2354 (n2015, n1752, n1066, n428, n260);
and  g2355 (n2362, n296, n237, n301, n395);
xnor g2356 (n2527, n1000, n188, n284, n388);
xor  g2357 (n2292, n958, n314, n1885, n1014);
xor  g2358 (n2245, n1862, n231, n1046, n1754);
xnor g2359 (n2065, n227, n202, n945, n1746);
xor  g2360 (n1924, n1745, n1734, n272, n1006);
nand g2361 (n2524, n218, n1851, n1033, n1864);
xnor g2362 (n2165, n1862, n365, n421, n283);
xor  g2363 (n2477, n1731, n371, n255, n200);
and  g2364 (n2486, n1047, n426, n405, n1805);
nand g2365 (n2306, n1883, n1823, n1005, n1830);
nand g2366 (n2407, n1861, n1076, n1835, n1770);
xor  g2367 (n2083, n386, n1824, n929, n358);
nor  g2368 (n1976, n373, n314, n409, n195);
xor  g2369 (n2397, n1731, n1860, n1730, n1018);
xnor g2370 (n1949, n349, n944, n1733, n1859);
and  g2371 (n2138, n369, n407, n1793, n1870);
nor  g2372 (n2186, n1828, n258, n945, n300);
xor  g2373 (n2325, n299, n1789, n340, n1050);
or   g2374 (n2334, n393, n433, n937, n959);
nand g2375 (n1906, n426, n1073, n281, n264);
and  g2376 (n2422, n278, n193, n402, n1730);
xor  g2377 (n1919, n1800, n1761, n290, n220);
xor  g2378 (n2445, n1804, n250, n933, n1825);
xnor g2379 (n2315, n1883, n420, n1860, n367);
or   g2380 (n2210, n1060, n1827, n378, n1037);
nor  g2381 (n2043, n1763, n306, n1023, n1811);
nand g2382 (n2189, n414, n1028, n1858, n421);
nor  g2383 (n2009, n1844, n977, n986, n293);
xor  g2384 (n2067, n1066, n199, n1884, n1805);
or   g2385 (n2150, n224, n347, n1777, n1769);
xnor g2386 (n2403, n1866, n1751, n293, n977);
or   g2387 (n2282, n1051, n942, n260, n307);
nand g2388 (n2363, n1830, n996, n967, n984);
or   g2389 (n2040, n411, n1001, n226, n1875);
nor  g2390 (n2291, n370, n1815, n1002, n223);
or   g2391 (n2230, n305, n1044, n1064, n318);
nand g2392 (n2167, n1017, n998, n1887, n217);
nor  g2393 (n2502, n258, n227, n1001, n1863);
or   g2394 (n2211, n209, n1771, n386, n1026);
and  g2395 (n2234, n423, n280, n291, n267);
and  g2396 (n2001, n1795, n933, n1792, n1854);
xor  g2397 (n2193, n1861, n1043, n310, n976);
or   g2398 (n2128, n306, n200, n1822, n1764);
or   g2399 (n2204, n199, n1050, n1779, n1793);
and  g2400 (n2528, n395, n1780, n964, n427);
and  g2401 (n2172, n412, n234, n1799, n1850);
or   g2402 (n2212, n1888, n1824, n420, n337);
or   g2403 (n2379, n329, n1042, n431, n406);
nor  g2404 (n2174, n1065, n1735, n1872, n333);
xnor g2405 (n2496, n949, n414, n1742, n1807);
nand g2406 (n2135, n298, n209, n1833, n335);
nand g2407 (n2287, n963, n1745, n1749, n1801);
nor  g2408 (n2125, n1023, n1855, n190, n257);
nor  g2409 (n2012, n1036, n1832, n1845, n275);
xor  g2410 (n1947, n1818, n312, n1038, n1807);
xnor g2411 (n2113, n272, n1798, n1067, n1778);
nand g2412 (n1952, n1782, n1049, n254, n1835);
xor  g2413 (n2277, n354, n971, n1781, n360);
xnor g2414 (n2491, n404, n1076, n1834, n421);
and  g2415 (n2272, n1048, n1050, n1880, n400);
xnor g2416 (n2010, n282, n1782, n247, n405);
or   g2417 (n2088, n343, n1842, n979, n271);
or   g2418 (n1965, n205, n954, n308, n1846);
xor  g2419 (n1980, n1024, n948, n200, n947);
and  g2420 (n1954, n1852, n246, n943, n375);
xor  g2421 (n1908, n226, n248, n1798, n311);
xor  g2422 (n2458, n993, n1018, n992, n342);
nor  g2423 (n2254, n1772, n1851, n1001, n1748);
xor  g2424 (n2381, n1062, n1757, n1783, n1775);
nor  g2425 (n2429, n1828, n422, n960, n973);
nand g2426 (n1922, n1746, n250, n1752, n981);
and  g2427 (n2307, n1838, n933, n434, n1767);
or   g2428 (n2011, n1882, n1829, n1840, n1791);
xor  g2429 (n1982, n197, n232, n210, n352);
nand g2430 (n1967, n1881, n1871, n993, n296);
nor  g2431 (n2016, n368, n983, n425, n264);
and  g2432 (n2141, n1887, n195, n386, n212);
xnor g2433 (n2215, n342, n1814, n987, n327);
xor  g2434 (n2261, n1059, n1838, n931, n1827);
nor  g2435 (n2080, n246, n1022, n302, n947);
xor  g2436 (n2251, n202, n1865, n331, n989);
xnor g2437 (n2388, n1809, n270, n227, n934);
or   g2438 (n2314, n1757, n1071, n358, n330);
and  g2439 (n2518, n1070, n1067, n1006, n187);
nand g2440 (n2192, n301, n383, n1795, n997);
or   g2441 (n2467, n271, n1047, n1068, n263);
xnor g2442 (n2142, n279, n1821, n1856, n1749);
nand g2443 (n2474, n418, n337, n1768, n387);
or   g2444 (n2345, n987, n243, n314, n1759);
xnor g2445 (n2095, n389, n271, n1737, n1884);
and  g2446 (n2161, n1736, n1783, n1044, n345);
xor  g2447 (n2201, n236, n415, n1839, n1007);
nor  g2448 (n2220, n198, n419, n927, n1857);
nor  g2449 (n1961, n1033, n364, n1040, n1002);
xor  g2450 (n2331, n962, n375, n354, n1810);
xor  g2451 (n2479, n231, n275, n242, n320);
nor  g2452 (n1992, n263, n244, n1778, n362);
nor  g2453 (n2433, n1794, n290, n317, n364);
xnor g2454 (n1926, n1790, n1879, n244, n1873);
or   g2455 (n2146, n1738, n357, n432, n355);
xnor g2456 (n2029, n998, n1023, n1871, n1832);
nand g2457 (n1970, n331, n285, n1061, n1734);
nand g2458 (n2241, n322, n999, n956, n1745);
xor  g2459 (n2013, n221, n984, n1753, n350);
nor  g2460 (n2278, n353, n214, n207, n1056);
nor  g2461 (n2475, n397, n1002, n306, n1757);
and  g2462 (n2464, n395, n362, n1874, n1785);
nor  g2463 (n2447, n278, n1770, n330, n378);
nand g2464 (n2444, n1762, n1855, n1002, n289);
or   g2465 (n2051, n401, n1013, n206, n994);
xor  g2466 (n1997, n968, n1765, n1775, n413);
xnor g2467 (n2139, n423, n340, n1857, n213);
nor  g2468 (n2387, n302, n361, n931, n242);
xor  g2469 (n2237, n1767, n1868, n1032, n1814);
nand g2470 (n2442, n392, n968, n1035, n990);
xnor g2471 (n2373, n330, n269, n1743, n305);
and  g2472 (n1932, n1771, n1874, n1861, n991);
xnor g2473 (n2053, n1788, n1835, n1843, n372);
or   g2474 (n1894, n1035, n983, n1073, n1817);
xor  g2475 (n2157, n993, n1765, n329, n1880);
and  g2476 (n2005, n389, n321, n1034, n1796);
xor  g2477 (n1890, n1816, n190, n1019, n1053);
xor  g2478 (n1910, n1867, n1780, n390, n274);
and  g2479 (n2337, n1759, n383, n1056, n1063);
nand g2480 (n2196, n208, n1873, n1741, n190);
and  g2481 (n2098, n366, n946, n1010, n942);
xor  g2482 (n2260, n399, n981, n204, n393);
nor  g2483 (n2504, n412, n996, n1780, n1755);
nor  g2484 (n1974, n409, n1053, n1742, n966);
and  g2485 (n2317, n328, n1847, n1746, n986);
xnor g2486 (n2103, n315, n951, n391, n1841);
xnor g2487 (n2392, n952, n1063, n410, n334);
xnor g2488 (n2022, n188, n1744, n383, n301);
nand g2489 (n1901, n385, n201, n252, n1826);
nor  g2490 (n2361, n209, n974, n364, n319);
nand g2491 (n2430, n997, n1742, n1872, n1852);
nor  g2492 (n2176, n1854, n1056, n1839, n1811);
xor  g2493 (n2062, n968, n304, n1823, n988);
nor  g2494 (n1939, n251, n392, n1759, n1772);
buf  g2495 (n2532, n2123);
buf  g2496 (n2612, n2258);
not  g2497 (n2560, n2211);
not  g2498 (n2541, n1977);
buf  g2499 (n2602, n2172);
not  g2500 (n2540, n2219);
not  g2501 (n2614, n1892);
or   g2502 (n2536, n2216, n2054);
nor  g2503 (n2551, n2114, n1955);
xnor g2504 (n2623, n2221, n2161);
or   g2505 (n2553, n2136, n2226, n2225);
or   g2506 (n2580, n2174, n2068, n1931, n2128);
xor  g2507 (n2628, n2141, n2087, n2235, n2013);
nor  g2508 (n2609, n2231, n2150, n2177, n1909);
xor  g2509 (n2533, n2155, n1997, n1959, n1976);
xnor g2510 (n2573, n2127, n2096, n2003, n2086);
or   g2511 (n2557, n2180, n2168, n1895, n2001);
xnor g2512 (n2547, n1994, n2183, n2027, n2237);
xnor g2513 (n2537, n2021, n2039, n2101, n1966);
xnor g2514 (n2606, n2181, n2018, n1915, n2124);
xor  g2515 (n2554, n1921, n2089, n1951, n2167);
nand g2516 (n2579, n2256, n1928, n2153, n1942);
nand g2517 (n2627, n2132, n2241, n2075, n1923);
xnor g2518 (n2577, n1963, n1904, n2073, n2193);
nand g2519 (n2564, n2061, n2196, n2179, n2232);
nand g2520 (n2535, n1933, n2159, n2148, n2255);
and  g2521 (n2556, n1988, n1967, n2130, n2240);
nor  g2522 (n2578, n2163, n2043, n2175, n2047);
nor  g2523 (n2566, n2212, n2137, n2229, n2165);
xor  g2524 (n2552, n1938, n2045, n2065, n2066);
and  g2525 (n2588, n2113, n1956, n1952, n1919);
or   g2526 (n2575, n2209, n2012, n2007, n2233);
nor  g2527 (n2561, n2058, n2122, n2037, n1910);
xor  g2528 (n2576, n2104, n2187, n2088, n1953);
and  g2529 (n2605, n2000, n1930, n1939, n2252);
xor  g2530 (n2545, n1890, n2204, n2248, n2035);
nand g2531 (n2574, n1949, n2217, n2200, n2227);
or   g2532 (n2617, n1929, n2042, n2249, n2195);
and  g2533 (n2546, n2059, n1926, n1984, n2169);
and  g2534 (n2589, n2069, n2213, n1999, n1993);
nand g2535 (n2583, n2092, n2011, n2030, n2090);
and  g2536 (n2597, n2034, n2071, n1987, n2245);
nand g2537 (n2601, n1960, n2072, n2103, n1990);
xor  g2538 (n2585, n1918, n2120, n1970, n2236);
nor  g2539 (n2549, n2015, n2033, n2182, n1980);
nor  g2540 (n2613, n1957, n2253, n2055, n2185);
nor  g2541 (n2600, n2040, n1981, n2057, n2228);
xor  g2542 (n2563, n1911, n2144, n2025, n2139);
xnor g2543 (n2569, n1900, n2108, n2170, n1925);
xor  g2544 (n2610, n2224, n2052, n2080, n2017);
xnor g2545 (n2570, n1934, n2105, n2234, n2138);
and  g2546 (n2587, n1944, n2184, n2145, n2063);
and  g2547 (n2544, n2186, n1924, n1896, n1917);
xor  g2548 (n2548, n1947, n2154, n2238, n1991);
nand g2549 (n2599, n2205, n2051, n2134, n1979);
nand g2550 (n2567, n1948, n1983, n2215, n1907);
and  g2551 (n2562, n2243, n1962, n2084, n2041);
xnor g2552 (n2571, n2083, n2020, n1901, n2214);
xor  g2553 (n2598, n2261, n1954, n1995, n1998);
xor  g2554 (n2539, n2060, n2106, n2147, n2028);
or   g2555 (n2584, n1898, n2121, n2085, n2110);
xnor g2556 (n2572, n2143, n1906, n2070, n2109);
xnor g2557 (n2555, n2010, n2005, n1908, n2115);
xor  g2558 (n2543, n1973, n2014, n2244, n2016);
xor  g2559 (n2582, n1958, n2220, n2146, n2162);
xor  g2560 (n2590, n2230, n1932, n1946, n2254);
nand g2561 (n2620, n2223, n2188, n2078, n2242);
or   g2562 (n2592, n1945, n2160, n1961, n2076);
xnor g2563 (n2534, n2157, n2156, n1943, n1996);
nor  g2564 (n2625, n2201, n2111, n2257, n2062);
xnor g2565 (n2568, n2032, n2094, n1975, n2194);
or   g2566 (n2619, n1971, n2202, n2191, n1920);
nand g2567 (n2530, n2119, n2079, n2091, n2189);
and  g2568 (n2607, n2117, n2097, n2098, n2158);
nand g2569 (n2595, n2250, n1986, n2081, n1985);
nand g2570 (n2581, n1912, n2029, n2151, n1902);
xnor g2571 (n2622, n2024, n2259, n2178, n1982);
xor  g2572 (n2550, n2152, n2023, n2207, n2046);
or   g2573 (n2626, n1922, n2192, n1940, n1894);
nor  g2574 (n2591, n1964, n2036, n2074, n2239);
xnor g2575 (n2624, n2056, n2002, n2133, n1897);
nand g2576 (n2565, n2198, n2142, n1905, n1935);
xnor g2577 (n2559, n1891, n2210, n2019, n2116);
xor  g2578 (n2603, n2208, n2164, n2260, n2206);
or   g2579 (n2629, n2218, n2140, n2093, n2006);
and  g2580 (n2558, n2067, n1969, n1893, n2118);
nand g2581 (n2611, n1899, n2149, n1914, n1972);
xnor g2582 (n2596, n2026, n1950, n1913, n2099);
and  g2583 (n2593, n2064, n2199, n2222, n2008);
xnor g2584 (n2604, n1968, n2049, n2166, n2171);
and  g2585 (n2608, n2004, n1937, n2131, n1936);
xnor g2586 (n2616, n1965, n1992, n2100, n1974);
or   g2587 (n2615, n2203, n2053, n2126, n2102);
nor  g2588 (n2586, n2135, n2190, n2050, n2095);
nand g2589 (n2531, n2031, n2044, n1941, n1989);
xor  g2590 (n2594, n2038, n2107, n1916, n2197);
nor  g2591 (n2542, n2009, n2022, n1903, n2048);
xnor g2592 (n2538, n2082, n1978, n2247, n2129);
xnor g2593 (n2618, n2112, n2176, n2251, n2246);
nor  g2594 (n2621, n2173, n1927, n2125, n2077);
nand g2595 (n2671, n2450, n2324, n2565, n2505);
xnor g2596 (n2680, n2592, n2358, n2364, n2521);
xor  g2597 (n2677, n2319, n2275, n2294, n2608);
or   g2598 (n2716, n2352, n2499, n2515, n2425);
nand g2599 (n2664, n2471, n2412, n2318, n2363);
nor  g2600 (n2714, n2397, n2479, n2292, n2287);
xnor g2601 (n2687, n2357, n2390, n2582, n2487);
nand g2602 (n2682, n2596, n2386, n2269, n2299);
xnor g2603 (n2659, n2456, n2559, n2551, n2411);
xnor g2604 (n2652, n2288, n2463, n2580, n2326);
and  g2605 (n2654, n2430, n2401, n2446, n2372);
nand g2606 (n2662, n2282, n2306, n2316, n2609);
xnor g2607 (n2670, n2460, n2360, n2455, n2549);
nor  g2608 (n2695, n2304, n2402, n2297, n2272);
nand g2609 (n2689, n2381, n2398, n2369, n2296);
xnor g2610 (n2685, n2518, n2510, n2418, n2492);
and  g2611 (n2713, n2268, n2554, n2420, n2616);
nand g2612 (n2694, n2498, n2553, n2507, n2391);
xor  g2613 (n2701, n2368, n2452, n2464, n2415);
xnor g2614 (n2640, n2388, n2396, n2544, n2522);
nand g2615 (n2678, n2338, n2378, n2373, n2508);
xor  g2616 (n2681, n2395, n2434, n2447, n2345);
and  g2617 (n2704, n2439, n2307, n2278, n2591);
and  g2618 (n2693, n2265, n2454, n2387, n2585);
and  g2619 (n2651, n2558, n2552, n2440, n2475);
and  g2620 (n2691, n2286, n2313, n2444, n2370);
xnor g2621 (n2641, n2276, n2274, n2422, n2538);
xor  g2622 (n2702, n2469, n2614, n2496, n2462);
or   g2623 (n2633, n2600, n2542, n2445, n2467);
and  g2624 (n2698, n2590, n2548, n2604, n2302);
xnor g2625 (n2692, n2281, n2605, n2533, n2556);
nand g2626 (n2655, n2485, n2394, n2470, n2343);
or   g2627 (n2660, n2502, n2607, n2303, n2419);
xnor g2628 (n2658, n2362, n2566, n2405, n2305);
xnor g2629 (n2648, n2375, n2428, n2380, n2482);
xor  g2630 (n2674, n2298, n2442, n2431, n2271);
xor  g2631 (n2647, n2356, n2555, n2325, n2584);
nand g2632 (n2634, n2270, n2277, n2513, n2483);
nor  g2633 (n2631, n2512, n2432, n2484, n2459);
and  g2634 (n2637, n2443, n2427, n2474, n2423);
xnor g2635 (n2683, n2346, n2535, n2441, n2476);
and  g2636 (n2668, n2611, n2490, n2290, n2336);
xor  g2637 (n2696, n2494, n2416, n2595, n2574);
or   g2638 (n2646, n2263, n2300, n2393, n2572);
and  g2639 (n2703, n2497, n2301, n2333, n2589);
xor  g2640 (n2669, n2573, n2530, n2337, n2560);
nand g2641 (n2663, n2328, n2340, n2339, n2361);
or   g2642 (n2643, n2561, n2291, n2517, n2355);
nor  g2643 (n2710, n2504, n2531, n2568, n2540);
xor  g2644 (n2688, n2283, n2327, n2501, n2519);
nor  g2645 (n2706, n2576, n2465, n2365, n2403);
xnor g2646 (n2656, n2543, n2341, n2266, n2334);
nand g2647 (n2630, n2457, n2366, n2400, n2408);
or   g2648 (n2642, n2367, n2516, n2478, n2262);
and  g2649 (n2709, n2347, n2541, n2433, n2267);
or   g2650 (n2673, n2308, n2311, n2448, n2389);
nor  g2651 (n2707, n2610, n2312, n2613, n2486);
nor  g2652 (n2636, n2284, n2488, n2451, n2532);
xnor g2653 (n2705, n2379, n2514, n2606, n2315);
or   g2654 (n2672, n2310, n2578, n2468, n2399);
nor  g2655 (n2632, n2285, n2453, n2493, n2371);
and  g2656 (n2635, n2342, n2438, n2537, n2279);
or   g2657 (n2712, n2567, n2314, n2376, n2598);
xnor g2658 (n2699, n2579, n2571, n2330, n2557);
nor  g2659 (n2686, n2500, n2383, n2534, n2382);
xnor g2660 (n2653, n2449, n2594, n2520, n2349);
nand g2661 (n2650, n2351, n2295, n2458, n2406);
nor  g2662 (n2700, n2385, n2563, n2593, n2583);
and  g2663 (n2639, n2581, n2417, n2359, n2350);
nor  g2664 (n2675, n2413, n2570, n2481, n2569);
nand g2665 (n2649, n2436, n2587, n2321, n2404);
xnor g2666 (n2708, n2472, n2599, n2564, n2562);
or   g2667 (n2638, n2601, n2575, n2421, n2506);
or   g2668 (n2711, n2409, n2545, n2491, n2603);
xnor g2669 (n2661, n2480, n2602, n2437, n2414);
xor  g2670 (n2684, n2329, n2509, n2473, n2615);
xor  g2671 (n2690, n2461, n2495, n2377, n2597);
and  g2672 (n2697, n2384, n2322, n2353, n2424);
or   g2673 (n2644, n2503, n2588, n2547, n2550);
or   g2674 (n2679, n2335, n2466, n2344, n2280);
nor  g2675 (n2676, n2332, n2331, n2577, n2392);
nand g2676 (n2665, n2293, n2323, n2320, n2536);
xor  g2677 (n2645, n2317, n2309, n2348, n2429);
and  g2678 (n2666, n2426, n2612, n2374, n2489);
nand g2679 (n2657, n2289, n2546, n2407, n2586);
nor  g2680 (n2715, n2477, n2539, n2410, n2435);
nor  g2681 (n2667, n2511, n2264, n2354, n2273);
not  g2682 (n2722, n2655);
buf  g2683 (n2717, n2661);
buf  g2684 (n2727, n2673);
not  g2685 (n2732, n2670);
buf  g2686 (n2741, n2649);
not  g2687 (n2726, n2641);
not  g2688 (n2729, n2679);
not  g2689 (n2718, n2667);
buf  g2690 (n2730, n2639);
not  g2691 (n2724, n2632);
buf  g2692 (n2721, n2648);
not  g2693 (n2739, n2650);
not  g2694 (n2735, n2663);
buf  g2695 (n2731, n2645);
not  g2696 (n2728, n2631);
not  g2697 (n2734, n2664);
nand g2698 (n2738, n2656, n2642);
or   g2699 (n2723, n2644, n2677, n2630, n2660);
or   g2700 (n2733, n2646, n2666, n2640, n2671);
and  g2701 (n2737, n2635, n2643, n2668, n2647);
nand g2702 (n2720, n2675, n2651, n2658, n2653);
xnor g2703 (n2740, n2662, n2636, n2674, n2654);
nand g2704 (n2725, n2665, n2657, n2637, n2634);
nand g2705 (n2736, n2672, n2652, n2633, n2669);
xnor g2706 (n2719, n2659, n2678, n2676, n2638);
xor  g2707 (n2742, n2717, n2683, n2691, n2689);
nor  g2708 (n2743, n2687, n2686, n2719, n2684);
or   g2709 (n2745, n2685, n2682, n2720, n2688);
nand g2710 (n2744, n2680, n2690, n2681, n2718);
buf  g2711 (n2746, n2742);
buf  g2712 (n2747, n2743);
or   g2713 (n2752, n1658, n2747, n1656);
nand g2714 (n2748, n1661, n2747, n1657);
and  g2715 (n2750, n2692, n2746, n1659);
nor  g2716 (n2751, n1662, n2744, n1654);
xnor g2717 (n2749, n1660, n2747, n1655);
not  g2718 (n2757, n2750);
buf  g2719 (n2754, n2749);
buf  g2720 (n2755, n2752);
buf  g2721 (n2756, n2751);
buf  g2722 (n2753, n2748);
or   g2723 (n2758, n2753, n1679);
and  g2724 (n2762, n33, n2758, n32);
and  g2725 (n2759, n33, n2758, n34);
nand g2726 (n2760, n32, n34);
or   g2727 (n2761, n33, n33, n32, n2758);
xor  g2728 (n2765, n117, n2759, n115, n2762);
xnor g2729 (n2766, n116, n117, n2761);
xor  g2730 (n2764, n116, n115, n118);
nor  g2731 (n2763, n115, n2762, n116, n2760);
or   g2732 (n2767, n118, n116, n115, n117);
not  g2733 (n2768, n2764);
and  g2734 (n2769, n2763, n436);
buf  g2735 (n2771, n2768);
not  g2736 (n2770, n2769);
not  g2737 (n2774, n2771);
not  g2738 (n2772, n2771);
not  g2739 (n2775, n2771);
not  g2740 (n2773, n2771);
buf  g2741 (n2779, n2773);
not  g2742 (n2778, n2774);
buf  g2743 (n2776, n2775);
nor  g2744 (n2777, n2772, n1077);
nor  g2745 (n2795, n2721, n2779, n2700, n2526);
and  g2746 (n2784, n2731, n2702, n2732, n2778);
nand g2747 (n2788, n2736, n2726, n2527, n2767);
xor  g2748 (n2789, n2524, n2696, n2523, n2727);
nand g2749 (n2793, n2703, n2707, n2765, n2778);
nand g2750 (n2780, n2778, n2695, n2741, n2724);
or   g2751 (n2787, n2722, n2735, n2733, n2698);
and  g2752 (n2794, n2728, n2699, n2740, n2697);
xnor g2753 (n2792, n2766, n2779, n2529, n2739);
xnor g2754 (n2786, n2693, n2704, n2777);
and  g2755 (n2783, n2777, n2779, n2737, n2723);
and  g2756 (n2782, n2694, n2741, n2777, n2525);
xor  g2757 (n2781, n2779, n2776, n2734);
xor  g2758 (n2785, n2706, n2701, n2776, n2730);
or   g2759 (n2790, n2725, n2705, n2776, n2778);
xor  g2760 (n2791, n2741, n2528, n2729, n2738);
xor  g2761 (n2810, n2795, n2788, n1108, n2780);
xor  g2762 (n2809, n2715, n1109, n2711, n1077);
nand g2763 (n2802, n2626, n1111, n1109, n2713);
xnor g2764 (n2806, n1077, n2627, n2629, n1111);
nand g2765 (n2797, n2792, n1108, n2782, n2790);
and  g2766 (n2814, n1110, n1112, n2789, n2714);
xor  g2767 (n2808, n2795, n2793, n2709, n2785);
or   g2768 (n2798, n2628, n1113, n1112, n2781);
nor  g2769 (n2811, n1112, n2784, n1109, n2790);
nor  g2770 (n2805, n2793, n2620, n1113, n2792);
xnor g2771 (n2796, n2621, n2617, n2787, n1107);
xnor g2772 (n2801, n2624, n1110, n2712, n1112);
and  g2773 (n2807, n2791, n1111, n1107, n2618);
nor  g2774 (n2800, n1110, n118, n2794, n2623);
xor  g2775 (n2804, n1077, n2625, n2795, n2794);
and  g2776 (n2799, n1113, n2783, n2716, n2793);
xnor g2777 (n2812, n2710, n2792, n2791, n2794);
and  g2778 (n2813, n1111, n1108, n1109, n2708);
xnor g2779 (n2803, n2622, n1110, n2790, n2791);
and  g2780 (n2815, n1113, n1108, n2619, n2786);
buf  g2781 (n2816, n2813);
not  g2782 (n2817, n2812);
or   g2783 (n2819, n2816, n2817, n437);
and  g2784 (n2822, n2815, n2817, n1183);
xnor g2785 (n2821, n1183, n2817, n438, n436);
and  g2786 (n2818, n2741, n438, n437);
nor  g2787 (n2820, n437, n438, n2814, n1183);
xnor g2788 (n2825, n2757, n1570, n1569, n2818);
xnor g2789 (n2828, n2756, n668, n2822, n1573);
nor  g2790 (n2827, n2819, n2822, n857);
or   g2791 (n2824, n2821, n2754, n2820, n1572);
or   g2792 (n2826, n670, n669, n2745, n2822);
and  g2793 (n2823, n671, n1568, n2755, n1571);
and  g2794 (n2832, n1575, n1578, n1582, n2823);
nand g2795 (n2830, n2824, n2825, n2826, n1583);
xnor g2796 (n2829, n1574, n1577, n2827, n2828);
and  g2797 (n2831, n1580, n1579, n1576, n1581);
nand g2798 (n2833, n2832, n2830, n2831, n2829);
endmodule
