// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_277_639 written by SynthGen on 2021/05/24 19:47:34
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_277_639 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21,
 n298, n293, n286, n291, n282, n294, n283, n296,
 n278, n287, n288, n279, n280, n276, n295, n277,
 n290, n281, n284, n285, n275, n289, n292, n297);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21;

output n298, n293, n286, n291, n282, n294, n283, n296,
 n278, n287, n288, n279, n280, n276, n295, n277,
 n290, n281, n284, n285, n275, n289, n292, n297;

wire n22, n23, n24, n25, n26, n27, n28, n29,
 n30, n31, n32, n33, n34, n35, n36, n37,
 n38, n39, n40, n41, n42, n43, n44, n45,
 n46, n47, n48, n49, n50, n51, n52, n53,
 n54, n55, n56, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n67, n68, n69,
 n70, n71, n72, n73, n74, n75, n76, n77,
 n78, n79, n80, n81, n82, n83, n84, n85,
 n86, n87, n88, n89, n90, n91, n92, n93,
 n94, n95, n96, n97, n98, n99, n100, n101,
 n102, n103, n104, n105, n106, n107, n108, n109,
 n110, n111, n112, n113, n114, n115, n116, n117,
 n118, n119, n120, n121, n122, n123, n124, n125,
 n126, n127, n128, n129, n130, n131, n132, n133,
 n134, n135, n136, n137, n138, n139, n140, n141,
 n142, n143, n144, n145, n146, n147, n148, n149,
 n150, n151, n152, n153, n154, n155, n156, n157,
 n158, n159, n160, n161, n162, n163, n164, n165,
 n166, n167, n168, n169, n170, n171, n172, n173,
 n174, n175, n176, n177, n178, n179, n180, n181,
 n182, n183, n184, n185, n186, n187, n188, n189,
 n190, n191, n192, n193, n194, n195, n196, n197,
 n198, n199, n200, n201, n202, n203, n204, n205,
 n206, n207, n208, n209, n210, n211, n212, n213,
 n214, n215, n216, n217, n218, n219, n220, n221,
 n222, n223, n224, n225, n226, n227, n228, n229,
 n230, n231, n232, n233, n234, n235, n236, n237,
 n238, n239, n240, n241, n242, n243, n244, n245,
 n246, n247, n248, n249, n250, n251, n252, n253,
 n254, n255, n256, n257, n258, n259, n260, n261,
 n262, n263, n264, n265, n266, n267, n268, n269,
 n270, n271, n272, n273, n274;

buf  g0 (n22, n5);
buf  g1 (n24, n2);
not  g2 (n25, n1);
not  g3 (n26, n4);
not  g4 (n23, n3);
not  g5 (n38, n25);
not  g6 (n39, n24);
not  g7 (n43, n23);
not  g8 (n37, n25);
buf  g9 (n32, n23);
buf  g10 (n36, n26);
not  g11 (n33, n26);
buf  g12 (n30, n24);
buf  g13 (n34, n23);
buf  g14 (n42, n26);
not  g15 (n29, n26);
buf  g16 (n35, n24);
not  g17 (n40, n25);
not  g18 (n28, n24);
not  g19 (n31, n23);
buf  g20 (n27, n25);
buf  g21 (n41, n22);
not  g22 (n62, n30);
not  g23 (n86, n32);
buf  g24 (n57, n39);
not  g25 (n88, n31);
buf  g26 (n69, n43);
buf  g27 (n102, n28);
buf  g28 (n50, n36);
buf  g29 (n96, n41);
buf  g30 (n58, n33);
not  g31 (n56, n42);
buf  g32 (n71, n39);
not  g33 (n98, n33);
not  g34 (n45, n29);
buf  g35 (n59, n42);
buf  g36 (n55, n28);
not  g37 (n68, n30);
buf  g38 (n66, n30);
buf  g39 (n78, n37);
not  g40 (n60, n43);
buf  g41 (n99, n43);
not  g42 (n95, n37);
not  g43 (n87, n33);
not  g44 (n63, n27);
buf  g45 (n67, n38);
buf  g46 (n80, n39);
buf  g47 (n101, n31);
not  g48 (n74, n29);
buf  g49 (n54, n33);
buf  g50 (n49, n38);
not  g51 (n64, n40);
not  g52 (n79, n32);
not  g53 (n44, n41);
not  g54 (n103, n35);
not  g55 (n92, n37);
not  g56 (n46, n38);
buf  g57 (n84, n37);
not  g58 (n82, n29);
buf  g59 (n97, n28);
not  g60 (n94, n34);
buf  g61 (n109, n41);
not  g62 (n53, n32);
buf  g63 (n51, n42);
buf  g64 (n85, n40);
not  g65 (n81, n34);
not  g66 (n72, n38);
not  g67 (n110, n39);
buf  g68 (n111, n34);
buf  g69 (n108, n27);
not  g70 (n104, n31);
not  g71 (n107, n28);
not  g72 (n100, n34);
buf  g73 (n89, n27);
not  g74 (n77, n40);
buf  g75 (n47, n35);
buf  g76 (n93, n30);
buf  g77 (n75, n29);
not  g78 (n83, n43);
buf  g79 (n52, n27);
buf  g80 (n73, n36);
not  g81 (n76, n41);
buf  g82 (n61, n35);
not  g83 (n65, n35);
not  g84 (n70, n40);
not  g85 (n48, n42);
buf  g86 (n106, n31);
buf  g87 (n90, n36);
not  g88 (n105, n32);
buf  g89 (n91, n36);
not  g90 (n181, n95);
buf  g91 (n189, n60);
buf  g92 (n180, n68);
not  g93 (n163, n76);
not  g94 (n178, n84);
not  g95 (n123, n65);
not  g96 (n187, n84);
buf  g97 (n193, n73);
buf  g98 (n179, n100);
buf  g99 (n125, n74);
not  g100 (n143, n19);
buf  g101 (n120, n10);
not  g102 (n167, n67);
nor  g103 (n130, n18, n51, n48);
and  g104 (n171, n82, n81, n51, n52);
nand g105 (n185, n67, n73, n106, n89);
and  g106 (n138, n17, n99, n60, n104);
nand g107 (n151, n87, n110, n55, n109);
and  g108 (n141, n56, n61, n82, n90);
nand g109 (n118, n101, n51, n61, n106);
nor  g110 (n152, n109, n75, n100);
xor  g111 (n160, n74, n111, n96);
xor  g112 (n135, n49, n56, n91, n97);
or   g113 (n186, n93, n84, n65, n85);
xor  g114 (n168, n46, n63, n75, n99);
and  g115 (n117, n102, n59, n64, n65);
or   g116 (n121, n83, n54, n76, n71);
and  g117 (n166, n106, n81, n104, n108);
xor  g118 (n124, n108, n53, n16, n11);
and  g119 (n164, n77, n54, n68, n21);
xnor g120 (n173, n45, n57, n44, n95);
and  g121 (n176, n82, n47, n44, n85);
nor  g122 (n153, n53, n69, n107, n68);
xor  g123 (n139, n58, n108, n52, n103);
and  g124 (n137, n51, n67, n110, n54);
and  g125 (n147, n80, n59, n53, n96);
xor  g126 (n128, n103, n93, n72, n84);
nand g127 (n155, n94, n55, n79, n49);
and  g128 (n184, n95, n57, n99, n105);
or   g129 (n142, n57, n89, n101, n88);
xnor g130 (n149, n94, n87, n95, n91);
xnor g131 (n182, n69, n66, n93, n92);
or   g132 (n136, n64, n100, n13, n54);
nand g133 (n114, n71, n111, n62, n58);
xnor g134 (n133, n97, n48, n109, n90);
and  g135 (n165, n64, n111, n50, n62);
xnor g136 (n190, n46, n75, n63, n66);
nand g137 (n144, n91, n49, n69, n87);
xnor g138 (n156, n62, n80, n73, n74);
nand g139 (n112, n98, n7, n105, n89);
or   g140 (n159, n109, n50, n70, n90);
and  g141 (n140, n102, n92, n48, n104);
xor  g142 (n175, n61, n68, n70, n97);
nand g143 (n132, n50, n98, n77, n96);
or   g144 (n177, n98, n107, n87, n81);
nand g145 (n131, n58, n79, n103, n45);
nand g146 (n174, n63, n8, n110, n60);
xnor g147 (n169, n88, n45, n102, n97);
or   g148 (n119, n103, n104, n83, n88);
or   g149 (n146, n46, n49, n71, n59);
xnor g150 (n154, n101, n12, n71, n85);
nand g151 (n129, n89, n60, n83, n86);
xnor g152 (n116, n52, n45, n98, n66);
xor  g153 (n192, n99, n44, n80, n77);
xor  g154 (n157, n70, n79, n107, n72);
nor  g155 (n191, n61, n108, n96, n107);
xor  g156 (n134, n56, n86, n64, n79);
xnor g157 (n158, n110, n105, n70, n48);
nor  g158 (n150, n6, n58, n102, n59);
or   g159 (n127, n77, n57, n55, n80);
nor  g160 (n148, n74, n56, n72, n50);
or   g161 (n172, n85, n55, n72, n106);
xnor g162 (n126, n78, n67, n47, n92);
and  g163 (n161, n78, n91, n92, n65);
xor  g164 (n113, n52, n82, n101, n90);
and  g165 (n183, n66, n86, n46, n76);
nand g166 (n188, n83, n9, n20, n47);
and  g167 (n145, n76, n44, n53, n78);
nand g168 (n115, n94, n78, n93, n62);
and  g169 (n162, n100, n105, n47, n94);
and  g170 (n170, n69, n15, n63, n81);
and  g171 (n122, n88, n86, n73, n14);
xor  g172 (n217, n134, n179, n148, n144);
nor  g173 (n212, n126, n124, n150, n136);
or   g174 (n218, n180, n112, n146, n182);
nand g175 (n258, n145, n123, n133);
and  g176 (n215, n129, n154, n190, n146);
nand g177 (n210, n114, n157, n128, n178);
and  g178 (n252, n182, n173, n162, n141);
xnor g179 (n268, n163, n166, n158, n134);
nand g180 (n220, n193, n172, n158, n177);
xnor g181 (n255, n174, n188, n159, n138);
xnor g182 (n260, n123, n168, n169);
or   g183 (n274, n168, n151, n164, n130);
and  g184 (n197, n156, n178, n190, n159);
nor  g185 (n233, n173, n152, n135, n141);
xor  g186 (n254, n126, n113, n130, n158);
or   g187 (n236, n141, n165, n183, n137);
xnor g188 (n227, n192, n124, n166, n119);
xor  g189 (n219, n120, n152, n142, n155);
and  g190 (n223, n170, n167, n136, n187);
xnor g191 (n239, n184, n118, n153, n120);
nand g192 (n246, n177, n188, n131, n141);
xor  g193 (n238, n176, n157, n114, n190);
nor  g194 (n213, n138, n127, n120, n152);
nor  g195 (n241, n176, n140, n118, n189);
nand g196 (n253, n185, n155, n179, n118);
nand g197 (n235, n155, n123, n163, n149);
and  g198 (n257, n191, n124, n116, n164);
and  g199 (n270, n174, n179, n125);
nor  g200 (n198, n161, n139, n174, n175);
or   g201 (n202, n192, n139, n134, n115);
or   g202 (n250, n177, n165, n147, n128);
xnor g203 (n249, n186, n164, n122, n157);
nand g204 (n229, n132, n186, n176, n169);
nor  g205 (n200, n177, n150, n162, n185);
nor  g206 (n206, n130, n136, n173, n134);
xnor g207 (n269, n116, n131, n150, n187);
xnor g208 (n194, n186, n183, n163, n148);
nand g209 (n266, n140, n138, n178, n121);
nand g210 (n195, n185, n140, n168, n143);
and  g211 (n271, n173, n132, n191, n167);
xnor g212 (n240, n135, n162, n159, n164);
and  g213 (n272, n147, n122, n145, n139);
xnor g214 (n261, n138, n157, n137, n156);
nor  g215 (n273, n151, n175, n149, n126);
and  g216 (n263, n137, n171, n121, n182);
xnor g217 (n211, n158, n130, n190, n170);
nor  g218 (n199, n113, n115, n125, n117);
or   g219 (n196, n142, n175, n181, n131);
nor  g220 (n248, n156, n128, n115, n132);
xor  g221 (n247, n153, n118, n182, n167);
and  g222 (n244, n115, n116, n117, n163);
or   g223 (n208, n144, n180, n187, n148);
or   g224 (n231, n161, n184, n127, n135);
and  g225 (n203, n125, n170, n127, n168);
xor  g226 (n265, n122, n181, n136, n189);
or   g227 (n242, n161, n176, n147, n124);
xnor g228 (n221, n191, n183, n154, n178);
nor  g229 (n256, n119, n133, n151, n117);
xor  g230 (n205, n171, n172, n142);
nor  g231 (n262, n160, n148, n152, n156);
xnor g232 (n204, n160, n169, n143, n180);
or   g233 (n226, n112, n189, n193, n174);
or   g234 (n224, n123, n145, n181, n140);
nand g235 (n214, n160, n116, n165, n143);
or   g236 (n232, n131, n150, n146, n132);
nor  g237 (n234, n129, n167, n153, n149);
nor  g238 (n245, n185, n137, n145, n192);
xnor g239 (n267, n122, n128, n184, n188);
nor  g240 (n230, n126, n186, n188, n159);
and  g241 (n222, n192, n135, n147, n149);
xnor g242 (n209, n144, n129, n121, n191);
xnor g243 (n251, n139, n143, n161, n119);
or   g244 (n259, n153, n187, n183, n142);
nor  g245 (n264, n184, n189, n170, n144);
nor  g246 (n228, n165, n119, n151, n114);
or   g247 (n237, n180, n146, n155, n166);
nor  g248 (n225, n162, n175, n121, n193);
xnor g249 (n207, n127, n171, n129, n133);
xnor g250 (n243, n193, n120, n154, n114);
and  g251 (n201, n181, n172, n171, n166);
xor  g252 (n216, n117, n160, n154, n125);
nand g253 (n289, n197, n245, n216, n223);
and  g254 (n276, n244, n208, n227, n273);
nand g255 (n293, n221, n203, n268, n194);
or   g256 (n298, n259, n254, n260, n246);
xor  g257 (n278, n226, n261, n270, n235);
xnor g258 (n294, n272, n270, n266, n198);
or   g259 (n282, n204, n220, n217, n239);
nor  g260 (n295, n222, n236, n256, n196);
xnor g261 (n290, n257, n232, n247, n274);
nand g262 (n286, n215, n274, n266, n269);
xnor g263 (n275, n234, n201, n274, n233);
xnor g264 (n291, n241, n264, n250, n253);
and  g265 (n285, n212, n238, n224, n248);
nor  g266 (n292, n249, n252, n210, n265);
xor  g267 (n296, n195, n240, n225, n205);
xor  g268 (n284, n264, n262, n219, n206);
xor  g269 (n287, n267, n237, n200, n271);
or   g270 (n288, n262, n230, n213, n263);
nor  g271 (n277, n229, n218, n265, n211);
xor  g272 (n280, n272, n268, n274, n271);
nand g273 (n281, n251, n202, n269, n267);
or   g274 (n283, n207, n228, n209, n214);
xnor g275 (n279, n255, n263, n258, n242);
and  g276 (n297, n199, n243, n231, n273);
endmodule
