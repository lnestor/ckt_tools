

module Stat_100_46
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n70,
  n69,
  n120,
  n102,
  n121,
  n106,
  n108,
  n112,
  n114,
  n109,
  n85,
  n83,
  n94,
  n111,
  n99,
  n115,
  n92,
  n116,
  n89,
  n86,
  n110,
  n119,
  n125,
  n123,
  n127,
  n131,
  n128,
  n126,
  n124,
  n132,
  n130,
  n129,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n70;
  output n69;
  output n120;
  output n102;
  output n121;
  output n106;
  output n108;
  output n112;
  output n114;
  output n109;
  output n85;
  output n83;
  output n94;
  output n111;
  output n99;
  output n115;
  output n92;
  output n116;
  output n89;
  output n86;
  output n110;
  output n119;
  output n125;
  output n123;
  output n127;
  output n131;
  output n128;
  output n126;
  output n124;
  output n132;
  output n130;
  output n129;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n84;
  wire n87;
  wire n88;
  wire n90;
  wire n91;
  wire n93;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n100;
  wire n101;
  wire n103;
  wire n104;
  wire n105;
  wire n107;
  wire n113;
  wire n117;
  wire n118;
  wire n122;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    KeyWire_0_34,
    n3
  );


  not
  g1
  (
    n35,
    n1
  );


  not
  g2
  (
    KeyWire_0_22,
    n10
  );


  not
  g3
  (
    n36,
    n5
  );


  buf
  g4
  (
    KeyWire_0_51,
    n4
  );


  buf
  g5
  (
    KeyWire_0_18,
    n9
  );


  buf
  g6
  (
    n33,
    n7
  );


  not
  g7
  (
    n41,
    n6
  );


  buf
  g8
  (
    KeyWire_0_20,
    n2
  );


  not
  g9
  (
    KeyWire_0_6,
    n11
  );


  not
  g10
  (
    n38,
    n8
  );


  not
  g11
  (
    KeyWire_0_26,
    n36
  );


  buf
  g12
  (
    n55,
    n35
  );


  buf
  g13
  (
    KeyWire_0_25,
    n37
  );


  not
  g14
  (
    n63,
    n36
  );


  buf
  g15
  (
    n71,
    n43
  );


  buf
  g16
  (
    n62,
    n41
  );


  buf
  g17
  (
    KeyWire_0_14,
    n41
  );


  not
  g18
  (
    KeyWire_0_32,
    n34
  );


  not
  g19
  (
    KeyWire_0_29,
    n42
  );


  buf
  g20
  (
    KeyWire_0_45,
    n38
  );


  not
  g21
  (
    KeyWire_0_0,
    n35
  );


  buf
  g22
  (
    KeyWire_0_13,
    n38
  );


  not
  g23
  (
    n47,
    n41
  );


  buf
  g24
  (
    KeyWire_0_3,
    n39
  );


  buf
  g25
  (
    KeyWire_0_48,
    n43
  );


  buf
  g26
  (
    KeyWire_0_23,
    n39
  );


  not
  g27
  (
    KeyWire_0_40,
    n36
  );


  not
  g28
  (
    KeyWire_0_43,
    n40
  );


  buf
  g29
  (
    KeyWire_0_10,
    n37
  );


  buf
  g30
  (
    KeyWire_0_36,
    n43
  );


  buf
  g31
  (
    KeyWire_0_9,
    n42
  );


  not
  g32
  (
    n61,
    n35
  );


  buf
  g33
  (
    KeyWire_0_8,
    n35
  );


  not
  g34
  (
    n51,
    n38
  );


  buf
  g35
  (
    KeyWire_0_59,
    n37
  );


  not
  g36
  (
    KeyWire_0_50,
    n34
  );


  not
  g37
  (
    n80,
    n38
  );


  buf
  g38
  (
    KeyWire_0_44,
    n34
  );


  not
  g39
  (
    KeyWire_0_49,
    n42
  );


  buf
  g40
  (
    KeyWire_0_4,
    n41
  );


  buf
  g41
  (
    n82,
    n36
  );


  buf
  g42
  (
    KeyWire_0_38,
    n39
  );


  buf
  g43
  (
    n72,
    n39
  );


  buf
  g44
  (
    KeyWire_0_35,
    n43
  );


  buf
  g45
  (
    KeyWire_0_1,
    n34
  );


  buf
  g46
  (
    KeyWire_0_47,
    n37
  );


  not
  g47
  (
    KeyWire_0_39,
    n40
  );


  buf
  g48
  (
    KeyWire_0_27,
    n42
  );


  buf
  g49
  (
    n53,
    n40
  );


  not
  g50
  (
    KeyWire_0_60,
    n70
  );


  buf
  g51
  (
    n91,
    n56
  );


  xor
  g52
  (
    KeyWire_0_31,
    n55,
    n72,
    n71
  );


  nor
  g53
  (
    n108,
    n77,
    n82,
    n69,
    n65
  );


  nor
  g54
  (
    n109,
    n46,
    n63,
    n60,
    n77
  );


  xor
  g55
  (
    n84,
    n46,
    n66,
    n58,
    n71
  );


  xnor
  g56
  (
    KeyWire_0_28,
    n78,
    n77,
    n50
  );


  or
  g57
  (
    KeyWire_0_12,
    n61,
    n47,
    n62,
    n68
  );


  or
  g58
  (
    n98,
    n79,
    n78,
    n55,
    n50
  );


  or
  g59
  (
    n104,
    n57,
    n81,
    n68
  );


  nor
  g60
  (
    n93,
    n78,
    n76,
    n79,
    n61
  );


  nor
  g61
  (
    KeyWire_0_54,
    n62,
    n73,
    n55,
    n57
  );


  xnor
  g62
  (
    n119,
    n70,
    n56,
    n49,
    n48
  );


  xor
  g63
  (
    n85,
    n59,
    n56,
    n80,
    n58
  );


  and
  g64
  (
    KeyWire_0_19,
    n67,
    n64,
    n81,
    n62
  );


  xnor
  g65
  (
    KeyWire_0_63,
    n75,
    n70,
    n60,
    n63
  );


  or
  g66
  (
    KeyWire_0_24,
    n79,
    n81,
    n51,
    n54
  );


  or
  g67
  (
    n117,
    n64,
    n59,
    n74,
    n82
  );


  or
  g68
  (
    KeyWire_0_42,
    n64,
    n76,
    n75,
    n73
  );


  xnor
  g69
  (
    KeyWire_0_61,
    n55,
    n75,
    n59,
    n64
  );


  nand
  g70
  (
    KeyWire_0_7,
    n48,
    n79,
    n71,
    n69
  );


  xor
  g71
  (
    KeyWire_0_16,
    n57,
    n45,
    n49,
    n73
  );


  or
  g72
  (
    KeyWire_0_2,
    n72,
    n80,
    n62,
    n74
  );


  xnor
  g73
  (
    KeyWire_0_37,
    n75,
    n60,
    n45,
    n69
  );


  or
  g74
  (
    KeyWire_0_57,
    n49,
    n51,
    n53
  );


  xor
  g75
  (
    KeyWire_0_41,
    n65,
    n47,
    n51,
    n66
  );


  nor
  g76
  (
    n89,
    n54,
    n54,
    n82,
    n50
  );


  and
  g77
  (
    n90,
    n80,
    n66,
    n57
  );


  xor
  g78
  (
    n106,
    n53,
    n50,
    n47,
    n12
  );


  xnor
  g79
  (
    n114,
    n72,
    n82,
    n61,
    n63
  );


  xor
  g80
  (
    n111,
    n65,
    n49,
    n76,
    n60
  );


  nand
  g81
  (
    n96,
    n45,
    n71,
    n48,
    n47
  );


  or
  g82
  (
    KeyWire_0_56,
    n58,
    n67,
    n53,
    n61
  );


  or
  g83
  (
    KeyWire_0_21,
    n67,
    n46,
    n69,
    n45
  );


  or
  g84
  (
    KeyWire_0_52,
    n76,
    n52,
    n73
  );


  nor
  g85
  (
    n115,
    n78,
    n56,
    n58,
    n68
  );


  nand
  g86
  (
    KeyWire_0_46,
    n59,
    n74,
    n80,
    n54
  );


  xnor
  g87
  (
    n87,
    n74,
    n65,
    n52,
    n70
  );


  xnor
  g88
  (
    KeyWire_0_30,
    n48,
    n68,
    n53,
    n67
  );


  nand
  g89
  (
    n103,
    n52,
    n72,
    n46,
    n63
  );


  xnor
  g90
  (
    KeyWire_0_62,
    n13,
    n105,
    n108,
    n110
  );


  nor
  g91
  (
    KeyWire_0_15,
    n115,
    n24,
    n119,
    n19
  );


  nand
  g92
  (
    KeyWire_0_33,
    n30,
    n113,
    n104,
    n28
  );


  nor
  g93
  (
    KeyWire_0_17,
    n114,
    n25,
    n111,
    n109
  );


  or
  g94
  (
    KeyWire_0_53,
    n122,
    n117,
    n29,
    n15
  );


  nand
  g95
  (
    KeyWire_0_11,
    n120,
    n14,
    n103,
    n16
  );


  or
  g96
  (
    n128,
    n112,
    n17,
    n26,
    n121
  );


  xor
  g97
  (
    KeyWire_0_58,
    n31,
    n20,
    n21,
    n23
  );


  or
  g98
  (
    KeyWire_0_55,
    n107,
    n116,
    n106,
    n118
  );


  and
  g99
  (
    KeyWire_0_5,
    n27,
    n22,
    n32,
    n18
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n59,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n77,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n116,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n74,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n46,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n125,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n34,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n112,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n49,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n69,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n78,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n131,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n83,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n75,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n70,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n129,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n121,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n123,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n40,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n105,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n39,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n107,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n43,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n73,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n100,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n56,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n48,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n52,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n86,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n68,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n94,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n95,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n57,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n124,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n42,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n54,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n79,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n118,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n66,
    keyIn_0_38,
    KeyWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n67,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n44,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    n92,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n122,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n81,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n65,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n64,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n102,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n58,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n45,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n50,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n60,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n37,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n88,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n130,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n101,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n132,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n97,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n113,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n127,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n76,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n110,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n99,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n126,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n120,
    KeyNOTWire_0_63
  );


endmodule

