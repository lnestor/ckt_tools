// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\6_15_large_circuits\Stat_1363_31_10 written by SynthGen on 2021/06/15 15:04:53
module Stat_1363_31_10( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n1117, n1123, n1116, n1121, n1110, n1124, n1122, n1119,
 n1118, n1128, n1409, n1407, n1403, n1401, n1410, n1408,
 n1405, n1411, n1402, n1406, n1404);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48;

output n1117, n1123, n1116, n1121, n1110, n1124, n1122, n1119,
 n1118, n1128, n1409, n1407, n1403, n1401, n1410, n1408,
 n1405, n1411, n1402, n1406, n1404;

wire n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1111, n1112, n1113,
 n1114, n1115, n1120, n1125, n1126, n1127, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400;

not  g0 (n178, n3);
buf  g1 (n58, n36);
buf  g2 (n196, n24);
buf  g3 (n208, n42);
not  g4 (n189, n1);
buf  g5 (n110, n4);
not  g6 (n120, n10);
buf  g7 (n215, n11);
not  g8 (n154, n9);
buf  g9 (n116, n36);
not  g10 (n114, n28);
not  g11 (n81, n24);
not  g12 (n49, n37);
buf  g13 (n216, n8);
buf  g14 (n129, n16);
not  g15 (n157, n21);
not  g16 (n199, n5);
not  g17 (n64, n41);
not  g18 (n94, n28);
buf  g19 (n193, n6);
buf  g20 (n141, n10);
buf  g21 (n174, n32);
buf  g22 (n133, n33);
buf  g23 (n186, n7);
buf  g24 (n105, n18);
buf  g25 (n102, n5);
not  g26 (n77, n8);
not  g27 (n175, n41);
not  g28 (n52, n2);
not  g29 (n185, n25);
buf  g30 (n167, n7);
not  g31 (n112, n23);
not  g32 (n184, n15);
buf  g33 (n214, n8);
not  g34 (n176, n14);
buf  g35 (n180, n26);
buf  g36 (n88, n4);
not  g37 (n137, n27);
not  g38 (n128, n6);
not  g39 (n104, n29);
buf  g40 (n205, n31);
buf  g41 (n50, n9);
not  g42 (n73, n33);
buf  g43 (n90, n29);
not  g44 (n107, n30);
buf  g45 (n111, n37);
buf  g46 (n158, n17);
buf  g47 (n192, n6);
not  g48 (n132, n13);
not  g49 (n86, n41);
buf  g50 (n82, n26);
not  g51 (n68, n17);
buf  g52 (n163, n33);
buf  g53 (n188, n23);
not  g54 (n70, n13);
not  g55 (n209, n29);
buf  g56 (n206, n12);
not  g57 (n170, n3);
not  g58 (n63, n41);
buf  g59 (n172, n24);
not  g60 (n165, n35);
buf  g61 (n67, n42);
buf  g62 (n181, n13);
not  g63 (n156, n7);
buf  g64 (n54, n10);
not  g65 (n144, n4);
not  g66 (n62, n2);
buf  g67 (n93, n15);
buf  g68 (n169, n20);
buf  g69 (n65, n25);
not  g70 (n145, n42);
buf  g71 (n113, n19);
buf  g72 (n127, n40);
not  g73 (n147, n23);
buf  g74 (n194, n20);
buf  g75 (n166, n10);
buf  g76 (n213, n34);
buf  g77 (n103, n28);
not  g78 (n123, n9);
buf  g79 (n210, n19);
buf  g80 (n198, n29);
not  g81 (n131, n22);
buf  g82 (n142, n17);
not  g83 (n191, n21);
buf  g84 (n56, n22);
buf  g85 (n152, n34);
not  g86 (n177, n11);
not  g87 (n97, n3);
buf  g88 (n190, n28);
buf  g89 (n161, n9);
buf  g90 (n99, n38);
buf  g91 (n117, n16);
buf  g92 (n160, n42);
not  g93 (n53, n30);
not  g94 (n85, n18);
not  g95 (n173, n35);
buf  g96 (n101, n34);
not  g97 (n149, n4);
not  g98 (n168, n35);
not  g99 (n211, n8);
not  g100 (n98, n20);
not  g101 (n138, n40);
buf  g102 (n153, n27);
buf  g103 (n202, n38);
buf  g104 (n92, n12);
buf  g105 (n79, n31);
buf  g106 (n171, n32);
not  g107 (n151, n14);
not  g108 (n162, n31);
not  g109 (n207, n21);
buf  g110 (n96, n5);
not  g111 (n115, n6);
not  g112 (n84, n24);
buf  g113 (n126, n26);
not  g114 (n95, n40);
not  g115 (n135, n30);
buf  g116 (n71, n19);
not  g117 (n91, n18);
not  g118 (n197, n16);
not  g119 (n183, n40);
not  g120 (n89, n12);
buf  g121 (n87, n2);
buf  g122 (n136, n37);
not  g123 (n143, n31);
buf  g124 (n80, n39);
buf  g125 (n130, n38);
buf  g126 (n60, n15);
not  g127 (n51, n27);
not  g128 (n134, n32);
not  g129 (n182, n32);
not  g130 (n108, n15);
not  g131 (n148, n27);
buf  g132 (n203, n14);
buf  g133 (n204, n25);
buf  g134 (n75, n5);
buf  g135 (n100, n21);
buf  g136 (n187, n22);
not  g137 (n72, n16);
not  g138 (n146, n13);
not  g139 (n109, n1);
buf  g140 (n125, n38);
not  g141 (n200, n1);
not  g142 (n179, n3);
not  g143 (n159, n36);
not  g144 (n106, n11);
not  g145 (n61, n20);
not  g146 (n124, n17);
not  g147 (n201, n26);
not  g148 (n212, n36);
not  g149 (n121, n35);
buf  g150 (n83, n39);
not  g151 (n155, n12);
not  g152 (n66, n1);
buf  g153 (n195, n33);
not  g154 (n139, n14);
buf  g155 (n164, n2);
not  g156 (n55, n34);
not  g157 (n78, n18);
not  g158 (n57, n25);
buf  g159 (n59, n11);
buf  g160 (n150, n39);
not  g161 (n74, n19);
not  g162 (n76, n39);
not  g163 (n118, n23);
not  g164 (n140, n22);
not  g165 (n119, n37);
not  g166 (n69, n30);
not  g167 (n122, n7);
not  g168 (n653, n137);
buf  g169 (n818, n125);
buf  g170 (n353, n178);
buf  g171 (n566, n150);
buf  g172 (n227, n135);
not  g173 (n218, n161);
buf  g174 (n248, n115);
not  g175 (n692, n131);
buf  g176 (n501, n125);
not  g177 (n698, n162);
buf  g178 (n365, n69);
not  g179 (n799, n115);
not  g180 (n350, n79);
buf  g181 (n622, n142);
buf  g182 (n803, n88);
not  g183 (n774, n143);
buf  g184 (n487, n187);
buf  g185 (n656, n112);
buf  g186 (n759, n153);
buf  g187 (n328, n167);
not  g188 (n804, n191);
not  g189 (n513, n137);
not  g190 (n287, n163);
not  g191 (n447, n112);
not  g192 (n289, n124);
buf  g193 (n363, n142);
not  g194 (n712, n189);
buf  g195 (n702, n192);
buf  g196 (n628, n100);
not  g197 (n836, n93);
not  g198 (n709, n147);
not  g199 (n681, n188);
not  g200 (n730, n87);
not  g201 (n242, n63);
not  g202 (n834, n73);
not  g203 (n543, n104);
not  g204 (n255, n121);
buf  g205 (n846, n91);
not  g206 (n439, n59);
buf  g207 (n641, n181);
not  g208 (n294, n191);
buf  g209 (n415, n84);
not  g210 (n408, n112);
not  g211 (n547, n115);
not  g212 (n637, n151);
not  g213 (n824, n68);
not  g214 (n463, n169);
buf  g215 (n417, n170);
buf  g216 (n428, n85);
not  g217 (n288, n128);
buf  g218 (n636, n64);
not  g219 (n310, n55);
not  g220 (n564, n145);
not  g221 (n259, n202);
not  g222 (n714, n50);
not  g223 (n745, n175);
buf  g224 (n652, n188);
not  g225 (n555, n65);
not  g226 (n472, n101);
not  g227 (n507, n175);
not  g228 (n768, n152);
buf  g229 (n512, n133);
not  g230 (n706, n132);
buf  g231 (n783, n148);
buf  g232 (n696, n75);
not  g233 (n635, n204);
not  g234 (n378, n112);
buf  g235 (n701, n66);
buf  g236 (n356, n49);
not  g237 (n568, n55);
not  g238 (n320, n120);
not  g239 (n838, n205);
not  g240 (n506, n104);
buf  g241 (n740, n127);
not  g242 (n282, n127);
not  g243 (n674, n66);
buf  g244 (n737, n113);
buf  g245 (n226, n127);
not  g246 (n843, n158);
buf  g247 (n492, n100);
not  g248 (n615, n92);
buf  g249 (n784, n106);
buf  g250 (n708, n180);
buf  g251 (n241, n160);
buf  g252 (n497, n85);
not  g253 (n291, n100);
buf  g254 (n546, n70);
buf  g255 (n277, n182);
not  g256 (n519, n173);
buf  g257 (n584, n113);
not  g258 (n822, n76);
buf  g259 (n461, n111);
buf  g260 (n411, n132);
buf  g261 (n613, n143);
buf  g262 (n420, n86);
buf  g263 (n359, n79);
buf  g264 (n658, n150);
buf  g265 (n526, n108);
buf  g266 (n751, n168);
buf  g267 (n357, n117);
buf  g268 (n471, n49);
buf  g269 (n811, n123);
not  g270 (n223, n180);
buf  g271 (n764, n76);
not  g272 (n738, n197);
not  g273 (n433, n207);
buf  g274 (n625, n124);
buf  g275 (n258, n155);
buf  g276 (n781, n152);
not  g277 (n264, n83);
not  g278 (n581, n169);
not  g279 (n779, n190);
not  g280 (n565, n109);
not  g281 (n302, n147);
not  g282 (n343, n199);
not  g283 (n261, n188);
not  g284 (n377, n164);
buf  g285 (n413, n107);
buf  g286 (n587, n206);
not  g287 (n435, n92);
buf  g288 (n247, n147);
buf  g289 (n621, n140);
buf  g290 (n796, n126);
not  g291 (n484, n137);
not  g292 (n713, n190);
not  g293 (n347, n80);
not  g294 (n369, n165);
buf  g295 (n711, n150);
buf  g296 (n485, n110);
buf  g297 (n829, n72);
not  g298 (n772, n122);
not  g299 (n493, n58);
buf  g300 (n807, n128);
not  g301 (n296, n188);
not  g302 (n518, n173);
buf  g303 (n601, n60);
not  g304 (n585, n171);
buf  g305 (n429, n183);
buf  g306 (n573, n161);
not  g307 (n780, n174);
buf  g308 (n797, n164);
not  g309 (n747, n50);
not  g310 (n726, n96);
not  g311 (n577, n49);
buf  g312 (n321, n62);
buf  g313 (n578, n126);
buf  g314 (n776, n88);
buf  g315 (n399, n72);
buf  g316 (n785, n189);
not  g317 (n693, n129);
buf  g318 (n596, n82);
buf  g319 (n643, n160);
buf  g320 (n603, n67);
buf  g321 (n375, n156);
not  g322 (n449, n167);
buf  g323 (n600, n176);
not  g324 (n389, n96);
not  g325 (n539, n114);
not  g326 (n246, n73);
buf  g327 (n267, n119);
buf  g328 (n406, n56);
buf  g329 (n346, n78);
buf  g330 (n669, n133);
not  g331 (n753, n63);
buf  g332 (n544, n76);
not  g333 (n503, n98);
buf  g334 (n739, n179);
buf  g335 (n680, n197);
buf  g336 (n474, n85);
buf  g337 (n450, n79);
buf  g338 (n252, n157);
buf  g339 (n763, n98);
not  g340 (n383, n133);
buf  g341 (n397, n138);
buf  g342 (n524, n96);
buf  g343 (n612, n107);
buf  g344 (n238, n197);
buf  g345 (n283, n168);
buf  g346 (n367, n142);
buf  g347 (n823, n158);
not  g348 (n298, n153);
not  g349 (n672, n194);
not  g350 (n315, n152);
not  g351 (n541, n151);
buf  g352 (n480, n174);
not  g353 (n830, n102);
buf  g354 (n390, n165);
not  g355 (n814, n85);
not  g356 (n683, n72);
not  g357 (n793, n93);
buf  g358 (n662, n87);
buf  g359 (n618, n67);
not  g360 (n736, n80);
not  g361 (n454, n199);
buf  g362 (n704, n154);
not  g363 (n778, n68);
buf  g364 (n404, n191);
not  g365 (n278, n65);
not  g366 (n393, n91);
not  g367 (n733, n167);
not  g368 (n514, n196);
buf  g369 (n465, n132);
not  g370 (n611, n157);
not  g371 (n540, n54);
not  g372 (n767, n139);
buf  g373 (n219, n68);
buf  g374 (n322, n156);
not  g375 (n668, n132);
buf  g376 (n409, n125);
not  g377 (n243, n149);
not  g378 (n607, n175);
buf  g379 (n624, n121);
buf  g380 (n281, n190);
buf  g381 (n634, n131);
not  g382 (n629, n53);
not  g383 (n679, n166);
not  g384 (n372, n51);
buf  g385 (n262, n93);
buf  g386 (n617, n69);
buf  g387 (n231, n179);
buf  g388 (n609, n141);
buf  g389 (n269, n69);
not  g390 (n334, n113);
buf  g391 (n639, n151);
not  g392 (n667, n199);
not  g393 (n659, n198);
not  g394 (n791, n111);
not  g395 (n813, n129);
not  g396 (n542, n110);
buf  g397 (n309, n90);
buf  g398 (n305, n162);
not  g399 (n469, n166);
buf  g400 (n695, n206);
not  g401 (n268, n193);
not  g402 (n563, n78);
buf  g403 (n230, n59);
buf  g404 (n689, n198);
not  g405 (n478, n121);
not  g406 (n479, n185);
not  g407 (n810, n144);
buf  g408 (n462, n52);
not  g409 (n286, n195);
buf  g410 (n528, n77);
buf  g411 (n339, n155);
buf  g412 (n762, n164);
not  g413 (n582, n56);
buf  g414 (n551, n116);
not  g415 (n424, n56);
not  g416 (n645, n205);
buf  g417 (n646, n148);
not  g418 (n591, n115);
not  g419 (n398, n58);
buf  g420 (n414, n200);
not  g421 (n719, n136);
not  g422 (n240, n134);
buf  g423 (n533, n189);
buf  g424 (n847, n99);
buf  g425 (n827, n67);
buf  g426 (n604, n172);
not  g427 (n486, n190);
not  g428 (n279, n136);
buf  g429 (n387, n106);
not  g430 (n438, n52);
not  g431 (n351, n140);
buf  g432 (n718, n95);
buf  g433 (n532, n203);
not  g434 (n329, n207);
buf  g435 (n537, n146);
not  g436 (n456, n70);
buf  g437 (n556, n160);
buf  g438 (n312, n50);
buf  g439 (n703, n186);
buf  g440 (n395, n170);
buf  g441 (n481, n87);
buf  g442 (n815, n80);
not  g443 (n729, n77);
buf  g444 (n642, n51);
not  g445 (n446, n89);
not  g446 (n835, n121);
buf  g447 (n598, n59);
not  g448 (n427, n74);
not  g449 (n345, n183);
not  g450 (n444, n184);
not  g451 (n661, n172);
not  g452 (n274, n177);
buf  g453 (n304, n136);
not  g454 (n549, n158);
buf  g455 (n579, n150);
not  g456 (n798, n134);
not  g457 (n314, n111);
not  g458 (n839, n106);
buf  g459 (n782, n145);
buf  g460 (n690, n154);
not  g461 (n233, n128);
buf  g462 (n300, n157);
not  g463 (n496, n80);
buf  g464 (n225, n141);
not  g465 (n816, n145);
buf  g466 (n728, n60);
not  g467 (n741, n193);
buf  g468 (n786, n181);
not  g469 (n384, n99);
buf  g470 (n284, n56);
not  g471 (n498, n167);
buf  g472 (n236, n202);
buf  g473 (n545, n77);
not  g474 (n657, n194);
not  g475 (n337, n94);
not  g476 (n280, n185);
not  g477 (n371, n53);
not  g478 (n531, n65);
buf  g479 (n677, n105);
not  g480 (n760, n170);
buf  g481 (n648, n164);
buf  g482 (n234, n181);
not  g483 (n841, n141);
buf  g484 (n299, n71);
buf  g485 (n732, n81);
buf  g486 (n473, n72);
not  g487 (n735, n124);
not  g488 (n567, n171);
buf  g489 (n686, n101);
not  g490 (n228, n182);
buf  g491 (n673, n61);
not  g492 (n602, n146);
not  g493 (n301, n109);
not  g494 (n335, n95);
not  g495 (n499, n86);
not  g496 (n491, n178);
buf  g497 (n220, n110);
not  g498 (n405, n204);
not  g499 (n520, n136);
buf  g500 (n434, n103);
not  g501 (n442, n198);
not  g502 (n569, n203);
not  g503 (n421, n103);
not  g504 (n235, n75);
not  g505 (n694, n159);
buf  g506 (n316, n172);
not  g507 (n410, n144);
buf  g508 (n344, n113);
buf  g509 (n597, n71);
not  g510 (n794, n192);
buf  g511 (n515, n91);
buf  g512 (n401, n195);
not  g513 (n251, n123);
buf  g514 (n423, n105);
not  g515 (n826, n97);
buf  g516 (n580, n123);
not  g517 (n670, n159);
buf  g518 (n821, n169);
buf  g519 (n691, n205);
buf  g520 (n654, n120);
not  g521 (n403, n96);
not  g522 (n361, n57);
buf  g523 (n490, n74);
buf  g524 (n769, n129);
buf  g525 (n483, n148);
buf  g526 (n400, n60);
not  g527 (n808, n205);
not  g528 (n529, n90);
buf  g529 (n755, n98);
not  g530 (n336, n82);
not  g531 (n527, n183);
not  g532 (n502, n201);
buf  g533 (n592, n62);
not  g534 (n352, n51);
not  g535 (n276, n97);
not  g536 (n575, n75);
not  g537 (n459, n54);
not  g538 (n599, n57);
buf  g539 (n222, n53);
buf  g540 (n663, n147);
buf  g541 (n746, n177);
not  g542 (n576, n58);
buf  g543 (n530, n71);
not  g544 (n623, n81);
buf  g545 (n265, n61);
buf  g546 (n303, n171);
not  g547 (n716, n186);
not  g548 (n705, n101);
buf  g549 (n844, n143);
buf  g550 (n470, n123);
not  g551 (n426, n66);
buf  g552 (n809, n182);
not  g553 (n761, n166);
not  g554 (n536, n117);
buf  g555 (n293, n204);
buf  g556 (n270, n187);
buf  g557 (n789, n81);
not  g558 (n458, n139);
not  g559 (n550, n206);
not  g560 (n752, n84);
buf  g561 (n845, n161);
buf  g562 (n440, n163);
not  g563 (n717, n77);
buf  g564 (n848, n78);
buf  g565 (n317, n53);
not  g566 (n833, n145);
buf  g567 (n297, n92);
buf  g568 (n432, n153);
buf  g569 (n430, n65);
buf  g570 (n385, n161);
not  g571 (n700, n75);
buf  g572 (n237, n49);
not  g573 (n801, n149);
buf  g574 (n720, n88);
buf  g575 (n460, n122);
buf  g576 (n381, n120);
buf  g577 (n368, n54);
buf  g578 (n306, n142);
buf  g579 (n311, n197);
not  g580 (n684, n172);
buf  g581 (n805, n187);
not  g582 (n825, n144);
buf  g583 (n562, n169);
buf  g584 (n790, n138);
not  g585 (n224, n168);
not  g586 (n425, n162);
buf  g587 (n715, n81);
not  g588 (n254, n203);
buf  g589 (n849, n98);
buf  g590 (n295, n195);
not  g591 (n837, n187);
not  g592 (n245, n126);
not  g593 (n391, n97);
not  g594 (n676, n183);
buf  g595 (n457, n118);
buf  g596 (n374, n66);
buf  g597 (n558, n107);
not  g598 (n724, n202);
buf  g599 (n557, n178);
buf  g600 (n734, n156);
not  g601 (n710, n149);
not  g602 (n272, n110);
not  g603 (n475, n69);
not  g604 (n436, n195);
buf  g605 (n742, n107);
buf  g606 (n770, n86);
not  g607 (n342, n118);
buf  g608 (n614, n73);
not  g609 (n416, n117);
buf  g610 (n412, n76);
buf  g611 (n232, n109);
not  g612 (n758, n191);
buf  g613 (n806, n63);
not  g614 (n535, n60);
not  g615 (n504, n201);
not  g616 (n360, n61);
buf  g617 (n553, n83);
buf  g618 (n508, n138);
buf  g619 (n370, n116);
not  g620 (n419, n189);
not  g621 (n627, n200);
buf  g622 (n616, n61);
not  g623 (n330, n87);
not  g624 (n355, n119);
not  g625 (n650, n140);
not  g626 (n548, n159);
not  g627 (n257, n184);
not  g628 (n271, n70);
buf  g629 (n748, n71);
buf  g630 (n773, n184);
buf  g631 (n244, n95);
buf  g632 (n586, n109);
buf  g633 (n757, n86);
buf  g634 (n831, n163);
buf  g635 (n338, n67);
buf  g636 (n756, n204);
not  g637 (n638, n151);
buf  g638 (n510, n58);
buf  g639 (n445, n54);
not  g640 (n290, n83);
buf  g641 (n500, n193);
buf  g642 (n792, n84);
buf  g643 (n422, n198);
not  g644 (n840, n180);
buf  g645 (n340, n146);
buf  g646 (n448, n68);
not  g647 (n590, n70);
buf  g648 (n464, n130);
not  g649 (n788, n148);
not  g650 (n812, n138);
not  g651 (n678, n114);
buf  g652 (n358, n128);
buf  g653 (n509, n55);
not  g654 (n292, n108);
not  g655 (n800, n141);
buf  g656 (n256, n120);
buf  g657 (n707, n158);
not  g658 (n561, n51);
not  g659 (n610, n135);
not  g660 (n386, n114);
not  g661 (n229, n140);
not  g662 (n402, n201);
buf  g663 (n495, n186);
buf  g664 (n766, n144);
not  g665 (n828, n192);
not  g666 (n333, n74);
buf  g667 (n332, n64);
buf  g668 (n494, n152);
not  g669 (n249, n101);
buf  g670 (n593, n196);
buf  g671 (n572, n179);
not  g672 (n687, n180);
not  g673 (n559, n55);
buf  g674 (n407, n117);
not  g675 (n731, n63);
not  g676 (n647, n94);
buf  g677 (n534, n124);
not  g678 (n795, n57);
buf  g679 (n285, n134);
buf  g680 (n476, n82);
buf  g681 (n632, n173);
not  g682 (n606, n83);
buf  g683 (n787, n199);
buf  g684 (n671, n116);
not  g685 (n522, n130);
not  g686 (n665, n182);
buf  g687 (n313, n89);
not  g688 (n777, n73);
not  g689 (n376, n122);
not  g690 (n239, n177);
buf  g691 (n323, n139);
not  g692 (n832, n106);
buf  g693 (n666, n157);
buf  g694 (n554, n59);
buf  g695 (n331, n185);
not  g696 (n688, n118);
buf  g697 (n754, n57);
not  g698 (n324, n166);
not  g699 (n517, n79);
buf  g700 (n588, n52);
buf  g701 (n660, n155);
not  g702 (n675, n91);
buf  g703 (n725, n181);
buf  g704 (n488, n194);
not  g705 (n468, n165);
not  g706 (n620, n162);
not  g707 (n765, n122);
not  g708 (n221, n108);
buf  g709 (n341, n130);
buf  g710 (n307, n89);
not  g711 (n354, n94);
not  g712 (n589, n116);
not  g713 (n552, n88);
not  g714 (n366, n108);
not  g715 (n452, n50);
buf  g716 (n364, n104);
buf  g717 (n253, n90);
buf  g718 (n505, n103);
buf  g719 (n318, n129);
not  g720 (n743, n104);
buf  g721 (n727, n168);
not  g722 (n392, n105);
buf  g723 (n583, n163);
not  g724 (n273, n103);
not  g725 (n850, n93);
not  g726 (n349, n178);
buf  g727 (n651, n194);
buf  g728 (n373, n64);
not  g729 (n466, n89);
buf  g730 (n560, n102);
not  g731 (n451, n196);
not  g732 (n489, n170);
buf  g733 (n266, n175);
buf  g734 (n594, n137);
buf  g735 (n263, n185);
buf  g736 (n388, n90);
not  g737 (n699, n154);
buf  g738 (n467, n62);
not  g739 (n644, n97);
not  g740 (n664, n203);
not  g741 (n626, n174);
buf  g742 (n308, n171);
not  g743 (n362, n119);
buf  g744 (n655, n206);
not  g745 (n418, n100);
buf  g746 (n453, n82);
not  g747 (n477, n94);
buf  g748 (n574, n102);
not  g749 (n379, n131);
not  g750 (n685, n186);
not  g751 (n721, n176);
not  g752 (n538, n99);
not  g753 (n217, n176);
buf  g754 (n851, n105);
buf  g755 (n749, n102);
buf  g756 (n608, n99);
not  g757 (n771, n92);
not  g758 (n649, n133);
buf  g759 (n441, n139);
buf  g760 (n640, n125);
not  g761 (n571, n78);
buf  g762 (n744, n177);
not  g763 (n380, n64);
not  g764 (n820, n179);
not  g765 (n443, n193);
not  g766 (n523, n160);
buf  g767 (n842, n149);
buf  g768 (n697, n84);
not  g769 (n817, n184);
not  g770 (n437, n156);
buf  g771 (n630, n207);
not  g772 (n605, n135);
buf  g773 (n631, n146);
buf  g774 (n802, n154);
buf  g775 (n525, n200);
not  g776 (n516, n131);
buf  g777 (n723, n134);
not  g778 (n250, n196);
not  g779 (n327, n62);
buf  g780 (n431, n95);
not  g781 (n750, n155);
buf  g782 (n260, n114);
buf  g783 (n325, n143);
buf  g784 (n396, n135);
buf  g785 (n382, n130);
not  g786 (n722, n118);
buf  g787 (n511, n127);
not  g788 (n570, n202);
not  g789 (n775, n165);
buf  g790 (n455, n74);
buf  g791 (n326, n119);
buf  g792 (n682, n153);
not  g793 (n275, n111);
not  g794 (n595, n159);
not  g795 (n319, n201);
not  g796 (n619, n176);
buf  g797 (n394, n173);
not  g798 (n482, n52);
not  g799 (n633, n200);
buf  g800 (n819, n192);
not  g801 (n521, n126);
buf  g802 (n348, n174);
xnor g803 (n949, n470, n290, n447, n420);
or   g804 (n948, n429, n387, n418, n445);
xor  g805 (n916, n441, n348, n584, n334);
or   g806 (n895, n656, n306, n323, n281);
or   g807 (n961, n226, n384, n315, n502);
nand g808 (n974, n625, n528, n375, n642);
nand g809 (n893, n761, n769, n771, n788);
and  g810 (n859, n758, n358, n262, n609);
nor  g811 (n878, n593, n278, n512, n777);
nor  g812 (n892, n643, n551, n293, n605);
nor  g813 (n942, n751, n602, n288, n545);
and  g814 (n889, n530, n667, n572, n564);
xnor g815 (n988, n388, n608, n604, n475);
and  g816 (n955, n220, n600, n424, n238);
xor  g817 (n900, n207, n535, n689, n465);
and  g818 (n968, n736, n303, n340, n362);
nor  g819 (n917, n663, n491, n742, n794);
xor  g820 (n918, n623, n639, n416, n511);
or   g821 (n959, n489, n628, n529, n498);
xor  g822 (n899, n360, n371, n433, n658);
nand g823 (n962, n403, n251, n611, n641);
or   g824 (n911, n634, n727, n257, n504);
xnor g825 (n934, n563, n582, n693, n601);
nor  g826 (n935, n701, n411, n263, n542);
or   g827 (n932, n786, n382, n485, n302);
nor  g828 (n869, n676, n330, n749, n737);
xnor g829 (n923, n482, n533, n432, n380);
or   g830 (n868, n633, n785, n274, n754);
xor  g831 (n958, n299, n507, n265, n366);
nor  g832 (n910, n450, n493, n280, n479);
nand g833 (n969, n789, n264, n253, n589);
xor  g834 (n896, n685, n467, n648, n506);
xnor g835 (n865, n614, n588, n461, n774);
xor  g836 (n928, n409, n252, n421, n718);
nand g837 (n936, n228, n569, n795, n574);
and  g838 (n901, n790, n462, n399, n760);
and  g839 (n913, n456, n515, n679, n219);
nand g840 (n960, n463, n596, n617, n494);
or   g841 (n938, n578, n223, n250, n546);
or   g842 (n866, n446, n335, n301, n757);
and  g843 (n951, n495, n417, n552, n367);
and  g844 (n920, n240, n540, n464, n566);
nor  g845 (n886, n733, n695, n653, n230);
nor  g846 (n981, n428, n256, n621, n324);
and  g847 (n941, n555, n597, n710, n668);
xnor g848 (n864, n361, n513, n332, n694);
nor  g849 (n979, n644, n365, n592, n452);
nor  g850 (n984, n556, n675, n791, n692);
nor  g851 (n929, n357, n442, n624, n469);
nand g852 (n983, n747, n410, n313, n570);
xor  g853 (n858, n729, n275, n440, n618);
nor  g854 (n905, n686, n327, n590, n347);
or   g855 (n952, n354, n460, n717, n522);
xor  g856 (n973, n339, n286, n239, n364);
xnor g857 (n922, n708, n343, n647, n294);
xor  g858 (n943, n422, n431, n224, n547);
and  g859 (n933, n383, n688, n379, n586);
xnor g860 (n867, n650, n743, n374, n405);
xor  g861 (n915, n439, n319, n603, n594);
xor  g862 (n987, n386, n671, n407, n517);
nor  g863 (n919, n395, n630, n300, n539);
xor  g864 (n975, n350, n778, n244, n304);
or   g865 (n853, n363, n497, n712, n328);
xor  g866 (n931, n599, n553, n295, n659);
or   g867 (n991, n261, n268, n472, n401);
or   g868 (n950, n558, n776, n466, n732);
xnor g869 (n921, n784, n780, n753, n707);
xnor g870 (n937, n703, n237, n698, n673);
nand g871 (n906, n412, n458, n247, n490);
xnor g872 (n927, n745, n266, n705, n775);
or   g873 (n926, n505, n400, n322, n437);
nand g874 (n863, n598, n550, n538, n503);
nand g875 (n884, n393, n724, n520, n782);
nand g876 (n872, n738, n474, n662, n516);
xor  g877 (n874, n756, n235, n255, n351);
xor  g878 (n857, n748, n763, n765, n344);
and  g879 (n982, n402, n587, n620, n514);
or   g880 (n940, n532, n459, n276, n660);
xor  g881 (n904, n414, n372, n764, n585);
xnor g882 (n887, n779, n486, n273, n355);
xor  g883 (n870, n752, n792, n687, n426);
xor  g884 (n956, n267, n483, n534, n787);
nor  g885 (n976, n723, n218, n557, n320);
xor  g886 (n971, n562, n269, n652, n773);
or   g887 (n882, n560, n317, n622, n312);
nand g888 (n989, n651, n677, n318, n523);
xor  g889 (n890, n443, n510, n316, n755);
and  g890 (n902, n481, n279, n619, n683);
and  g891 (n912, n283, n715, n739, n271);
xor  g892 (n860, n478, n666, n720, n356);
xor  g893 (n925, n419, n436, n455, n616);
nor  g894 (n966, n728, n338, n245, n635);
nand g895 (n992, n243, n607, n632, n438);
nor  g896 (n894, n649, n242, n711, n772);
xnor g897 (n881, n484, n285, n615, n329);
nand g898 (n862, n249, n565, n413, n548);
and  g899 (n970, n398, n561, n337, n292);
xor  g900 (n898, n770, n640, n581, n225);
nor  g901 (n963, n744, n352, n654, n699);
and  g902 (n897, n759, n377, n521, n314);
xor  g903 (n994, n310, n369, n353, n696);
or   g904 (n891, n454, n722, n719, n378);
and  g905 (n930, n227, n576, n451, n298);
xnor g906 (n875, n783, n746, n396, n741);
nand g907 (n985, n704, n793, n571, n691);
xnor g908 (n965, n473, n305, n277, n735);
nand g909 (n852, n331, n381, n270, n664);
or   g910 (n888, n716, n449, n488, n246);
or   g911 (n996, n681, n341, n531, n453);
xnor g912 (n856, n536, n404, n713, n579);
nor  g913 (n972, n518, n231, n731, n389);
xnor g914 (n967, n645, n448, n241, n670);
xnor g915 (n903, n349, n415, n333, n346);
and  g916 (n855, n629, n359, n509, n408);
nand g917 (n964, n549, n610, n222, n326);
nor  g918 (n879, n457, n730, n311, n248);
and  g919 (n873, n373, n376, n740, n684);
or   g920 (n990, n568, n697, n307, n537);
xor  g921 (n885, n613, n674, n526, n544);
nor  g922 (n947, n406, n519, n287, n527);
and  g923 (n907, n427, n236, n390, n525);
xor  g924 (n908, n444, n471, n233, n750);
and  g925 (n909, n487, n342, n725, n655);
xor  g926 (n861, n309, n259, n700, n591);
or   g927 (n953, n284, n612, n595, n260);
xor  g928 (n939, n657, n682, n468, n661);
xnor g929 (n978, n709, n423, n606, n234);
and  g930 (n986, n706, n480, n714, n282);
nand g931 (n944, n325, n781, n258, n434);
or   g932 (n924, n768, n678, n492, n627);
and  g933 (n946, n345, n541, n336, n680);
or   g934 (n954, n577, n297, n291, n477);
nor  g935 (n854, n394, n646, n500, n573);
xor  g936 (n876, n397, n499, n496, n554);
or   g937 (n883, n232, n626, n476, n721);
xnor g938 (n880, n669, n665, n289, n726);
or   g939 (n993, n229, n767, n690, n296);
nor  g940 (n877, n580, n430, n524, n637);
and  g941 (n957, n559, n308, n501, n391);
and  g942 (n914, n370, n272, n385, n368);
and  g943 (n945, n636, n567, n435, n702);
xor  g944 (n995, n254, n672, n221, n321);
or   g945 (n980, n631, n508, n762, n217);
and  g946 (n871, n425, n734, n543, n583);
xor  g947 (n977, n766, n638, n575, n392);
xnor g948 (n1001, n852, n864);
nor  g949 (n1004, n869, n874);
xnor g950 (n1003, n879, n881);
nor  g951 (n1005, n878, n883);
or   g952 (n999, n872, n859);
xor  g953 (n1007, n871, n876);
xor  g954 (n1002, n863, n868);
nand g955 (n1008, n877, n856);
or   g956 (n1009, n882, n860);
xnor g957 (n1000, n853, n854);
nor  g958 (n997, n867, n865);
nand g959 (n998, n857, n873);
and  g960 (n1011, n858, n862);
xor  g961 (n1006, n866, n880);
and  g962 (n1012, n855, n875);
and  g963 (n1010, n870, n861);
buf  g964 (n1013, n998);
buf  g965 (n1014, n997);
buf  g966 (n1018, n1013);
not  g967 (n1017, n1013);
not  g968 (n1016, n1013);
not  g969 (n1015, n1013);
xor  g970 (n1019, n900, n1001, n1015, n1003);
xor  g971 (n1025, n906, n1004, n887, n902);
xnor g972 (n1022, n1015, n1001, n911, n999);
xnor g973 (n1024, n1001, n1016, n897, n905);
nand g974 (n1021, n889, n1017, n899, n1002);
and  g975 (n1020, n884, n891, n1015, n910);
nor  g976 (n1027, n1016, n1000, n907, n901);
nand g977 (n1032, n1004, n1017, n1002, n898);
nor  g978 (n1033, n1000, n894, n1017, n1016);
nor  g979 (n1023, n1018, n1018, n890, n1001);
or   g980 (n1031, n912, n904, n1018, n1015);
xor  g981 (n1034, n903, n1017, n886, n1002);
and  g982 (n1029, n1018, n888, n1003);
nand g983 (n1028, n1016, n1003, n885, n895);
nor  g984 (n1030, n909, n893, n1004, n892);
or   g985 (n1026, n896, n1000, n908, n1002);
or   g986 (n1037, n46, n47, n48);
xor  g987 (n1041, n43, n1023, n45, n44);
xnor g988 (n1042, n43, n1026, n48, n45);
xor  g989 (n1040, n1022, n43, n47, n44);
nand g990 (n1038, n43, n46, n1020, n1025);
nand g991 (n1036, n44, n45, n48, n1021);
nor  g992 (n1039, n45, n48, n1019, n46);
or   g993 (n1035, n46, n47, n1024, n44);
not  g994 (n1063, n1040);
not  g995 (n1050, n210);
buf  g996 (n1060, n1038);
buf  g997 (n1052, n1039);
not  g998 (n1051, n1037);
buf  g999 (n1061, n210);
not  g1000 (n1047, n209);
not  g1001 (n1059, n209);
buf  g1002 (n1057, n208);
not  g1003 (n1043, n208);
not  g1004 (n1056, n1042);
buf  g1005 (n1046, n1036);
buf  g1006 (n1048, n208);
not  g1007 (n1044, n1035);
buf  g1008 (n1058, n1042);
not  g1009 (n1062, n1041);
not  g1010 (n1045, n1036);
xor  g1011 (n1053, n1037, n1041, n1038);
or   g1012 (n1054, n1041, n210, n209, n1040);
and  g1013 (n1049, n1039, n209, n1040, n1042);
xor  g1014 (n1055, n1040, n1035, n208, n1041);
not  g1015 (n1075, n1043);
buf  g1016 (n1067, n1043);
buf  g1017 (n1065, n1043);
not  g1018 (n1074, n796);
buf  g1019 (n1071, n1044);
buf  g1020 (n1070, n1044);
buf  g1021 (n1064, n1045);
buf  g1022 (n1072, n1045);
not  g1023 (n1066, n1044);
buf  g1024 (n1073, n1044);
and  g1025 (n1068, n1043, n798);
and  g1026 (n1069, n797, n1045, n799);
buf  g1027 (n1085, n1064);
not  g1028 (n1077, n1066);
not  g1029 (n1089, n1067);
not  g1030 (n1081, n1067);
not  g1031 (n1080, n1067);
not  g1032 (n1087, n1067);
buf  g1033 (n1079, n1064);
not  g1034 (n1090, n1066);
not  g1035 (n1082, n1065);
buf  g1036 (n1088, n1064);
buf  g1037 (n1076, n1066);
not  g1038 (n1078, n1065);
buf  g1039 (n1084, n1066);
buf  g1040 (n1086, n1064);
buf  g1041 (n1083, n1065);
buf  g1042 (n1091, n1065);
not  g1043 (n1105, n1079);
not  g1044 (n1108, n1077);
not  g1045 (n1107, n1076);
not  g1046 (n1093, n1079);
buf  g1047 (n1103, n1080);
not  g1048 (n1095, n1078);
buf  g1049 (n1106, n1079);
buf  g1050 (n1098, n1077);
not  g1051 (n1096, n1076);
buf  g1052 (n1099, n1078);
buf  g1053 (n1094, n1080);
not  g1054 (n1100, n1077);
buf  g1055 (n1104, n1078);
buf  g1056 (n1109, n1077);
not  g1057 (n1092, n1076);
buf  g1058 (n1101, n1078);
not  g1059 (n1097, n1076);
not  g1060 (n1102, n1079);
not  g1061 (n1115, n918);
not  g1062 (n1119, n1094);
buf  g1063 (n1117, n1092);
not  g1064 (n1123, n914);
not  g1065 (n1111, n1095);
not  g1066 (n1126, n1094);
not  g1067 (n1121, n1092);
not  g1068 (n1127, n1014);
not  g1069 (n1112, n1093);
buf  g1070 (n1118, n1096);
not  g1071 (n1122, n1014);
not  g1072 (n1113, n1095);
buf  g1073 (n1124, n1096);
not  g1074 (n1116, n1014);
buf  g1075 (n1110, n1095);
xnor g1076 (n1128, n915, n913);
or   g1077 (n1114, n916, n917, n1093, n1096);
and  g1078 (n1125, n1014, n1094, n1093);
and  g1079 (n1120, n1094, n1092, n1095);
xnor g1080 (n1136, n214, n1122, n215);
and  g1081 (n1131, n1121, n1120, n216, n210);
nor  g1082 (n1137, n216, n1124, n919, n211);
or   g1083 (n1129, n211, n214, n920, n1127);
xnor g1084 (n1130, n1125, n216, n212);
xor  g1085 (n1132, n213, n213, n211, n1128);
nor  g1086 (n1133, n211, n214, n212);
and  g1087 (n1134, n1126, n213, n214);
xnor g1088 (n1135, n216, n215, n1123);
nor  g1089 (n1149, n805, n808, n811, n801);
xor  g1090 (n1144, n1028, n1031, n802, n1132);
or   g1091 (n1145, n1132, n1133, n807, n814);
xor  g1092 (n1146, n820, n804, n825, n824);
xor  g1093 (n1147, n809, n1033, n1029, n1129);
or   g1094 (n1141, n803, n812, n1133, n1131);
nor  g1095 (n1148, n821, n1134, n1130, n1129);
or   g1096 (n1140, n806, n1134, n819, n827);
nor  g1097 (n1138, n813, n1130, n818, n1032);
nor  g1098 (n1139, n816, n822, n817, n1131);
nand g1099 (n1143, n800, n810, n815, n1034);
xnor g1100 (n1142, n826, n1027, n1030, n823);
not  g1101 (n1155, n1138);
not  g1102 (n1150, n1138);
not  g1103 (n1151, n1139);
not  g1104 (n1154, n1139);
not  g1105 (n1153, n1139);
not  g1106 (n1152, n1139);
nor  g1107 (n1158, n1057, n1152, n1062, n1054);
nor  g1108 (n1175, n1058, n1153, n1055, n1061);
and  g1109 (n1160, n1063, n1154, n1057);
xor  g1110 (n1167, n1051, n1150, n1060, n1059);
xor  g1111 (n1177, n1153, n1052, n1154, n1051);
xor  g1112 (n1168, n1059, n1056, n1050, n1063);
xor  g1113 (n1165, n1150, n1155, n1053);
or   g1114 (n1171, n1063, n1152, n1047, n1051);
and  g1115 (n1161, n1062, n1059, n1053, n1054);
nor  g1116 (n1159, n1052, n1051, n1153, n1055);
nor  g1117 (n1178, n1054, n1055, n1151, n1153);
or   g1118 (n1173, n1154, n1049, n1152, n1050);
nor  g1119 (n1170, n1060, n1060, n1049, n1055);
nand g1120 (n1156, n1151, n1048, n1047, n1046);
nor  g1121 (n1176, n1155, n1151, n1054, n1058);
or   g1122 (n1169, n1059, n1150, n1152, n1060);
xor  g1123 (n1172, n1155, n1049, n1056);
xor  g1124 (n1163, n1056, n1155, n1151, n1063);
xor  g1125 (n1162, n1046, n1048, n1150);
and  g1126 (n1164, n1047, n1053, n1046, n1061);
and  g1127 (n1166, n1047, n1062, n1061);
xnor g1128 (n1174, n1050, n1057, n1052, n1049);
nor  g1129 (n1157, n1154, n1058, n1061, n1050);
nor  g1130 (n1179, n1058, n1052, n1046, n1048);
buf  g1131 (n1183, n1156);
buf  g1132 (n1181, n1158);
not  g1133 (n1182, n1157);
buf  g1134 (n1180, n1157);
nand g1135 (n1187, n1086, n1090, n1087, n1182);
nand g1136 (n1190, n1183, n1091, n1087, n1084);
xor  g1137 (n1188, n1085, n1183, n1086, n1090);
xnor g1138 (n1186, n1089, n1088, n1083, n1082);
or   g1139 (n1192, n1088, n1090, n1180, n1081);
xor  g1140 (n1184, n1089, n1087, n1083, n1086);
xnor g1141 (n1185, n921, n1085, n1180, n1089);
or   g1142 (n1197, n1182, n1181, n1088, n1080);
xor  g1143 (n1198, n1084, n1086, n1091);
nand g1144 (n1193, n1088, n1084, n1083, n1180);
or   g1145 (n1196, n1084, n1082, n1181);
nor  g1146 (n1199, n1080, n1083, n1085, n1183);
xnor g1147 (n1195, n922, n1081, n1091);
and  g1148 (n1194, n1180, n1181, n1085, n1090);
and  g1149 (n1191, n1089, n1087, n1081, n1183);
nor  g1150 (n1189, n1082, n1182, n1181);
xor  g1151 (n1204, n1195, n1099, n1100, n1005);
nand g1152 (n1219, n1195, n1196, n1158, n1097);
nand g1153 (n1203, n1006, n1007, n1102, n1191);
and  g1154 (n1221, n1196, n1159, n1107, n1008);
xor  g1155 (n1208, n1103, n1187, n1098, n1188);
xnor g1156 (n1224, n1101, n1186, n1160, n1105);
nor  g1157 (n1228, n1105, n1109, n1103, n1100);
nand g1158 (n1225, n1104, n1097, n1193, n1160);
and  g1159 (n1220, n1190, n1161, n1109, n1007);
nor  g1160 (n1216, n1195, n1134, n1161, n1106);
or   g1161 (n1217, n1098, n1163, n1107, n1193);
nor  g1162 (n1222, n1107, n1005, n1162, n1159);
nand g1163 (n1211, n1007, n1106, n1005);
or   g1164 (n1213, n1194, n1004, n1105, n1187);
nand g1165 (n1212, n1100, n1190, n1105, n1108);
or   g1166 (n1201, n1194, n1194, n1101, n1102);
or   g1167 (n1200, n1163, n1096, n1101, n1109);
or   g1168 (n1226, n1163, n1108, n1097);
and  g1169 (n1206, n1104, n1102, n1160, n1101);
nand g1170 (n1209, n1008, n1108, n1007, n1005);
and  g1171 (n1218, n1184, n1099, n1192, n1104);
nor  g1172 (n1214, n1162, n1103, n1189, n1163);
and  g1173 (n1210, n1189, n1109, n1191, n1162);
or   g1174 (n1223, n1100, n1192, n1104, n1006);
nand g1175 (n1202, n1008, n1097, n1006, n1193);
xnor g1176 (n1229, n1161, n1188, n1103, n1099);
nor  g1177 (n1215, n1102, n1160, n1194, n1186);
xnor g1178 (n1227, n1161, n1195, n1162, n1193);
nand g1179 (n1205, n1106, n1098, n1008, n1099);
nand g1180 (n1207, n1185, n1006, n1098, n1107);
not  g1181 (n1230, n1212);
buf  g1182 (n1234, n1211);
not  g1183 (n1235, n1216);
buf  g1184 (n1242, n1202);
not  g1185 (n1233, n1214);
buf  g1186 (n1245, n1207);
buf  g1187 (n1244, n1203);
not  g1188 (n1240, n1210);
not  g1189 (n1243, n1204);
buf  g1190 (n1237, n1200);
buf  g1191 (n1247, n1205);
buf  g1192 (n1239, n1208);
not  g1193 (n1236, n1217);
buf  g1194 (n1238, n1209);
buf  g1195 (n1231, n1213);
not  g1196 (n1246, n1206);
not  g1197 (n1232, n1201);
not  g1198 (n1241, n1215);
not  g1199 (n1250, n1230);
not  g1200 (n1249, n1230);
not  g1201 (n1248, n1230);
nand g1202 (n1256, n1248, n1144, n1146, n1140);
xor  g1203 (n1254, n1148, n1147, n1249, n1145);
xnor g1204 (n1259, n1147, n1144, n1145);
or   g1205 (n1262, n1143, n1249, n1141, n1250);
nor  g1206 (n1258, n1140, n1249, n1143);
xor  g1207 (n1257, n1148, n1146, n1142);
xnor g1208 (n1253, n1147, n1248, n1141, n1146);
nand g1209 (n1251, n1144, n1143, n1248, n1145);
xor  g1210 (n1260, n1148, n1145, n1248, n1140);
or   g1211 (n1255, n1148, n1142, n1250);
nand g1212 (n1261, n1146, n1141, n1140);
nor  g1213 (n1252, n1250, n1147, n1249, n1142);
buf  g1214 (n1275, n1252);
buf  g1215 (n1277, n956);
not  g1216 (n1274, n933);
nand g1217 (n1278, n1254, n940, n936);
or   g1218 (n1264, n1257, n953, n957, n1251);
nand g1219 (n1271, n951, n943, n925, n960);
xor  g1220 (n1268, n1254, n934, n1252, n939);
or   g1221 (n1266, n954, n944, n930, n937);
or   g1222 (n1265, n927, n1257, n942, n1256);
or   g1223 (n1276, n952, n1258, n924, n931);
xnor g1224 (n1269, n1253, n965, n947, n962);
xnor g1225 (n1280, n945, n932, n1251, n948);
xnor g1226 (n1267, n964, n1258, n941, n963);
or   g1227 (n1263, n935, n926, n946, n1255);
xnor g1228 (n1272, n938, n961, n928, n949);
and  g1229 (n1273, n923, n955, n1255, n1258);
nor  g1230 (n1279, n966, n950, n929, n1259);
or   g1231 (n1270, n1256, n1253, n958, n959);
or   g1232 (n1282, n1263, n1166, n1164);
or   g1233 (n1284, n1167, n1166, n1165, n1168);
nor  g1234 (n1285, n1264, n1165);
nor  g1235 (n1283, n1167, n1166, n1265, n1164);
or   g1236 (n1286, n1167, n1267, n1268, n1168);
nand g1237 (n1281, n1266, n1167, n1164, n1166);
buf  g1238 (n1287, n1281);
buf  g1239 (n1288, n1283);
not  g1240 (n1289, n1282);
xor  g1241 (n1293, n1198, n1196, n1199, n1197);
and  g1242 (n1291, n1197, n1198, n1289);
or   g1243 (n1290, n1288, n1197, n1289, n1287);
xnor g1244 (n1292, n1199, n1199, n1269, n1288);
or   g1245 (n1294, n1199, n1198, n1196, n1197);
nand g1246 (n1296, n1279, n1136, n1226, n1219);
xor  g1247 (n1312, n1276, n1291, n1290, n1136);
xnor g1248 (n1310, n1277, n1226, n1224);
and  g1249 (n1306, n1294, n1293, n1292);
xnor g1250 (n1299, n1135, n1229, n1222, n1225);
xnor g1251 (n1311, n1275, n1136, n1227);
nand g1252 (n1300, n1290, n1228, n1292, n1291);
xor  g1253 (n1297, n1223, n1273, n1272, n1274);
nor  g1254 (n1304, n1229, n1294, n1137, n1278);
or   g1255 (n1303, n1278, n1291, n1273, n1226);
and  g1256 (n1305, n1227, n1228, n1134, n1229);
nor  g1257 (n1314, n1276, n1221, n1275, n1293);
or   g1258 (n1298, n1277, n1270, n1220, n1135);
and  g1259 (n1307, n1277, n1292, n1135, n1290);
xnor g1260 (n1295, n1218, n1225, n1293, n1229);
nand g1261 (n1301, n1225, n1277, n1227, n1224);
nand g1262 (n1309, n1135, n1223, n1271, n1292);
nand g1263 (n1308, n1228, n1272, n1290, n1278);
or   g1264 (n1302, n1291, n1225, n1227, n1278);
xnor g1265 (n1313, n1228, n1294, n1274);
and  g1266 (n1350, n842, n1245, n1313, n1312);
xnor g1267 (n1361, n1242, n1069, n844, n1238);
or   g1268 (n1335, n829, n1011, n1238, n1074);
nor  g1269 (n1318, n1010, n1285, n834, n1311);
and  g1270 (n1322, n1300, n1233, n1231, n1235);
or   g1271 (n1352, n1072, n848, n1240, n1010);
or   g1272 (n1347, n1069, n1012, n1305, n1301);
nor  g1273 (n1344, n1244, n1314, n1243, n1012);
or   g1274 (n1328, n1241, n846, n1071, n828);
nor  g1275 (n1343, n1069, n850, n1239);
xor  g1276 (n1366, n1071, n1239, n847, n1074);
or   g1277 (n1354, n1075, n839, n1302, n1073);
and  g1278 (n1327, n1245, n830, n1242, n1244);
nor  g1279 (n1333, n1073, n1259, n1075, n1307);
xnor g1280 (n1341, n1308, n1247, n1305, n1231);
nor  g1281 (n1356, n1231, n1071, n1306, n1009);
or   g1282 (n1359, n837, n1243, n840, n1070);
xor  g1283 (n1321, n1236, n838, n831, n1012);
xor  g1284 (n1357, n1240, n1235, n841, n1236);
nand g1285 (n1355, n1011, n1299, n1309, n1298);
nand g1286 (n1365, n1234, n1241, n1069, n845);
nand g1287 (n1362, n1149, n1279, n1313, n1247);
nand g1288 (n1358, n1075, n1305, n1149, n1231);
or   g1289 (n1342, n843, n1308, n1299, n1071);
and  g1290 (n1340, n967, n1074, n1312, n1313);
xnor g1291 (n1338, n1073, n1312, n1070, n1244);
nor  g1292 (n1353, n1238, n1070, n1230, n1297);
or   g1293 (n1316, n1072, n1297, n1240, n1241);
and  g1294 (n1324, n1009, n1308, n1242, n1307);
xor  g1295 (n1364, n1279, n1235, n1302, n1296);
and  g1296 (n1351, n1068, n1243, n1244, n1234);
or   g1297 (n1325, n1310, n1303, n1237, n1011);
nand g1298 (n1348, n1314, n1234, n1309, n1295);
xor  g1299 (n1326, n1237, n1068, n1304, n836);
xor  g1300 (n1329, n1070, n1072, n1296, n832);
xnor g1301 (n1363, n1068, n1236, n1075, n1072);
and  g1302 (n1337, n968, n1284, n1246, n1237);
xnor g1303 (n1339, n1241, n1295, n1238, n1304);
xnor g1304 (n1319, n1242, n1012, n1232, n1313);
nor  g1305 (n1345, n1237, n1246, n969, n1234);
xnor g1306 (n1317, n1309, n1232, n1042, n1233);
or   g1307 (n1360, n1149, n851, n1009, n1010);
nor  g1308 (n1346, n1235, n1286, n1314, n1307);
or   g1309 (n1315, n1247, n1301, n1243, n1068);
nor  g1310 (n1349, n1314, n835, n1310, n1233);
xor  g1311 (n1331, n1311, n1011, n1310, n849);
nor  g1312 (n1336, n1311, n1279, n1239, n1306);
or   g1313 (n1334, n1009, n1246, n1010, n1232);
or   g1314 (n1320, n1298, n1245, n1074, n1236);
nand g1315 (n1332, n1245, n1306, n1303, n1149);
xnor g1316 (n1323, n1233, n1232, n1300, n1246);
xor  g1317 (n1330, n1247, n1073, n1240, n833);
xor  g1318 (n1378, n1178, n1168, n1320, n1335);
xor  g1319 (n1375, n1177, n1171, n992, n989);
nor  g1320 (n1382, n1170, n1360, n1365, n1327);
xnor g1321 (n1385, n1329, n1179, n990, n1259);
xnor g1322 (n1389, n1325, n1352, n1350, n1174);
and  g1323 (n1390, n1361, n1322, n1174, n1171);
or   g1324 (n1371, n1176, n1179, n1362, n1354);
xnor g1325 (n1377, n1355, n1315, n1280, n974);
xnor g1326 (n1374, n1364, n1178, n1324, n1176);
xnor g1327 (n1397, n1363, n1340, n993, n1260);
xor  g1328 (n1381, n1137, n1172, n1168);
xnor g1329 (n1391, n1280, n1323, n971, n1177);
nor  g1330 (n1368, n1353, n1346, n1333, n1137);
xnor g1331 (n1370, n978, n1170, n1280, n1356);
and  g1332 (n1398, n1172, n1345, n984, n982);
nand g1333 (n1379, n1169, n1177, n1171, n1178);
xnor g1334 (n1395, n1326, n979, n1173, n1316);
xnor g1335 (n1367, n1321, n1178, n1169, n1343);
nor  g1336 (n1386, n1179, n994, n1170, n973);
and  g1337 (n1388, n1338, n1179, n1357, n1366);
nand g1338 (n1394, n1334, n1331, n1342, n1344);
xor  g1339 (n1369, n1259, n1349, n1339, n1359);
nand g1340 (n1396, n991, n983, n1319, n1170);
xnor g1341 (n1393, n986, n1348, n975, n1260);
and  g1342 (n1383, n995, n1328, n976, n970);
nand g1343 (n1392, n1171, n1175, n987, n1358);
and  g1344 (n1384, n1175, n1351, n1173, n1318);
xor  g1345 (n1372, n977, n1169, n981, n1175);
nand g1346 (n1376, n1330, n1174, n1137, n972);
xnor g1347 (n1400, n1280, n1337, n1173, n985);
and  g1348 (n1373, n996, n1177, n1317, n980);
or   g1349 (n1387, n1174, n1332, n1169, n1172);
nor  g1350 (n1380, n988, n1176, n1341);
xnor g1351 (n1399, n1336, n1175, n1173, n1347);
or   g1352 (n1401, n1384, n1372, n1400, n1376);
xor  g1353 (n1403, n1379, n1371, n1390, n1260);
or   g1354 (n1405, n1262, n1388, n1398, n1374);
and  g1355 (n1410, n1375, n1399, n1261, n1394);
nand g1356 (n1409, n1262, n1387, n1261, n1395);
nor  g1357 (n1411, n1369, n1389, n1261, n1380);
and  g1358 (n1402, n1377, n1370, n1397, n1383);
xor  g1359 (n1406, n1373, n1378, n1260, n1381);
nand g1360 (n1404, n1367, n1393, n1368, n1386);
nand g1361 (n1407, n1382, n1261, n1392, n1391);
xor  g1362 (n1408, n1385, n1396, n1262);
endmodule
