// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_803_2716 written by SynthGen on 2021/05/24 19:48:30
module Stat_803_2716( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27,
 n698, n701, n689, n693, n794, n830, n820, n828,
 n819, n821, n825, n824, n823, n829, n827, n822,
 n826);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27;

output n698, n701, n689, n693, n794, n830, n820, n828,
 n819, n821, n825, n824, n823, n829, n827, n822,
 n826;

wire n28, n29, n30, n31, n32, n33, n34, n35,
 n36, n37, n38, n39, n40, n41, n42, n43,
 n44, n45, n46, n47, n48, n49, n50, n51,
 n52, n53, n54, n55, n56, n57, n58, n59,
 n60, n61, n62, n63, n64, n65, n66, n67,
 n68, n69, n70, n71, n72, n73, n74, n75,
 n76, n77, n78, n79, n80, n81, n82, n83,
 n84, n85, n86, n87, n88, n89, n90, n91,
 n92, n93, n94, n95, n96, n97, n98, n99,
 n100, n101, n102, n103, n104, n105, n106, n107,
 n108, n109, n110, n111, n112, n113, n114, n115,
 n116, n117, n118, n119, n120, n121, n122, n123,
 n124, n125, n126, n127, n128, n129, n130, n131,
 n132, n133, n134, n135, n136, n137, n138, n139,
 n140, n141, n142, n143, n144, n145, n146, n147,
 n148, n149, n150, n151, n152, n153, n154, n155,
 n156, n157, n158, n159, n160, n161, n162, n163,
 n164, n165, n166, n167, n168, n169, n170, n171,
 n172, n173, n174, n175, n176, n177, n178, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n189, n190, n191, n192, n193, n194, n195,
 n196, n197, n198, n199, n200, n201, n202, n203,
 n204, n205, n206, n207, n208, n209, n210, n211,
 n212, n213, n214, n215, n216, n217, n218, n219,
 n220, n221, n222, n223, n224, n225, n226, n227,
 n228, n229, n230, n231, n232, n233, n234, n235,
 n236, n237, n238, n239, n240, n241, n242, n243,
 n244, n245, n246, n247, n248, n249, n250, n251,
 n252, n253, n254, n255, n256, n257, n258, n259,
 n260, n261, n262, n263, n264, n265, n266, n267,
 n268, n269, n270, n271, n272, n273, n274, n275,
 n276, n277, n278, n279, n280, n281, n282, n283,
 n284, n285, n286, n287, n288, n289, n290, n291,
 n292, n293, n294, n295, n296, n297, n298, n299,
 n300, n301, n302, n303, n304, n305, n306, n307,
 n308, n309, n310, n311, n312, n313, n314, n315,
 n316, n317, n318, n319, n320, n321, n322, n323,
 n324, n325, n326, n327, n328, n329, n330, n331,
 n332, n333, n334, n335, n336, n337, n338, n339,
 n340, n341, n342, n343, n344, n345, n346, n347,
 n348, n349, n350, n351, n352, n353, n354, n355,
 n356, n357, n358, n359, n360, n361, n362, n363,
 n364, n365, n366, n367, n368, n369, n370, n371,
 n372, n373, n374, n375, n376, n377, n378, n379,
 n380, n381, n382, n383, n384, n385, n386, n387,
 n388, n389, n390, n391, n392, n393, n394, n395,
 n396, n397, n398, n399, n400, n401, n402, n403,
 n404, n405, n406, n407, n408, n409, n410, n411,
 n412, n413, n414, n415, n416, n417, n418, n419,
 n420, n421, n422, n423, n424, n425, n426, n427,
 n428, n429, n430, n431, n432, n433, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n571,
 n572, n573, n574, n575, n576, n577, n578, n579,
 n580, n581, n582, n583, n584, n585, n586, n587,
 n588, n589, n590, n591, n592, n593, n594, n595,
 n596, n597, n598, n599, n600, n601, n602, n603,
 n604, n605, n606, n607, n608, n609, n610, n611,
 n612, n613, n614, n615, n616, n617, n618, n619,
 n620, n621, n622, n623, n624, n625, n626, n627,
 n628, n629, n630, n631, n632, n633, n634, n635,
 n636, n637, n638, n639, n640, n641, n642, n643,
 n644, n645, n646, n647, n648, n649, n650, n651,
 n652, n653, n654, n655, n656, n657, n658, n659,
 n660, n661, n662, n663, n664, n665, n666, n667,
 n668, n669, n670, n671, n672, n673, n674, n675,
 n676, n677, n678, n679, n680, n681, n682, n683,
 n684, n685, n686, n687, n688, n690, n691, n692,
 n694, n695, n696, n697, n699, n700, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735,
 n736, n737, n738, n739, n740, n741, n742, n743,
 n744, n745, n746, n747, n748, n749, n750, n751,
 n752, n753, n754, n755, n756, n757, n758, n759,
 n760, n761, n762, n763, n764, n765, n766, n767,
 n768, n769, n770, n771, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818;

not  g0 (n80, n8);
buf  g1 (n119, n16);
not  g2 (n123, n5);
not  g3 (n74, n23);
buf  g4 (n88, n8);
not  g5 (n77, n9);
not  g6 (n107, n12);
not  g7 (n47, n5);
buf  g8 (n70, n18);
buf  g9 (n65, n4);
not  g10 (n97, n3);
not  g11 (n46, n12);
buf  g12 (n98, n6);
buf  g13 (n109, n24);
buf  g14 (n55, n14);
not  g15 (n35, n7);
buf  g16 (n89, n10);
buf  g17 (n58, n2);
buf  g18 (n45, n6);
not  g19 (n114, n22);
not  g20 (n39, n2);
buf  g21 (n76, n21);
buf  g22 (n108, n8);
not  g23 (n78, n6);
not  g24 (n53, n14);
not  g25 (n103, n15);
buf  g26 (n106, n14);
buf  g27 (n44, n2);
not  g28 (n82, n6);
not  g29 (n68, n10);
buf  g30 (n41, n1);
buf  g31 (n50, n11);
not  g32 (n96, n13);
not  g33 (n36, n7);
not  g34 (n59, n10);
not  g35 (n75, n13);
not  g36 (n126, n22);
not  g37 (n85, n25);
not  g38 (n64, n16);
buf  g39 (n63, n17);
not  g40 (n118, n9);
buf  g41 (n71, n15);
not  g42 (n81, n23);
buf  g43 (n51, n21);
buf  g44 (n124, n12);
not  g45 (n69, n18);
not  g46 (n56, n24);
buf  g47 (n60, n12);
buf  g48 (n113, n2);
not  g49 (n62, n23);
buf  g50 (n94, n19);
buf  g51 (n30, n1);
not  g52 (n110, n21);
buf  g53 (n48, n20);
not  g54 (n117, n4);
buf  g55 (n112, n10);
buf  g56 (n105, n1);
not  g57 (n66, n13);
not  g58 (n52, n20);
not  g59 (n57, n4);
buf  g60 (n91, n17);
buf  g61 (n61, n4);
buf  g62 (n84, n19);
buf  g63 (n54, n13);
not  g64 (n121, n16);
buf  g65 (n125, n17);
buf  g66 (n33, n7);
buf  g67 (n42, n7);
buf  g68 (n86, n9);
not  g69 (n83, n18);
not  g70 (n40, n3);
not  g71 (n31, n5);
buf  g72 (n73, n19);
buf  g73 (n95, n3);
buf  g74 (n90, n11);
not  g75 (n122, n20);
buf  g76 (n92, n25);
not  g77 (n93, n15);
buf  g78 (n120, n19);
not  g79 (n34, n17);
not  g80 (n115, n8);
not  g81 (n37, n21);
buf  g82 (n87, n20);
buf  g83 (n67, n15);
not  g84 (n43, n23);
buf  g85 (n100, n11);
buf  g86 (n72, n14);
buf  g87 (n101, n24);
buf  g88 (n29, n16);
not  g89 (n99, n1);
not  g90 (n104, n24);
buf  g91 (n32, n9);
not  g92 (n116, n11);
buf  g93 (n111, n3);
not  g94 (n49, n5);
not  g95 (n28, n22);
not  g96 (n79, n18);
buf  g97 (n102, n25);
buf  g98 (n38, n22);
buf  g99 (n169, n29);
buf  g100 (n394, n30);
buf  g101 (n207, n43);
buf  g102 (n349, n67);
buf  g103 (n320, n54);
buf  g104 (n202, n50);
buf  g105 (n257, n40);
not  g106 (n290, n55);
not  g107 (n385, n84);
buf  g108 (n301, n89);
not  g109 (n263, n97);
not  g110 (n162, n32);
buf  g111 (n293, n42);
not  g112 (n152, n97);
buf  g113 (n265, n44);
buf  g114 (n194, n40);
not  g115 (n363, n60);
not  g116 (n333, n79);
buf  g117 (n184, n64);
buf  g118 (n392, n96);
not  g119 (n187, n36);
not  g120 (n221, n93);
buf  g121 (n168, n89);
buf  g122 (n277, n38);
not  g123 (n155, n71);
buf  g124 (n182, n93);
not  g125 (n241, n88);
buf  g126 (n356, n30);
buf  g127 (n147, n82);
buf  g128 (n315, n79);
buf  g129 (n188, n67);
buf  g130 (n171, n72);
not  g131 (n195, n43);
buf  g132 (n170, n59);
buf  g133 (n238, n38);
buf  g134 (n179, n82);
buf  g135 (n323, n34);
not  g136 (n208, n73);
buf  g137 (n218, n32);
buf  g138 (n390, n68);
not  g139 (n410, n44);
not  g140 (n236, n48);
not  g141 (n283, n56);
not  g142 (n159, n76);
not  g143 (n373, n37);
buf  g144 (n177, n29);
buf  g145 (n205, n92);
buf  g146 (n346, n31);
buf  g147 (n369, n57);
buf  g148 (n300, n79);
not  g149 (n381, n99);
buf  g150 (n371, n67);
not  g151 (n364, n57);
buf  g152 (n255, n75);
buf  g153 (n359, n60);
not  g154 (n312, n83);
not  g155 (n294, n55);
buf  g156 (n134, n74);
not  g157 (n271, n31);
not  g158 (n180, n42);
buf  g159 (n299, n95);
buf  g160 (n386, n78);
not  g161 (n302, n40);
buf  g162 (n193, n72);
buf  g163 (n225, n80);
not  g164 (n228, n87);
buf  g165 (n328, n54);
buf  g166 (n166, n37);
buf  g167 (n370, n65);
buf  g168 (n259, n57);
not  g169 (n274, n45);
not  g170 (n230, n92);
buf  g171 (n137, n52);
buf  g172 (n128, n99);
not  g173 (n192, n58);
not  g174 (n148, n88);
buf  g175 (n295, n72);
not  g176 (n181, n32);
buf  g177 (n269, n61);
buf  g178 (n209, n30);
not  g179 (n270, n46);
buf  g180 (n331, n40);
buf  g181 (n150, n33);
not  g182 (n136, n94);
not  g183 (n264, n96);
buf  g184 (n345, n69);
not  g185 (n232, n53);
buf  g186 (n223, n88);
buf  g187 (n324, n58);
buf  g188 (n282, n48);
buf  g189 (n336, n62);
buf  g190 (n178, n98);
not  g191 (n298, n69);
not  g192 (n142, n39);
not  g193 (n332, n80);
not  g194 (n379, n78);
buf  g195 (n201, n28);
not  g196 (n376, n73);
not  g197 (n189, n63);
buf  g198 (n206, n35);
buf  g199 (n245, n66);
buf  g200 (n297, n87);
buf  g201 (n317, n61);
buf  g202 (n341, n87);
buf  g203 (n243, n54);
buf  g204 (n186, n33);
buf  g205 (n174, n67);
buf  g206 (n337, n35);
not  g207 (n139, n49);
not  g208 (n304, n97);
buf  g209 (n289, n29);
buf  g210 (n404, n86);
buf  g211 (n260, n65);
buf  g212 (n343, n95);
buf  g213 (n327, n77);
not  g214 (n316, n83);
not  g215 (n211, n37);
not  g216 (n391, n32);
buf  g217 (n130, n70);
buf  g218 (n388, n46);
not  g219 (n144, n82);
buf  g220 (n314, n56);
buf  g221 (n351, n91);
buf  g222 (n262, n37);
buf  g223 (n239, n63);
buf  g224 (n254, n92);
buf  g225 (n272, n55);
buf  g226 (n131, n50);
buf  g227 (n335, n91);
not  g228 (n368, n84);
buf  g229 (n252, n47);
buf  g230 (n402, n96);
not  g231 (n354, n74);
not  g232 (n309, n46);
buf  g233 (n384, n33);
buf  g234 (n286, n77);
not  g235 (n242, n85);
not  g236 (n375, n28);
not  g237 (n244, n63);
buf  g238 (n352, n91);
not  g239 (n382, n47);
buf  g240 (n220, n90);
buf  g241 (n306, n80);
buf  g242 (n378, n78);
not  g243 (n361, n85);
buf  g244 (n258, n34);
buf  g245 (n129, n49);
not  g246 (n231, n98);
buf  g247 (n200, n75);
buf  g248 (n401, n99);
not  g249 (n127, n45);
not  g250 (n279, n86);
not  g251 (n350, n41);
buf  g252 (n355, n66);
buf  g253 (n338, n45);
buf  g254 (n342, n96);
buf  g255 (n387, n34);
buf  g256 (n374, n51);
buf  g257 (n226, n63);
buf  g258 (n339, n42);
buf  g259 (n308, n60);
not  g260 (n393, n36);
not  g261 (n249, n45);
not  g262 (n358, n82);
buf  g263 (n311, n60);
buf  g264 (n197, n71);
not  g265 (n222, n53);
not  g266 (n367, n59);
buf  g267 (n268, n38);
buf  g268 (n141, n94);
not  g269 (n247, n41);
buf  g270 (n140, n34);
buf  g271 (n348, n66);
buf  g272 (n353, n39);
buf  g273 (n253, n69);
not  g274 (n227, n90);
not  g275 (n303, n64);
not  g276 (n413, n95);
not  g277 (n248, n98);
buf  g278 (n234, n68);
buf  g279 (n411, n81);
buf  g280 (n143, n52);
not  g281 (n377, n92);
buf  g282 (n278, n64);
buf  g283 (n344, n79);
buf  g284 (n198, n84);
not  g285 (n204, n93);
buf  g286 (n276, n81);
not  g287 (n224, n85);
not  g288 (n291, n56);
buf  g289 (n135, n59);
buf  g290 (n365, n66);
not  g291 (n360, n71);
not  g292 (n172, n33);
buf  g293 (n305, n81);
buf  g294 (n214, n53);
not  g295 (n215, n70);
not  g296 (n176, n65);
buf  g297 (n330, n89);
buf  g298 (n389, n51);
not  g299 (n213, n77);
not  g300 (n167, n86);
not  g301 (n199, n52);
buf  g302 (n149, n43);
not  g303 (n267, n28);
buf  g304 (n372, n38);
buf  g305 (n325, n89);
not  g306 (n395, n98);
buf  g307 (n326, n83);
not  g308 (n321, n83);
not  g309 (n292, n46);
buf  g310 (n400, n95);
not  g311 (n318, n47);
not  g312 (n246, n36);
buf  g313 (n133, n30);
buf  g314 (n396, n44);
not  g315 (n157, n74);
not  g316 (n217, n58);
not  g317 (n319, n50);
buf  g318 (n409, n76);
buf  g319 (n240, n55);
not  g320 (n380, n76);
not  g321 (n307, n29);
not  g322 (n407, n31);
buf  g323 (n256, n41);
buf  g324 (n160, n64);
buf  g325 (n273, n70);
buf  g326 (n158, n77);
buf  g327 (n237, n36);
buf  g328 (n163, n80);
buf  g329 (n313, n62);
not  g330 (n196, n58);
buf  g331 (n164, n59);
buf  g332 (n357, n97);
not  g333 (n412, n73);
buf  g334 (n183, n93);
not  g335 (n347, n49);
buf  g336 (n175, n81);
not  g337 (n132, n68);
not  g338 (n296, n88);
not  g339 (n154, n90);
buf  g340 (n173, n90);
not  g341 (n287, n91);
buf  g342 (n190, n28);
not  g343 (n185, n68);
not  g344 (n405, n73);
buf  g345 (n281, n48);
buf  g346 (n310, n51);
buf  g347 (n146, n53);
not  g348 (n235, n85);
not  g349 (n250, n44);
not  g350 (n251, n69);
buf  g351 (n153, n54);
not  g352 (n329, n78);
not  g353 (n275, n94);
buf  g354 (n340, n31);
not  g355 (n156, n75);
buf  g356 (n399, n94);
not  g357 (n145, n41);
buf  g358 (n216, n61);
not  g359 (n151, n86);
not  g360 (n233, n65);
not  g361 (n261, n43);
buf  g362 (n219, n39);
buf  g363 (n266, n35);
buf  g364 (n408, n70);
not  g365 (n285, n47);
buf  g366 (n229, n49);
not  g367 (n210, n57);
not  g368 (n203, n84);
buf  g369 (n288, n74);
buf  g370 (n334, n52);
not  g371 (n280, n50);
not  g372 (n138, n56);
buf  g373 (n322, n51);
not  g374 (n284, n35);
not  g375 (n406, n76);
buf  g376 (n191, n75);
buf  g377 (n165, n61);
not  g378 (n212, n62);
not  g379 (n362, n71);
buf  g380 (n366, n62);
buf  g381 (n398, n72);
buf  g382 (n383, n48);
buf  g383 (n397, n87);
not  g384 (n161, n39);
buf  g385 (n403, n42);
not  g386 (n430, n146);
not  g387 (n423, n135);
not  g388 (n431, n147);
buf  g389 (n429, n151);
not  g390 (n433, n152);
buf  g391 (n421, n150);
buf  g392 (n434, n145);
buf  g393 (n426, n133);
buf  g394 (n422, n130);
buf  g395 (n424, n134);
not  g396 (n436, n140);
not  g397 (n419, n144);
buf  g398 (n427, n138);
buf  g399 (n414, n132);
buf  g400 (n420, n129);
not  g401 (n435, n128);
buf  g402 (n428, n137);
not  g403 (n432, n131);
not  g404 (n416, n142);
not  g405 (n417, n136);
buf  g406 (n439, n149);
not  g407 (n425, n143);
buf  g408 (n418, n141);
buf  g409 (n437, n127);
buf  g410 (n438, n148);
buf  g411 (n415, n139);
nand g412 (n474, n260, n177, n174, n197);
xnor g413 (n452, n239, n195, n266, n262);
xnor g414 (n533, n416, n155, n275, n425);
nand g415 (n524, n194, n284, n298, n430);
nor  g416 (n503, n314, n183, n180, n298);
or   g417 (n527, n269, n208, n251, n415);
xor  g418 (n455, n237, n244, n204, n270);
nor  g419 (n448, n295, n242, n250, n189);
xnor g420 (n479, n314, n429, n425, n439);
xor  g421 (n523, n253, n424, n265);
nor  g422 (n511, n302, n437, n428, n198);
xor  g423 (n493, n286, n291, n236, n312);
and  g424 (n463, n437, n249, n303, n438);
xor  g425 (n505, n272, n190, n431, n280);
nand g426 (n506, n309, n426, n157, n219);
xor  g427 (n520, n222, n434, n303, n240);
xnor g428 (n515, n256, n214, n185, n300);
nor  g429 (n532, n229, n289, n206, n249);
nand g430 (n528, n436, n275, n420, n418);
and  g431 (n489, n223, n247, n189, n284);
xor  g432 (n540, n311, n156, n435, n287);
or   g433 (n497, n420, n239, n294, n283);
xor  g434 (n501, n228, n261, n205, n252);
xor  g435 (n539, n216, n260, n419, n425);
nor  g436 (n480, n267, n301, n203, n432);
xor  g437 (n478, n273, n261, n299, n256);
and  g438 (n471, n271, n282, n428, n186);
nand g439 (n459, n422, n164, n304, n424);
and  g440 (n472, n431, n163, n423, n427);
xor  g441 (n457, n418, n417, n192, n421);
and  g442 (n498, n421, n251, n434, n230);
and  g443 (n488, n192, n435, n224, n198);
or   g444 (n473, n180, n272, n226, n199);
nand g445 (n494, n181, n268, n175, n211);
or   g446 (n442, n209, n212, n219, n439);
nor  g447 (n504, n221, n201, n278, n257);
xor  g448 (n484, n305, n211, n214, n171);
or   g449 (n451, n286, n264, n296, n419);
nand g450 (n537, n215, n193, n207, n288);
xnor g451 (n464, n308, n292, n429, n433);
or   g452 (n477, n308, n416, n306, n297);
nor  g453 (n519, n184, n154, n310, n199);
xor  g454 (n440, n184, n257, n422, n235);
xnor g455 (n486, n414, n196, n438, n417);
and  g456 (n460, n233, n267, n208, n244);
xnor g457 (n514, n283, n417, n234, n217);
xor  g458 (n444, n315, n188, n187, n289);
xor  g459 (n453, n414, n243, n161, n202);
nand g460 (n535, n241, n427, n309, n224);
nand g461 (n462, n271, n282, n218, n212);
nand g462 (n482, n246, n248, n238, n172);
and  g463 (n443, n312, n229, n253, n436);
or   g464 (n513, n299, n302, n158, n430);
xor  g465 (n529, n194, n420, n285, n290);
and  g466 (n526, n296, n434, n414, n221);
xnor g467 (n500, n162, n170, n429, n255);
nand g468 (n490, n281, n245, n231, n220);
xnor g469 (n456, n218, n174, n277, n424);
xor  g470 (n491, n231, n259, n238, n290);
xor  g471 (n447, n181, n175, n255, n429);
xnor g472 (n485, n297, n268, n422, n307);
or   g473 (n475, n300, n213, n421, n227);
nor  g474 (n454, n292, n311, n258, n165);
nand g475 (n517, n226, n263, n415, n168);
xor  g476 (n522, n177, n414, n423, n313);
nor  g477 (n487, n438, n430, n188, n160);
nand g478 (n458, n201, n243, n195, n313);
xor  g479 (n510, n416, n439, n274, n437);
or   g480 (n468, n295, n420, n426, n173);
xor  g481 (n534, n310, n285, n276, n258);
nand g482 (n446, n179, n437, n436, n259);
nand g483 (n481, n287, n232, n432, n204);
xor  g484 (n538, n305, n430, n190, n423);
xor  g485 (n507, n217, n176, n433, n419);
xnor g486 (n465, n193, n222, n435, n307);
xnor g487 (n469, n171, n247, n206, n438);
nand g488 (n441, n209, n215, n252, n235);
xnor g489 (n450, n236, n182, n187, n197);
xor  g490 (n525, n233, n280, n225);
xnor g491 (n512, n270, n200, n427, n168);
nand g492 (n449, n248, n419, n428, n427);
xnor g493 (n516, n418, n265, n254, n220);
and  g494 (n461, n207, n263, n281, n415);
xor  g495 (n483, n432, n433, n426, n173);
nor  g496 (n508, n200, n432, n277, n227);
nand g497 (n530, n279, n417, n264, n433);
nor  g498 (n531, n416, n273, n304, n237);
nor  g499 (n496, n415, n216, n223, n178);
nand g500 (n521, n316, n426, n170, n254);
nand g501 (n541, n288, n202, n182, n436);
xnor g502 (n467, n279, n178, n291, n191);
nor  g503 (n542, n269, n210, n169, n153);
or   g504 (n470, n274, n439, n431, n230);
nand g505 (n518, n418, n262, n250, n306);
nor  g506 (n543, n205, n213, n293, n241);
xnor g507 (n492, n431, n266, n293, n245);
xor  g508 (n466, n242, n176, n191, n435);
nand g509 (n495, n172, n232, n315, n159);
nand g510 (n445, n183, n246, n278, n425);
xor  g511 (n476, n434, n179, n196, n240);
nor  g512 (n499, n203, n186, n234, n167);
xor  g513 (n536, n423, n428, n185, n166);
nor  g514 (n509, n210, n421, n422, n301);
xor  g515 (n502, n276, n294, n228, n169);
xnor g516 (n555, n354, n352, n344, n391);
nor  g517 (n582, n354, n515, n377, n364);
or   g518 (n561, n376, n383, n351, n346);
nor  g519 (n571, n368, n106, n350, n324);
xor  g520 (n605, n497, n319, n512, n378);
and  g521 (n576, n443, n375, n385, n387);
xor  g522 (n595, n485, n363, n110, n530);
xor  g523 (n622, n338, n471, n362, n389);
nand g524 (n577, n379, n331, n455, n366);
nand g525 (n620, n382, n101, n339, n104);
xnor g526 (n628, n349, n518, n331, n453);
xnor g527 (n592, n357, n488, n379, n343);
xnor g528 (n560, n344, n531, n350, n353);
xnor g529 (n544, n441, n475, n109, n354);
nand g530 (n631, n384, n360, n377, n380);
and  g531 (n606, n342, n377, n393, n379);
xor  g532 (n642, n395, n338, n348, n26);
xnor g533 (n565, n365, n322, n492, n347);
xnor g534 (n645, n348, n371, n355, n326);
xor  g535 (n636, n364, n371, n365, n388);
nor  g536 (n640, n496, n318, n105, n389);
or   g537 (n545, n337, n337, n26, n528);
nor  g538 (n619, n508, n370, n527, n449);
nor  g539 (n617, n447, n369, n103, n363);
or   g540 (n648, n457, n330, n339, n483);
nand g541 (n625, n371, n387, n341, n110);
and  g542 (n610, n394, n327, n108, n516);
nand g543 (n553, n395, n359, n342);
xor  g544 (n623, n456, n459, n26, n350);
xnor g545 (n575, n392, n340, n376, n393);
xnor g546 (n566, n516, n349, n332, n345);
xnor g547 (n594, n355, n355, n372, n526);
or   g548 (n638, n329, n317, n476, n370);
xnor g549 (n562, n506, n386, n390, n323);
xor  g550 (n643, n364, n382, n336, n387);
xor  g551 (n614, n366, n332, n358, n464);
nand g552 (n556, n369, n329, n375, n491);
xor  g553 (n651, n100, n463, n384, n520);
nand g554 (n599, n367, n525, n379, n460);
nand g555 (n586, n360, n102, n372, n345);
xnor g556 (n591, n451, n502, n360, n322);
nand g557 (n564, n361, n321, n27, n100);
or   g558 (n615, n111, n509, n360, n378);
xor  g559 (n548, n477, n347, n353, n361);
and  g560 (n621, n388, n524, n325, n101);
nor  g561 (n583, n388, n376, n389, n366);
nor  g562 (n629, n381, n103, n521, n442);
and  g563 (n585, n380, n383, n320, n343);
xor  g564 (n587, n374, n378, n371, n394);
nor  g565 (n637, n351, n501, n390, n367);
or   g566 (n641, n481, n390, n363, n366);
xor  g567 (n616, n529, n107, n462, n368);
and  g568 (n611, n106, n469, n356, n522);
nor  g569 (n581, n498, n350, n394, n367);
nor  g570 (n633, n385, n383, n382, n102);
xor  g571 (n563, n334, n104, n386, n482);
nand g572 (n613, n520, n103, n359, n109);
nand g573 (n546, n103, n369, n109, n110);
or   g574 (n653, n357, n487, n110, n356);
and  g575 (n632, n364, n474, n374, n381);
nor  g576 (n549, n368, n374, n479, n104);
and  g577 (n644, n107, n109, n522, n333);
xnor g578 (n590, n383, n388, n466, n344);
xor  g579 (n574, n510, n27, n472, n377);
or   g580 (n552, n486, n100, n105, n529);
xnor g581 (n607, n374, n448, n523, n384);
xnor g582 (n551, n393, n357, n367, n362);
and  g583 (n650, n27, n323, n320, n339);
and  g584 (n600, n351, n505, n528, n499);
xor  g585 (n646, n369, n445, n342, n348);
and  g586 (n593, n381, n467, n99, n25);
or   g587 (n559, n345, n317, n513, n484);
nor  g588 (n627, n465, n111, n328, n341);
nand g589 (n649, n444, n100, n343, n346);
or   g590 (n626, n385, n517, n380, n500);
nand g591 (n580, n382, n511, n515, n346);
xnor g592 (n608, n328, n391, n346, n375);
and  g593 (n579, n373, n358, n504, n490);
and  g594 (n618, n394, n321, n334, n513);
xnor g595 (n654, n461, n108, n386, n530);
xnor g596 (n567, n356, n495, n335, n378);
nand g597 (n647, n519, n106, n478, n503);
and  g598 (n630, n392, n108, n390, n352);
and  g599 (n554, n395, n348, n393, n102);
and  g600 (n558, n341, n343, n26, n318);
xnor g601 (n550, n362, n365, n470, n458);
nor  g602 (n609, n356, n27, n353, n384);
nor  g603 (n584, n494, n370, n440);
and  g604 (n604, n101, n373, n518, n514);
and  g605 (n603, n352, n396, n480, n108);
xor  g606 (n588, n392, n351, n361, n347);
nor  g607 (n547, n523, n316, n368, n373);
and  g608 (n573, n473, n330, n358, n333);
or   g609 (n568, n362, n335, n373, n391);
nand g610 (n602, n326, n372, n489, n386);
nand g611 (n639, n358, n363, n340, n519);
nand g612 (n570, n454, n507, n359, n396);
xnor g613 (n598, n352, n353, n385, n517);
xnor g614 (n589, n340, n375, n395, n355);
and  g615 (n652, n327, n349, n340, n101);
xor  g616 (n578, n372, n347, n102, n106);
xor  g617 (n557, n514, n446, n392, n338);
and  g618 (n601, n468, n349, n380, n341);
xor  g619 (n597, n105, n450, n339, n493);
nor  g620 (n569, n357, n521, n525, n107);
nor  g621 (n612, n381, n361, n526, n325);
xnor g622 (n596, n512, n345, n111, n365);
xor  g623 (n572, n376, n319, n391, n336);
xnor g624 (n634, n387, n105, n524, n104);
xnor g625 (n624, n107, n359, n324, n354);
or   g626 (n635, n344, n452, n389, n527);
not  g627 (n658, n531);
not  g628 (n661, n548);
buf  g629 (n657, n546);
buf  g630 (n656, n549);
buf  g631 (n660, n532);
not  g632 (n659, n547);
nand g633 (n655, n550, n545, n544);
and  g634 (n681, n597, n556, n575, n587);
or   g635 (n679, n631, n623, n574, n657);
or   g636 (n676, n613, n571, n581, n582);
xnor g637 (n684, n660, n658, n661, n553);
nor  g638 (n685, n551, n660, n594, n656);
nor  g639 (n678, n656, n555, n657, n585);
nor  g640 (n675, n554, n628, n611, n626);
xnor g641 (n669, n624, n655, n615, n608);
or   g642 (n677, n593, n614, n592, n603);
xnor g643 (n687, n604, n589, n620, n625);
nor  g644 (n664, n655, n606, n661, n612);
nor  g645 (n667, n568, n569, n618, n591);
nor  g646 (n672, n610, n605, n659, n599);
nand g647 (n662, n588, n561, n564, n590);
nor  g648 (n673, n629, n570, n661, n659);
nor  g649 (n682, n622, n660, n563, n627);
nor  g650 (n668, n562, n572, n578, n558);
nor  g651 (n674, n583, n657, n566, n658);
nor  g652 (n671, n621, n576, n602, n586);
nor  g653 (n688, n661, n552, n658, n573);
nor  g654 (n680, n656, n560, n617, n616);
nor  g655 (n666, n565, n658, n584, n656);
or   g656 (n670, n657, n601, n659, n579);
xor  g657 (n686, n609, n596, n580, n660);
xnor g658 (n663, n655, n607, n577, n630);
and  g659 (n665, n595, n619, n600, n598);
nand g660 (n683, n559, n557, n659, n567);
or   g661 (n692, n119, n121, n115, n117);
or   g662 (n707, n113, n116, n124, n125);
nor  g663 (n703, n663, n117, n673, n675);
and  g664 (n701, n664, n118, n122);
or   g665 (n697, n114, n669, n119, n112);
or   g666 (n696, n114, n668, n676, n124);
nand g667 (n689, n121, n125, n117, n111);
or   g668 (n700, n676, n120, n118);
nor  g669 (n690, n676, n113, n122, n123);
xnor g670 (n698, n674, n119, n662, n123);
or   g671 (n704, n121, n671, n675, n126);
and  g672 (n693, n123, n118, n121, n122);
nand g673 (n705, n115, n113, n125);
nor  g674 (n691, n124, n114, n675, n115);
xor  g675 (n702, n120, n113, n666, n124);
nor  g676 (n708, n118, n114, n119, n672);
and  g677 (n694, n670, n675, n126, n120);
or   g678 (n699, n123, n116, n665, n112);
nand g679 (n706, n117, n116, n115);
xor  g680 (n695, n667, n126, n112);
xor  g681 (n721, n397, n402, n406, n696);
xor  g682 (n722, n404, n407, n400, n697);
xor  g683 (n710, n399, n397, n404, n401);
nand g684 (n718, n703, n398, n400);
or   g685 (n712, n405, n396, n403, n401);
or   g686 (n717, n702, n397, n407, n398);
nor  g687 (n719, n399, n706, n701, n407);
nand g688 (n711, n406, n707, n705, n397);
and  g689 (n724, n400, n398, n403);
or   g690 (n723, n694, n399, n396, n402);
nor  g691 (n716, n402, n693, n403, n404);
nand g692 (n713, n708, n408, n699);
xor  g693 (n714, n399, n401, n406, n700);
xor  g694 (n720, n406, n698, n405);
and  g695 (n709, n407, n404, n402, n405);
xor  g696 (n715, n695, n401, n704, n403);
nor  g697 (n726, n649, n648, n640, n652);
nor  g698 (n725, n635, n710, n643);
nor  g699 (n727, n642, n710, n709);
nand g700 (n729, n632, n650, n637, n647);
or   g701 (n728, n645, n646, n641, n638);
or   g702 (n730, n636, n644, n709);
nand g703 (n731, n634, n651, n633, n639);
nand g704 (n741, n717, n718, n728, n713);
xnor g705 (n742, n713, n716, n711, n712);
nand g706 (n733, n717, n716, n729, n712);
nand g707 (n734, n717, n711, n712, n728);
xnor g708 (n732, n714, n717, n715, n716);
xor  g709 (n737, n718, n714, n729);
nand g710 (n735, n718, n713, n719, n726);
nand g711 (n739, n715, n725, n727, n714);
nand g712 (n738, n712, n715, n711, n718);
nor  g713 (n740, n711, n727, n728);
nand g714 (n736, n713, n715, n728, n716);
and  g715 (n743, n680, n409, n734, n679);
xor  g716 (n749, n680, n678, n677);
nand g717 (n748, n678, n408, n679);
xnor g718 (n747, n737, n680, n677);
and  g719 (n745, n735, n678, n733, n732);
xor  g720 (n746, n677, n681, n676, n738);
or   g721 (n744, n736, n679, n408, n680);
nand g722 (n753, n744, n739, n748, n533);
xnor g723 (n752, n742, n721, n740, n720);
xnor g724 (n751, n746, n719, n721);
xnor g725 (n750, n533, n743, n720, n719);
xnor g726 (n755, n741, n720, n745, n747);
and  g727 (n754, n721, n719, n720, n532);
xor  g728 (n758, n681, n682, n752);
nor  g729 (n756, n750, n681, n722);
nand g730 (n757, n683, n751, n682);
and  g731 (n760, n757, n730);
xnor g732 (n759, n729, n729, n730, n756);
xnor g733 (n762, n723, n723, n760, n722);
nor  g734 (n761, n722, n759, n760, n723);
nor  g735 (n763, n722, n724, n723);
buf  g736 (n770, n761);
not  g737 (n766, n731);
not  g738 (n764, n762);
buf  g739 (n769, n731);
buf  g740 (n768, n731);
buf  g741 (n773, n762);
not  g742 (n772, n749);
and  g743 (n765, n683, n763, n731);
xnor g744 (n767, n763, n761, n762);
nor  g745 (n771, n762, n763);
not  g746 (n775, n764);
not  g747 (n774, n764);
xnor g748 (n779, n774, n765, n764, n769);
xnor g749 (n776, n766, n766, n775, n768);
or   g750 (n783, n768, n766, n765, n774);
nor  g751 (n778, n765, n766, n768, n764);
xnor g752 (n780, n774, n724, n767, n775);
nand g753 (n781, n767, n767, n768, n774);
or   g754 (n782, n775, n769, n767);
nor  g755 (n777, n769, n765, n775, n724);
not  g756 (n791, n410);
not  g757 (n792, n410);
not  g758 (n786, n412);
buf  g759 (n790, n779);
nand g760 (n785, n778, n776, n409, n410);
or   g761 (n788, n412, n411, n780, n409);
or   g762 (n789, n781, n411, n779);
nand g763 (n787, n778, n410, n412, n777);
nand g764 (n784, n780, n409, n412, n411);
buf  g765 (n793, n784);
not  g766 (n794, n784);
or   g767 (n795, n794, n413);
xnor g768 (n796, n755, n654, n795, n753);
nor  g769 (n797, n653, n795, n758, n754);
xnor g770 (n798, n796, n770);
or   g771 (n799, n798, n786, n787);
xnor g772 (n801, n787, n788, n798, n786);
nand g773 (n800, n787, n786, n785);
nor  g774 (n802, n797, n798, n788);
or   g775 (n816, n536, n802, n535, n543);
nand g776 (n803, n540, n771, n537, n782);
and  g777 (n813, n538, n772, n801);
nand g778 (n804, n802, n773, n684, n800);
xor  g779 (n814, n772, n799, n800);
and  g780 (n818, n537, n536, n540, n800);
nand g781 (n805, n541, n773, n126, n535);
nor  g782 (n808, n801, n685, n772, n534);
nand g783 (n812, n771, n802, n801, n799);
nand g784 (n806, n771, n538, n683, n782);
xor  g785 (n809, n781, n542, n771);
xor  g786 (n815, n772, n543, n539, n773);
or   g787 (n817, n413, n684);
xor  g788 (n810, n683, n800, n799, n770);
and  g789 (n807, n534, n802, n685, n539);
xnor g790 (n811, n685, n541, n783);
or   g791 (n820, n810, n773, n807, n804);
and  g792 (n819, n811, n791, n688, n790);
nor  g793 (n826, n688, n685, n791, n818);
nand g794 (n821, n803, n790, n686, n687);
xnor g795 (n829, n792, n687, n791);
xnor g796 (n828, n815, n817, n788, n790);
or   g797 (n822, n790, n688, n687, n792);
xnor g798 (n830, n805, n816, n789, n791);
nor  g799 (n827, n808, n686, n789, n792);
or   g800 (n824, n792, n813, n812, n789);
or   g801 (n823, n688, n788, n789, n809);
nand g802 (n825, n686, n686, n814, n806);
endmodule
