

module Stat_1443_32_4
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n947,
  n950,
  n940,
  n948,
  n949,
  n941,
  n945,
  n942,
  n939,
  n943,
  n946,
  n958,
  n1461,
  n1465,
  n1471,
  n1468,
  n1469,
  n1470,
  n1459,
  n1466,
  n1457,
  n1463,
  n1464,
  n1458,
  n1467,
  n1472,
  n1460,
  n1462,
  n1473
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n947;output n950;output n940;output n948;output n949;output n941;output n945;output n942;output n939;output n943;output n946;output n958;output n1461;output n1465;output n1471;output n1468;output n1469;output n1470;output n1459;output n1466;output n1457;output n1463;output n1464;output n1458;output n1467;output n1472;output n1460;output n1462;output n1473;
  wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n944;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyNOTWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyNOTWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyNOTWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyNOTWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyNOTWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    n52,
    n21
  );


  buf
  g1
  (
    n88,
    n23
  );


  buf
  g2
  (
    n100,
    n28
  );


  not
  g3
  (
    n65,
    n27
  );


  buf
  g4
  (
    n113,
    n1
  );


  not
  g5
  (
    n61,
    n5
  );


  not
  g6
  (
    n83,
    n22
  );


  not
  g7
  (
    n59,
    n7
  );


  not
  g8
  (
    n120,
    n6
  );


  not
  g9
  (
    n45,
    n14
  );


  buf
  g10
  (
    n69,
    n9
  );


  not
  g11
  (
    n44,
    n11
  );


  not
  g12
  (
    n121,
    n11
  );


  not
  g13
  (
    n87,
    n21
  );


  buf
  g14
  (
    n105,
    n8
  );


  not
  g15
  (
    n108,
    n29
  );


  buf
  g16
  (
    n99,
    n30
  );


  buf
  g17
  (
    KeyWire_0_25,
    n29
  );


  not
  g18
  (
    n118,
    n1
  );


  buf
  g19
  (
    n126,
    n18
  );


  not
  g20
  (
    n149,
    n6
  );


  buf
  g21
  (
    n48,
    n26
  );


  not
  g22
  (
    n36,
    n1
  );


  buf
  g23
  (
    n39,
    n10
  );


  buf
  g24
  (
    n33,
    n9
  );


  not
  g25
  (
    n147,
    n26
  );


  not
  g26
  (
    n43,
    n2
  );


  not
  g27
  (
    n103,
    n12
  );


  not
  g28
  (
    n68,
    n12
  );


  not
  g29
  (
    n95,
    n5
  );


  buf
  g30
  (
    n35,
    n27
  );


  buf
  g31
  (
    n58,
    n23
  );


  buf
  g32
  (
    n146,
    n3
  );


  buf
  g33
  (
    n123,
    n23
  );


  not
  g34
  (
    n122,
    n28
  );


  not
  g35
  (
    n101,
    n24
  );


  not
  g36
  (
    n49,
    n4
  );


  not
  g37
  (
    n50,
    n16
  );


  not
  g38
  (
    n137,
    n24
  );


  buf
  g39
  (
    n150,
    n8
  );


  not
  g40
  (
    n74,
    n18
  );


  not
  g41
  (
    n96,
    n10
  );


  buf
  g42
  (
    n90,
    n13
  );


  buf
  g43
  (
    n38,
    n19
  );


  not
  g44
  (
    n53,
    n29
  );


  not
  g45
  (
    n144,
    n5
  );


  buf
  g46
  (
    n63,
    n1
  );


  not
  g47
  (
    n62,
    n25
  );


  buf
  g48
  (
    n111,
    n10
  );


  not
  g49
  (
    n117,
    n15
  );


  buf
  g50
  (
    n93,
    n2
  );


  not
  g51
  (
    n42,
    n8
  );


  not
  g52
  (
    n116,
    n11
  );


  not
  g53
  (
    KeyWire_0_9,
    n19
  );


  not
  g54
  (
    n91,
    n25
  );


  not
  g55
  (
    n78,
    n9
  );


  not
  g56
  (
    n141,
    n7
  );


  not
  g57
  (
    n136,
    n22
  );


  not
  g58
  (
    n31,
    n7
  );


  not
  g59
  (
    n106,
    n4
  );


  buf
  g60
  (
    n37,
    n22
  );


  not
  g61
  (
    n55,
    n13
  );


  not
  g62
  (
    n133,
    n3
  );


  not
  g63
  (
    KeyWire_0_8,
    n16
  );


  buf
  g64
  (
    n86,
    n12
  );


  not
  g65
  (
    n75,
    n14
  );


  not
  g66
  (
    n72,
    n2
  );


  not
  g67
  (
    n110,
    n4
  );


  not
  g68
  (
    n40,
    n13
  );


  not
  g69
  (
    n77,
    n17
  );


  not
  g70
  (
    n85,
    n16
  );


  buf
  g71
  (
    n109,
    n30
  );


  buf
  g72
  (
    n47,
    n6
  );


  buf
  g73
  (
    KeyWire_0_60,
    n28
  );


  buf
  g74
  (
    n128,
    n26
  );


  buf
  g75
  (
    n92,
    n24
  );


  buf
  g76
  (
    n81,
    n3
  );


  buf
  g77
  (
    n80,
    n14
  );


  buf
  g78
  (
    n51,
    n4
  );


  not
  g79
  (
    n97,
    n27
  );


  not
  g80
  (
    n71,
    n19
  );


  not
  g81
  (
    n56,
    n8
  );


  not
  g82
  (
    n139,
    n26
  );


  not
  g83
  (
    n41,
    n9
  );


  buf
  g84
  (
    n34,
    n10
  );


  not
  g85
  (
    n32,
    n20
  );


  not
  g86
  (
    n127,
    n7
  );


  buf
  g87
  (
    n89,
    n11
  );


  buf
  g88
  (
    n54,
    n27
  );


  buf
  g89
  (
    KeyWire_0_18,
    n18
  );


  not
  g90
  (
    n143,
    n22
  );


  not
  g91
  (
    n64,
    n21
  );


  buf
  g92
  (
    KeyWire_0_42,
    n5
  );


  not
  g93
  (
    n132,
    n30
  );


  not
  g94
  (
    n131,
    n25
  );


  not
  g95
  (
    n107,
    n23
  );


  not
  g96
  (
    n148,
    n13
  );


  not
  g97
  (
    n57,
    n17
  );


  not
  g98
  (
    n119,
    n3
  );


  not
  g99
  (
    n98,
    n18
  );


  buf
  g100
  (
    KeyWire_0_54,
    n25
  );


  not
  g101
  (
    n130,
    n15
  );


  buf
  g102
  (
    n66,
    n20
  );


  not
  g103
  (
    n73,
    n20
  );


  not
  g104
  (
    n76,
    n17
  );


  not
  g105
  (
    n114,
    n15
  );


  buf
  g106
  (
    n145,
    n17
  );


  not
  g107
  (
    n94,
    n12
  );


  buf
  g108
  (
    n60,
    n30
  );


  buf
  g109
  (
    n124,
    n16
  );


  not
  g110
  (
    n82,
    n19
  );


  buf
  g111
  (
    n140,
    n20
  );


  not
  g112
  (
    n104,
    n21
  );


  not
  g113
  (
    n138,
    n14
  );


  buf
  g114
  (
    KeyWire_0_58,
    n28
  );


  buf
  g115
  (
    n134,
    n15
  );


  not
  g116
  (
    n112,
    n29
  );


  buf
  g117
  (
    n129,
    n6
  );


  buf
  g118
  (
    n102,
    n2
  );


  not
  g119
  (
    n67,
    n24
  );


  not
  g120
  (
    n396,
    n91
  );


  buf
  g121
  (
    n195,
    n45
  );


  buf
  g122
  (
    n244,
    n57
  );


  buf
  g123
  (
    n331,
    n75
  );


  buf
  g124
  (
    n276,
    n136
  );


  not
  g125
  (
    n500,
    n45
  );


  buf
  g126
  (
    n463,
    n87
  );


  buf
  g127
  (
    n362,
    n116
  );


  buf
  g128
  (
    n531,
    n77
  );


  buf
  g129
  (
    n451,
    n113
  );


  buf
  g130
  (
    n273,
    n140
  );


  buf
  g131
  (
    n335,
    n53
  );


  not
  g132
  (
    n548,
    n138
  );


  buf
  g133
  (
    n208,
    n90
  );


  not
  g134
  (
    n570,
    n70
  );


  buf
  g135
  (
    n435,
    n63
  );


  not
  g136
  (
    n374,
    n43
  );


  not
  g137
  (
    n155,
    n87
  );


  buf
  g138
  (
    n163,
    n121
  );


  buf
  g139
  (
    n579,
    n142
  );


  not
  g140
  (
    KeyWire_0_11,
    n102
  );


  not
  g141
  (
    n459,
    n94
  );


  not
  g142
  (
    n348,
    n147
  );


  not
  g143
  (
    n324,
    n31
  );


  not
  g144
  (
    n466,
    n81
  );


  buf
  g145
  (
    n234,
    n95
  );


  not
  g146
  (
    n578,
    n125
  );


  buf
  g147
  (
    n478,
    n44
  );


  not
  g148
  (
    n555,
    n137
  );


  buf
  g149
  (
    n165,
    n136
  );


  buf
  g150
  (
    n593,
    n98
  );


  not
  g151
  (
    n328,
    n48
  );


  buf
  g152
  (
    n426,
    n149
  );


  not
  g153
  (
    n268,
    n31
  );


  not
  g154
  (
    n588,
    n62
  );


  not
  g155
  (
    n461,
    n134
  );


  buf
  g156
  (
    n176,
    n130
  );


  buf
  g157
  (
    n563,
    n79
  );


  not
  g158
  (
    n158,
    n108
  );


  not
  g159
  (
    KeyWire_0_23,
    n89
  );


  buf
  g160
  (
    n402,
    n99
  );


  not
  g161
  (
    n380,
    n129
  );


  not
  g162
  (
    n439,
    n45
  );


  buf
  g163
  (
    n289,
    n112
  );


  buf
  g164
  (
    n377,
    n70
  );


  buf
  g165
  (
    n498,
    n40
  );


  not
  g166
  (
    n455,
    n93
  );


  not
  g167
  (
    n510,
    n33
  );


  buf
  g168
  (
    n428,
    n123
  );


  buf
  g169
  (
    n390,
    n132
  );


  buf
  g170
  (
    n318,
    n45
  );


  buf
  g171
  (
    n198,
    n128
  );


  buf
  g172
  (
    n352,
    n116
  );


  not
  g173
  (
    n201,
    n82
  );


  not
  g174
  (
    n308,
    n57
  );


  not
  g175
  (
    n481,
    n97
  );


  not
  g176
  (
    n577,
    n103
  );


  not
  g177
  (
    n366,
    n35
  );


  buf
  g178
  (
    n256,
    n132
  );


  not
  g179
  (
    n556,
    n105
  );


  not
  g180
  (
    n334,
    n69
  );


  not
  g181
  (
    n355,
    n90
  );


  not
  g182
  (
    n499,
    n148
  );


  not
  g183
  (
    n238,
    n71
  );


  buf
  g184
  (
    KeyWire_0_50,
    n31
  );


  not
  g185
  (
    n544,
    n113
  );


  not
  g186
  (
    n248,
    n111
  );


  not
  g187
  (
    n271,
    n114
  );


  not
  g188
  (
    n370,
    n59
  );


  not
  g189
  (
    n230,
    n123
  );


  buf
  g190
  (
    n381,
    n100
  );


  not
  g191
  (
    n560,
    n146
  );


  buf
  g192
  (
    n539,
    n108
  );


  not
  g193
  (
    n433,
    n44
  );


  not
  g194
  (
    n407,
    n38
  );


  buf
  g195
  (
    n185,
    n96
  );


  not
  g196
  (
    n501,
    n47
  );


  not
  g197
  (
    n462,
    n107
  );


  not
  g198
  (
    n496,
    n127
  );


  not
  g199
  (
    n387,
    n125
  );


  not
  g200
  (
    n251,
    n136
  );


  not
  g201
  (
    KeyWire_0_35,
    n135
  );


  buf
  g202
  (
    n558,
    n107
  );


  buf
  g203
  (
    n359,
    n46
  );


  buf
  g204
  (
    n250,
    n105
  );


  not
  g205
  (
    n412,
    n139
  );


  buf
  g206
  (
    n225,
    n100
  );


  buf
  g207
  (
    n495,
    n96
  );


  not
  g208
  (
    n533,
    n149
  );


  buf
  g209
  (
    n564,
    n55
  );


  not
  g210
  (
    n247,
    n134
  );


  buf
  g211
  (
    n421,
    n69
  );


  buf
  g212
  (
    n333,
    n67
  );


  buf
  g213
  (
    n399,
    n46
  );


  buf
  g214
  (
    n442,
    n55
  );


  not
  g215
  (
    n403,
    n60
  );


  buf
  g216
  (
    n192,
    n103
  );


  not
  g217
  (
    n460,
    n66
  );


  not
  g218
  (
    n206,
    n66
  );


  not
  g219
  (
    KeyWire_0_62,
    n101
  );


  not
  g220
  (
    n162,
    n71
  );


  buf
  g221
  (
    n154,
    n66
  );


  buf
  g222
  (
    n423,
    n96
  );


  buf
  g223
  (
    n221,
    n80
  );


  buf
  g224
  (
    n411,
    n108
  );


  not
  g225
  (
    n446,
    n115
  );


  not
  g226
  (
    n493,
    n39
  );


  buf
  g227
  (
    n180,
    n96
  );


  buf
  g228
  (
    KeyWire_0_61,
    n118
  );


  buf
  g229
  (
    n311,
    n65
  );


  not
  g230
  (
    n263,
    n34
  );


  buf
  g231
  (
    n346,
    n68
  );


  not
  g232
  (
    n282,
    n106
  );


  buf
  g233
  (
    n332,
    n98
  );


  not
  g234
  (
    n571,
    n85
  );


  buf
  g235
  (
    n384,
    n60
  );


  not
  g236
  (
    n281,
    n54
  );


  buf
  g237
  (
    n521,
    n88
  );


  not
  g238
  (
    n508,
    n135
  );


  buf
  g239
  (
    n522,
    n54
  );


  buf
  g240
  (
    n371,
    n65
  );


  buf
  g241
  (
    n364,
    n106
  );


  buf
  g242
  (
    n541,
    n97
  );


  buf
  g243
  (
    n231,
    n138
  );


  not
  g244
  (
    n336,
    n76
  );


  buf
  g245
  (
    n589,
    n89
  );


  buf
  g246
  (
    n404,
    n64
  );


  not
  g247
  (
    n188,
    n115
  );


  buf
  g248
  (
    n279,
    n121
  );


  not
  g249
  (
    KeyWire_0_19,
    n147
  );


  buf
  g250
  (
    n193,
    n144
  );


  buf
  g251
  (
    n400,
    n68
  );


  buf
  g252
  (
    KeyWire_0_38,
    n105
  );


  buf
  g253
  (
    n302,
    n67
  );


  not
  g254
  (
    n235,
    n142
  );


  buf
  g255
  (
    KeyWire_0_59,
    n99
  );


  buf
  g256
  (
    n452,
    n83
  );


  not
  g257
  (
    n479,
    n124
  );


  buf
  g258
  (
    n431,
    n126
  );


  buf
  g259
  (
    n365,
    n62
  );


  not
  g260
  (
    n349,
    n123
  );


  not
  g261
  (
    n434,
    n117
  );


  buf
  g262
  (
    n554,
    n56
  );


  not
  g263
  (
    n291,
    n50
  );


  not
  g264
  (
    n216,
    n114
  );


  not
  g265
  (
    n388,
    n114
  );


  buf
  g266
  (
    n204,
    n130
  );


  not
  g267
  (
    n223,
    n115
  );


  not
  g268
  (
    n534,
    n49
  );


  buf
  g269
  (
    n559,
    n111
  );


  buf
  g270
  (
    n327,
    n42
  );


  not
  g271
  (
    n186,
    n89
  );


  buf
  g272
  (
    n361,
    n94
  );


  buf
  g273
  (
    n547,
    n104
  );


  not
  g274
  (
    n267,
    n98
  );


  buf
  g275
  (
    n591,
    n106
  );


  buf
  g276
  (
    n528,
    n53
  );


  not
  g277
  (
    n317,
    n108
  );


  buf
  g278
  (
    n294,
    n121
  );


  buf
  g279
  (
    n545,
    n78
  );


  not
  g280
  (
    n574,
    n131
  );


  buf
  g281
  (
    n406,
    n92
  );


  not
  g282
  (
    n464,
    n141
  );


  not
  g283
  (
    n546,
    n38
  );


  buf
  g284
  (
    n448,
    n103
  );


  not
  g285
  (
    n450,
    n74
  );


  not
  g286
  (
    n269,
    n63
  );


  not
  g287
  (
    n425,
    n129
  );


  not
  g288
  (
    n303,
    n115
  );


  buf
  g289
  (
    n550,
    n80
  );


  not
  g290
  (
    n520,
    n117
  );


  not
  g291
  (
    n492,
    n148
  );


  buf
  g292
  (
    n167,
    n82
  );


  not
  g293
  (
    n511,
    n91
  );


  buf
  g294
  (
    n487,
    n85
  );


  buf
  g295
  (
    n491,
    n131
  );


  buf
  g296
  (
    n474,
    n71
  );


  not
  g297
  (
    n417,
    n82
  );


  buf
  g298
  (
    n212,
    n48
  );


  not
  g299
  (
    n429,
    n88
  );


  not
  g300
  (
    n242,
    n93
  );


  not
  g301
  (
    n392,
    n104
  );


  buf
  g302
  (
    n304,
    n146
  );


  buf
  g303
  (
    n529,
    n83
  );


  buf
  g304
  (
    n241,
    n95
  );


  not
  g305
  (
    KeyWire_0_39,
    n86
  );


  buf
  g306
  (
    n194,
    n54
  );


  buf
  g307
  (
    n350,
    n71
  );


  buf
  g308
  (
    KeyWire_0_1,
    n33
  );


  buf
  g309
  (
    n486,
    n92
  );


  buf
  g310
  (
    n530,
    n85
  );


  buf
  g311
  (
    n465,
    n36
  );


  not
  g312
  (
    n319,
    n70
  );


  not
  g313
  (
    n477,
    n124
  );


  not
  g314
  (
    n488,
    n90
  );


  buf
  g315
  (
    n284,
    n132
  );


  not
  g316
  (
    n264,
    n59
  );


  buf
  g317
  (
    n383,
    n42
  );


  buf
  g318
  (
    n594,
    n56
  );


  buf
  g319
  (
    n200,
    n64
  );


  buf
  g320
  (
    n257,
    n110
  );


  buf
  g321
  (
    n543,
    n33
  );


  buf
  g322
  (
    n509,
    n117
  );


  buf
  g323
  (
    n287,
    n140
  );


  buf
  g324
  (
    n405,
    n128
  );


  not
  g325
  (
    n181,
    n74
  );


  buf
  g326
  (
    n504,
    n147
  );


  not
  g327
  (
    n443,
    n52
  );


  buf
  g328
  (
    n345,
    n149
  );


  buf
  g329
  (
    n196,
    n68
  );


  buf
  g330
  (
    n280,
    n118
  );


  buf
  g331
  (
    n572,
    n34
  );


  not
  g332
  (
    n270,
    n39
  );


  not
  g333
  (
    n265,
    n35
  );


  buf
  g334
  (
    n398,
    n44
  );


  buf
  g335
  (
    n447,
    n84
  );


  buf
  g336
  (
    n414,
    n102
  );


  buf
  g337
  (
    n581,
    n60
  );


  buf
  g338
  (
    n449,
    n94
  );


  buf
  g339
  (
    n151,
    n143
  );


  not
  g340
  (
    n199,
    n42
  );


  not
  g341
  (
    n557,
    n135
  );


  not
  g342
  (
    n299,
    n97
  );


  buf
  g343
  (
    n240,
    n76
  );


  not
  g344
  (
    n567,
    n138
  );


  buf
  g345
  (
    n306,
    n101
  );


  buf
  g346
  (
    n358,
    n41
  );


  buf
  g347
  (
    n183,
    n75
  );


  not
  g348
  (
    n540,
    n125
  );


  not
  g349
  (
    n475,
    n119
  );


  buf
  g350
  (
    n395,
    n43
  );


  not
  g351
  (
    n369,
    n75
  );


  buf
  g352
  (
    n353,
    n44
  );


  buf
  g353
  (
    n249,
    n49
  );


  buf
  g354
  (
    n322,
    n61
  );


  not
  g355
  (
    n523,
    n99
  );


  not
  g356
  (
    n214,
    n109
  );


  not
  g357
  (
    n340,
    n122
  );


  not
  g358
  (
    n323,
    n82
  );


  not
  g359
  (
    n285,
    n116
  );


  not
  g360
  (
    n297,
    n114
  );


  buf
  g361
  (
    n168,
    n141
  );


  not
  g362
  (
    n532,
    n51
  );


  buf
  g363
  (
    n440,
    n105
  );


  not
  g364
  (
    n413,
    n120
  );


  not
  g365
  (
    n347,
    n38
  );


  buf
  g366
  (
    n290,
    n79
  );


  buf
  g367
  (
    n171,
    n86
  );


  not
  g368
  (
    n561,
    n50
  );


  buf
  g369
  (
    n397,
    n48
  );


  not
  g370
  (
    n469,
    n131
  );


  not
  g371
  (
    n401,
    n109
  );


  not
  g372
  (
    n224,
    n113
  );


  buf
  g373
  (
    n159,
    n101
  );


  not
  g374
  (
    n432,
    n81
  );


  buf
  g375
  (
    n473,
    n79
  );


  buf
  g376
  (
    n471,
    n64
  );


  buf
  g377
  (
    n515,
    n120
  );


  not
  g378
  (
    n228,
    n145
  );


  buf
  g379
  (
    n552,
    n134
  );


  not
  g380
  (
    n503,
    n57
  );


  buf
  g381
  (
    n261,
    n148
  );


  buf
  g382
  (
    n368,
    n119
  );


  buf
  g383
  (
    n226,
    n150
  );


  buf
  g384
  (
    n456,
    n150
  );


  not
  g385
  (
    n191,
    n107
  );


  not
  g386
  (
    n507,
    n113
  );


  not
  g387
  (
    n236,
    n135
  );


  buf
  g388
  (
    n325,
    n41
  );


  not
  g389
  (
    n326,
    n141
  );


  buf
  g390
  (
    n445,
    n37
  );


  buf
  g391
  (
    n438,
    n143
  );


  not
  g392
  (
    n215,
    n62
  );


  not
  g393
  (
    n386,
    n66
  );


  not
  g394
  (
    n293,
    n124
  );


  not
  g395
  (
    n419,
    n133
  );


  buf
  g396
  (
    n255,
    n31
  );


  not
  g397
  (
    n153,
    n126
  );


  not
  g398
  (
    n343,
    n47
  );


  not
  g399
  (
    n375,
    n78
  );


  buf
  g400
  (
    n382,
    n119
  );


  buf
  g401
  (
    n490,
    n100
  );


  not
  g402
  (
    n389,
    n127
  );


  not
  g403
  (
    n275,
    n58
  );


  buf
  g404
  (
    n542,
    n110
  );


  not
  g405
  (
    n483,
    n92
  );


  buf
  g406
  (
    n305,
    n142
  );


  not
  g407
  (
    n569,
    n50
  );


  buf
  g408
  (
    n203,
    n32
  );


  buf
  g409
  (
    n222,
    n131
  );


  not
  g410
  (
    n157,
    n40
  );


  buf
  g411
  (
    n517,
    n134
  );


  not
  g412
  (
    n217,
    n72
  );


  buf
  g413
  (
    n182,
    n92
  );


  not
  g414
  (
    n177,
    n123
  );


  not
  g415
  (
    n516,
    n32
  );


  not
  g416
  (
    n262,
    n84
  );


  not
  g417
  (
    n524,
    n46
  );


  not
  g418
  (
    n526,
    n48
  );


  not
  g419
  (
    n489,
    n121
  );


  buf
  g420
  (
    n277,
    n143
  );


  not
  g421
  (
    n424,
    n122
  );


  buf
  g422
  (
    n367,
    n83
  );


  buf
  g423
  (
    n436,
    n49
  );


  buf
  g424
  (
    n506,
    n59
  );


  buf
  g425
  (
    n295,
    n118
  );


  not
  g426
  (
    n258,
    n112
  );


  buf
  g427
  (
    n394,
    n95
  );


  buf
  g428
  (
    n537,
    n53
  );


  not
  g429
  (
    KeyWire_0_12,
    n58
  );


  not
  g430
  (
    n566,
    n52
  );


  buf
  g431
  (
    n378,
    n56
  );


  buf
  g432
  (
    n274,
    n43
  );


  not
  g433
  (
    n184,
    n61
  );


  buf
  g434
  (
    n341,
    n119
  );


  buf
  g435
  (
    n160,
    n55
  );


  not
  g436
  (
    n468,
    n148
  );


  not
  g437
  (
    n309,
    n127
  );


  not
  g438
  (
    n512,
    n88
  );


  not
  g439
  (
    n170,
    n81
  );


  buf
  g440
  (
    n253,
    n69
  );


  buf
  g441
  (
    KeyWire_0_34,
    n72
  );


  buf
  g442
  (
    n441,
    n34
  );


  buf
  g443
  (
    n197,
    n37
  );


  not
  g444
  (
    n245,
    n107
  );


  buf
  g445
  (
    n283,
    n78
  );


  not
  g446
  (
    n320,
    n38
  );


  buf
  g447
  (
    n373,
    n86
  );


  not
  g448
  (
    n164,
    n40
  );


  buf
  g449
  (
    n219,
    n73
  );


  not
  g450
  (
    n519,
    n93
  );


  not
  g451
  (
    n233,
    n116
  );


  buf
  g452
  (
    n286,
    n94
  );


  not
  g453
  (
    n416,
    n34
  );


  buf
  g454
  (
    n587,
    n126
  );


  buf
  g455
  (
    n298,
    n138
  );


  buf
  g456
  (
    KeyWire_0_36,
    n125
  );


  not
  g457
  (
    n497,
    n128
  );


  buf
  g458
  (
    n209,
    n142
  );


  not
  g459
  (
    n344,
    n56
  );


  buf
  g460
  (
    n453,
    n80
  );


  buf
  g461
  (
    n391,
    n150
  );


  buf
  g462
  (
    n301,
    n83
  );


  not
  g463
  (
    n166,
    n33
  );


  not
  g464
  (
    n538,
    n91
  );


  not
  g465
  (
    KeyWire_0_15,
    n132
  );


  not
  g466
  (
    n376,
    n32
  );


  not
  g467
  (
    n213,
    n39
  );


  buf
  g468
  (
    n568,
    n62
  );


  buf
  g469
  (
    n329,
    n109
  );


  buf
  g470
  (
    n300,
    n58
  );


  buf
  g471
  (
    n457,
    n106
  );


  not
  g472
  (
    n174,
    n102
  );


  not
  g473
  (
    n580,
    n91
  );


  buf
  g474
  (
    n272,
    n137
  );


  not
  g475
  (
    n229,
    n49
  );


  buf
  g476
  (
    n549,
    n84
  );


  buf
  g477
  (
    n339,
    n133
  );


  not
  g478
  (
    n467,
    n50
  );


  not
  g479
  (
    n239,
    n51
  );


  not
  g480
  (
    n357,
    n55
  );


  not
  g481
  (
    n513,
    n77
  );


  not
  g482
  (
    n385,
    n76
  );


  buf
  g483
  (
    n356,
    n137
  );


  buf
  g484
  (
    n260,
    n111
  );


  buf
  g485
  (
    n485,
    n37
  );


  buf
  g486
  (
    n207,
    n36
  );


  buf
  g487
  (
    KeyWire_0_31,
    n120
  );


  not
  g488
  (
    n592,
    n143
  );


  not
  g489
  (
    n484,
    n139
  );


  buf
  g490
  (
    n205,
    n103
  );


  buf
  g491
  (
    n393,
    n64
  );


  not
  g492
  (
    n254,
    n53
  );


  buf
  g493
  (
    n227,
    n87
  );


  buf
  g494
  (
    n292,
    n73
  );


  buf
  g495
  (
    n470,
    n35
  );


  not
  g496
  (
    n175,
    n77
  );


  not
  g497
  (
    n211,
    n149
  );


  not
  g498
  (
    n189,
    n109
  );


  buf
  g499
  (
    n232,
    n145
  );


  buf
  g500
  (
    n278,
    n117
  );


  buf
  g501
  (
    n218,
    n145
  );


  buf
  g502
  (
    n472,
    n144
  );


  not
  g503
  (
    n321,
    n78
  );


  buf
  g504
  (
    n315,
    n100
  );


  not
  g505
  (
    n565,
    n130
  );


  buf
  g506
  (
    n220,
    n137
  );


  buf
  g507
  (
    n476,
    n70
  );


  not
  g508
  (
    n152,
    n51
  );


  not
  g509
  (
    n179,
    n140
  );


  not
  g510
  (
    n422,
    n99
  );


  buf
  g511
  (
    n502,
    n79
  );


  buf
  g512
  (
    n527,
    n144
  );


  not
  g513
  (
    n161,
    n90
  );


  not
  g514
  (
    n296,
    n145
  );


  not
  g515
  (
    n307,
    n147
  );


  buf
  g516
  (
    n237,
    n47
  );


  not
  g517
  (
    n202,
    n95
  );


  not
  g518
  (
    n525,
    n39
  );


  not
  g519
  (
    n430,
    n61
  );


  buf
  g520
  (
    n259,
    n72
  );


  buf
  g521
  (
    n156,
    n36
  );


  buf
  g522
  (
    n575,
    n73
  );


  not
  g523
  (
    n437,
    n72
  );


  buf
  g524
  (
    n190,
    n101
  );


  buf
  g525
  (
    n427,
    n139
  );


  not
  g526
  (
    n583,
    n136
  );


  buf
  g527
  (
    KeyWire_0_51,
    n88
  );


  not
  g528
  (
    n553,
    n122
  );


  buf
  g529
  (
    n409,
    n146
  );


  buf
  g530
  (
    n480,
    n46
  );


  buf
  g531
  (
    n351,
    n122
  );


  buf
  g532
  (
    n562,
    n41
  );


  not
  g533
  (
    n420,
    n37
  );


  buf
  g534
  (
    n514,
    n73
  );


  buf
  g535
  (
    n354,
    n63
  );


  buf
  g536
  (
    n372,
    n40
  );


  buf
  g537
  (
    KeyWire_0_21,
    n102
  );


  buf
  g538
  (
    n573,
    n127
  );


  buf
  g539
  (
    n535,
    n120
  );


  not
  g540
  (
    n178,
    n43
  );


  buf
  g541
  (
    n494,
    n54
  );


  buf
  g542
  (
    n586,
    n104
  );


  buf
  g543
  (
    n172,
    n141
  );


  buf
  g544
  (
    n252,
    n93
  );


  not
  g545
  (
    n458,
    n74
  );


  not
  g546
  (
    n444,
    n68
  );


  buf
  g547
  (
    n454,
    n80
  );


  nor
  g548
  (
    n288,
    n126,
    n118,
    n52
  );


  or
  g549
  (
    n310,
    n133,
    n76,
    n112
  );


  xnor
  g550
  (
    KeyWire_0_47,
    n74,
    n52,
    n124
  );


  or
  g551
  (
    n518,
    n139,
    n130,
    n69
  );


  and
  g552
  (
    n360,
    n61,
    n65,
    n77
  );


  nor
  g553
  (
    n313,
    n144,
    n42,
    n110
  );


  xnor
  g554
  (
    n379,
    n81,
    n41,
    n75
  );


  or
  g555
  (
    n312,
    n129,
    n65,
    n140
  );


  or
  g556
  (
    n210,
    n36,
    n63,
    n89
  );


  nor
  g557
  (
    n582,
    n133,
    n111,
    n84
  );


  and
  g558
  (
    n576,
    n51,
    n87,
    n129
  );


  nor
  g559
  (
    n187,
    n67,
    n98,
    n85
  );


  or
  g560
  (
    n551,
    n35,
    n60,
    n97
  );


  and
  g561
  (
    n173,
    n58,
    n104,
    n32
  );


  xnor
  g562
  (
    n595,
    n59,
    n86,
    n110
  );


  xor
  g563
  (
    n585,
    n57,
    n146,
    n47
  );


  nand
  g564
  (
    n342,
    n112,
    n67,
    n128
  );


  or
  g565
  (
    n686,
    n252,
    n460
  );


  xnor
  g566
  (
    n639,
    n244,
    n516
  );


  xnor
  g567
  (
    n683,
    n275,
    n334
  );


  xor
  g568
  (
    n680,
    n206,
    n423
  );


  xor
  g569
  (
    n641,
    n344,
    n170,
    n407,
    n479
  );


  nor
  g570
  (
    n608,
    n475,
    n514,
    n516,
    n506
  );


  and
  g571
  (
    n609,
    n298,
    n436,
    n513,
    n372
  );


  or
  g572
  (
    n668,
    n483,
    n283,
    n326,
    n409
  );


  xnor
  g573
  (
    n694,
    n383,
    n245,
    n166,
    n373
  );


  xor
  g574
  (
    n688,
    n513,
    n207,
    n359,
    n367
  );


  nand
  g575
  (
    n670,
    n255,
    n476,
    n178,
    n189
  );


  xor
  g576
  (
    n648,
    n439,
    n312,
    n485,
    n159
  );


  nor
  g577
  (
    n674,
    n256,
    n214,
    n402,
    n273
  );


  nor
  g578
  (
    n602,
    n309,
    n265,
    n495,
    n432
  );


  nand
  g579
  (
    n692,
    n461,
    n263,
    n472,
    n175
  );


  nor
  g580
  (
    n678,
    n321,
    n360,
    n365,
    n464
  );


  or
  g581
  (
    n657,
    n468,
    n492,
    n240,
    n156
  );


  xor
  g582
  (
    n606,
    n433,
    n497,
    n427,
    n151
  );


  nand
  g583
  (
    n682,
    n164,
    n318,
    n430,
    n517
  );


  nand
  g584
  (
    n669,
    n336,
    n271,
    n512,
    n504
  );


  nor
  g585
  (
    n619,
    n354,
    n316,
    n229,
    n233
  );


  nor
  g586
  (
    n666,
    n442,
    n418,
    n301,
    n313
  );


  and
  g587
  (
    n650,
    n511,
    n474,
    n153,
    n364
  );


  or
  g588
  (
    n656,
    n201,
    n486,
    n500,
    n203
  );


  or
  g589
  (
    n638,
    n390,
    n329,
    n225,
    n362
  );


  or
  g590
  (
    n695,
    n174,
    n266,
    n465,
    n481
  );


  xor
  g591
  (
    n614,
    n305,
    n351,
    n406,
    n243
  );


  and
  g592
  (
    n689,
    n394,
    n511,
    n399,
    n458
  );


  and
  g593
  (
    n655,
    n215,
    n302,
    n403,
    n180
  );


  nor
  g594
  (
    n631,
    n400,
    n519,
    n469,
    n210
  );


  xnor
  g595
  (
    n625,
    n332,
    n199,
    n342,
    n269
  );


  xor
  g596
  (
    n637,
    n186,
    n404,
    n197,
    n218
  );


  nor
  g597
  (
    n649,
    n381,
    n514,
    n454,
    n513
  );


  xor
  g598
  (
    n662,
    n398,
    n235,
    n155,
    n177
  );


  or
  g599
  (
    n618,
    n347,
    n484,
    n194,
    n236
  );


  nor
  g600
  (
    KeyWire_0_33,
    n438,
    n322,
    n279,
    n437
  );


  or
  g601
  (
    n634,
    n384,
    n196,
    n370,
    n154
  );


  nand
  g602
  (
    n617,
    n284,
    n282,
    n323,
    n232
  );


  and
  g603
  (
    n643,
    n386,
    n357,
    n290,
    n341
  );


  nor
  g604
  (
    n633,
    n519,
    n493,
    n325,
    n517
  );


  xor
  g605
  (
    n604,
    n511,
    n505,
    n172,
    n519
  );


  xnor
  g606
  (
    KeyWire_0_4,
    n258,
    n230,
    n509,
    n328
  );


  xnor
  g607
  (
    n663,
    n397,
    n227,
    n408,
    n338
  );


  nor
  g608
  (
    n598,
    n482,
    n508,
    n366,
    n499
  );


  or
  g609
  (
    n658,
    n160,
    n356,
    n324,
    n451
  );


  nor
  g610
  (
    n660,
    n158,
    n231,
    n424,
    n228
  );


  xor
  g611
  (
    n635,
    n202,
    n515,
    n507,
    n462
  );


  xor
  g612
  (
    n615,
    n339,
    n268,
    n152,
    n488
  );


  xor
  g613
  (
    n675,
    n264,
    n463,
    n453,
    n498
  );


  xor
  g614
  (
    n623,
    n456,
    n369,
    n452,
    n379
  );


  and
  g615
  (
    KeyWire_0_44,
    n297,
    n183,
    n165,
    n181
  );


  or
  g616
  (
    n672,
    n415,
    n270,
    n518,
    n314
  );


  nand
  g617
  (
    KeyWire_0_16,
    n272,
    n376,
    n512,
    n393
  );


  xnor
  g618
  (
    n626,
    n250,
    n274,
    n185,
    n299
  );


  nor
  g619
  (
    n630,
    n368,
    n502,
    n184,
    n517
  );


  nor
  g620
  (
    n628,
    n510,
    n459,
    n306,
    n191
  );


  and
  g621
  (
    n621,
    n392,
    n285,
    n278,
    n288
  );


  or
  g622
  (
    KeyWire_0_22,
    n176,
    n286,
    n434,
    n251
  );


  nor
  g623
  (
    n636,
    n287,
    n308,
    n320,
    n350
  );


  or
  g624
  (
    n616,
    n173,
    n470,
    n234,
    n337
  );


  nand
  g625
  (
    n597,
    n190,
    n204,
    n371,
    n248
  );


  nand
  g626
  (
    n681,
    n448,
    n277,
    n307,
    n496
  );


  or
  g627
  (
    n661,
    n444,
    n200,
    n167,
    n241
  );


  nor
  g628
  (
    n679,
    n249,
    n217,
    n348,
    n445
  );


  nand
  g629
  (
    n690,
    n161,
    n391,
    n510,
    n513
  );


  or
  g630
  (
    n624,
    n515,
    n171,
    n471,
    n220
  );


  xor
  g631
  (
    n691,
    n396,
    n515,
    n226,
    n519
  );


  and
  g632
  (
    KeyWire_0_32,
    n431,
    n327,
    n192,
    n440
  );


  and
  g633
  (
    n665,
    n512,
    n512,
    n361,
    n411
  );


  and
  g634
  (
    n645,
    n417,
    n216,
    n262,
    n426
  );


  nor
  g635
  (
    n620,
    n317,
    n450,
    n428,
    n447
  );


  or
  g636
  (
    n644,
    n375,
    n501,
    n518,
    n343
  );


  xor
  g637
  (
    n632,
    n385,
    n224,
    n242,
    n246
  );


  or
  g638
  (
    n651,
    n510,
    n413,
    n416,
    n518
  );


  or
  g639
  (
    n629,
    n310,
    n296,
    n198,
    n412
  );


  and
  g640
  (
    n693,
    n466,
    n304,
    n380,
    n374
  );


  nand
  g641
  (
    n654,
    n331,
    n422,
    n188,
    n377
  );


  or
  g642
  (
    n646,
    n494,
    n414,
    n520,
    n213
  );


  xnor
  g643
  (
    n687,
    n435,
    n388,
    n345,
    n300
  );


  nor
  g644
  (
    n685,
    n378,
    n169,
    n446,
    n294
  );


  xor
  g645
  (
    n696,
    n489,
    n247,
    n187,
    n335
  );


  xor
  g646
  (
    n610,
    n349,
    n293,
    n352,
    n315
  );


  and
  g647
  (
    n601,
    n455,
    n449,
    n222,
    n267
  );


  and
  g648
  (
    n653,
    n179,
    n358,
    n295,
    n443
  );


  xnor
  g649
  (
    n659,
    n212,
    n363,
    n219,
    n223
  );


  nand
  g650
  (
    KeyWire_0_46,
    n515,
    n387,
    n163,
    n395
  );


  nand
  g651
  (
    n622,
    n261,
    n517,
    n289,
    n340
  );


  or
  g652
  (
    n599,
    n157,
    n291,
    n410,
    n311
  );


  or
  g653
  (
    n652,
    n511,
    n195,
    n516,
    n209
  );


  or
  g654
  (
    n697,
    n421,
    n382,
    n389,
    n205
  );


  nand
  g655
  (
    n611,
    n473,
    n238,
    n514,
    n333
  );


  or
  g656
  (
    n664,
    n257,
    n346,
    n303,
    n276
  );


  nand
  g657
  (
    n607,
    n237,
    n260,
    n477,
    n193
  );


  nand
  g658
  (
    n671,
    n292,
    n330,
    n253,
    n239
  );


  nand
  g659
  (
    n642,
    n280,
    n429,
    n254,
    n510
  );


  and
  g660
  (
    n612,
    n353,
    n425,
    n491,
    n162
  );


  nor
  g661
  (
    n596,
    n208,
    n281,
    n211,
    n405
  );


  nor
  g662
  (
    n673,
    n516,
    n514,
    n420,
    n401
  );


  or
  g663
  (
    n667,
    n441,
    n490,
    n518,
    n478
  );


  xor
  g664
  (
    n603,
    n487,
    n419,
    n259,
    n480
  );


  nor
  g665
  (
    n647,
    n182,
    n319,
    n503,
    n457
  );


  xor
  g666
  (
    n684,
    n168,
    n355,
    n467,
    n221
  );


  buf
  g667
  (
    n727,
    n656
  );


  not
  g668
  (
    n724,
    n621
  );


  buf
  g669
  (
    n709,
    n596
  );


  buf
  g670
  (
    n721,
    n620
  );


  not
  g671
  (
    n703,
    n605
  );


  not
  g672
  (
    n700,
    n609
  );


  buf
  g673
  (
    n723,
    n639
  );


  not
  g674
  (
    n705,
    n648
  );


  not
  g675
  (
    n707,
    n622
  );


  buf
  g676
  (
    n711,
    n599
  );


  not
  g677
  (
    n728,
    n657
  );


  not
  g678
  (
    n726,
    n611
  );


  buf
  g679
  (
    n720,
    n649
  );


  not
  g680
  (
    n699,
    n600
  );


  buf
  g681
  (
    n708,
    n627
  );


  not
  g682
  (
    n698,
    n636
  );


  not
  g683
  (
    n713,
    n608
  );


  not
  g684
  (
    n704,
    n598
  );


  not
  g685
  (
    n718,
    n618
  );


  not
  g686
  (
    n710,
    n604
  );


  buf
  g687
  (
    n719,
    n633
  );


  or
  g688
  (
    n712,
    n642,
    n641,
    n652
  );


  and
  g689
  (
    n717,
    n655,
    n631,
    n606,
    n597
  );


  xor
  g690
  (
    n716,
    n607,
    n614,
    n628,
    n635
  );


  xnor
  g691
  (
    n725,
    n616,
    n640,
    n615,
    n651
  );


  or
  g692
  (
    n729,
    n630,
    n625,
    n645,
    n629
  );


  xor
  g693
  (
    n701,
    n602,
    n646,
    n656,
    n603
  );


  nand
  g694
  (
    n706,
    n647,
    n613,
    n632,
    n610
  );


  or
  g695
  (
    n715,
    n617,
    n634,
    n654,
    n626
  );


  and
  g696
  (
    n702,
    n612,
    n637,
    n643,
    n624
  );


  xnor
  g697
  (
    n714,
    n601,
    n656,
    n650,
    n623
  );


  nor
  g698
  (
    n722,
    n619,
    n644,
    n638,
    n653
  );


  buf
  g699
  (
    n730,
    n699
  );


  not
  g700
  (
    n735,
    n698
  );


  not
  g701
  (
    n732,
    n698
  );


  not
  g702
  (
    n736,
    n700
  );


  buf
  g703
  (
    n737,
    n698
  );


  and
  g704
  (
    n738,
    n699,
    n701,
    n702
  );


  xnor
  g705
  (
    n739,
    n699,
    n700
  );


  or
  g706
  (
    n733,
    n702,
    n701,
    n700
  );


  xnor
  g707
  (
    n731,
    n701,
    n702
  );


  and
  g708
  (
    n734,
    n698,
    n701,
    n699
  );


  buf
  g709
  (
    n745,
    n737
  );


  not
  g710
  (
    n742,
    n735
  );


  nand
  g711
  (
    n740,
    n704,
    n733,
    n703,
    n730
  );


  nand
  g712
  (
    n746,
    n704,
    n703,
    n705
  );


  and
  g713
  (
    n743,
    n739,
    n731,
    n705
  );


  xor
  g714
  (
    n741,
    n704,
    n738,
    n703
  );


  nor
  g715
  (
    n744,
    n736,
    n704,
    n732,
    n734
  );


  buf
  g716
  (
    n747,
    n520
  );


  and
  g717
  (
    n750,
    n522,
    n706,
    n746
  );


  or
  g718
  (
    n752,
    n746,
    n520,
    n741
  );


  and
  g719
  (
    n749,
    n742,
    n743,
    n521,
    n740
  );


  or
  g720
  (
    n748,
    n746,
    n744,
    n521
  );


  or
  g721
  (
    n751,
    n745,
    n521,
    n746,
    n706
  );


  buf
  g722
  (
    n759,
    n751
  );


  not
  g723
  (
    n768,
    n711
  );


  buf
  g724
  (
    n758,
    n713
  );


  buf
  g725
  (
    n755,
    n711
  );


  buf
  g726
  (
    n776,
    n748
  );


  buf
  g727
  (
    n757,
    n712
  );


  buf
  g728
  (
    n773,
    n706
  );


  not
  g729
  (
    n774,
    n750
  );


  buf
  g730
  (
    n756,
    n749
  );


  buf
  g731
  (
    n764,
    n706
  );


  buf
  g732
  (
    n766,
    n712
  );


  not
  g733
  (
    n754,
    n711
  );


  or
  g734
  (
    n760,
    n709,
    n749
  );


  nor
  g735
  (
    n767,
    n752,
    n749,
    n751,
    n709
  );


  nor
  g736
  (
    n761,
    n713,
    n714,
    n711,
    n749
  );


  xor
  g737
  (
    n769,
    n750,
    n707,
    n748,
    n713
  );


  xnor
  g738
  (
    n765,
    n707,
    n707,
    n709,
    n748
  );


  and
  g739
  (
    n772,
    n710,
    n710,
    n708,
    n752
  );


  and
  g740
  (
    n775,
    n748,
    n710,
    n747,
    n714
  );


  nand
  g741
  (
    n763,
    n750,
    n713,
    n751,
    n714
  );


  xnor
  g742
  (
    n753,
    n708,
    n712,
    n709
  );


  xnor
  g743
  (
    n770,
    n708,
    n747,
    n710
  );


  xor
  g744
  (
    n771,
    n708,
    n751,
    n747,
    n752
  );


  or
  g745
  (
    n762,
    n707,
    n714,
    n750,
    n752
  );


  buf
  g746
  (
    n781,
    n753
  );


  not
  g747
  (
    n782,
    n753
  );


  buf
  g748
  (
    n784,
    n758
  );


  not
  g749
  (
    n790,
    n757
  );


  not
  g750
  (
    n785,
    n756
  );


  not
  g751
  (
    n789,
    n758
  );


  buf
  g752
  (
    n792,
    n758
  );


  not
  g753
  (
    n778,
    n754
  );


  not
  g754
  (
    n791,
    n755
  );


  and
  g755
  (
    n783,
    n757,
    n754
  );


  xnor
  g756
  (
    n780,
    n757,
    n756
  );


  and
  g757
  (
    n788,
    n756,
    n753
  );


  or
  g758
  (
    n787,
    n757,
    n754
  );


  nor
  g759
  (
    n779,
    n756,
    n754
  );


  xnor
  g760
  (
    n777,
    n755,
    n753
  );


  nand
  g761
  (
    n786,
    n755,
    n758
  );


  xnor
  g762
  (
    n799,
    n792,
    n530,
    n791,
    n531
  );


  xnor
  g763
  (
    n811,
    n790,
    n778,
    n531,
    n716
  );


  nand
  g764
  (
    n794,
    n525,
    n715,
    n528
  );


  nor
  g765
  (
    n801,
    n790,
    n532,
    n784
  );


  nand
  g766
  (
    n802,
    n525,
    n779,
    n781,
    n523
  );


  xor
  g767
  (
    n818,
    n530,
    n788,
    n533,
    n789
  );


  or
  g768
  (
    n812,
    n525,
    n531,
    n791,
    n789
  );


  xor
  g769
  (
    n815,
    n792,
    n523,
    n718
  );


  xor
  g770
  (
    n796,
    n533,
    n718,
    n789,
    n522
  );


  and
  g771
  (
    n816,
    n524,
    n527,
    n715,
    n525
  );


  and
  g772
  (
    n797,
    n777,
    n717,
    n535,
    n533
  );


  xnor
  g773
  (
    n800,
    n789,
    n782,
    n792,
    n716
  );


  nor
  g774
  (
    n798,
    n786,
    n718,
    n717,
    n535
  );


  or
  g775
  (
    n808,
    n785,
    n528,
    n780,
    n790
  );


  xnor
  g776
  (
    n807,
    n527,
    n657,
    n787,
    n715
  );


  or
  g777
  (
    n805,
    n523,
    n522,
    n528,
    n716
  );


  nor
  g778
  (
    n793,
    n527,
    n527,
    n526,
    n534
  );


  and
  g779
  (
    n817,
    n529,
    n526,
    n532,
    n534
  );


  xor
  g780
  (
    n795,
    n657,
    n534,
    n530
  );


  nor
  g781
  (
    n813,
    n535,
    n535,
    n791,
    n526
  );


  xnor
  g782
  (
    n814,
    n524,
    n532,
    n792,
    n536
  );


  xnor
  g783
  (
    n803,
    n717,
    n718,
    n791,
    n790
  );


  xnor
  g784
  (
    KeyWire_0_48,
    n526,
    n529,
    n522,
    n717
  );


  nor
  g785
  (
    n809,
    n783,
    n531,
    n533,
    n529
  );


  xnor
  g786
  (
    n810,
    n524,
    n716,
    n536,
    n530
  );


  nor
  g787
  (
    n806,
    n715,
    n524,
    n536,
    n529
  );


  not
  g788
  (
    n826,
    n793
  );


  buf
  g789
  (
    n828,
    n798
  );


  not
  g790
  (
    n819,
    n793
  );


  buf
  g791
  (
    n822,
    n797
  );


  buf
  g792
  (
    n827,
    n797
  );


  not
  g793
  (
    n821,
    n795
  );


  buf
  g794
  (
    n829,
    n796
  );


  xnor
  g795
  (
    n820,
    n795,
    n793
  );


  and
  g796
  (
    n824,
    n795,
    n798,
    n794,
    n797
  );


  xor
  g797
  (
    n823,
    n797,
    n795,
    n794,
    n793
  );


  xor
  g798
  (
    n825,
    n796,
    n794
  );


  buf
  g799
  (
    n836,
    n822
  );


  not
  g800
  (
    n831,
    n719
  );


  not
  g801
  (
    n834,
    n826
  );


  buf
  g802
  (
    n833,
    n820
  );


  or
  g803
  (
    n835,
    n819,
    n825
  );


  xor
  g804
  (
    n832,
    n829,
    n719,
    n823,
    n828
  );


  xnor
  g805
  (
    n830,
    n827,
    n824,
    n821,
    n719
  );


  nand
  g806
  (
    n839,
    n831,
    n762,
    n833,
    n832
  );


  xor
  g807
  (
    n858,
    n761,
    n719,
    n764,
    n720
  );


  nor
  g808
  (
    n843,
    n832,
    n767,
    n764,
    n769
  );


  and
  g809
  (
    n842,
    n834,
    n772,
    n771,
    n773
  );


  xnor
  g810
  (
    KeyWire_0_41,
    n721,
    n771,
    n772
  );


  nand
  g811
  (
    n863,
    n759,
    n766,
    n769
  );


  and
  g812
  (
    n840,
    n833,
    n830,
    n722,
    n768
  );


  and
  g813
  (
    n853,
    n832,
    n759,
    n836,
    n831
  );


  nand
  g814
  (
    n848,
    n761,
    n720,
    n759,
    n767
  );


  nand
  g815
  (
    n856,
    n767,
    n836,
    n835,
    n720
  );


  nand
  g816
  (
    n857,
    n723,
    n763,
    n724,
    n760
  );


  xnor
  g817
  (
    n849,
    n830,
    n764,
    n767,
    n723
  );


  and
  g818
  (
    n862,
    n836,
    n773,
    n721,
    n765
  );


  and
  g819
  (
    n852,
    n761,
    n763,
    n770,
    n723
  );


  xnor
  g820
  (
    n860,
    n836,
    n761,
    n835,
    n833
  );


  and
  g821
  (
    n837,
    n834,
    n771,
    n765,
    n770
  );


  and
  g822
  (
    n841,
    n835,
    n768,
    n764
  );


  and
  g823
  (
    n861,
    n835,
    n724,
    n831,
    n721
  );


  or
  g824
  (
    n855,
    n832,
    n766,
    n763,
    n760
  );


  xnor
  g825
  (
    n854,
    n760,
    n833,
    n721,
    n834
  );


  xnor
  g826
  (
    n847,
    n773,
    n765,
    n724,
    n766
  );


  and
  g827
  (
    n844,
    n722,
    n762,
    n770
  );


  or
  g828
  (
    n845,
    n720,
    n770,
    n763,
    n769
  );


  nand
  g829
  (
    n851,
    n769,
    n723,
    n762,
    n834
  );


  nand
  g830
  (
    KeyWire_0_37,
    n771,
    n831,
    n536,
    n773
  );


  nand
  g831
  (
    n838,
    n722,
    n768,
    n772,
    n760
  );


  or
  g832
  (
    n846,
    n759,
    n765,
    n830,
    n722
  );


  buf
  g833
  (
    KeyWire_0_5,
    n853
  );


  not
  g834
  (
    n904,
    n809
  );


  buf
  g835
  (
    n899,
    n659
  );


  buf
  g836
  (
    n912,
    n846
  );


  buf
  g837
  (
    n914,
    n857
  );


  not
  g838
  (
    n910,
    n800
  );


  not
  g839
  (
    n890,
    n805
  );


  not
  g840
  (
    n877,
    n861
  );


  not
  g841
  (
    n889,
    n863
  );


  not
  g842
  (
    n892,
    n726
  );


  buf
  g843
  (
    n868,
    n848
  );


  not
  g844
  (
    n883,
    n658
  );


  not
  g845
  (
    n881,
    n802
  );


  not
  g846
  (
    n876,
    n851
  );


  and
  g847
  (
    n882,
    n810,
    n861,
    n849,
    n726
  );


  or
  g848
  (
    n896,
    n852,
    n855,
    n807
  );


  xor
  g849
  (
    n865,
    n809,
    n809,
    n813,
    n806
  );


  nor
  g850
  (
    n873,
    n725,
    n725,
    n858,
    n847
  );


  or
  g851
  (
    n902,
    n854,
    n803,
    n537,
    n847
  );


  nor
  g852
  (
    KeyWire_0_56,
    n799,
    n801,
    n811,
    n857
  );


  nor
  g853
  (
    n898,
    n841,
    n804,
    n855,
    n847
  );


  and
  g854
  (
    n887,
    n803,
    n852,
    n842,
    n854
  );


  xnor
  g855
  (
    n888,
    n802,
    n854,
    n853,
    n858
  );


  and
  g856
  (
    n908,
    n812,
    n856,
    n843,
    n657
  );


  xor
  g857
  (
    n900,
    n806,
    n855,
    n808,
    n860
  );


  nor
  g858
  (
    n894,
    n846,
    n852,
    n860,
    n844
  );


  nor
  g859
  (
    n878,
    n859,
    n726,
    n806,
    n724
  );


  and
  g860
  (
    n907,
    n725,
    n659
  );


  or
  g861
  (
    n874,
    n537,
    n862,
    n850,
    n807
  );


  xnor
  g862
  (
    n906,
    n808,
    n850,
    n838,
    n849
  );


  nand
  g863
  (
    n879,
    n798,
    n851,
    n804,
    n856
  );


  xor
  g864
  (
    n897,
    n862,
    n801,
    n658,
    n800
  );


  nor
  g865
  (
    KeyWire_0_52,
    n800,
    n863,
    n860,
    n850
  );


  and
  g866
  (
    n895,
    n858,
    n862,
    n854,
    n801
  );


  or
  g867
  (
    n880,
    n803,
    n849,
    n805,
    n808
  );


  or
  g868
  (
    n867,
    n857,
    n850,
    n859,
    n811
  );


  or
  g869
  (
    n911,
    n860,
    n658,
    n812,
    n853
  );


  xor
  g870
  (
    n875,
    n805,
    n810,
    n804,
    n839
  );


  xnor
  g871
  (
    n901,
    n847,
    n837,
    n660,
    n799
  );


  xnor
  g872
  (
    n913,
    n848,
    n808,
    n856,
    n846
  );


  xor
  g873
  (
    n893,
    n802,
    n859,
    n658,
    n805
  );


  or
  g874
  (
    n866,
    n799,
    n812,
    n811,
    n807
  );


  and
  g875
  (
    n872,
    n802,
    n810,
    n538,
    n859
  );


  xnor
  g876
  (
    n903,
    n811,
    n848,
    n803,
    n861
  );


  nand
  g877
  (
    n869,
    n852,
    n863,
    n798,
    n537
  );


  or
  g878
  (
    n885,
    n856,
    n858,
    n804,
    n809
  );


  nand
  g879
  (
    n891,
    n810,
    n800,
    n845,
    n863
  );


  and
  g880
  (
    n864,
    n801,
    n659,
    n807,
    n861
  );


  nand
  g881
  (
    n905,
    n851,
    n812,
    n848,
    n806
  );


  xnor
  g882
  (
    n886,
    n849,
    n853,
    n857,
    n862
  );


  or
  g883
  (
    n909,
    n840,
    n851,
    n537,
    n799
  );


  or
  g884
  (
    n922,
    n882,
    n899,
    n906,
    n874
  );


  xnor
  g885
  (
    n927,
    n902,
    n909,
    n906,
    n867
  );


  and
  g886
  (
    n918,
    n894,
    n898,
    n875,
    n893
  );


  nor
  g887
  (
    n915,
    n880,
    n904,
    n866
  );


  nand
  g888
  (
    n920,
    n908,
    n870,
    n904,
    n865
  );


  and
  g889
  (
    n923,
    n903,
    n869,
    n873,
    n881
  );


  xnor
  g890
  (
    n928,
    n877,
    n907,
    n906
  );


  xor
  g891
  (
    n917,
    n908,
    n906,
    n905,
    n868
  );


  and
  g892
  (
    n925,
    n888,
    n907,
    n883,
    n879
  );


  and
  g893
  (
    n921,
    n909,
    n878,
    n887,
    n876
  );


  and
  g894
  (
    n929,
    n889,
    n891,
    n872,
    n885
  );


  nand
  g895
  (
    n916,
    n908,
    n905,
    n904
  );


  nor
  g896
  (
    n924,
    n905,
    n900,
    n897,
    n892
  );


  nand
  g897
  (
    n930,
    n907,
    n886,
    n864,
    n884
  );


  and
  g898
  (
    KeyWire_0_13,
    n871,
    n895,
    n909,
    n896
  );


  and
  g899
  (
    n919,
    n890,
    n909,
    n901,
    n908
  );


  not
  g900
  (
    n934,
    n919
  );


  not
  g901
  (
    n931,
    n921
  );


  buf
  g902
  (
    n935,
    n920
  );


  not
  g903
  (
    n937,
    n915
  );


  buf
  g904
  (
    n933,
    n923
  );


  not
  g905
  (
    n932,
    n923
  );


  buf
  g906
  (
    n936,
    n922
  );


  and
  g907
  (
    n938,
    n918,
    n916,
    n917
  );


  xor
  g908
  (
    n939,
    n935,
    n937,
    n936,
    n814
  );


  nor
  g909
  (
    n944,
    n933,
    n931,
    n936,
    n938
  );


  xnor
  g910
  (
    n950,
    n936,
    n937,
    n910
  );


  nor
  g911
  (
    n946,
    n910,
    n934,
    n935
  );


  and
  g912
  (
    n948,
    n936,
    n933,
    n938
  );


  or
  g913
  (
    n942,
    n813,
    n813,
    n934,
    n935
  );


  or
  g914
  (
    n940,
    n815,
    n911
  );


  or
  g915
  (
    KeyWire_0_24,
    n938,
    n814,
    n934
  );


  or
  g916
  (
    n947,
    n938,
    n813,
    n910,
    n932
  );


  nor
  g917
  (
    n945,
    n815,
    n932,
    n911
  );


  xor
  g918
  (
    n949,
    n814,
    n937,
    n931
  );


  and
  g919
  (
    n941,
    n933,
    n935,
    n932,
    n910
  );


  or
  g920
  (
    n951,
    n924,
    n950,
    n923
  );


  not
  g921
  (
    n954,
    n951
  );


  not
  g922
  (
    n952,
    n951
  );


  buf
  g923
  (
    n953,
    n951
  );


  buf
  g924
  (
    n955,
    n951
  );


  buf
  g925
  (
    n956,
    n952
  );


  buf
  g926
  (
    n958,
    n956
  );


  not
  g927
  (
    n957,
    n956
  );


  xor
  g928
  (
    n959,
    n924,
    n958
  );


  or
  g929
  (
    n962,
    n925,
    n924
  );


  and
  g930
  (
    n960,
    n927,
    n926,
    n959
  );


  or
  g931
  (
    n961,
    n926,
    n959,
    n925
  );


  xor
  g932
  (
    n963,
    n959,
    n926,
    n927,
    n925
  );


  or
  g933
  (
    n967,
    n548,
    n541,
    n962,
    n960
  );


  or
  g934
  (
    n964,
    n544,
    n547,
    n538
  );


  nand
  g935
  (
    n969,
    n543,
    n726,
    n542,
    n544
  );


  and
  g936
  (
    n974,
    n546,
    n962,
    n541,
    n542
  );


  xor
  g937
  (
    n971,
    n541,
    n545,
    n961
  );


  xnor
  g938
  (
    n968,
    n547,
    n544,
    n540,
    n963
  );


  xnor
  g939
  (
    n973,
    n960,
    n545,
    n962,
    n549
  );


  or
  g940
  (
    n977,
    n548,
    n545,
    n540,
    n547
  );


  and
  g941
  (
    n970,
    n542,
    n548,
    n961,
    n541
  );


  xnor
  g942
  (
    n965,
    n540,
    n539,
    n543,
    n538
  );


  nor
  g943
  (
    n975,
    n546,
    n548,
    n539
  );


  xor
  g944
  (
    n978,
    n543,
    n961,
    n546,
    n539
  );


  xnor
  g945
  (
    n972,
    n549,
    n727,
    n543,
    n960
  );


  xnor
  g946
  (
    n966,
    n727,
    n540,
    n544,
    n963
  );


  xnor
  g947
  (
    n976,
    n546,
    n963,
    n545,
    n547
  );


  nor
  g948
  (
    n979,
    n962,
    n542,
    n960,
    n963
  );


  buf
  g949
  (
    n998,
    n964
  );


  buf
  g950
  (
    KeyWire_0_55,
    n968
  );


  buf
  g951
  (
    n996,
    n967
  );


  buf
  g952
  (
    n995,
    n965
  );


  not
  g953
  (
    n993,
    n968
  );


  not
  g954
  (
    n992,
    n967
  );


  buf
  g955
  (
    n983,
    n968
  );


  buf
  g956
  (
    n988,
    n965
  );


  buf
  g957
  (
    n987,
    n966
  );


  not
  g958
  (
    n997,
    n966
  );


  not
  g959
  (
    n985,
    n969
  );


  buf
  g960
  (
    n999,
    n964
  );


  buf
  g961
  (
    n989,
    n967
  );


  not
  g962
  (
    n1000,
    n964
  );


  buf
  g963
  (
    n990,
    n967
  );


  not
  g964
  (
    n981,
    n965
  );


  buf
  g965
  (
    n994,
    n965
  );


  not
  g966
  (
    n980,
    n966
  );


  buf
  g967
  (
    n982,
    n966
  );


  buf
  g968
  (
    n1001,
    n969
  );


  not
  g969
  (
    n984,
    n968
  );


  buf
  g970
  (
    n986,
    n964
  );


  xnor
  g971
  (
    KeyWire_0_63,
    n980,
    n981,
    n982
  );


  nor
  g972
  (
    n1002,
    n988,
    n984,
    n983
  );


  and
  g973
  (
    n1010,
    n988,
    n989,
    n981,
    n985
  );


  nor
  g974
  (
    n1005,
    n982,
    n987,
    n980,
    n983
  );


  nand
  g975
  (
    KeyWire_0_28,
    n986,
    n983,
    n982,
    n988
  );


  nor
  g976
  (
    n1004,
    n987,
    n990,
    n986,
    n989
  );


  nor
  g977
  (
    n1006,
    n980,
    n982,
    n989,
    n990
  );


  nand
  g978
  (
    n1012,
    n986,
    n980,
    n990,
    n985
  );


  xor
  g979
  (
    n1008,
    n985,
    n985,
    n984,
    n987
  );


  xnor
  g980
  (
    n1007,
    n989,
    n988,
    n987,
    n981
  );


  xnor
  g981
  (
    n1009,
    n986,
    n990,
    n984,
    n983
  );


  and
  g982
  (
    n1021,
    n815,
    n817,
    n816
  );


  or
  g983
  (
    n1015,
    n815,
    n816,
    n729
  );


  nor
  g984
  (
    n1020,
    n956,
    n1011,
    n727,
    n728
  );


  nand
  g985
  (
    n1016,
    n928,
    n818,
    n1002
  );


  or
  g986
  (
    n1019,
    n928,
    n1003,
    n729,
    n927
  );


  and
  g987
  (
    n1022,
    n1005,
    n928,
    n818,
    n728
  );


  xor
  g988
  (
    n1013,
    n1006,
    n927,
    n817,
    n1007
  );


  xor
  g989
  (
    n1017,
    n817,
    n727,
    n1010,
    n1008
  );


  xnor
  g990
  (
    n1018,
    n816,
    n728,
    n1004,
    n729
  );


  or
  g991
  (
    n1014,
    n1012,
    n956,
    n1009,
    n728
  );


  not
  g992
  (
    n1036,
    n928
  );


  buf
  g993
  (
    n1040,
    n912
  );


  buf
  g994
  (
    n1031,
    n1015
  );


  not
  g995
  (
    n1038,
    n913
  );


  not
  g996
  (
    n1033,
    n914
  );


  buf
  g997
  (
    n1034,
    n1022
  );


  not
  g998
  (
    n1029,
    n1018
  );


  buf
  g999
  (
    n1039,
    n1021
  );


  buf
  g1000
  (
    n1027,
    n1016
  );


  buf
  g1001
  (
    n1024,
    n929
  );


  not
  g1002
  (
    n1026,
    n914
  );


  buf
  g1003
  (
    n1030,
    n1020
  );


  or
  g1004
  (
    n1037,
    n1014,
    n1020
  );


  xor
  g1005
  (
    n1028,
    n929,
    n929,
    n1017,
    n930
  );


  or
  g1006
  (
    n1035,
    n913,
    n914,
    n1013,
    n930
  );


  xor
  g1007
  (
    n1032,
    n912,
    n818,
    n1022,
    n1020
  );


  nor
  g1008
  (
    n1023,
    n1020,
    n913,
    n1022
  );


  xnor
  g1009
  (
    n1025,
    n1022,
    n1021,
    n912
  );


  or
  g1010
  (
    n1041,
    n929,
    n1019,
    n1021
  );


  xor
  g1011
  (
    n1055,
    n590,
    n574,
    n1035,
    n975
  );


  nor
  g1012
  (
    n1076,
    n1039,
    n587,
    n595,
    n559
  );


  nor
  g1013
  (
    n1094,
    n572,
    n593,
    n569,
    n1033
  );


  nand
  g1014
  (
    n1091,
    n595,
    n559,
    n1037,
    n1027
  );


  xnor
  g1015
  (
    n1086,
    n581,
    n970,
    n1028,
    n554
  );


  nand
  g1016
  (
    n1048,
    n557,
    n591,
    n1026,
    n977
  );


  and
  g1017
  (
    n1087,
    n561,
    n570,
    n1023,
    n1035
  );


  nand
  g1018
  (
    n1063,
    n1031,
    n595,
    n552,
    n1032
  );


  xnor
  g1019
  (
    n1107,
    n971,
    n973,
    n555,
    n1027
  );


  xnor
  g1020
  (
    n1089,
    n549,
    n572,
    n589,
    n585
  );


  nor
  g1021
  (
    n1077,
    n578,
    n971,
    n1029,
    n1030
  );


  xnor
  g1022
  (
    n1080,
    n556,
    n563,
    n1039,
    n1026
  );


  and
  g1023
  (
    n1113,
    n583,
    n974,
    n977,
    n586
  );


  nor
  g1024
  (
    n1054,
    n972,
    n552,
    n1039,
    n556
  );


  xnor
  g1025
  (
    n1104,
    n555,
    n973,
    n573,
    n589
  );


  nand
  g1026
  (
    n1062,
    n553,
    n551,
    n581,
    n575
  );


  xnor
  g1027
  (
    KeyWire_0_40,
    n572,
    n568,
    n1040,
    n570
  );


  or
  g1028
  (
    n1070,
    n557,
    n558,
    n552,
    n563
  );


  or
  g1029
  (
    n1057,
    n566,
    n571,
    n975,
    n1041
  );


  xor
  g1030
  (
    n1106,
    n573,
    n581,
    n1038,
    n580
  );


  xnor
  g1031
  (
    n1044,
    n588,
    n579,
    n969,
    n1035
  );


  xnor
  g1032
  (
    n1112,
    n568,
    n584,
    n561,
    n564
  );


  nand
  g1033
  (
    n1042,
    n1031,
    n579,
    n1038,
    n976
  );


  and
  g1034
  (
    n1098,
    n1036,
    n1032,
    n575,
    n977
  );


  nand
  g1035
  (
    n1046,
    n974,
    n566,
    n978,
    n558
  );


  and
  g1036
  (
    n1067,
    n1034,
    n565,
    n584,
    n560
  );


  nand
  g1037
  (
    n1078,
    n594,
    n979,
    n590,
    n975
  );


  nor
  g1038
  (
    n1109,
    n553,
    n554,
    n1027,
    n584
  );


  nand
  g1039
  (
    n1071,
    n593,
    n586,
    n1037,
    n562
  );


  nor
  g1040
  (
    n1051,
    n594,
    n560,
    n562,
    n550
  );


  and
  g1041
  (
    n1090,
    n582,
    n579,
    n974,
    n592
  );


  nand
  g1042
  (
    n1116,
    n1037,
    n1024,
    n592,
    n580
  );


  xor
  g1043
  (
    n1075,
    n974,
    n586,
    n1034,
    n970
  );


  nor
  g1044
  (
    n1114,
    n560,
    n1028,
    n593
  );


  xnor
  g1045
  (
    n1052,
    n574,
    n576,
    n578,
    n554
  );


  xnor
  g1046
  (
    n1072,
    n970,
    n570,
    n1033
  );


  xor
  g1047
  (
    n1060,
    n556,
    n567,
    n976,
    n579
  );


  nand
  g1048
  (
    n1102,
    n582,
    n571,
    n567,
    n583
  );


  nand
  g1049
  (
    n1117,
    n590,
    n555,
    n1023,
    n588
  );


  or
  g1050
  (
    n1100,
    n1025,
    n553,
    n1031,
    n1036
  );


  xor
  g1051
  (
    n1081,
    n577,
    n972,
    n1034,
    n1026
  );


  or
  g1052
  (
    n1045,
    n551,
    n586,
    n587,
    n577
  );


  nand
  g1053
  (
    n1065,
    n1023,
    n565,
    n1030,
    n1041
  );


  xnor
  g1054
  (
    n1053,
    n565,
    n588,
    n1032,
    n1033
  );


  and
  g1055
  (
    n1047,
    n576,
    n561,
    n1032,
    n1031
  );


  xnor
  g1056
  (
    n1088,
    n561,
    n568,
    n972,
    n580
  );


  xnor
  g1057
  (
    KeyWire_0_10,
    n1026,
    n594,
    n1024
  );


  xor
  g1058
  (
    n1111,
    n552,
    n557,
    n589,
    n1036
  );


  nor
  g1059
  (
    n1096,
    n550,
    n1039,
    n563,
    n569
  );


  xor
  g1060
  (
    n1066,
    n567,
    n578,
    n1029,
    n550
  );


  and
  g1061
  (
    KeyWire_0_49,
    n589,
    n1041,
    n581
  );


  nand
  g1062
  (
    n1099,
    n969,
    n564,
    n978,
    n566
  );


  xnor
  g1063
  (
    n1101,
    n554,
    n978,
    n558,
    n557
  );


  xnor
  g1064
  (
    n1085,
    n563,
    n587,
    n979,
    n566
  );


  xor
  g1065
  (
    KeyWire_0_45,
    n1029,
    n551,
    n1025,
    n582
  );


  xor
  g1066
  (
    n1110,
    n1025,
    n1038,
    n1040,
    n573
  );


  or
  g1067
  (
    n1083,
    n575,
    n1035,
    n1038,
    n558
  );


  and
  g1068
  (
    KeyWire_0_30,
    n580,
    n551,
    n577,
    n590
  );


  xnor
  g1069
  (
    n1050,
    n585,
    n592,
    n1037,
    n1029
  );


  and
  g1070
  (
    n1061,
    n973,
    n568,
    n587,
    n1024
  );


  xnor
  g1071
  (
    n1058,
    n578,
    n559,
    n549,
    n978
  );


  xor
  g1072
  (
    n1092,
    n565,
    n973,
    n591,
    n575
  );


  and
  g1073
  (
    n1093,
    n1023,
    n970,
    n560,
    n1024
  );


  xnor
  g1074
  (
    n1082,
    n1040,
    n593,
    n550,
    n556
  );


  nand
  g1075
  (
    n1068,
    n583,
    n576,
    n1025
  );


  and
  g1076
  (
    n1097,
    n567,
    n559,
    n583,
    n574
  );


  or
  g1077
  (
    n1095,
    n588,
    n562,
    n976,
    n569
  );


  xnor
  g1078
  (
    n1059,
    n570,
    n1034,
    n572,
    n1027
  );


  nor
  g1079
  (
    n1105,
    n585,
    n971,
    n1028,
    n591
  );


  xnor
  g1080
  (
    n1079,
    n595,
    n584,
    n564
  );


  nor
  g1081
  (
    n1084,
    n972,
    n1036,
    n569,
    n577
  );


  xor
  g1082
  (
    n1115,
    n553,
    n976,
    n1030,
    n573
  );


  or
  g1083
  (
    n1064,
    n975,
    n562,
    n1030,
    n574
  );


  xnor
  g1084
  (
    n1108,
    n571,
    n977,
    n585,
    n1040
  );


  and
  g1085
  (
    n1049,
    n979,
    n571,
    n591,
    n971
  );


  or
  g1086
  (
    n1069,
    n979,
    n555,
    n592,
    n582
  );


  buf
  g1087
  (
    KeyWire_0_7,
    n1088
  );


  buf
  g1088
  (
    n1227,
    n729
  );


  not
  g1089
  (
    n1379,
    n688
  );


  buf
  g1090
  (
    n1157,
    n1109
  );


  buf
  g1091
  (
    n1127,
    n697
  );


  buf
  g1092
  (
    n1352,
    n1084
  );


  buf
  g1093
  (
    n1185,
    n1110
  );


  buf
  g1094
  (
    n1241,
    n1072
  );


  buf
  g1095
  (
    n1229,
    n1095
  );


  buf
  g1096
  (
    n1258,
    n1111
  );


  not
  g1097
  (
    n1167,
    n1062
  );


  buf
  g1098
  (
    n1270,
    n1000
  );


  not
  g1099
  (
    n1184,
    n1107
  );


  not
  g1100
  (
    n1187,
    n1058
  );


  buf
  g1101
  (
    n1336,
    n684
  );


  not
  g1102
  (
    n1234,
    n1070
  );


  not
  g1103
  (
    n1307,
    n670
  );


  not
  g1104
  (
    n1326,
    n1098
  );


  not
  g1105
  (
    n1226,
    n677
  );


  buf
  g1106
  (
    n1286,
    n1051
  );


  buf
  g1107
  (
    n1249,
    n681
  );


  buf
  g1108
  (
    n1180,
    n682
  );


  not
  g1109
  (
    n1351,
    n1108
  );


  not
  g1110
  (
    n1150,
    n991
  );


  not
  g1111
  (
    n1289,
    n1104
  );


  buf
  g1112
  (
    n1164,
    n671
  );


  buf
  g1113
  (
    n1162,
    n1117
  );


  buf
  g1114
  (
    n1370,
    n1094
  );


  buf
  g1115
  (
    n1342,
    n681
  );


  buf
  g1116
  (
    n1321,
    n682
  );


  buf
  g1117
  (
    n1269,
    n1046
  );


  not
  g1118
  (
    n1135,
    n1075
  );


  not
  g1119
  (
    n1247,
    n1079
  );


  not
  g1120
  (
    n1260,
    n993
  );


  buf
  g1121
  (
    n1278,
    n1098
  );


  buf
  g1122
  (
    KeyWire_0_17,
    n687
  );


  not
  g1123
  (
    n1219,
    n696
  );


  not
  g1124
  (
    n1338,
    n1099
  );


  not
  g1125
  (
    n1188,
    n995
  );


  buf
  g1126
  (
    n1346,
    n1066
  );


  buf
  g1127
  (
    n1299,
    n1087
  );


  not
  g1128
  (
    n1333,
    n1051
  );


  not
  g1129
  (
    n1385,
    n660
  );


  buf
  g1130
  (
    n1197,
    n1096
  );


  not
  g1131
  (
    n1172,
    n669
  );


  buf
  g1132
  (
    n1181,
    n1046
  );


  buf
  g1133
  (
    n1281,
    n1091
  );


  not
  g1134
  (
    n1268,
    n696
  );


  buf
  g1135
  (
    n1144,
    n1043
  );


  not
  g1136
  (
    n1245,
    n694
  );


  buf
  g1137
  (
    n1355,
    n668
  );


  not
  g1138
  (
    n1308,
    n678
  );


  buf
  g1139
  (
    n1210,
    n672
  );


  buf
  g1140
  (
    n1147,
    n1087
  );


  not
  g1141
  (
    n1262,
    n1050
  );


  not
  g1142
  (
    n1153,
    n1076
  );


  buf
  g1143
  (
    n1298,
    n1117
  );


  not
  g1144
  (
    n1177,
    n1077
  );


  buf
  g1145
  (
    n1128,
    n662
  );


  buf
  g1146
  (
    n1133,
    n954
  );


  not
  g1147
  (
    n1216,
    n1083
  );


  not
  g1148
  (
    n1345,
    n1073
  );


  buf
  g1149
  (
    n1366,
    n676
  );


  buf
  g1150
  (
    n1192,
    n1044
  );


  not
  g1151
  (
    n1330,
    n1060
  );


  buf
  g1152
  (
    n1146,
    n1115
  );


  buf
  g1153
  (
    n1118,
    n1058
  );


  buf
  g1154
  (
    n1228,
    n1102
  );


  buf
  g1155
  (
    n1362,
    n996
  );


  buf
  g1156
  (
    n1313,
    n1092
  );


  buf
  g1157
  (
    n1317,
    n1085
  );


  not
  g1158
  (
    n1374,
    n1114
  );


  not
  g1159
  (
    n1203,
    n1095
  );


  buf
  g1160
  (
    n1222,
    n1100
  );


  not
  g1161
  (
    n1137,
    n695
  );


  buf
  g1162
  (
    n1384,
    n1097
  );


  not
  g1163
  (
    n1334,
    n1086
  );


  not
  g1164
  (
    KeyWire_0_14,
    n993
  );


  not
  g1165
  (
    n1253,
    n1106
  );


  buf
  g1166
  (
    KeyWire_0_6,
    n996
  );


  buf
  g1167
  (
    n1266,
    n1080
  );


  not
  g1168
  (
    n1246,
    n1074
  );


  buf
  g1169
  (
    n1288,
    n1089
  );


  not
  g1170
  (
    KeyWire_0_26,
    n1104
  );


  not
  g1171
  (
    n1305,
    n1102
  );


  buf
  g1172
  (
    n1272,
    n1042
  );


  buf
  g1173
  (
    n1230,
    n669
  );


  buf
  g1174
  (
    n1332,
    n1052
  );


  buf
  g1175
  (
    n1171,
    n1084
  );


  buf
  g1176
  (
    n1295,
    n668
  );


  not
  g1177
  (
    n1138,
    n1075
  );


  buf
  g1178
  (
    n1195,
    n1067
  );


  buf
  g1179
  (
    n1207,
    n681
  );


  buf
  g1180
  (
    n1275,
    n1057
  );


  buf
  g1181
  (
    n1339,
    n1090
  );


  buf
  g1182
  (
    n1261,
    n1057
  );


  buf
  g1183
  (
    n1340,
    n1048
  );


  buf
  g1184
  (
    n1263,
    n914
  );


  not
  g1185
  (
    n1240,
    n1043
  );


  buf
  g1186
  (
    n1347,
    n686
  );


  not
  g1187
  (
    n1237,
    n999
  );


  buf
  g1188
  (
    n1169,
    n1108
  );


  buf
  g1189
  (
    n1165,
    n678
  );


  buf
  g1190
  (
    n1232,
    n1103
  );


  buf
  g1191
  (
    n1218,
    n1092
  );


  buf
  g1192
  (
    n1327,
    n693
  );


  buf
  g1193
  (
    n1163,
    n1103
  );


  buf
  g1194
  (
    n1325,
    n955
  );


  buf
  g1195
  (
    n1357,
    n676
  );


  buf
  g1196
  (
    n1208,
    n1053
  );


  buf
  g1197
  (
    n1331,
    n953
  );


  not
  g1198
  (
    n1130,
    n1078
  );


  buf
  g1199
  (
    n1296,
    n1063
  );


  not
  g1200
  (
    n1145,
    n677
  );


  not
  g1201
  (
    n1126,
    n1075
  );


  buf
  g1202
  (
    n1361,
    n1093
  );


  not
  g1203
  (
    n1178,
    n680
  );


  not
  g1204
  (
    n1283,
    n1042
  );


  buf
  g1205
  (
    n1182,
    n1113
  );


  not
  g1206
  (
    n1372,
    n1112
  );


  not
  g1207
  (
    n1318,
    n1112
  );


  not
  g1208
  (
    n1309,
    n661
  );


  buf
  g1209
  (
    n1252,
    n1107
  );


  not
  g1210
  (
    n1194,
    n672
  );


  buf
  g1211
  (
    n1320,
    n683
  );


  not
  g1212
  (
    n1174,
    n1049
  );


  not
  g1213
  (
    n1319,
    n1081
  );


  not
  g1214
  (
    n1121,
    n1084
  );


  not
  g1215
  (
    n1280,
    n997
  );


  not
  g1216
  (
    n1265,
    n991
  );


  not
  g1217
  (
    n1363,
    n689
  );


  buf
  g1218
  (
    n1122,
    n1094
  );


  not
  g1219
  (
    KeyWire_0_57,
    n1077
  );


  not
  g1220
  (
    n1154,
    n1109
  );


  buf
  g1221
  (
    n1139,
    n1054
  );


  not
  g1222
  (
    n1156,
    n672
  );


  buf
  g1223
  (
    n1143,
    n1056
  );


  buf
  g1224
  (
    n1380,
    n1116
  );


  not
  g1225
  (
    n1236,
    n930
  );


  buf
  g1226
  (
    n1291,
    n1067
  );


  not
  g1227
  (
    n1123,
    n1110
  );


  not
  g1228
  (
    n1341,
    n1000
  );


  not
  g1229
  (
    n1134,
    n660
  );


  buf
  g1230
  (
    n1344,
    n1090
  );


  buf
  g1231
  (
    n1142,
    n1087
  );


  not
  g1232
  (
    n1239,
    n1047
  );


  buf
  g1233
  (
    n1255,
    n667
  );


  buf
  g1234
  (
    n1206,
    n674
  );


  not
  g1235
  (
    n1383,
    n690
  );


  not
  g1236
  (
    n1368,
    n687
  );


  not
  g1237
  (
    n1186,
    n1081
  );


  not
  g1238
  (
    n1175,
    n954
  );


  buf
  g1239
  (
    n1259,
    n1093
  );


  buf
  g1240
  (
    n1140,
    n1064
  );


  buf
  g1241
  (
    n1251,
    n1072
  );


  buf
  g1242
  (
    n1354,
    n685
  );


  not
  g1243
  (
    n1277,
    n1087
  );


  not
  g1244
  (
    n1214,
    n1066
  );


  not
  g1245
  (
    n1300,
    n685
  );


  buf
  g1246
  (
    n1369,
    n1117
  );


  buf
  g1247
  (
    n1287,
    n1085
  );


  buf
  g1248
  (
    n1310,
    n679
  );


  not
  g1249
  (
    n1202,
    n1083
  );


  not
  g1250
  (
    n1364,
    n661
  );


  buf
  g1251
  (
    n1221,
    n1097
  );


  not
  g1252
  (
    n1271,
    n1105
  );


  not
  g1253
  (
    KeyWire_0_27,
    n1067
  );


  buf
  g1254
  (
    n1284,
    n999
  );


  buf
  g1255
  (
    n1170,
    n696
  );


  not
  g1256
  (
    n1224,
    n994
  );


  not
  g1257
  (
    n1302,
    n1081
  );


  buf
  g1258
  (
    KeyWire_0_0,
    n684
  );


  not
  g1259
  (
    n1343,
    n1106
  );


  not
  g1260
  (
    n1282,
    n697
  );


  buf
  g1261
  (
    n1314,
    n673
  );


  not
  g1262
  (
    n1242,
    n1094
  );


  not
  g1263
  (
    n1297,
    n1089
  );


  not
  g1264
  (
    n1276,
    n1105
  );


  buf
  g1265
  (
    n1179,
    n993
  );


  buf
  g1266
  (
    n1367,
    n1079
  );


  buf
  g1267
  (
    n1190,
    n1111
  );


  not
  g1268
  (
    n1119,
    n1094
  );


  not
  g1269
  (
    n1231,
    n1071
  );


  not
  g1270
  (
    n1131,
    n1074
  );


  buf
  g1271
  (
    n1211,
    n1100
  );


  nor
  g1272
  (
    n1204,
    n995,
    n668,
    n1063,
    n1078
  );


  xnor
  g1273
  (
    n1217,
    n1051,
    n1114,
    n1061,
    n1093
  );


  nor
  g1274
  (
    n1183,
    n999,
    n1092,
    n663,
    n1076
  );


  nor
  g1275
  (
    n1264,
    n1086,
    n775,
    n1116,
    n1077
  );


  xnor
  g1276
  (
    n1205,
    n1080,
    n693,
    n1088,
    n686
  );


  xor
  g1277
  (
    n1220,
    n676,
    n1096,
    n1099,
    n669
  );


  xnor
  g1278
  (
    n1151,
    n691,
    n1065,
    n1060
  );


  xnor
  g1279
  (
    n1293,
    n1001,
    n1051,
    n671,
    n680
  );


  or
  g1280
  (
    n1168,
    n1001,
    n1043,
    n995,
    n1068
  );


  xor
  g1281
  (
    n1301,
    n690,
    n1082,
    n693,
    n1101
  );


  and
  g1282
  (
    n1387,
    n1061,
    n1050,
    n686
  );


  nor
  g1283
  (
    n1159,
    n992,
    n685,
    n1074,
    n673
  );


  nor
  g1284
  (
    n1124,
    n687,
    n1113,
    n997,
    n678
  );


  or
  g1285
  (
    n1201,
    n688,
    n1042,
    n692,
    n1063
  );


  xnor
  g1286
  (
    n1248,
    n1079,
    n1096,
    n675,
    n685
  );


  and
  g1287
  (
    n1348,
    n1082,
    n1086,
    n693,
    n688
  );


  or
  g1288
  (
    n1199,
    n695,
    n678,
    n1081,
    n1085
  );


  or
  g1289
  (
    n1292,
    n1071,
    n691,
    n661,
    n1068
  );


  xor
  g1290
  (
    n1148,
    n1091,
    n1047,
    n697,
    n1109
  );


  and
  g1291
  (
    n1244,
    n774,
    n1055,
    n1078
  );


  xnor
  g1292
  (
    n1316,
    n1112,
    n1064,
    n1092,
    n1091
  );


  or
  g1293
  (
    n1256,
    n1063,
    n664,
    n1050,
    n992
  );


  or
  g1294
  (
    n1323,
    n1046,
    n996,
    n662,
    n1104
  );


  and
  g1295
  (
    n1267,
    n667,
    n1065,
    n1077,
    n994
  );


  nor
  g1296
  (
    n1290,
    n994,
    n1044,
    n1057,
    n954
  );


  nand
  g1297
  (
    n1322,
    n999,
    n1069,
    n664,
    n1047
  );


  xnor
  g1298
  (
    n1125,
    n694,
    n1044,
    n1053,
    n1056
  );


  xnor
  g1299
  (
    n1200,
    n1083,
    n692,
    n682,
    n1062
  );


  or
  g1300
  (
    n1233,
    n1101,
    n675,
    n776,
    n1082
  );


  xnor
  g1301
  (
    n1376,
    n694,
    n662,
    n670,
    n1073
  );


  nand
  g1302
  (
    n1196,
    n1068,
    n663,
    n992
  );


  and
  g1303
  (
    n1350,
    n683,
    n1103,
    n1076,
    n776
  );


  nand
  g1304
  (
    n1279,
    n672,
    n1045,
    n1059,
    n1115
  );


  nor
  g1305
  (
    n1315,
    n1116,
    n1059,
    n1070,
    n683
  );


  or
  g1306
  (
    n1382,
    n673,
    n680,
    n1105,
    n930
  );


  nor
  g1307
  (
    n1365,
    n1078,
    n669,
    n774,
    n991
  );


  and
  g1308
  (
    n1209,
    n1101,
    n1074,
    n1097,
    n665
  );


  nor
  g1309
  (
    n1120,
    n1062,
    n1086,
    n1073,
    n674
  );


  xnor
  g1310
  (
    n1378,
    n1045,
    n689,
    n1117,
    n668
  );


  xor
  g1311
  (
    n1257,
    n1060,
    n665,
    n1102,
    n1083
  );


  nor
  g1312
  (
    n1294,
    n1109,
    n1054,
    n660,
    n679
  );


  xor
  g1313
  (
    n1353,
    n697,
    n1042,
    n690,
    n997
  );


  nand
  g1314
  (
    n1388,
    n1114,
    n674,
    n1069,
    n775
  );


  nand
  g1315
  (
    n1176,
    n1054,
    n1115,
    n1071
  );


  nor
  g1316
  (
    n1198,
    n1049,
    n1052,
    n1090,
    n682
  );


  and
  g1317
  (
    n1193,
    n1088,
    n1099,
    n662,
    n1048
  );


  or
  g1318
  (
    n1381,
    n1088,
    n666,
    n1089,
    n695
  );


  and
  g1319
  (
    n1129,
    n1107,
    n663,
    n775,
    n1057
  );


  xnor
  g1320
  (
    n1160,
    n689,
    n671,
    n1073,
    n1116
  );


  and
  g1321
  (
    KeyWire_0_20,
    n1068,
    n955,
    n687,
    n954
  );


  or
  g1322
  (
    n1356,
    n991,
    n1100,
    n670,
    n1113
  );


  xor
  g1323
  (
    n1225,
    n1058,
    n1049,
    n1106,
    n684
  );


  nor
  g1324
  (
    n1273,
    n666,
    n1093,
    n1000,
    n1098
  );


  xor
  g1325
  (
    n1329,
    n1066,
    n775,
    n673,
    n1001
  );


  nor
  g1326
  (
    KeyWire_0_3,
    n776,
    n1070,
    n1066,
    n1106
  );


  or
  g1327
  (
    n1324,
    n1046,
    n677,
    n661,
    n1084
  );


  xor
  g1328
  (
    n1235,
    n1065,
    n679,
    n1112,
    n692
  );


  and
  g1329
  (
    n1360,
    n670,
    n1000,
    n774,
    n1053
  );


  xnor
  g1330
  (
    n1306,
    n680,
    n953,
    n1079,
    n675
  );


  xnor
  g1331
  (
    n1285,
    n679,
    n1001,
    n665,
    n1114
  );


  xor
  g1332
  (
    n1215,
    n1099,
    n996,
    n665,
    n1070
  );


  and
  g1333
  (
    n1223,
    n1100,
    n674,
    n696,
    n694
  );


  nand
  g1334
  (
    n1274,
    n1095,
    n1053,
    n955,
    n1104
  );


  or
  g1335
  (
    n1337,
    n691,
    n1055,
    n994,
    n1108
  );


  xnor
  g1336
  (
    n1132,
    n1069,
    n955,
    n1095,
    n1054
  );


  or
  g1337
  (
    n1303,
    n998,
    n1043,
    n1064,
    n1102
  );


  and
  g1338
  (
    n1238,
    n1048,
    n1044,
    n1069,
    n997
  );


  or
  g1339
  (
    n1152,
    n993,
    n1059,
    n1111,
    n1097
  );


  or
  g1340
  (
    n1189,
    n1061,
    n666,
    n1052,
    n1091
  );


  xor
  g1341
  (
    n1304,
    n683,
    n1050,
    n953,
    n1045
  );


  xnor
  g1342
  (
    n1335,
    n1108,
    n664,
    n1085,
    n1113
  );


  nand
  g1343
  (
    n1311,
    n692,
    n1110,
    n1075,
    n1090
  );


  xor
  g1344
  (
    n1373,
    n1048,
    n998,
    n688,
    n1060
  );


  xor
  g1345
  (
    n1371,
    n1072,
    n1067,
    n676,
    n684
  );


  xnor
  g1346
  (
    n1328,
    n1049,
    n677,
    n689,
    n1056
  );


  xor
  g1347
  (
    n1358,
    n1062,
    n681,
    n1101,
    n1061
  );


  and
  g1348
  (
    n1250,
    n1071,
    n1098,
    n1059,
    n992
  );


  and
  g1349
  (
    n1312,
    n952,
    n774,
    n1047,
    n691
  );


  or
  g1350
  (
    n1213,
    n1064,
    n1080,
    n1058
  );


  nand
  g1351
  (
    n1191,
    n1052,
    n1082,
    n1076,
    n776
  );


  nor
  g1352
  (
    n1141,
    n1105,
    n667,
    n1072,
    n1096
  );


  and
  g1353
  (
    n1161,
    n1107,
    n1055,
    n952,
    n695
  );


  nor
  g1354
  (
    n1243,
    n998,
    n1056,
    n667,
    n671
  );


  nor
  g1355
  (
    n1166,
    n1110,
    n664,
    n1089,
    n1045
  );


  nor
  g1356
  (
    n1158,
    n690,
    n953,
    n995,
    n666
  );


  and
  g1357
  (
    n1212,
    n675,
    n1103,
    n998,
    n1111
  );


  nor
  g1358
  (
    n1441,
    n1354,
    n1205,
    n1129,
    n1216
  );


  nand
  g1359
  (
    n1416,
    n1188,
    n1192,
    n1118,
    n1139
  );


  and
  g1360
  (
    n1406,
    n1258,
    n1120,
    n1374,
    n1283
  );


  xnor
  g1361
  (
    n1442,
    n1232,
    n1353,
    n1328,
    n1274
  );


  nand
  g1362
  (
    n1411,
    n1160,
    n1231,
    n1256,
    n1313
  );


  or
  g1363
  (
    n1430,
    n1127,
    n1380,
    n1195,
    n1329
  );


  xor
  g1364
  (
    n1440,
    n1336,
    n1255,
    n1164,
    n1133
  );


  nor
  g1365
  (
    n1447,
    n1292,
    n1306,
    n1239,
    n1135
  );


  or
  g1366
  (
    n1446,
    n1257,
    n1279,
    n1251,
    n1348
  );


  nand
  g1367
  (
    n1432,
    n1125,
    n1370,
    n1134,
    n1181
  );


  xor
  g1368
  (
    n1395,
    n1153,
    n1298,
    n1140,
    n1335
  );


  xor
  g1369
  (
    n1434,
    n1371,
    n1237,
    n1322,
    n1361
  );


  nand
  g1370
  (
    n1410,
    n1185,
    n1148,
    n1282,
    n1357
  );


  xnor
  g1371
  (
    n1427,
    n1327,
    n1286,
    n1199,
    n1377
  );


  nand
  g1372
  (
    n1445,
    n1180,
    n1310,
    n1303,
    n1320
  );


  xnor
  g1373
  (
    n1423,
    n1356,
    n1280,
    n1271,
    n1152
  );


  and
  g1374
  (
    n1452,
    n1189,
    n1291,
    n1200,
    n1247
  );


  nor
  g1375
  (
    n1415,
    n1159,
    n1224,
    n1318,
    n1171
  );


  nand
  g1376
  (
    n1394,
    n1349,
    n1208,
    n1337,
    n1317
  );


  xnor
  g1377
  (
    n1397,
    n1342,
    n1272,
    n1381,
    n1379
  );


  nor
  g1378
  (
    n1437,
    n1131,
    n1254,
    n1297,
    n1220
  );


  or
  g1379
  (
    n1409,
    n1301,
    n1369,
    n1172,
    n1176
  );


  nand
  g1380
  (
    n1436,
    n1333,
    n1136,
    n1215,
    n1162
  );


  xnor
  g1381
  (
    n1439,
    n1157,
    n1229,
    n1124,
    n1248
  );


  xnor
  g1382
  (
    n1396,
    n1341,
    n1163,
    n1223,
    n1260
  );


  xnor
  g1383
  (
    n1408,
    n1352,
    n1177,
    n1193,
    n1363
  );


  xor
  g1384
  (
    n1421,
    n1326,
    n1373,
    n1230,
    n1305
  );


  xor
  g1385
  (
    n1438,
    n1145,
    n1222,
    n1187,
    n1197
  );


  and
  g1386
  (
    n1431,
    n1285,
    n1364,
    n1347,
    n1156
  );


  nor
  g1387
  (
    n1425,
    n1267,
    n1319,
    n1170,
    n1375
  );


  and
  g1388
  (
    n1414,
    n1385,
    n1281,
    n1179,
    n1138
  );


  or
  g1389
  (
    n1404,
    n1294,
    n1144,
    n1234,
    n1128
  );


  xnor
  g1390
  (
    n1435,
    n1201,
    n1288,
    n1266,
    n1209
  );


  nor
  g1391
  (
    n1407,
    n1250,
    n1241,
    n1240,
    n1167
  );


  nand
  g1392
  (
    n1398,
    n1372,
    n1264,
    n1228,
    n1242
  );


  and
  g1393
  (
    n1412,
    n1293,
    n1270,
    n1206,
    n1307
  );


  or
  g1394
  (
    n1399,
    n1233,
    n1161,
    n1304,
    n1277
  );


  xor
  g1395
  (
    n1402,
    n1225,
    n1296,
    n1269,
    n1386
  );


  nor
  g1396
  (
    n1455,
    n1299,
    n1360,
    n1121,
    n1236
  );


  xor
  g1397
  (
    n1420,
    n1150,
    n1166,
    n1122,
    n1249
  );


  nor
  g1398
  (
    n1391,
    n1334,
    n1142,
    n1343,
    n1244
  );


  xnor
  g1399
  (
    n1433,
    n1202,
    n1173,
    n1332,
    n1366
  );


  nand
  g1400
  (
    n1392,
    n1323,
    n1265,
    n1221,
    n1194
  );


  xor
  g1401
  (
    n1405,
    n1315,
    n1155,
    n1132,
    n1126
  );


  nor
  g1402
  (
    n1389,
    n1227,
    n1316,
    n1289,
    n1290
  );


  xnor
  g1403
  (
    n1429,
    n1218,
    n1190,
    n1183,
    n1235
  );


  or
  g1404
  (
    KeyWire_0_29,
    n1308,
    n1219,
    n1330,
    n1245
  );


  xnor
  g1405
  (
    n1403,
    n1340,
    n1154,
    n1324,
    n1355
  );


  and
  g1406
  (
    n1450,
    n1149,
    n1368,
    n1212,
    n1226
  );


  nand
  g1407
  (
    KeyWire_0_53,
    n1275,
    n1210,
    n1146,
    n1273
  );


  nor
  g1408
  (
    n1443,
    n1262,
    n1376,
    n1178,
    n1169
  );


  xor
  g1409
  (
    n1451,
    n1268,
    n1331,
    n1350,
    n1174
  );


  nand
  g1410
  (
    n1456,
    n1309,
    n1191,
    n1362,
    n1182
  );


  xor
  g1411
  (
    n1393,
    n1147,
    n1253,
    n1312,
    n1278
  );


  nand
  g1412
  (
    n1390,
    n1238,
    n1158,
    n1339,
    n1365
  );


  or
  g1413
  (
    n1424,
    n1211,
    n1314,
    n1203,
    n1130
  );


  xor
  g1414
  (
    n1448,
    n1261,
    n1143,
    n1338,
    n1311
  );


  xnor
  g1415
  (
    KeyWire_0_2,
    n1123,
    n1378,
    n1213,
    n1263
  );


  and
  g1416
  (
    n1454,
    n1246,
    n1367,
    n1302,
    n1186
  );


  and
  g1417
  (
    n1413,
    n1295,
    n150,
    n1325,
    n1276
  );


  nand
  g1418
  (
    n1422,
    n1252,
    n1346,
    n1184,
    n1284
  );


  xor
  g1419
  (
    n1417,
    n1137,
    n1198,
    n1345,
    n1141
  );


  nand
  g1420
  (
    n1444,
    n1214,
    n1119,
    n1175,
    n1382
  );


  xor
  g1421
  (
    n1453,
    n1204,
    n1344,
    n1217,
    n1387
  );


  and
  g1422
  (
    n1428,
    n1287,
    n1243,
    n1165,
    n1383
  );


  xnor
  g1423
  (
    n1401,
    n1351,
    n1388,
    n1168,
    n1196
  );


  xnor
  g1424
  (
    n1419,
    n1259,
    n1358,
    n1384,
    n1321
  );


  and
  g1425
  (
    n1426,
    n1359,
    n1300,
    n1207,
    n1151
  );


  or
  g1426
  (
    n1463,
    n1402,
    n1389,
    n1409,
    n1449
  );


  and
  g1427
  (
    n1470,
    n1424,
    n1455,
    n1407,
    n1440
  );


  nand
  g1428
  (
    n1459,
    n1448,
    n1435,
    n1410,
    n1419
  );


  xnor
  g1429
  (
    n1464,
    n1427,
    n1416,
    n1450,
    n1403
  );


  xnor
  g1430
  (
    n1458,
    n1444,
    n1453,
    n1446,
    n1436
  );


  xor
  g1431
  (
    n1467,
    n1443,
    n1406,
    n1415,
    n1445
  );


  or
  g1432
  (
    n1472,
    n1456,
    n1439,
    n1441,
    n1428
  );


  or
  g1433
  (
    n1460,
    n1417,
    n1425,
    n1411,
    n1392
  );


  nor
  g1434
  (
    n1469,
    n1447,
    n1399,
    n1432,
    n1414
  );


  and
  g1435
  (
    n1466,
    n1400,
    n1405,
    n1434,
    n1430
  );


  xnor
  g1436
  (
    n1473,
    n1390,
    n1426,
    n1396,
    n1404
  );


  and
  g1437
  (
    n1471,
    n1442,
    n1420,
    n1429,
    n1452
  );


  xor
  g1438
  (
    KeyWire_0_43,
    n1401,
    n1423,
    n1437,
    n1433
  );


  nor
  g1439
  (
    n1468,
    n1438,
    n1408,
    n1393,
    n1413
  );


  nand
  g1440
  (
    n1457,
    n1451,
    n1431,
    n1397,
    n1422
  );


  xor
  g1441
  (
    n1461,
    n1412,
    n1391,
    n1395,
    n1394
  );


  nor
  g1442
  (
    n1462,
    n1421,
    n1454,
    n1418,
    n1398
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1377,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n408,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1418,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n1149,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n640,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n884,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1155,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1173,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n142,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n135,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1074,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n314,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n316,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n926,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1375,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n590,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n600,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n1136,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n79,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n169,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1349,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n505,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n627,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n410,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n943,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n70,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1254,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1386,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1003,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n1449,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1103,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n338,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n613,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n605,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n246,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n482,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n536,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n859,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n363,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n330,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n1073,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n850,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n46,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n1465,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n677,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n1043,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n676,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n266,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n804,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n1056,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n415,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n418,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n870,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n1400,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n84,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n991,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n871,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n1359,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n125,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n584,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n115,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n337,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n243,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n1011,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


