// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_164_430 written by SynthGen on 2021/05/24 19:45:41
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_164_430 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31,
 n181, n193, n178, n189, n179, n184, n183, n182,
 n194, n186, n188, n192, n190, n191, n180, n195,
 n187, n185);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31;

output n181, n193, n178, n189, n179, n184, n183, n182,
 n194, n186, n188, n192, n190, n191, n180, n195,
 n187, n185;

wire n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177;

not  g0 (n53, n12);
buf  g1 (n43, n10);
buf  g2 (n85, n30);
not  g3 (n113, n3);
buf  g4 (n46, n5);
buf  g5 (n66, n22);
buf  g6 (n82, n21);
not  g7 (n130, n20);
not  g8 (n68, n22);
buf  g9 (n126, n11);
not  g10 (n119, n4);
not  g11 (n98, n18);
not  g12 (n110, n9);
buf  g13 (n77, n28);
buf  g14 (n79, n4);
buf  g15 (n102, n30);
not  g16 (n76, n12);
not  g17 (n57, n1);
not  g18 (n78, n20);
not  g19 (n33, n22);
buf  g20 (n70, n8);
buf  g21 (n47, n29);
not  g22 (n115, n2);
not  g23 (n95, n1);
buf  g24 (n106, n29);
not  g25 (n51, n27);
buf  g26 (n101, n17);
not  g27 (n59, n31);
buf  g28 (n122, n13);
not  g29 (n92, n27);
buf  g30 (n75, n19);
not  g31 (n73, n1);
not  g32 (n114, n17);
buf  g33 (n36, n6);
buf  g34 (n118, n11);
not  g35 (n135, n21);
not  g36 (n134, n24);
not  g37 (n72, n26);
buf  g38 (n49, n19);
buf  g39 (n67, n7);
not  g40 (n54, n23);
buf  g41 (n50, n6);
not  g42 (n99, n29);
buf  g43 (n87, n23);
not  g44 (n38, n16);
not  g45 (n121, n14);
not  g46 (n133, n23);
buf  g47 (n40, n28);
buf  g48 (n91, n2);
not  g49 (n80, n26);
buf  g50 (n63, n26);
buf  g51 (n90, n28);
not  g52 (n55, n25);
buf  g53 (n105, n7);
buf  g54 (n127, n24);
not  g55 (n35, n8);
buf  g56 (n52, n28);
buf  g57 (n56, n21);
buf  g58 (n132, n2);
not  g59 (n88, n30);
not  g60 (n74, n13);
buf  g61 (n111, n26);
buf  g62 (n93, n24);
buf  g63 (n97, n30);
buf  g64 (n64, n25);
buf  g65 (n83, n19);
buf  g66 (n103, n22);
not  g67 (n58, n31);
not  g68 (n107, n12);
not  g69 (n125, n4);
not  g70 (n104, n8);
not  g71 (n116, n21);
not  g72 (n128, n5);
buf  g73 (n108, n19);
buf  g74 (n34, n9);
buf  g75 (n136, n27);
not  g76 (n44, n3);
buf  g77 (n62, n9);
buf  g78 (n42, n17);
not  g79 (n112, n7);
not  g80 (n100, n3);
buf  g81 (n45, n20);
buf  g82 (n81, n10);
buf  g83 (n60, n10);
buf  g84 (n32, n13);
not  g85 (n41, n16);
buf  g86 (n65, n6);
buf  g87 (n69, n24);
not  g88 (n137, n15);
not  g89 (n123, n14);
buf  g90 (n48, n5);
not  g91 (n129, n15);
buf  g92 (n124, n25);
not  g93 (n71, n18);
buf  g94 (n89, n31);
buf  g95 (n37, n11);
buf  g96 (n86, n20);
buf  g97 (n131, n31);
not  g98 (n96, n16);
buf  g99 (n109, n23);
not  g100 (n84, n18);
buf  g101 (n39, n25);
buf  g102 (n117, n29);
not  g103 (n120, n14);
not  g104 (n61, n15);
not  g105 (n94, n27);
buf  g106 (n140, n44);
buf  g107 (n149, n43);
not  g108 (n142, n48);
not  g109 (n148, n49);
buf  g110 (n155, n47);
not  g111 (n139, n32);
not  g112 (n153, n53);
buf  g113 (n151, n36);
not  g114 (n141, n38);
buf  g115 (n152, n46);
buf  g116 (n145, n37);
not  g117 (n150, n33);
not  g118 (n154, n34);
not  g119 (n144, n41);
buf  g120 (n147, n51);
buf  g121 (n143, n52);
buf  g122 (n156, n40);
not  g123 (n138, n42);
not  g124 (n157, n39);
buf  g125 (n158, n45);
nand g126 (n146, n50, n35);
not  g127 (n163, n54);
buf  g128 (n159, n55);
not  g129 (n167, n148);
not  g130 (n162, n69);
buf  g131 (n160, n84);
not  g132 (n164, n146);
and  g133 (n172, n71, n153);
xnor g134 (n165, n85, n67);
nor  g135 (n174, n142, n86);
nor  g136 (n169, n73, n81, n143, n64);
and  g137 (n168, n61, n140, n78, n80);
and  g138 (n175, n145, n141, n151, n72);
xor  g139 (n161, n77, n65, n62, n144);
xnor g140 (n171, n138, n68, n83, n156);
xnor g141 (n170, n63, n57, n139, n60);
and  g142 (n166, n70, n149, n154, n58);
or   g143 (n176, n66, n74, n76, n155);
nand g144 (n173, n56, n75, n147, n150);
and  g145 (n177, n152, n82, n59, n79);
xnor g146 (n195, n103, n134, n176, n177);
and  g147 (n188, n137, n93, n112, n92);
or   g148 (n190, n124, n115, n88, n131);
nand g149 (n184, n104, n135, n173, n105);
and  g150 (n194, n163, n161, n175, n128);
xor  g151 (n189, n167, n127, n117, n174);
xnor g152 (n192, n97, n106, n125, n120);
or   g153 (n180, n90, n101, n165, n116);
and  g154 (n179, n94, n87, n126, n136);
or   g155 (n193, n133, n102, n108, n157);
xnor g156 (n186, n166, n118, n164, n119);
or   g157 (n183, n99, n114, n98, n121);
and  g158 (n182, n169, n111, n162, n168);
nor  g159 (n191, n113, n130, n123, n107);
and  g160 (n187, n122, n160, n170, n96);
xnor g161 (n185, n132, n110, n159, n172);
and  g162 (n178, n100, n171, n95, n129);
nand g163 (n181, n158, n91, n109, n89);
endmodule
