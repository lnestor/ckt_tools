

module Stat_834_381
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n177,
  n183,
  n175,
  n176,
  n192,
  n194,
  n181,
  n186,
  n196,
  n189,
  n590,
  n597,
  n587,
  n840,
  n852,
  n854,
  n860,
  n861,
  n865
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n177;output n183;output n175;output n176;output n192;output n194;output n181;output n186;output n196;output n189;output n590;output n597;output n587;output n840;output n852;output n854;output n860;output n861;output n865;
  wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n178;wire n179;wire n180;wire n182;wire n184;wire n185;wire n187;wire n188;wire n190;wire n191;wire n193;wire n195;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n588;wire n589;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n853;wire n855;wire n856;wire n857;wire n858;wire n859;wire n862;wire n863;wire n864;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n64,
    n9
  );


  not
  g1
  (
    n33,
    n25
  );


  not
  g2
  (
    n47,
    n23
  );


  not
  g3
  (
    n83,
    n3
  );


  not
  g4
  (
    KeyWire_0_3,
    n8
  );


  buf
  g5
  (
    n74,
    n12
  );


  not
  g6
  (
    n77,
    n27
  );


  buf
  g7
  (
    n49,
    n30
  );


  not
  g8
  (
    n93,
    n25
  );


  not
  g9
  (
    n34,
    n10
  );


  buf
  g10
  (
    n106,
    n14
  );


  buf
  g11
  (
    n105,
    n5
  );


  buf
  g12
  (
    KeyWire_0_18,
    n10
  );


  not
  g13
  (
    n78,
    n15
  );


  not
  g14
  (
    n109,
    n13
  );


  not
  g15
  (
    n69,
    n6
  );


  not
  g16
  (
    n118,
    n10
  );


  buf
  g17
  (
    n44,
    n20
  );


  not
  g18
  (
    n97,
    n31
  );


  not
  g19
  (
    n68,
    n30
  );


  not
  g20
  (
    n96,
    n14
  );


  buf
  g21
  (
    n115,
    n5
  );


  buf
  g22
  (
    n98,
    n27
  );


  buf
  g23
  (
    n42,
    n18
  );


  buf
  g24
  (
    n95,
    n19
  );


  buf
  g25
  (
    n41,
    n12
  );


  buf
  g26
  (
    n123,
    n5
  );


  not
  g27
  (
    n122,
    n6
  );


  buf
  g28
  (
    n54,
    n21
  );


  buf
  g29
  (
    n50,
    n26
  );


  buf
  g30
  (
    n103,
    n15
  );


  buf
  g31
  (
    n101,
    n16
  );


  not
  g32
  (
    n121,
    n20
  );


  buf
  g33
  (
    n84,
    n4
  );


  buf
  g34
  (
    n38,
    n11
  );


  buf
  g35
  (
    n37,
    n29
  );


  not
  g36
  (
    n85,
    n24
  );


  buf
  g37
  (
    n51,
    n16
  );


  not
  g38
  (
    n46,
    n31
  );


  buf
  g39
  (
    n32,
    n3
  );


  not
  g40
  (
    n53,
    n1
  );


  not
  g41
  (
    n90,
    n18
  );


  not
  g42
  (
    n110,
    n17
  );


  not
  g43
  (
    n35,
    n27
  );


  buf
  g44
  (
    n89,
    n7
  );


  not
  g45
  (
    n56,
    n28
  );


  buf
  g46
  (
    n111,
    n2
  );


  buf
  g47
  (
    n102,
    n30
  );


  not
  g48
  (
    n100,
    n31
  );


  not
  g49
  (
    n72,
    n6
  );


  not
  g50
  (
    n71,
    n2
  );


  not
  g51
  (
    n60,
    n4
  );


  not
  g52
  (
    n79,
    n13
  );


  not
  g53
  (
    n108,
    n7
  );


  not
  g54
  (
    n65,
    n9
  );


  buf
  g55
  (
    n91,
    n1
  );


  buf
  g56
  (
    n63,
    n17
  );


  buf
  g57
  (
    n99,
    n26
  );


  buf
  g58
  (
    n66,
    n8
  );


  buf
  g59
  (
    n45,
    n13
  );


  not
  g60
  (
    n57,
    n28
  );


  buf
  g61
  (
    n82,
    n25
  );


  buf
  g62
  (
    n70,
    n4
  );


  buf
  g63
  (
    n39,
    n1
  );


  buf
  g64
  (
    n117,
    n21
  );


  buf
  g65
  (
    n58,
    n17
  );


  not
  g66
  (
    n59,
    n7
  );


  buf
  g67
  (
    n114,
    n24
  );


  not
  g68
  (
    n107,
    n19
  );


  not
  g69
  (
    n86,
    n22
  );


  buf
  g70
  (
    n67,
    n22
  );


  buf
  g71
  (
    n76,
    n23
  );


  buf
  g72
  (
    n52,
    n16
  );


  buf
  g73
  (
    n62,
    n21
  );


  not
  g74
  (
    n113,
    n11
  );


  not
  g75
  (
    n55,
    n3
  );


  not
  g76
  (
    n104,
    n20
  );


  buf
  g77
  (
    n81,
    n19
  );


  buf
  g78
  (
    n119,
    n22
  );


  buf
  g79
  (
    n40,
    n12
  );


  buf
  g80
  (
    n87,
    n2
  );


  not
  g81
  (
    n112,
    n18
  );


  not
  g82
  (
    n94,
    n8
  );


  not
  g83
  (
    KeyWire_0_14,
    n28
  );


  buf
  g84
  (
    n120,
    n26
  );


  buf
  g85
  (
    n73,
    n15
  );


  not
  g86
  (
    n124,
    n29
  );


  not
  g87
  (
    n75,
    n29
  );


  buf
  g88
  (
    n48,
    n24
  );


  not
  g89
  (
    n116,
    n11
  );


  not
  g90
  (
    n80,
    n14
  );


  buf
  g91
  (
    n88,
    n9
  );


  not
  g92
  (
    n43,
    n23
  );


  buf
  g93
  (
    n170,
    n41
  );


  not
  g94
  (
    n145,
    n59
  );


  not
  g95
  (
    n160,
    n79
  );


  buf
  g96
  (
    n159,
    n55
  );


  not
  g97
  (
    n136,
    n49
  );


  buf
  g98
  (
    n167,
    n59
  );


  not
  g99
  (
    n157,
    n44
  );


  buf
  g100
  (
    n152,
    n73
  );


  buf
  g101
  (
    n132,
    n76
  );


  nand
  g102
  (
    n137,
    n60,
    n62
  );


  or
  g103
  (
    n171,
    n58,
    n62,
    n84,
    n80
  );


  nand
  g104
  (
    n133,
    n77,
    n51,
    n74
  );


  xnor
  g105
  (
    KeyWire_0_10,
    n44,
    n52,
    n58,
    n87
  );


  nor
  g106
  (
    n166,
    n76,
    n32,
    n68,
    n81
  );


  xnor
  g107
  (
    n150,
    n61,
    n32,
    n46,
    n54
  );


  xnor
  g108
  (
    n165,
    n37,
    n86,
    n36,
    n87
  );


  and
  g109
  (
    n155,
    n43,
    n69,
    n64,
    n40
  );


  xor
  g110
  (
    n172,
    n51,
    n64,
    n63,
    n86
  );


  xor
  g111
  (
    n144,
    n49,
    n70,
    n45,
    n60
  );


  xor
  g112
  (
    n128,
    n80,
    n75,
    n50
  );


  nand
  g113
  (
    n158,
    n57,
    n43,
    n42,
    n66
  );


  xnor
  g114
  (
    n127,
    n41,
    n72,
    n83,
    n74
  );


  xor
  g115
  (
    n139,
    n35,
    n72,
    n85,
    n67
  );


  nor
  g116
  (
    n151,
    n67,
    n85,
    n77,
    n65
  );


  xor
  g117
  (
    n129,
    n73,
    n78,
    n50,
    n39
  );


  and
  g118
  (
    n135,
    n71,
    n66,
    n36,
    n62
  );


  xor
  g119
  (
    n156,
    n44,
    n40,
    n79,
    n33
  );


  or
  g120
  (
    n126,
    n63,
    n85,
    n71,
    n84
  );


  nor
  g121
  (
    n163,
    n82,
    n48,
    n46,
    n84
  );


  and
  g122
  (
    n148,
    n48,
    n35,
    n82,
    n56
  );


  xnor
  g123
  (
    n162,
    n69,
    n64,
    n53,
    n49
  );


  and
  g124
  (
    n154,
    n61,
    n55,
    n72,
    n78
  );


  or
  g125
  (
    n169,
    n71,
    n39,
    n37,
    n35
  );


  xnor
  g126
  (
    n168,
    n83,
    n55,
    n33,
    n76
  );


  nand
  g127
  (
    n141,
    n47,
    n81,
    n51,
    n50
  );


  or
  g128
  (
    n164,
    n48,
    n38
  );


  and
  g129
  (
    n138,
    n37,
    n56,
    n34,
    n79
  );


  or
  g130
  (
    n134,
    n39,
    n61,
    n34,
    n57
  );


  nand
  g131
  (
    n173,
    n33,
    n69,
    n36,
    n60
  );


  xor
  g132
  (
    n146,
    n47,
    n65,
    n45,
    n56
  );


  xnor
  g133
  (
    n143,
    n57,
    n83,
    n54,
    n80
  );


  or
  g134
  (
    n142,
    n43,
    n75,
    n86,
    n59
  );


  xor
  g135
  (
    n130,
    n82,
    n52,
    n70
  );


  or
  g136
  (
    n161,
    n70,
    n77,
    n67,
    n66
  );


  or
  g137
  (
    n125,
    n41,
    n46,
    n42
  );


  xor
  g138
  (
    n153,
    n40,
    n78,
    n65,
    n32
  );


  and
  g139
  (
    n147,
    n47,
    n58,
    n53,
    n68
  );


  nand
  g140
  (
    n140,
    n53,
    n45,
    n81,
    n54
  );


  or
  g141
  (
    n131,
    n73,
    n68,
    n34,
    n63
  );


  not
  g142
  (
    n197,
    n126
  );


  not
  g143
  (
    n194,
    n140
  );


  buf
  g144
  (
    n195,
    n133
  );


  buf
  g145
  (
    n174,
    n152
  );


  not
  g146
  (
    n181,
    n128
  );


  buf
  g147
  (
    n200,
    n146
  );


  buf
  g148
  (
    n180,
    n138
  );


  buf
  g149
  (
    n182,
    n127
  );


  not
  g150
  (
    n198,
    n145
  );


  not
  g151
  (
    n183,
    n141
  );


  not
  g152
  (
    KeyWire_0_13,
    n139
  );


  buf
  g153
  (
    n189,
    n137
  );


  not
  g154
  (
    n185,
    n142
  );


  buf
  g155
  (
    n201,
    n136
  );


  buf
  g156
  (
    n190,
    n149
  );


  buf
  g157
  (
    n184,
    n129
  );


  buf
  g158
  (
    n193,
    n125
  );


  buf
  g159
  (
    n177,
    n144
  );


  not
  g160
  (
    KeyWire_0_30,
    n130
  );


  buf
  g161
  (
    n187,
    n143
  );


  buf
  g162
  (
    n186,
    n134
  );


  buf
  g163
  (
    n196,
    n132
  );


  not
  g164
  (
    n199,
    n151
  );


  buf
  g165
  (
    n176,
    n148
  );


  buf
  g166
  (
    n192,
    n147
  );


  not
  g167
  (
    n188,
    n131
  );


  not
  g168
  (
    n191,
    n135
  );


  buf
  g169
  (
    n175,
    n150
  );


  not
  g170
  (
    n205,
    n89
  );


  not
  g171
  (
    n210,
    n89
  );


  buf
  g172
  (
    n213,
    n197
  );


  buf
  g173
  (
    n206,
    n198
  );


  not
  g174
  (
    n216,
    n190
  );


  buf
  g175
  (
    n207,
    n192
  );


  not
  g176
  (
    KeyWire_0_25,
    n191
  );


  not
  g177
  (
    n204,
    n193
  );


  not
  g178
  (
    n212,
    n186
  );


  buf
  g179
  (
    n203,
    n187
  );


  buf
  g180
  (
    n219,
    n201
  );


  not
  g181
  (
    n209,
    n194
  );


  buf
  g182
  (
    n208,
    n195
  );


  not
  g183
  (
    n214,
    n199
  );


  nor
  g184
  (
    n218,
    n89,
    n88
  );


  nor
  g185
  (
    n211,
    n196,
    n88,
    n188,
    n90
  );


  nand
  g186
  (
    n217,
    n184,
    n200,
    n90,
    n88
  );


  and
  g187
  (
    n202,
    n189,
    n87,
    n185,
    n90
  );


  buf
  g188
  (
    n223,
    n208
  );


  not
  g189
  (
    n222,
    n202
  );


  and
  g190
  (
    n220,
    n206,
    n209
  );


  xnor
  g191
  (
    n227,
    n203,
    n210
  );


  and
  g192
  (
    n228,
    n209,
    n206,
    n204,
    n205
  );


  and
  g193
  (
    n226,
    n203,
    n205,
    n209,
    n210
  );


  nor
  g194
  (
    n225,
    n208,
    n211,
    n210,
    n202
  );


  xor
  g195
  (
    n229,
    n207,
    n206,
    n211,
    n208
  );


  xnor
  g196
  (
    n221,
    n204,
    n202,
    n207,
    n211
  );


  nor
  g197
  (
    n224,
    n203,
    n205,
    n204,
    n207
  );


  buf
  g198
  (
    n236,
    n226
  );


  buf
  g199
  (
    n231,
    n227
  );


  not
  g200
  (
    n234,
    n225
  );


  not
  g201
  (
    n230,
    n222
  );


  buf
  g202
  (
    n232,
    n221
  );


  buf
  g203
  (
    n238,
    n224
  );


  buf
  g204
  (
    n237,
    n223
  );


  not
  g205
  (
    n235,
    n228
  );


  not
  g206
  (
    n233,
    n220
  );


  not
  g207
  (
    n240,
    n235
  );


  not
  g208
  (
    n241,
    n236
  );


  not
  g209
  (
    n247,
    n232
  );


  not
  g210
  (
    n239,
    n231
  );


  not
  g211
  (
    n254,
    n232
  );


  not
  g212
  (
    n257,
    n235
  );


  buf
  g213
  (
    n255,
    n236
  );


  buf
  g214
  (
    n243,
    n234
  );


  not
  g215
  (
    n251,
    n233
  );


  buf
  g216
  (
    n242,
    n233
  );


  buf
  g217
  (
    n244,
    n232
  );


  buf
  g218
  (
    KeyWire_0_8,
    n230
  );


  not
  g219
  (
    n246,
    n234
  );


  not
  g220
  (
    n250,
    n230
  );


  not
  g221
  (
    n248,
    n231
  );


  buf
  g222
  (
    n256,
    n231
  );


  buf
  g223
  (
    n249,
    n234
  );


  not
  g224
  (
    n252,
    n233
  );


  buf
  g225
  (
    n253,
    n235
  );


  buf
  g226
  (
    n258,
    n230
  );


  buf
  g227
  (
    n272,
    n244
  );


  not
  g228
  (
    n264,
    n212
  );


  not
  g229
  (
    n285,
    n216
  );


  not
  g230
  (
    n283,
    n251
  );


  not
  g231
  (
    n280,
    n246
  );


  buf
  g232
  (
    n259,
    n242
  );


  buf
  g233
  (
    n282,
    n258
  );


  not
  g234
  (
    n278,
    n249
  );


  not
  g235
  (
    n267,
    n213
  );


  not
  g236
  (
    n274,
    n243
  );


  buf
  g237
  (
    n269,
    n249
  );


  not
  g238
  (
    n270,
    n153
  );


  xor
  g239
  (
    n276,
    n216,
    n255,
    n239,
    n248
  );


  xor
  g240
  (
    n260,
    n244,
    n256,
    n240,
    n248
  );


  xor
  g241
  (
    n281,
    n215,
    n241,
    n250,
    n252
  );


  xnor
  g242
  (
    n265,
    n154,
    n241,
    n250,
    n156
  );


  or
  g243
  (
    n262,
    n215,
    n253,
    n244,
    n251
  );


  nor
  g244
  (
    n273,
    n243,
    n248,
    n241,
    n254
  );


  or
  g245
  (
    KeyWire_0_16,
    n254,
    n245,
    n216,
    n257
  );


  and
  g246
  (
    n266,
    n247,
    n252,
    n251,
    n249
  );


  nand
  g247
  (
    n287,
    n213,
    n213,
    n246,
    n240
  );


  xnor
  g248
  (
    n275,
    n157,
    n215,
    n256,
    n254
  );


  xnor
  g249
  (
    n279,
    n214,
    n155,
    n239,
    n258
  );


  nor
  g250
  (
    n263,
    n252,
    n258,
    n214,
    n250
  );


  or
  g251
  (
    n277,
    n257,
    n257,
    n242,
    n253
  );


  nand
  g252
  (
    n284,
    n253,
    n245,
    n242,
    n214
  );


  and
  g253
  (
    n261,
    n246,
    n256,
    n255,
    n245
  );


  and
  g254
  (
    n286,
    n239,
    n247,
    n243,
    n212
  );


  xor
  g255
  (
    n268,
    n212,
    n247,
    n240,
    n255
  );


  buf
  g256
  (
    n302,
    n264
  );


  buf
  g257
  (
    n308,
    n263
  );


  buf
  g258
  (
    n301,
    n271
  );


  not
  g259
  (
    n298,
    n277
  );


  not
  g260
  (
    n289,
    n275
  );


  buf
  g261
  (
    n290,
    n276
  );


  not
  g262
  (
    n294,
    n273
  );


  buf
  g263
  (
    n300,
    n274
  );


  not
  g264
  (
    n297,
    n265
  );


  not
  g265
  (
    n309,
    n266
  );


  not
  g266
  (
    n292,
    n261
  );


  not
  g267
  (
    n304,
    n260
  );


  not
  g268
  (
    n296,
    n270
  );


  buf
  g269
  (
    KeyWire_0_29,
    n278
  );


  not
  g270
  (
    n305,
    n276
  );


  buf
  g271
  (
    n306,
    n277
  );


  buf
  g272
  (
    n307,
    n267
  );


  not
  g273
  (
    n295,
    n272
  );


  buf
  g274
  (
    KeyWire_0_15,
    n268
  );


  buf
  g275
  (
    n299,
    n275
  );


  not
  g276
  (
    n310,
    n262
  );


  buf
  g277
  (
    n291,
    n259
  );


  buf
  g278
  (
    n288,
    n278
  );


  buf
  g279
  (
    n311,
    n269
  );


  not
  g280
  (
    KeyWire_0_31,
    n288
  );


  not
  g281
  (
    n325,
    n290
  );


  buf
  g282
  (
    n320,
    n289
  );


  not
  g283
  (
    n326,
    n292
  );


  buf
  g284
  (
    n313,
    n290
  );


  not
  g285
  (
    n321,
    n295
  );


  buf
  g286
  (
    n312,
    n289
  );


  buf
  g287
  (
    n317,
    n288
  );


  not
  g288
  (
    n323,
    n290
  );


  not
  g289
  (
    n316,
    n296
  );


  nor
  g290
  (
    n318,
    n294,
    n293,
    n295
  );


  xnor
  g291
  (
    n322,
    n294,
    n296,
    n292,
    n295
  );


  xnor
  g292
  (
    n324,
    n291,
    n293,
    n288,
    n297
  );


  xnor
  g293
  (
    n315,
    n291,
    n289,
    n296,
    n292
  );


  nor
  g294
  (
    KeyWire_0_0,
    n291,
    n294,
    n297
  );


  not
  g295
  (
    n331,
    n322
  );


  buf
  g296
  (
    KeyWire_0_23,
    n312
  );


  buf
  g297
  (
    n342,
    n316
  );


  buf
  g298
  (
    n338,
    n321
  );


  buf
  g299
  (
    n335,
    n313
  );


  not
  g300
  (
    n343,
    n324
  );


  buf
  g301
  (
    n328,
    n321
  );


  buf
  g302
  (
    n339,
    n318
  );


  buf
  g303
  (
    n337,
    n323
  );


  buf
  g304
  (
    n340,
    n323
  );


  not
  g305
  (
    n344,
    n325
  );


  not
  g306
  (
    n332,
    n325
  );


  not
  g307
  (
    n327,
    n317
  );


  not
  g308
  (
    n336,
    n326
  );


  not
  g309
  (
    n330,
    n314
  );


  buf
  g310
  (
    n329,
    n315
  );


  buf
  g311
  (
    n333,
    n324
  );


  buf
  g312
  (
    n341,
    n320
  );


  buf
  g313
  (
    n334,
    n322
  );


  buf
  g314
  (
    n346,
    n319
  );


  buf
  g315
  (
    n359,
    n346
  );


  buf
  g316
  (
    n362,
    n343
  );


  not
  g317
  (
    n361,
    n93
  );


  buf
  g318
  (
    KeyWire_0_6,
    n95
  );


  not
  g319
  (
    n368,
    n238
  );


  buf
  g320
  (
    n352,
    n100
  );


  buf
  g321
  (
    n353,
    n94
  );


  not
  g322
  (
    n369,
    n96
  );


  buf
  g323
  (
    n351,
    n101
  );


  buf
  g324
  (
    n364,
    n328
  );


  nor
  g325
  (
    n355,
    n342,
    n237
  );


  and
  g326
  (
    n354,
    n336,
    n329,
    n99,
    n327
  );


  nor
  g327
  (
    n366,
    n94,
    n99,
    n339,
    n344
  );


  and
  g328
  (
    n370,
    n331,
    n330,
    n101,
    n237
  );


  xnor
  g329
  (
    n365,
    n96,
    n333,
    n100,
    n101
  );


  xnor
  g330
  (
    n349,
    n345,
    n103,
    n97,
    n343
  );


  nor
  g331
  (
    n367,
    n338,
    n99,
    n92,
    n102
  );


  or
  g332
  (
    n357,
    n332,
    n96,
    n92,
    n97
  );


  and
  g333
  (
    n347,
    n340,
    n91,
    n102,
    n97
  );


  nor
  g334
  (
    n372,
    n236,
    n103,
    n93,
    n238
  );


  or
  g335
  (
    n363,
    n94,
    n335,
    n346,
    n342
  );


  nand
  g336
  (
    n371,
    n344,
    n334,
    n98,
    n95
  );


  nor
  g337
  (
    n360,
    n93,
    n237,
    n103,
    n238
  );


  or
  g338
  (
    n356,
    n98,
    n95,
    n341,
    n102
  );


  nand
  g339
  (
    n350,
    n345,
    n91,
    n337
  );


  and
  g340
  (
    n358,
    n98,
    n92,
    n100,
    n341
  );


  buf
  g341
  (
    n373,
    n301
  );


  not
  g342
  (
    n375,
    n303
  );


  buf
  g343
  (
    n393,
    n299
  );


  buf
  g344
  (
    n418,
    n368
  );


  not
  g345
  (
    n415,
    n302
  );


  not
  g346
  (
    n403,
    n302
  );


  not
  g347
  (
    KeyWire_0_24,
    n104
  );


  buf
  g348
  (
    n376,
    n350
  );


  buf
  g349
  (
    n387,
    n302
  );


  not
  g350
  (
    n402,
    n355
  );


  buf
  g351
  (
    n416,
    n349
  );


  buf
  g352
  (
    n411,
    n218
  );


  buf
  g353
  (
    n392,
    n362
  );


  not
  g354
  (
    n413,
    n367
  );


  buf
  g355
  (
    n412,
    n303
  );


  buf
  g356
  (
    n381,
    n300
  );


  not
  g357
  (
    n408,
    n219
  );


  buf
  g358
  (
    n386,
    n363
  );


  not
  g359
  (
    n390,
    n219
  );


  buf
  g360
  (
    n400,
    n359
  );


  not
  g361
  (
    n420,
    n303
  );


  not
  g362
  (
    n417,
    n358
  );


  buf
  g363
  (
    n394,
    n105
  );


  not
  g364
  (
    KeyWire_0_27,
    n354
  );


  not
  g365
  (
    KeyWire_0_5,
    n368
  );


  buf
  g366
  (
    KeyWire_0_28,
    n298
  );


  not
  g367
  (
    n391,
    n218
  );


  buf
  g368
  (
    n406,
    n356
  );


  not
  g369
  (
    n384,
    n369
  );


  not
  g370
  (
    n401,
    n370
  );


  nand
  g371
  (
    n424,
    n217,
    n351,
    n106
  );


  nor
  g372
  (
    n383,
    n371,
    n347,
    n108
  );


  and
  g373
  (
    n385,
    n217,
    n105,
    n360
  );


  nor
  g374
  (
    n374,
    n219,
    n108,
    n369
  );


  xnor
  g375
  (
    n422,
    n357,
    n352,
    n300
  );


  xnor
  g376
  (
    n419,
    n356,
    n106,
    n347
  );


  nor
  g377
  (
    n379,
    n107,
    n364
  );


  and
  g378
  (
    n410,
    n298,
    n355,
    n371
  );


  nand
  g379
  (
    n397,
    n353,
    n107,
    n108
  );


  or
  g380
  (
    n396,
    n360,
    n300,
    n217
  );


  nor
  g381
  (
    n398,
    n104,
    n354,
    n366
  );


  xor
  g382
  (
    n388,
    n106,
    n365,
    n362
  );


  nand
  g383
  (
    n395,
    n351,
    n104,
    n348
  );


  xnor
  g384
  (
    n409,
    n105,
    n361,
    n218
  );


  nor
  g385
  (
    n423,
    n357,
    n298,
    n109
  );


  nor
  g386
  (
    n399,
    n301,
    n358,
    n367
  );


  and
  g387
  (
    n407,
    n301,
    n361,
    n372
  );


  nand
  g388
  (
    n421,
    n299,
    n107,
    n359
  );


  and
  g389
  (
    n380,
    n370,
    n352,
    n372
  );


  and
  g390
  (
    n377,
    n365,
    n363,
    n366
  );


  nor
  g391
  (
    n404,
    n349,
    n350,
    n299
  );


  xor
  g392
  (
    n405,
    n353,
    n348,
    n109
  );


  buf
  g393
  (
    n468,
    n390
  );


  not
  g394
  (
    n427,
    n413
  );


  buf
  g395
  (
    n443,
    n404
  );


  buf
  g396
  (
    n511,
    n380
  );


  not
  g397
  (
    n448,
    n380
  );


  buf
  g398
  (
    n469,
    n410
  );


  not
  g399
  (
    n487,
    n390
  );


  buf
  g400
  (
    n545,
    n385
  );


  buf
  g401
  (
    n445,
    n401
  );


  buf
  g402
  (
    n562,
    n379
  );


  buf
  g403
  (
    n461,
    n389
  );


  buf
  g404
  (
    n464,
    n391
  );


  not
  g405
  (
    n442,
    n399
  );


  not
  g406
  (
    n564,
    n399
  );


  not
  g407
  (
    n539,
    n393
  );


  not
  g408
  (
    n538,
    n409
  );


  not
  g409
  (
    n555,
    n417
  );


  buf
  g410
  (
    n561,
    n379
  );


  not
  g411
  (
    n536,
    n403
  );


  not
  g412
  (
    n513,
    n408
  );


  not
  g413
  (
    n466,
    n381
  );


  buf
  g414
  (
    n432,
    n415
  );


  not
  g415
  (
    n475,
    n382
  );


  not
  g416
  (
    n566,
    n400
  );


  buf
  g417
  (
    n472,
    n415
  );


  not
  g418
  (
    n494,
    n402
  );


  buf
  g419
  (
    n485,
    n417
  );


  not
  g420
  (
    n527,
    n398
  );


  not
  g421
  (
    n535,
    n407
  );


  not
  g422
  (
    n517,
    n400
  );


  buf
  g423
  (
    n462,
    n397
  );


  buf
  g424
  (
    n565,
    n392
  );


  not
  g425
  (
    n433,
    n413
  );


  not
  g426
  (
    n543,
    n397
  );


  not
  g427
  (
    KeyWire_0_22,
    n406
  );


  not
  g428
  (
    n456,
    n406
  );


  not
  g429
  (
    n471,
    n376
  );


  buf
  g430
  (
    n467,
    n416
  );


  buf
  g431
  (
    n457,
    n404
  );


  buf
  g432
  (
    n495,
    n394
  );


  not
  g433
  (
    n544,
    n378
  );


  buf
  g434
  (
    n516,
    n414
  );


  not
  g435
  (
    n463,
    n409
  );


  not
  g436
  (
    n453,
    n384
  );


  not
  g437
  (
    n506,
    n389
  );


  not
  g438
  (
    n431,
    n393
  );


  buf
  g439
  (
    KeyWire_0_17,
    n396
  );


  not
  g440
  (
    n434,
    n376
  );


  not
  g441
  (
    n512,
    n383
  );


  not
  g442
  (
    n437,
    n402
  );


  not
  g443
  (
    n482,
    n375
  );


  not
  g444
  (
    n502,
    n410
  );


  buf
  g445
  (
    n438,
    n396
  );


  not
  g446
  (
    n473,
    n381
  );


  buf
  g447
  (
    n440,
    n412
  );


  buf
  g448
  (
    n515,
    n373
  );


  buf
  g449
  (
    n501,
    n404
  );


  buf
  g450
  (
    n531,
    n411
  );


  not
  g451
  (
    n558,
    n417
  );


  buf
  g452
  (
    n490,
    n398
  );


  not
  g453
  (
    n533,
    n419
  );


  not
  g454
  (
    n550,
    n377
  );


  buf
  g455
  (
    n508,
    n373
  );


  not
  g456
  (
    n521,
    n405
  );


  not
  g457
  (
    n559,
    n401
  );


  not
  g458
  (
    KeyWire_0_21,
    n382
  );


  buf
  g459
  (
    n476,
    n403
  );


  buf
  g460
  (
    n478,
    n403
  );


  not
  g461
  (
    n548,
    n387
  );


  not
  g462
  (
    n451,
    n384
  );


  buf
  g463
  (
    n509,
    n418
  );


  not
  g464
  (
    n481,
    n391
  );


  buf
  g465
  (
    n557,
    n397
  );


  not
  g466
  (
    n452,
    n411
  );


  not
  g467
  (
    n454,
    n374
  );


  buf
  g468
  (
    n522,
    n378
  );


  buf
  g469
  (
    n524,
    n405
  );


  not
  g470
  (
    n503,
    n416
  );


  buf
  g471
  (
    n491,
    n392
  );


  buf
  g472
  (
    n430,
    n398
  );


  not
  g473
  (
    n534,
    n395
  );


  buf
  g474
  (
    n514,
    n418
  );


  not
  g475
  (
    n529,
    n386
  );


  buf
  g476
  (
    n426,
    n412
  );


  buf
  g477
  (
    n542,
    n419
  );


  buf
  g478
  (
    n553,
    n380
  );


  not
  g479
  (
    n504,
    n413
  );


  buf
  g480
  (
    n450,
    n393
  );


  not
  g481
  (
    n435,
    n420
  );


  not
  g482
  (
    n460,
    n374
  );


  buf
  g483
  (
    n519,
    n375
  );


  not
  g484
  (
    n439,
    n399
  );


  not
  g485
  (
    n477,
    n394
  );


  buf
  g486
  (
    n540,
    n388
  );


  buf
  g487
  (
    n479,
    n412
  );


  not
  g488
  (
    n441,
    n386
  );


  buf
  g489
  (
    n554,
    n389
  );


  not
  g490
  (
    n486,
    n382
  );


  buf
  g491
  (
    n549,
    n383
  );


  buf
  g492
  (
    n458,
    n406
  );


  buf
  g493
  (
    n520,
    n414
  );


  not
  g494
  (
    n560,
    n401
  );


  not
  g495
  (
    n470,
    n390
  );


  not
  g496
  (
    n444,
    n375
  );


  buf
  g497
  (
    KeyWire_0_26,
    n408
  );


  not
  g498
  (
    n541,
    n388
  );


  buf
  g499
  (
    n447,
    n387
  );


  not
  g500
  (
    n551,
    n416
  );


  buf
  g501
  (
    n455,
    n411
  );


  not
  g502
  (
    n489,
    n376
  );


  not
  g503
  (
    n499,
    n407
  );


  buf
  g504
  (
    n429,
    n415
  );


  not
  g505
  (
    n507,
    n419
  );


  buf
  g506
  (
    n525,
    n379
  );


  not
  g507
  (
    n497,
    n384
  );


  buf
  g508
  (
    n484,
    n395
  );


  not
  g509
  (
    n492,
    n378
  );


  buf
  g510
  (
    n459,
    n374
  );


  buf
  g511
  (
    n563,
    n396
  );


  not
  g512
  (
    n537,
    n385
  );


  buf
  g513
  (
    n474,
    n402
  );


  not
  g514
  (
    n552,
    n418
  );


  buf
  g515
  (
    n523,
    n383
  );


  not
  g516
  (
    n500,
    n409
  );


  not
  g517
  (
    n547,
    n377
  );


  not
  g518
  (
    n480,
    n386
  );


  not
  g519
  (
    n532,
    n385
  );


  not
  g520
  (
    n546,
    n407
  );


  buf
  g521
  (
    n526,
    n395
  );


  buf
  g522
  (
    n496,
    n373
  );


  buf
  g523
  (
    n465,
    n408
  );


  not
  g524
  (
    n518,
    n387
  );


  not
  g525
  (
    n528,
    n410
  );


  buf
  g526
  (
    n493,
    n381
  );


  buf
  g527
  (
    n498,
    n391
  );


  buf
  g528
  (
    n488,
    n394
  );


  not
  g529
  (
    n425,
    n377
  );


  not
  g530
  (
    n556,
    n400
  );


  not
  g531
  (
    n446,
    n388
  );


  buf
  g532
  (
    n428,
    n414
  );


  buf
  g533
  (
    n483,
    n392
  );


  buf
  g534
  (
    n510,
    n405
  );


  buf
  g535
  (
    n578,
    n436
  );


  not
  g536
  (
    n568,
    n427
  );


  buf
  g537
  (
    n574,
    n435
  );


  not
  g538
  (
    n576,
    n428
  );


  not
  g539
  (
    n572,
    n438
  );


  not
  g540
  (
    n577,
    n434
  );


  buf
  g541
  (
    n570,
    n432
  );


  not
  g542
  (
    n575,
    n430
  );


  buf
  g543
  (
    n571,
    n437
  );


  nor
  g544
  (
    n580,
    n426,
    n437,
    n429
  );


  nand
  g545
  (
    n573,
    n434,
    n429,
    n433,
    n431
  );


  xnor
  g546
  (
    n579,
    n428,
    n438,
    n430,
    n432
  );


  nor
  g547
  (
    n567,
    n426,
    n427,
    n436,
    n431
  );


  or
  g548
  (
    n569,
    n425,
    n425,
    n433,
    n435
  );


  xor
  g549
  (
    n597,
    n446,
    n443,
    n579
  );


  or
  g550
  (
    n591,
    n578,
    n571,
    n439,
    n569
  );


  nand
  g551
  (
    n594,
    n447,
    n574,
    n567,
    n445
  );


  and
  g552
  (
    n593,
    n568,
    n571,
    n572,
    n569
  );


  xnor
  g553
  (
    n595,
    n578,
    n568,
    n577
  );


  and
  g554
  (
    n598,
    n569,
    n576,
    n570,
    n446
  );


  or
  g555
  (
    n586,
    n567,
    n574,
    n439
  );


  or
  g556
  (
    n584,
    n110,
    n579,
    n567,
    n444
  );


  nor
  g557
  (
    n583,
    n580,
    n578,
    n577,
    n576
  );


  nand
  g558
  (
    n581,
    n579,
    n573,
    n110,
    n440
  );


  or
  g559
  (
    n582,
    n447,
    n575,
    n576
  );


  nor
  g560
  (
    n590,
    n448,
    n572,
    n570,
    n580
  );


  xnor
  g561
  (
    n585,
    n109,
    n579,
    n578,
    n575
  );


  xnor
  g562
  (
    n592,
    n576,
    n442,
    n440,
    n570
  );


  xnor
  g563
  (
    n587,
    n441,
    n442,
    n444,
    n580
  );


  xor
  g564
  (
    n596,
    n575,
    n111,
    n573
  );


  xnor
  g565
  (
    n589,
    n445,
    n580,
    n577
  );


  and
  g566
  (
    n588,
    n572,
    n571,
    n110,
    n441
  );


  buf
  g567
  (
    n602,
    n592
  );


  not
  g568
  (
    n613,
    n587
  );


  not
  g569
  (
    n601,
    n590
  );


  buf
  g570
  (
    n611,
    n596
  );


  not
  g571
  (
    n609,
    n597
  );


  buf
  g572
  (
    n612,
    n585
  );


  not
  g573
  (
    n608,
    n593
  );


  buf
  g574
  (
    n610,
    n584
  );


  not
  g575
  (
    n599,
    n589
  );


  not
  g576
  (
    KeyWire_0_9,
    n588
  );


  not
  g577
  (
    n604,
    n586
  );


  buf
  g578
  (
    n607,
    n591
  );


  not
  g579
  (
    n605,
    n595
  );


  not
  g580
  (
    n603,
    n111
  );


  or
  g581
  (
    n606,
    n594,
    n598
  );


  xor
  g582
  (
    n652,
    n466,
    n498,
    n487
  );


  nand
  g583
  (
    n662,
    n599,
    n483,
    n456,
    n601
  );


  and
  g584
  (
    n638,
    n612,
    n472,
    n606,
    n502
  );


  nand
  g585
  (
    n620,
    n478,
    n492,
    n509,
    n493
  );


  and
  g586
  (
    n621,
    n485,
    n448,
    n606,
    n601
  );


  nor
  g587
  (
    n635,
    n609,
    n495,
    n490,
    n610
  );


  nand
  g588
  (
    n632,
    n458,
    n602,
    n506,
    n607
  );


  nand
  g589
  (
    n616,
    n471,
    n602,
    n603,
    n501
  );


  xor
  g590
  (
    n648,
    n613,
    n497,
    n304,
    n599
  );


  or
  g591
  (
    n642,
    n457,
    n473,
    n496,
    n604
  );


  xor
  g592
  (
    n647,
    n482,
    n456,
    n612,
    n304
  );


  xnor
  g593
  (
    n637,
    n453,
    n499,
    n493,
    n506
  );


  nand
  g594
  (
    n660,
    n304,
    n500,
    n484,
    n476
  );


  nand
  g595
  (
    n619,
    n492,
    n496,
    n477,
    n475
  );


  and
  g596
  (
    n655,
    n611,
    n491,
    n490,
    n487
  );


  or
  g597
  (
    n640,
    n478,
    n472,
    n508,
    n449
  );


  nand
  g598
  (
    n653,
    n305,
    n504,
    n454,
    n505
  );


  nand
  g599
  (
    n624,
    n607,
    n449,
    n450,
    n600
  );


  nor
  g600
  (
    n631,
    n455,
    n603,
    n479,
    n488
  );


  xor
  g601
  (
    n644,
    n494,
    n475,
    n465,
    n605
  );


  or
  g602
  (
    n622,
    n604,
    n502,
    n613,
    n496
  );


  and
  g603
  (
    n649,
    n610,
    n458,
    n509,
    n499
  );


  nor
  g604
  (
    n651,
    n450,
    n468,
    n501,
    n504
  );


  xnor
  g605
  (
    n643,
    n474,
    n451,
    n459,
    n489
  );


  or
  g606
  (
    n656,
    n493,
    n457,
    n507,
    n506
  );


  nand
  g607
  (
    n614,
    n491,
    n503,
    n602,
    n467
  );


  xor
  g608
  (
    n615,
    n611,
    n486,
    n489,
    n607
  );


  nand
  g609
  (
    n636,
    n495,
    n500,
    n507,
    n461
  );


  xnor
  g610
  (
    n623,
    n476,
    n494,
    n468,
    n500
  );


  nor
  g611
  (
    n626,
    n611,
    n505,
    n600,
    n601
  );


  xor
  g612
  (
    n654,
    n471,
    n499,
    n610,
    n606
  );


  and
  g613
  (
    n630,
    n599,
    n613,
    n484,
    n464
  );


  xor
  g614
  (
    n625,
    n609,
    n466,
    n463,
    n477
  );


  and
  g615
  (
    n659,
    n507,
    n480,
    n470,
    n464
  );


  or
  g616
  (
    n645,
    n503,
    n454,
    n467,
    n460
  );


  and
  g617
  (
    n646,
    n608,
    n462,
    n501,
    n612
  );


  nor
  g618
  (
    n641,
    n603,
    n460,
    n605,
    n498
  );


  or
  g619
  (
    n633,
    n459,
    n504,
    n488,
    n495
  );


  xnor
  g620
  (
    n618,
    n481,
    n485,
    n469,
    n608
  );


  and
  g621
  (
    n657,
    n452,
    n481,
    n473,
    n502
  );


  xnor
  g622
  (
    n639,
    n470,
    n489,
    n455,
    n505
  );


  or
  g623
  (
    n658,
    n451,
    n482,
    n483,
    n611
  );


  nand
  g624
  (
    n634,
    n604,
    n508,
    n474,
    n453
  );


  xor
  g625
  (
    n650,
    n605,
    n508,
    n490,
    n612
  );


  nor
  g626
  (
    n617,
    n465,
    n461,
    n463,
    n479
  );


  xnor
  g627
  (
    n627,
    n480,
    n494,
    n497,
    n452
  );


  nand
  g628
  (
    n628,
    n469,
    n609,
    n491,
    n462
  );


  xnor
  g629
  (
    n629,
    n608,
    n497,
    n492,
    n610
  );


  nand
  g630
  (
    n661,
    n486,
    n503,
    n613,
    n600
  );


  or
  g631
  (
    n700,
    n645,
    n531,
    n117,
    n617
  );


  xor
  g632
  (
    n717,
    n539,
    n555,
    n650,
    n111
  );


  or
  g633
  (
    n698,
    n518,
    n662,
    n658,
    n529
  );


  nand
  g634
  (
    n670,
    n625,
    n639,
    n647,
    n517
  );


  or
  g635
  (
    n694,
    n538,
    n546,
    n639,
    n541
  );


  and
  g636
  (
    n709,
    n537,
    n654,
    n633,
    n645
  );


  xor
  g637
  (
    n676,
    n622,
    n531,
    n114,
    n519
  );


  xnor
  g638
  (
    n715,
    n626,
    n513,
    n115,
    n116
  );


  nand
  g639
  (
    KeyWire_0_20,
    n620,
    n648,
    n531,
    n638
  );


  nand
  g640
  (
    n739,
    n545,
    n646,
    n533,
    n523
  );


  nor
  g641
  (
    n663,
    n521,
    n620,
    n510,
    n549
  );


  xnor
  g642
  (
    n678,
    n513,
    n619,
    n541,
    n642
  );


  xnor
  g643
  (
    n691,
    n637,
    n638,
    n520,
    n646
  );


  or
  g644
  (
    n701,
    n556,
    n656,
    n555
  );


  and
  g645
  (
    n683,
    n642,
    n420,
    n651,
    n614
  );


  xnor
  g646
  (
    n696,
    n634,
    n524,
    n512,
    n616
  );


  xor
  g647
  (
    n667,
    n641,
    n525,
    n650,
    n516
  );


  or
  g648
  (
    n737,
    n615,
    n618,
    n113,
    n625
  );


  nor
  g649
  (
    n723,
    n546,
    n621,
    n533,
    n515
  );


  nor
  g650
  (
    n679,
    n661,
    n545,
    n112,
    n641
  );


  or
  g651
  (
    n689,
    n659,
    n550,
    n622,
    n657
  );


  and
  g652
  (
    n680,
    n654,
    n615,
    n634,
    n625
  );


  xnor
  g653
  (
    n684,
    n516,
    n550,
    n545,
    n636
  );


  nor
  g654
  (
    n703,
    n534,
    n420,
    n547,
    n523
  );


  nand
  g655
  (
    n695,
    n629,
    n525,
    n535
  );


  and
  g656
  (
    n736,
    n618,
    n624,
    n650,
    n631
  );


  xor
  g657
  (
    n688,
    n540,
    n643,
    n554,
    n543
  );


  xor
  g658
  (
    n735,
    n624,
    n635,
    n645,
    n513
  );


  xor
  g659
  (
    n732,
    n113,
    n647,
    n619,
    n511
  );


  nor
  g660
  (
    n674,
    n656,
    n644,
    n623,
    n528
  );


  nor
  g661
  (
    KeyWire_0_12,
    n522,
    n547,
    n516,
    n633
  );


  nor
  g662
  (
    n675,
    n116,
    n552,
    n640,
    n626
  );


  or
  g663
  (
    n666,
    n640,
    n114,
    n536,
    n526
  );


  nor
  g664
  (
    n693,
    n653,
    n511,
    n518,
    n548
  );


  nor
  g665
  (
    n710,
    n529,
    n655,
    n617,
    n648
  );


  nor
  g666
  (
    n681,
    n551,
    n651,
    n547,
    n660
  );


  xor
  g667
  (
    n721,
    n649,
    n542,
    n662
  );


  nor
  g668
  (
    n692,
    n636,
    n662,
    n525,
    n551
  );


  nand
  g669
  (
    n685,
    n649,
    n517,
    n514,
    n526
  );


  xnor
  g670
  (
    n707,
    n652,
    n115,
    n616,
    n628
  );


  nand
  g671
  (
    n724,
    n661,
    n628,
    n634,
    n631
  );


  and
  g672
  (
    n690,
    n522,
    n655,
    n627,
    n537
  );


  xnor
  g673
  (
    n708,
    n540,
    n532,
    n112,
    n549
  );


  xor
  g674
  (
    n699,
    n517,
    n658,
    n524,
    n530
  );


  and
  g675
  (
    n719,
    n648,
    n640,
    n512,
    n553
  );


  and
  g676
  (
    n671,
    n550,
    n637,
    n642,
    n655
  );


  xor
  g677
  (
    n726,
    n643,
    n512,
    n631,
    n515
  );


  and
  g678
  (
    n668,
    n532,
    n552,
    n548,
    n649
  );


  xnor
  g679
  (
    n714,
    n526,
    n115,
    n623,
    n549
  );


  or
  g680
  (
    n665,
    n538,
    n534,
    n639,
    n515
  );


  nor
  g681
  (
    n702,
    n537,
    n519,
    n615,
    n632
  );


  nand
  g682
  (
    n704,
    n657,
    n544,
    n541,
    n546
  );


  nor
  g683
  (
    n677,
    n646,
    n659,
    n621,
    n653
  );


  nor
  g684
  (
    n731,
    n527,
    n536,
    n618,
    n651
  );


  nand
  g685
  (
    n728,
    n520,
    n556,
    n533,
    n626
  );


  xor
  g686
  (
    n682,
    n629,
    n654,
    n658,
    n511
  );


  or
  g687
  (
    n738,
    n628,
    n622,
    n112,
    n530
  );


  and
  g688
  (
    n725,
    n551,
    n629,
    n630,
    n616
  );


  xnor
  g689
  (
    n673,
    n114,
    n528,
    n553,
    n635
  );


  nor
  g690
  (
    n686,
    n633,
    n535,
    n552,
    n527
  );


  xor
  g691
  (
    n734,
    n621,
    n544,
    n528,
    n521
  );


  nor
  g692
  (
    n669,
    n614,
    n620,
    n518,
    n660
  );


  nor
  g693
  (
    n687,
    n532,
    n540,
    n659,
    n638
  );


  nor
  g694
  (
    n697,
    n660,
    n644,
    n627,
    n519
  );


  xor
  g695
  (
    n727,
    n636,
    n637,
    n530,
    n553
  );


  nor
  g696
  (
    n711,
    n539,
    n521,
    n623,
    n617
  );


  xor
  g697
  (
    n733,
    n632,
    n635,
    n661,
    n652
  );


  and
  g698
  (
    n722,
    n643,
    n630,
    n527
  );


  nor
  g699
  (
    n706,
    n544,
    n652,
    n641,
    n644
  );


  and
  g700
  (
    n705,
    n627,
    n534,
    n556,
    n523
  );


  xnor
  g701
  (
    n720,
    n619,
    n624,
    n522,
    n554
  );


  nor
  g702
  (
    n730,
    n520,
    n539,
    n647,
    n632
  );


  xor
  g703
  (
    n664,
    n554,
    n509,
    n548,
    n538
  );


  and
  g704
  (
    n718,
    n510,
    n542,
    n555,
    n113
  );


  xor
  g705
  (
    n713,
    n657,
    n543,
    n614,
    n653
  );


  or
  g706
  (
    n716,
    n529,
    n543,
    n116,
    n536
  );


  nand
  g707
  (
    n712,
    n524,
    n514,
    n510
  );


  or
  g708
  (
    n744,
    n683,
    n676,
    n665,
    n685
  );


  nand
  g709
  (
    n743,
    n672,
    n673,
    n670,
    n666
  );


  or
  g710
  (
    n741,
    n667,
    n674,
    n664,
    n677
  );


  and
  g711
  (
    n742,
    n668,
    n691,
    n679,
    n684
  );


  nor
  g712
  (
    KeyWire_0_1,
    n678,
    n688,
    n681,
    n689
  );


  nand
  g713
  (
    n747,
    n663,
    n686,
    n671,
    n692
  );


  xor
  g714
  (
    n746,
    n669,
    n680,
    n682,
    n690
  );


  xnor
  g715
  (
    n740,
    n694,
    n675,
    n687,
    n693
  );


  buf
  g716
  (
    n758,
    n743
  );


  buf
  g717
  (
    n750,
    n743
  );


  not
  g718
  (
    n748,
    n741
  );


  not
  g719
  (
    n751,
    n746
  );


  not
  g720
  (
    n757,
    n746
  );


  not
  g721
  (
    n753,
    n742
  );


  not
  g722
  (
    n766,
    n741
  );


  buf
  g723
  (
    n759,
    n740
  );


  buf
  g724
  (
    n755,
    n742
  );


  not
  g725
  (
    n760,
    n743
  );


  not
  g726
  (
    n765,
    n741
  );


  not
  g727
  (
    n764,
    n744
  );


  not
  g728
  (
    n752,
    n159
  );


  buf
  g729
  (
    n754,
    n745
  );


  and
  g730
  (
    n768,
    n745,
    n118
  );


  xnor
  g731
  (
    n767,
    n119,
    n743,
    n118,
    n747
  );


  xnor
  g732
  (
    n756,
    n695,
    n696,
    n747,
    n746
  );


  xnor
  g733
  (
    n761,
    n117,
    n744,
    n747,
    n742
  );


  xor
  g734
  (
    KeyWire_0_7,
    n744,
    n747,
    n746,
    n119
  );


  nor
  g735
  (
    n749,
    n745,
    n158,
    n740,
    n117
  );


  or
  g736
  (
    n769,
    n744,
    n742,
    n741,
    n119
  );


  nand
  g737
  (
    n762,
    n745,
    n740,
    n697,
    n118
  );


  buf
  g738
  (
    n790,
    n768
  );


  not
  g739
  (
    KeyWire_0_19,
    n769
  );


  buf
  g740
  (
    n774,
    n285
  );


  buf
  g741
  (
    n788,
    n560
  );


  buf
  g742
  (
    n784,
    n761
  );


  buf
  g743
  (
    n771,
    n759
  );


  and
  g744
  (
    n792,
    n284,
    n120,
    n559,
    n749
  );


  xnor
  g745
  (
    n782,
    n758,
    n120,
    n422,
    n757
  );


  and
  g746
  (
    n779,
    n765,
    n283,
    n120,
    n423
  );


  and
  g747
  (
    n791,
    n759,
    n422,
    n760
  );


  xnor
  g748
  (
    n776,
    n754,
    n557,
    n763,
    n285
  );


  nand
  g749
  (
    n786,
    n558,
    n766,
    n762
  );


  or
  g750
  (
    n777,
    n750,
    n559,
    n560,
    n765
  );


  xnor
  g751
  (
    n787,
    n557,
    n422,
    n558,
    n282
  );


  nand
  g752
  (
    n775,
    n762,
    n286,
    n748,
    n421
  );


  xor
  g753
  (
    n770,
    n283,
    n764,
    n121,
    n768
  );


  xor
  g754
  (
    n783,
    n764,
    n761,
    n763,
    n561
  );


  xnor
  g755
  (
    n780,
    n769,
    n280,
    n281,
    n279
  );


  and
  g756
  (
    n773,
    n755,
    n557,
    n558,
    n286
  );


  nor
  g757
  (
    n772,
    n752,
    n281,
    n756,
    n767
  );


  nand
  g758
  (
    n789,
    n280,
    n282,
    n305,
    n421
  );


  nor
  g759
  (
    n781,
    n767,
    n279,
    n284,
    n560
  );


  nor
  g760
  (
    n778,
    n753,
    n751,
    n421,
    n559
  );


  buf
  g761
  (
    n799,
    n770
  );


  buf
  g762
  (
    n802,
    n779
  );


  buf
  g763
  (
    n797,
    n776
  );


  buf
  g764
  (
    n798,
    n777
  );


  not
  g765
  (
    n800,
    n774
  );


  buf
  g766
  (
    n795,
    n775
  );


  buf
  g767
  (
    n794,
    n773
  );


  buf
  g768
  (
    n793,
    n772
  );


  not
  g769
  (
    n796,
    n778
  );


  buf
  g770
  (
    n801,
    n771
  );


  nor
  g771
  (
    n806,
    n793,
    n712,
    n160,
    n306
  );


  xnor
  g772
  (
    n818,
    n729,
    n800,
    n715,
    n727
  );


  or
  g773
  (
    n821,
    n307,
    n792,
    n121,
    n802
  );


  xor
  g774
  (
    n809,
    n795,
    n170,
    n736,
    n229
  );


  and
  g775
  (
    n824,
    n561,
    n121,
    n308,
    n725
  );


  or
  g776
  (
    n822,
    n166,
    n788,
    n800,
    n306
  );


  or
  g777
  (
    n810,
    n739,
    n796,
    n167,
    n562
  );


  nor
  g778
  (
    n815,
    n798,
    n782,
    n307,
    n733
  );


  and
  g779
  (
    n805,
    n307,
    n801,
    n797
  );


  and
  g780
  (
    n811,
    n171,
    n711,
    n699,
    n722
  );


  nor
  g781
  (
    KeyWire_0_4,
    n306,
    n787,
    n789,
    n802
  );


  xnor
  g782
  (
    n820,
    n793,
    n717,
    n703,
    n563
  );


  or
  g783
  (
    n827,
    n709,
    n802,
    n737,
    n162
  );


  nor
  g784
  (
    n819,
    n735,
    n308,
    n704,
    n706
  );


  xor
  g785
  (
    n828,
    n718,
    n783,
    n786,
    n796
  );


  nor
  g786
  (
    n817,
    n172,
    n720,
    n702,
    n705
  );


  or
  g787
  (
    n804,
    n563,
    n710,
    n780,
    n790
  );


  or
  g788
  (
    n832,
    n561,
    n799,
    n796,
    n173
  );


  xnor
  g789
  (
    n813,
    n714,
    n700,
    n164,
    n728
  );


  nand
  g790
  (
    n829,
    n784,
    n721,
    n708,
    n799
  );


  nand
  g791
  (
    n830,
    n781,
    n795,
    n169,
    n732
  );


  or
  g792
  (
    n807,
    n161,
    n793,
    n798,
    n785
  );


  and
  g793
  (
    n816,
    n730,
    n724,
    n738,
    n726
  );


  and
  g794
  (
    n808,
    n562,
    n168,
    n163,
    n698
  );


  xor
  g795
  (
    n825,
    n308,
    n701,
    n562,
    n723
  );


  nand
  g796
  (
    n823,
    n794,
    n563,
    n801,
    n305
  );


  nor
  g797
  (
    n814,
    n800,
    n165,
    n731,
    n713
  );


  nand
  g798
  (
    n831,
    n719,
    n716,
    n795,
    n794
  );


  or
  g799
  (
    n803,
    n707,
    n797,
    n794,
    n734
  );


  and
  g800
  (
    n826,
    n791,
    n799,
    n798,
    n797
  );


  not
  g801
  (
    n834,
    n804
  );


  not
  g802
  (
    KeyWire_0_11,
    n803
  );


  and
  g803
  (
    n837,
    n807,
    n812,
    n806,
    n805
  );


  or
  g804
  (
    n836,
    n808,
    n809,
    n810,
    n813
  );


  xnor
  g805
  (
    n835,
    n811,
    n833,
    n834
  );


  not
  g806
  (
    KeyWire_0_2,
    n836
  );


  nand
  g807
  (
    n842,
    n122,
    n836,
    n837
  );


  or
  g808
  (
    n841,
    n424,
    n564,
    n836,
    n837
  );


  xor
  g809
  (
    n839,
    n835,
    n564,
    n814
  );


  or
  g810
  (
    n838,
    n815,
    n835,
    n565,
    n423
  );


  xnor
  g811
  (
    n843,
    n835,
    n423,
    n837,
    n816
  );


  nand
  g812
  (
    n844,
    n122,
    n839,
    n819,
    n817
  );


  and
  g813
  (
    n846,
    n818,
    n841,
    n824,
    n565
  );


  and
  g814
  (
    n845,
    n843,
    n820,
    n821,
    n122
  );


  and
  g815
  (
    n847,
    n822,
    n823,
    n840,
    n842
  );


  or
  g816
  (
    n849,
    n825,
    n847
  );


  xor
  g817
  (
    n848,
    n845,
    n826,
    n123,
    n828
  );


  and
  g818
  (
    n850,
    n846,
    n123,
    n827,
    n844
  );


  buf
  g819
  (
    n851,
    n829
  );


  or
  g820
  (
    n852,
    n848,
    n849,
    n124,
    n123
  );


  or
  g821
  (
    n853,
    n852,
    n309
  );


  and
  g822
  (
    n855,
    n853,
    n124,
    n424
  );


  or
  g823
  (
    n854,
    n853,
    n287,
    n124
  );


  nand
  g824
  (
    n856,
    n855,
    n310
  );


  xnor
  g825
  (
    n858,
    n856,
    n326,
    n311
  );


  xor
  g826
  (
    n857,
    n856,
    n311
  );


  buf
  g827
  (
    n859,
    n850
  );


  buf
  g828
  (
    n860,
    n858
  );


  or
  g829
  (
    n861,
    n858,
    n857
  );


  and
  g830
  (
    n862,
    n566,
    n566,
    n861,
    n565
  );


  buf
  g831
  (
    n863,
    n862
  );


  and
  g832
  (
    n864,
    n830,
    n862,
    n831
  );


  xor
  g833
  (
    n865,
    n832,
    n566,
    n864,
    n863
  );


  xnor
  KeyGate_0_0
  (
    n314,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n745,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n840,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n61,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n812,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n382,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n348,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n763,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n245,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n600,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n149,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n833,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n729,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n178,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n36,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n303,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n271,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n449,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n92,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n785,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n672,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n505,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n530,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n345,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n389,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n215,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n436,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n414,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n378,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n293,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n179,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n319,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


