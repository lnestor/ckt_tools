

module Stat_1000_107
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n988,
  n1010,
  n1012,
  n990,
  n986,
  n1000,
  n997,
  n991,
  n1013,
  n1016,
  n1002,
  n993,
  n1001,
  n989,
  n992,
  n985,
  n1015,
  n1005,
  n1026,
  n1022,
  n1023,
  n1021,
  n1025,
  n1030,
  n1031,
  n1020,
  n1032,
  n1019,
  n1024,
  n1029,
  n1027,
  n1028,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n988;
  output n1010;
  output n1012;
  output n990;
  output n986;
  output n1000;
  output n997;
  output n991;
  output n1013;
  output n1016;
  output n1002;
  output n993;
  output n1001;
  output n989;
  output n992;
  output n985;
  output n1015;
  output n1005;
  output n1026;
  output n1022;
  output n1023;
  output n1021;
  output n1025;
  output n1030;
  output n1031;
  output n1020;
  output n1032;
  output n1019;
  output n1024;
  output n1029;
  output n1027;
  output n1028;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n987;
  wire n994;
  wire n995;
  wire n996;
  wire n998;
  wire n999;
  wire n1003;
  wire n1004;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1011;
  wire n1014;
  wire n1017;
  wire n1018;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n107,
    n6
  );


  not
  g1
  (
    n43,
    n22
  );


  buf
  g2
  (
    n44,
    n19
  );


  not
  g3
  (
    n83,
    n6
  );


  buf
  g4
  (
    n102,
    n21
  );


  buf
  g5
  (
    n110,
    n11
  );


  buf
  g6
  (
    n69,
    n16
  );


  not
  g7
  (
    n95,
    n5
  );


  not
  g8
  (
    n51,
    n16
  );


  not
  g9
  (
    n97,
    n7
  );


  not
  g10
  (
    n81,
    n12
  );


  buf
  g11
  (
    n74,
    n5
  );


  buf
  g12
  (
    n70,
    n3
  );


  buf
  g13
  (
    n36,
    n17
  );


  buf
  g14
  (
    n72,
    n4
  );


  buf
  g15
  (
    n80,
    n20
  );


  not
  g16
  (
    n67,
    n3
  );


  not
  g17
  (
    n94,
    n17
  );


  not
  g18
  (
    n50,
    n17
  );


  buf
  g19
  (
    n86,
    n13
  );


  buf
  g20
  (
    n47,
    n9
  );


  buf
  g21
  (
    n82,
    n7
  );


  buf
  g22
  (
    n106,
    n8
  );


  buf
  g23
  (
    n90,
    n20
  );


  not
  g24
  (
    n104,
    n9
  );


  buf
  g25
  (
    n37,
    n5
  );


  buf
  g26
  (
    n103,
    n18
  );


  not
  g27
  (
    n59,
    n16
  );


  buf
  g28
  (
    n76,
    n7
  );


  buf
  g29
  (
    n91,
    n13
  );


  buf
  g30
  (
    n66,
    n19
  );


  not
  g31
  (
    n46,
    n14
  );


  buf
  g32
  (
    n105,
    n4
  );


  buf
  g33
  (
    n96,
    n14
  );


  buf
  g34
  (
    n39,
    n15
  );


  not
  g35
  (
    n57,
    n14
  );


  not
  g36
  (
    n49,
    n19
  );


  not
  g37
  (
    n100,
    n18
  );


  buf
  g38
  (
    n101,
    n14
  );


  not
  g39
  (
    n71,
    n21
  );


  not
  g40
  (
    n40,
    n20
  );


  buf
  g41
  (
    n93,
    n7
  );


  not
  g42
  (
    n75,
    n12
  );


  not
  g43
  (
    n62,
    n17
  );


  buf
  g44
  (
    n79,
    n10
  );


  not
  g45
  (
    n33,
    n1
  );


  not
  g46
  (
    n108,
    n9
  );


  not
  g47
  (
    n73,
    n11
  );


  not
  g48
  (
    n68,
    n10
  );


  not
  g49
  (
    KeyWire_0_6,
    n3
  );


  not
  g50
  (
    n53,
    n18
  );


  buf
  g51
  (
    n38,
    n8
  );


  buf
  g52
  (
    n88,
    n10
  );


  buf
  g53
  (
    n52,
    n15
  );


  buf
  g54
  (
    n35,
    n6
  );


  not
  g55
  (
    n99,
    n21
  );


  buf
  g56
  (
    n55,
    n13
  );


  buf
  g57
  (
    KeyWire_0_15,
    n18
  );


  not
  g58
  (
    n85,
    n19
  );


  not
  g59
  (
    n109,
    n11
  );


  not
  g60
  (
    n61,
    n21
  );


  not
  g61
  (
    n87,
    n3
  );


  buf
  g62
  (
    n60,
    n4
  );


  not
  g63
  (
    n65,
    n11
  );


  not
  g64
  (
    n54,
    n10
  );


  not
  g65
  (
    n41,
    n6
  );


  buf
  g66
  (
    n89,
    n22
  );


  buf
  g67
  (
    n56,
    n15
  );


  not
  g68
  (
    n112,
    n5
  );


  not
  g69
  (
    n45,
    n13
  );


  not
  g70
  (
    n92,
    n4
  );


  buf
  g71
  (
    n111,
    n15
  );


  not
  g72
  (
    n77,
    n16
  );


  not
  g73
  (
    n98,
    n20
  );


  buf
  g74
  (
    n58,
    n2
  );


  not
  g75
  (
    n64,
    n8
  );


  buf
  g76
  (
    n63,
    n9
  );


  not
  g77
  (
    n42,
    n12
  );


  buf
  g78
  (
    n34,
    n12
  );


  buf
  g79
  (
    n48,
    n8
  );


  not
  g80
  (
    n228,
    n60
  );


  buf
  g81
  (
    n254,
    n60
  );


  buf
  g82
  (
    n159,
    n58
  );


  not
  g83
  (
    n160,
    n45
  );


  not
  g84
  (
    n267,
    n41
  );


  not
  g85
  (
    n259,
    n67
  );


  not
  g86
  (
    n165,
    n55
  );


  buf
  g87
  (
    n256,
    n66
  );


  buf
  g88
  (
    KeyWire_0_14,
    n38
  );


  not
  g89
  (
    n276,
    n40
  );


  not
  g90
  (
    n154,
    n34
  );


  buf
  g91
  (
    n173,
    n47
  );


  not
  g92
  (
    n118,
    n46
  );


  not
  g93
  (
    n146,
    n64
  );


  buf
  g94
  (
    n137,
    n64
  );


  not
  g95
  (
    n216,
    n73
  );


  buf
  g96
  (
    n136,
    n42
  );


  buf
  g97
  (
    n208,
    n48
  );


  not
  g98
  (
    n127,
    n42
  );


  not
  g99
  (
    n266,
    n54
  );


  not
  g100
  (
    n141,
    n48
  );


  not
  g101
  (
    n144,
    n60
  );


  buf
  g102
  (
    n152,
    n51
  );


  not
  g103
  (
    n130,
    n55
  );


  buf
  g104
  (
    n156,
    n73
  );


  not
  g105
  (
    n148,
    n43
  );


  buf
  g106
  (
    n178,
    n43
  );


  buf
  g107
  (
    n187,
    n71
  );


  not
  g108
  (
    n197,
    n39
  );


  buf
  g109
  (
    n205,
    n47
  );


  not
  g110
  (
    n221,
    n43
  );


  buf
  g111
  (
    n206,
    n40
  );


  buf
  g112
  (
    n237,
    n63
  );


  buf
  g113
  (
    n211,
    n37
  );


  buf
  g114
  (
    n196,
    n67
  );


  not
  g115
  (
    n224,
    n42
  );


  not
  g116
  (
    n210,
    n53
  );


  not
  g117
  (
    n193,
    n38
  );


  buf
  g118
  (
    n180,
    n70
  );


  buf
  g119
  (
    n183,
    n65
  );


  not
  g120
  (
    n195,
    n62
  );


  buf
  g121
  (
    n273,
    n36
  );


  buf
  g122
  (
    n149,
    n57
  );


  buf
  g123
  (
    n263,
    n46
  );


  not
  g124
  (
    n181,
    n52
  );


  buf
  g125
  (
    n203,
    n49
  );


  buf
  g126
  (
    n269,
    n50
  );


  not
  g127
  (
    n214,
    n37
  );


  not
  g128
  (
    n200,
    n63
  );


  not
  g129
  (
    n257,
    n35
  );


  not
  g130
  (
    n172,
    n44
  );


  buf
  g131
  (
    n161,
    n65
  );


  not
  g132
  (
    n151,
    n48
  );


  not
  g133
  (
    n139,
    n57
  );


  buf
  g134
  (
    KeyWire_0_10,
    n33
  );


  buf
  g135
  (
    n143,
    n61
  );


  not
  g136
  (
    n184,
    n51
  );


  not
  g137
  (
    n252,
    n46
  );


  not
  g138
  (
    n247,
    n50
  );


  buf
  g139
  (
    n125,
    n49
  );


  not
  g140
  (
    KeyWire_0_18,
    n68
  );


  buf
  g141
  (
    n215,
    n34
  );


  not
  g142
  (
    n231,
    n36
  );


  buf
  g143
  (
    n190,
    n73
  );


  not
  g144
  (
    n167,
    n56
  );


  buf
  g145
  (
    n201,
    n70
  );


  not
  g146
  (
    n171,
    n56
  );


  buf
  g147
  (
    n240,
    n35
  );


  not
  g148
  (
    n245,
    n66
  );


  not
  g149
  (
    n189,
    n62
  );


  buf
  g150
  (
    n272,
    n37
  );


  buf
  g151
  (
    KeyWire_0_13,
    n54
  );


  not
  g152
  (
    n233,
    n33
  );


  buf
  g153
  (
    n209,
    n36
  );


  buf
  g154
  (
    n163,
    n45
  );


  not
  g155
  (
    n198,
    n43
  );


  buf
  g156
  (
    n229,
    n56
  );


  not
  g157
  (
    n249,
    n48
  );


  not
  g158
  (
    n170,
    n72
  );


  not
  g159
  (
    n115,
    n33
  );


  buf
  g160
  (
    n232,
    n49
  );


  buf
  g161
  (
    n212,
    n47
  );


  buf
  g162
  (
    n114,
    n67
  );


  buf
  g163
  (
    n243,
    n58
  );


  buf
  g164
  (
    n227,
    n70
  );


  buf
  g165
  (
    n133,
    n62
  );


  buf
  g166
  (
    n220,
    n68
  );


  buf
  g167
  (
    n138,
    n42
  );


  buf
  g168
  (
    n120,
    n46
  );


  not
  g169
  (
    n261,
    n57
  );


  buf
  g170
  (
    n140,
    n64
  );


  not
  g171
  (
    n244,
    n49
  );


  not
  g172
  (
    n202,
    n65
  );


  not
  g173
  (
    n119,
    n39
  );


  buf
  g174
  (
    n204,
    n53
  );


  buf
  g175
  (
    n135,
    n69
  );


  not
  g176
  (
    n157,
    n39
  );


  not
  g177
  (
    n177,
    n67
  );


  not
  g178
  (
    n168,
    n57
  );


  buf
  g179
  (
    n121,
    n71
  );


  buf
  g180
  (
    n213,
    n44
  );


  buf
  g181
  (
    n124,
    n39
  );


  buf
  g182
  (
    KeyWire_0_19,
    n68
  );


  not
  g183
  (
    n142,
    n69
  );


  not
  g184
  (
    n162,
    n50
  );


  buf
  g185
  (
    n199,
    n69
  );


  not
  g186
  (
    n248,
    n35
  );


  buf
  g187
  (
    n271,
    n40
  );


  buf
  g188
  (
    n147,
    n65
  );


  buf
  g189
  (
    n113,
    n73
  );


  not
  g190
  (
    n166,
    n51
  );


  buf
  g191
  (
    n264,
    n35
  );


  not
  g192
  (
    n238,
    n34
  );


  not
  g193
  (
    KeyWire_0_9,
    n37
  );


  not
  g194
  (
    n275,
    n70
  );


  not
  g195
  (
    n175,
    n59
  );


  not
  g196
  (
    n242,
    n55
  );


  buf
  g197
  (
    n217,
    n44
  );


  not
  g198
  (
    n255,
    n36
  );


  buf
  g199
  (
    n174,
    n72
  );


  not
  g200
  (
    n191,
    n41
  );


  not
  g201
  (
    n251,
    n34
  );


  not
  g202
  (
    KeyWire_0_29,
    n71
  );


  buf
  g203
  (
    n236,
    n58
  );


  buf
  g204
  (
    n218,
    n58
  );


  not
  g205
  (
    n164,
    n38
  );


  buf
  g206
  (
    n122,
    n38
  );


  not
  g207
  (
    n188,
    n64
  );


  buf
  g208
  (
    n239,
    n52
  );


  buf
  g209
  (
    n126,
    n33
  );


  buf
  g210
  (
    n185,
    n59
  );


  buf
  g211
  (
    n222,
    n63
  );


  not
  g212
  (
    n123,
    n63
  );


  buf
  g213
  (
    n145,
    n45
  );


  buf
  g214
  (
    n182,
    n40
  );


  not
  g215
  (
    n234,
    n51
  );


  not
  g216
  (
    n223,
    n45
  );


  buf
  g217
  (
    n274,
    n61
  );


  buf
  g218
  (
    n235,
    n56
  );


  not
  g219
  (
    n117,
    n69
  );


  not
  g220
  (
    n131,
    n41
  );


  not
  g221
  (
    n158,
    n53
  );


  not
  g222
  (
    n176,
    n71
  );


  not
  g223
  (
    n241,
    n47
  );


  buf
  g224
  (
    n153,
    n54
  );


  not
  g225
  (
    n129,
    n50
  );


  not
  g226
  (
    n132,
    n55
  );


  not
  g227
  (
    n262,
    n41
  );


  not
  g228
  (
    n207,
    n62
  );


  buf
  g229
  (
    KeyWire_0_7,
    n59
  );


  buf
  g230
  (
    n194,
    n72
  );


  not
  g231
  (
    n116,
    n68
  );


  not
  g232
  (
    n226,
    n72
  );


  not
  g233
  (
    n268,
    n66
  );


  buf
  g234
  (
    n179,
    n60
  );


  buf
  g235
  (
    n134,
    n61
  );


  buf
  g236
  (
    n270,
    n52
  );


  buf
  g237
  (
    n150,
    n61
  );


  buf
  g238
  (
    n230,
    n44
  );


  buf
  g239
  (
    n250,
    n52
  );


  buf
  g240
  (
    n128,
    n66
  );


  not
  g241
  (
    n253,
    n54
  );


  not
  g242
  (
    n246,
    n59
  );


  buf
  g243
  (
    n265,
    n53
  );


  not
  g244
  (
    n291,
    n122
  );


  buf
  g245
  (
    n339,
    n75
  );


  buf
  g246
  (
    n299,
    n117
  );


  not
  g247
  (
    n293,
    n114
  );


  buf
  g248
  (
    n323,
    n127
  );


  buf
  g249
  (
    n318,
    n113
  );


  not
  g250
  (
    n335,
    n118
  );


  not
  g251
  (
    n305,
    n75
  );


  buf
  g252
  (
    n342,
    n127
  );


  not
  g253
  (
    n289,
    n113
  );


  buf
  g254
  (
    n295,
    n120
  );


  not
  g255
  (
    n325,
    n122
  );


  not
  g256
  (
    n333,
    n122
  );


  buf
  g257
  (
    n313,
    n116
  );


  buf
  g258
  (
    n279,
    n74
  );


  not
  g259
  (
    n334,
    n125
  );


  buf
  g260
  (
    n294,
    n128
  );


  not
  g261
  (
    n329,
    n74
  );


  buf
  g262
  (
    n297,
    n116
  );


  buf
  g263
  (
    n328,
    n120
  );


  not
  g264
  (
    n282,
    n117
  );


  buf
  g265
  (
    n277,
    n115
  );


  not
  g266
  (
    n302,
    n123
  );


  buf
  g267
  (
    n324,
    n115
  );


  buf
  g268
  (
    n326,
    n119
  );


  not
  g269
  (
    n341,
    n127
  );


  buf
  g270
  (
    n306,
    n121
  );


  buf
  g271
  (
    n321,
    n120
  );


  not
  g272
  (
    n280,
    n123
  );


  not
  g273
  (
    n301,
    n123
  );


  not
  g274
  (
    n310,
    n74
  );


  not
  g275
  (
    n343,
    n120
  );


  not
  g276
  (
    n303,
    n123
  );


  buf
  g277
  (
    n330,
    n114
  );


  not
  g278
  (
    n332,
    n129
  );


  buf
  g279
  (
    n315,
    n126
  );


  buf
  g280
  (
    n311,
    n129
  );


  not
  g281
  (
    n320,
    n128
  );


  not
  g282
  (
    n286,
    n126
  );


  not
  g283
  (
    n307,
    n113
  );


  not
  g284
  (
    n340,
    n118
  );


  buf
  g285
  (
    n312,
    n121
  );


  buf
  g286
  (
    n287,
    n118
  );


  not
  g287
  (
    n316,
    n125
  );


  buf
  g288
  (
    n319,
    n115
  );


  not
  g289
  (
    n331,
    n117
  );


  not
  g290
  (
    n308,
    n121
  );


  not
  g291
  (
    n296,
    n129
  );


  not
  g292
  (
    KeyWire_0_24,
    n125
  );


  not
  g293
  (
    n284,
    n116
  );


  not
  g294
  (
    n309,
    n128
  );


  not
  g295
  (
    n278,
    n125
  );


  buf
  g296
  (
    n314,
    n122
  );


  buf
  g297
  (
    n283,
    n113
  );


  buf
  g298
  (
    n298,
    n127
  );


  not
  g299
  (
    n300,
    n126
  );


  buf
  g300
  (
    n281,
    n117
  );


  buf
  g301
  (
    n285,
    n74
  );


  buf
  g302
  (
    n304,
    n124
  );


  not
  g303
  (
    n336,
    n118
  );


  buf
  g304
  (
    n327,
    n115
  );


  not
  g305
  (
    n292,
    n121
  );


  not
  g306
  (
    n288,
    n116
  );


  not
  g307
  (
    n290,
    n119
  );


  buf
  g308
  (
    n338,
    n124
  );


  xor
  g309
  (
    n317,
    n75,
    n119,
    n114,
    n128
  );


  xor
  g310
  (
    n322,
    n119,
    n126,
    n114,
    n124
  );


  xor
  g311
  (
    n437,
    n149,
    n331,
    n181,
    n283
  );


  nand
  g312
  (
    n508,
    n248,
    n29,
    n172
  );


  and
  g313
  (
    n565,
    n80,
    n309,
    n204,
    n197
  );


  or
  g314
  (
    n512,
    n312,
    n208,
    n286,
    n254
  );


  xor
  g315
  (
    n539,
    n314,
    n131,
    n259,
    n166
  );


  and
  g316
  (
    n488,
    n242,
    n159,
    n165,
    n256
  );


  nand
  g317
  (
    n414,
    n289,
    n224,
    n247,
    n202
  );


  nand
  g318
  (
    n453,
    n294,
    n270,
    n224,
    n217
  );


  xnor
  g319
  (
    n397,
    n224,
    n267,
    n277,
    n148
  );


  nand
  g320
  (
    KeyWire_0_4,
    n176,
    n181,
    n255,
    n285
  );


  or
  g321
  (
    n558,
    n305,
    n26,
    n273,
    n248
  );


  xor
  g322
  (
    n441,
    n192,
    n253,
    n210,
    n136
  );


  xor
  g323
  (
    n416,
    n24,
    n192,
    n290,
    n249
  );


  nand
  g324
  (
    n349,
    n311,
    n141,
    n282,
    n330
  );


  nand
  g325
  (
    n454,
    n299,
    n322,
    n265,
    n314
  );


  xnor
  g326
  (
    n474,
    n326,
    n299,
    n286,
    n239
  );


  nand
  g327
  (
    n363,
    n151,
    n250,
    n305,
    n82
  );


  and
  g328
  (
    n447,
    n318,
    n30,
    n197,
    n23
  );


  nor
  g329
  (
    n464,
    n149,
    n164,
    n313,
    n258
  );


  xor
  g330
  (
    n419,
    n311,
    n199,
    n171,
    n27
  );


  xnor
  g331
  (
    n350,
    n219,
    n141,
    n237,
    n274
  );


  nor
  g332
  (
    n456,
    n327,
    n333,
    n250,
    n308
  );


  xor
  g333
  (
    n470,
    n236,
    n175,
    n244,
    n155
  );


  nand
  g334
  (
    n404,
    n178,
    n147,
    n255,
    n136
  );


  nand
  g335
  (
    n442,
    n82,
    n235,
    n269,
    n134
  );


  xor
  g336
  (
    n415,
    n290,
    n177,
    n301,
    n209
  );


  and
  g337
  (
    n457,
    n214,
    n173,
    n288,
    n142
  );


  nand
  g338
  (
    n503,
    n176,
    n257,
    n160,
    n134
  );


  xnor
  g339
  (
    n461,
    n236,
    n283,
    n329,
    n326
  );


  or
  g340
  (
    n510,
    n145,
    n200,
    n178,
    n194
  );


  and
  g341
  (
    n514,
    n246,
    n310,
    n214,
    n139
  );


  nand
  g342
  (
    n466,
    n218,
    n270,
    n130,
    n81
  );


  and
  g343
  (
    n505,
    n247,
    n215,
    n29,
    n233
  );


  and
  g344
  (
    n557,
    n295,
    n239,
    n332,
    n260
  );


  or
  g345
  (
    n483,
    n239,
    n310,
    n205,
    n294
  );


  xor
  g346
  (
    n484,
    n281,
    n161,
    n249,
    n229
  );


  or
  g347
  (
    n430,
    n309,
    n247,
    n288
  );


  xor
  g348
  (
    n384,
    n176,
    n334,
    n264,
    n333
  );


  or
  g349
  (
    n480,
    n157,
    n184,
    n140,
    n320
  );


  and
  g350
  (
    n538,
    n156,
    n314,
    n228,
    n330
  );


  or
  g351
  (
    n489,
    n145,
    n251,
    n163,
    n151
  );


  xnor
  g352
  (
    n395,
    n327,
    n177,
    n28,
    n226
  );


  nand
  g353
  (
    n523,
    n289,
    n24,
    n234,
    n231
  );


  nand
  g354
  (
    n463,
    n175,
    n260,
    n329,
    n181
  );


  xnor
  g355
  (
    n353,
    n261,
    n237,
    n137,
    n134
  );


  or
  g356
  (
    n344,
    n206,
    n212,
    n175,
    n311
  );


  and
  g357
  (
    n405,
    n218,
    n272,
    n204,
    n165
  );


  and
  g358
  (
    n385,
    n271,
    n133,
    n222,
    n285
  );


  and
  g359
  (
    n533,
    n244,
    n291,
    n286,
    n189
  );


  nand
  g360
  (
    n532,
    n173,
    n82,
    n169,
    n164
  );


  and
  g361
  (
    n418,
    n153,
    n170,
    n85,
    n133
  );


  and
  g362
  (
    n511,
    n255,
    n240,
    n296,
    n242
  );


  xor
  g363
  (
    n548,
    n221,
    n293,
    n205,
    n266
  );


  or
  g364
  (
    n401,
    n156,
    n177,
    n166,
    n307
  );


  xnor
  g365
  (
    n455,
    n77,
    n274,
    n135,
    n241
  );


  xor
  g366
  (
    n517,
    n159,
    n179,
    n250,
    n132
  );


  or
  g367
  (
    n377,
    n186,
    n298,
    n214,
    n259
  );


  nand
  g368
  (
    n346,
    n135,
    n280,
    n220,
    n195
  );


  and
  g369
  (
    n536,
    n86,
    n260,
    n301,
    n299
  );


  or
  g370
  (
    n481,
    n31,
    n202,
    n177,
    n315
  );


  nand
  g371
  (
    n406,
    n154,
    n205,
    n185,
    n27
  );


  xor
  g372
  (
    n542,
    n172,
    n297,
    n79,
    n331
  );


  nand
  g373
  (
    n535,
    n264,
    n277,
    n130,
    n131
  );


  or
  g374
  (
    n562,
    n253,
    n163,
    n281,
    n213
  );


  xor
  g375
  (
    n378,
    n157,
    n129,
    n22,
    n155
  );


  nand
  g376
  (
    n379,
    n137,
    n203,
    n266,
    n188
  );


  nor
  g377
  (
    n396,
    n141,
    n238,
    n158,
    n331
  );


  nor
  g378
  (
    n452,
    n324,
    n220,
    n211,
    n133
  );


  and
  g379
  (
    n446,
    n190,
    n230,
    n221,
    n335
  );


  and
  g380
  (
    n360,
    n25,
    n182,
    n132,
    n245
  );


  xnor
  g381
  (
    n370,
    n276,
    n180,
    n317,
    n323
  );


  xor
  g382
  (
    n450,
    n161,
    n176,
    n199,
    n281
  );


  nand
  g383
  (
    n388,
    n306,
    n308,
    n219,
    n23
  );


  xnor
  g384
  (
    n439,
    n282,
    n249,
    n199,
    n168
  );


  and
  g385
  (
    n567,
    n226,
    n312,
    n165,
    n179
  );


  xnor
  g386
  (
    n554,
    n317,
    n229,
    n152,
    n25
  );


  xor
  g387
  (
    n352,
    n216,
    n300,
    n268,
    n143
  );


  nand
  g388
  (
    KeyWire_0_23,
    n275,
    n207,
    n198,
    n155
  );


  xnor
  g389
  (
    n424,
    n259,
    n240,
    n193,
    n160
  );


  nand
  g390
  (
    n513,
    n233,
    n301,
    n182,
    n311
  );


  nand
  g391
  (
    n528,
    n159,
    n232,
    n174,
    n284
  );


  nand
  g392
  (
    n389,
    n328,
    n182,
    n278,
    n170
  );


  or
  g393
  (
    n383,
    n313,
    n190,
    n131,
    n144
  );


  nor
  g394
  (
    n478,
    n319,
    n274,
    n328,
    n81
  );


  nor
  g395
  (
    n364,
    n186,
    n196,
    n321,
    n294
  );


  xnor
  g396
  (
    n403,
    n136,
    n285,
    n169,
    n243
  );


  nor
  g397
  (
    n440,
    n198,
    n316,
    n196,
    n302
  );


  nor
  g398
  (
    n398,
    n146,
    n76,
    n234,
    n140
  );


  xor
  g399
  (
    n375,
    n151,
    n257,
    n319,
    n165
  );


  nand
  g400
  (
    n537,
    n222,
    n321,
    n261,
    n215
  );


  and
  g401
  (
    n436,
    n202,
    n227,
    n167,
    n326
  );


  or
  g402
  (
    n553,
    n261,
    n151,
    n246,
    n325
  );


  nand
  g403
  (
    n345,
    n304,
    n272,
    n174,
    n83
  );


  or
  g404
  (
    n357,
    n142,
    n84,
    n229,
    n28
  );


  nor
  g405
  (
    n520,
    n30,
    n159,
    n180,
    n300
  );


  or
  g406
  (
    n556,
    n326,
    n268,
    n225,
    n241
  );


  and
  g407
  (
    n506,
    n319,
    n147,
    n296,
    n298
  );


  xnor
  g408
  (
    n497,
    n229,
    n85,
    n150,
    n328
  );


  and
  g409
  (
    n555,
    n302,
    n241,
    n284,
    n318
  );


  xor
  g410
  (
    n391,
    n32,
    n280,
    n306,
    n225
  );


  xnor
  g411
  (
    n449,
    n222,
    n192,
    n208,
    n154
  );


  xor
  g412
  (
    n382,
    n153,
    n131,
    n180,
    n216
  );


  xnor
  g413
  (
    n423,
    n262,
    n206,
    n279,
    n323
  );


  or
  g414
  (
    n550,
    n145,
    n169,
    n147,
    n191
  );


  and
  g415
  (
    n515,
    n32,
    n213,
    n263,
    n318
  );


  xnor
  g416
  (
    n545,
    n307,
    n221,
    n202,
    n83
  );


  xnor
  g417
  (
    n568,
    n188,
    n85,
    n185,
    n246
  );


  xor
  g418
  (
    n410,
    n322,
    n219,
    n324,
    n76
  );


  or
  g419
  (
    n407,
    n184,
    n30,
    n319,
    n212
  );


  xor
  g420
  (
    n356,
    n236,
    n320,
    n172,
    n277
  );


  and
  g421
  (
    n492,
    n292,
    n164,
    n201,
    n268
  );


  xnor
  g422
  (
    n429,
    n220,
    n26,
    n242,
    n226
  );


  nand
  g423
  (
    n465,
    n305,
    n80,
    n146,
    n332
  );


  and
  g424
  (
    n438,
    n230,
    n244,
    n84,
    n135
  );


  and
  g425
  (
    n354,
    n184,
    n275,
    n263,
    n287
  );


  or
  g426
  (
    n460,
    n237,
    n234,
    n304,
    n25
  );


  or
  g427
  (
    n501,
    n204,
    n153,
    n135,
    n149
  );


  xnor
  g428
  (
    n496,
    n232,
    n210,
    n77,
    n140
  );


  nand
  g429
  (
    n551,
    n160,
    n180,
    n200,
    n278
  );


  xor
  g430
  (
    n380,
    n223,
    n291,
    n22,
    n268
  );


  xnor
  g431
  (
    n373,
    n79,
    n185,
    n31,
    n196
  );


  xor
  g432
  (
    n444,
    n190,
    n193,
    n174,
    n187
  );


  or
  g433
  (
    n534,
    n216,
    n84,
    n232,
    n30
  );


  xnor
  g434
  (
    n500,
    n196,
    n259,
    n304,
    n269
  );


  nor
  g435
  (
    n507,
    n208,
    n303,
    n171,
    n142
  );


  nand
  g436
  (
    n431,
    n213,
    n251,
    n327,
    n148
  );


  xor
  g437
  (
    n358,
    n313,
    n312,
    n292,
    n258
  );


  or
  g438
  (
    n521,
    n153,
    n152,
    n288,
    n322
  );


  nor
  g439
  (
    n413,
    n186,
    n206,
    n238,
    n265
  );


  nand
  g440
  (
    n408,
    n191,
    n152,
    n31,
    n78
  );


  xnor
  g441
  (
    n409,
    n327,
    n317,
    n198,
    n282
  );


  nand
  g442
  (
    n458,
    n185,
    n271,
    n217,
    n234
  );


  xnor
  g443
  (
    n529,
    n243,
    n280,
    n183,
    n249
  );


  xor
  g444
  (
    n469,
    n158,
    n162,
    n279,
    n323
  );


  xnor
  g445
  (
    n428,
    n150,
    n212,
    n164,
    n324
  );


  nor
  g446
  (
    n549,
    n83,
    n188,
    n138,
    n269
  );


  xnor
  g447
  (
    n371,
    n297,
    n295,
    n31,
    n207
  );


  nor
  g448
  (
    n476,
    n266,
    n201,
    n263,
    n198
  );


  xnor
  g449
  (
    n531,
    n292,
    n261,
    n132,
    n162
  );


  nor
  g450
  (
    n546,
    n272,
    n208,
    n187,
    n199
  );


  and
  g451
  (
    n530,
    n316,
    n300,
    n293,
    n156
  );


  or
  g452
  (
    n499,
    n201,
    n138,
    n86
  );


  xnor
  g453
  (
    n462,
    n256,
    n152,
    n240,
    n272
  );


  nand
  g454
  (
    n504,
    n255,
    n27,
    n143,
    n77
  );


  nand
  g455
  (
    n495,
    n24,
    n257,
    n174,
    n146
  );


  xor
  g456
  (
    n390,
    n320,
    n145,
    n291,
    n303
  );


  and
  g457
  (
    n386,
    n298,
    n144,
    n287,
    n312
  );


  xor
  g458
  (
    n490,
    n287,
    n333,
    n187,
    n76
  );


  nand
  g459
  (
    n566,
    n134,
    n179,
    n170,
    n166
  );


  xor
  g460
  (
    n491,
    n204,
    n325,
    n209,
    n187
  );


  xor
  g461
  (
    n411,
    n140,
    n139,
    n245,
    n298
  );


  xor
  g462
  (
    n399,
    n306,
    n239,
    n267,
    n194
  );


  xnor
  g463
  (
    n351,
    n191,
    n77,
    n289,
    n279
  );


  xor
  g464
  (
    n544,
    n143,
    n235,
    n209,
    n258
  );


  and
  g465
  (
    n524,
    n28,
    n226,
    n147,
    n263
  );


  or
  g466
  (
    n369,
    n330,
    n29,
    n262,
    n282
  );


  xnor
  g467
  (
    n365,
    n32,
    n306,
    n205,
    n252
  );


  nand
  g468
  (
    n559,
    n23,
    n332,
    n183,
    n227
  );


  or
  g469
  (
    n420,
    n167,
    n310,
    n251,
    n290
  );


  xnor
  g470
  (
    n475,
    n146,
    n320,
    n228,
    n25
  );


  or
  g471
  (
    n448,
    n211,
    n225,
    n216,
    n150
  );


  xor
  g472
  (
    n348,
    n221,
    n233,
    n175,
    n295
  );


  nor
  g473
  (
    n564,
    n295,
    n253,
    n137,
    n333
  );


  nand
  g474
  (
    n569,
    n217,
    n81,
    n210,
    n162
  );


  or
  g475
  (
    n498,
    n328,
    n218,
    n264,
    n168
  );


  nor
  g476
  (
    n427,
    n188,
    n267,
    n163,
    n323
  );


  or
  g477
  (
    n400,
    n200,
    n154,
    n283,
    n160
  );


  and
  g478
  (
    n355,
    n195,
    n211,
    n296,
    n223
  );


  xor
  g479
  (
    n426,
    n284,
    n189,
    n197,
    n274
  );


  or
  g480
  (
    n367,
    n23,
    n193,
    n276,
    n84
  );


  nand
  g481
  (
    n486,
    n250,
    n252,
    n273
  );


  and
  g482
  (
    n393,
    n173,
    n168,
    n157,
    n76
  );


  xnor
  g483
  (
    KeyWire_0_16,
    n233,
    n218,
    n316,
    n137
  );


  xor
  g484
  (
    n361,
    n172,
    n256,
    n314,
    n227
  );


  and
  g485
  (
    n482,
    n75,
    n270,
    n236,
    n243
  );


  and
  g486
  (
    n526,
    n253,
    n265,
    n192,
    n215
  );


  nand
  g487
  (
    n471,
    n231,
    n184,
    n308,
    n222
  );


  xor
  g488
  (
    n434,
    n28,
    n315,
    n223,
    n130
  );


  and
  g489
  (
    n552,
    n212,
    n245,
    n301,
    n148
  );


  and
  g490
  (
    n494,
    n215,
    n200,
    n331,
    n161
  );


  and
  g491
  (
    n412,
    n232,
    n293,
    n330,
    n310
  );


  and
  g492
  (
    n563,
    n225,
    n189,
    n315,
    n148
  );


  and
  g493
  (
    n443,
    n329,
    n210,
    n265,
    n194
  );


  and
  g494
  (
    n502,
    n82,
    n275,
    n133,
    n83
  );


  xor
  g495
  (
    n433,
    n80,
    n139,
    n241,
    n186
  );


  xor
  g496
  (
    n392,
    n302,
    n224,
    n26,
    n141
  );


  nor
  g497
  (
    n560,
    n203,
    n270,
    n271,
    n325
  );


  nand
  g498
  (
    n570,
    n286,
    n273,
    n161,
    n158
  );


  nor
  g499
  (
    n368,
    n201,
    n228,
    n157,
    n136
  );


  nor
  g500
  (
    n509,
    n209,
    n285,
    n142,
    n290
  );


  nor
  g501
  (
    n435,
    n262,
    n139,
    n173,
    n321
  );


  nand
  g502
  (
    n518,
    n79,
    n171,
    n163,
    n143
  );


  xnor
  g503
  (
    KeyWire_0_26,
    n183,
    n203,
    n292,
    n303
  );


  and
  g504
  (
    n422,
    n207,
    n329,
    n238,
    n26
  );


  xnor
  g505
  (
    n421,
    n279,
    n264,
    n162,
    n138
  );


  or
  g506
  (
    n372,
    n130,
    n230,
    n220,
    n317
  );


  xnor
  g507
  (
    n522,
    n254,
    n297,
    n244,
    n235
  );


  xnor
  g508
  (
    n417,
    n144,
    n315,
    n211,
    n171
  );


  xor
  g509
  (
    n374,
    n254,
    n213,
    n322,
    n195
  );


  xnor
  g510
  (
    n425,
    n78,
    n325,
    n150,
    n243
  );


  nor
  g511
  (
    n541,
    n280,
    n223,
    n299,
    n149
  );


  and
  g512
  (
    n402,
    n278,
    n283,
    n276,
    n324
  );


  or
  g513
  (
    n547,
    n195,
    n230,
    n307,
    n296
  );


  or
  g514
  (
    n347,
    n334,
    n167,
    n156,
    n277
  );


  xnor
  g515
  (
    n362,
    n191,
    n267,
    n228,
    n284
  );


  xor
  g516
  (
    n366,
    n276,
    n304,
    n269,
    n27
  );


  xnor
  g517
  (
    n472,
    n194,
    n251,
    n303,
    n242
  );


  nor
  g518
  (
    KeyWire_0_22,
    n307,
    n318,
    n248,
    n305
  );


  nand
  g519
  (
    n468,
    n335,
    n203,
    n178,
    n169
  );


  nor
  g520
  (
    n487,
    n197,
    n227,
    n24,
    n80
  );


  and
  g521
  (
    n543,
    n334,
    n252,
    n178
  );


  xnor
  g522
  (
    n432,
    n167,
    n217,
    n231,
    n154
  );


  or
  g523
  (
    n387,
    n132,
    n238,
    n32,
    n254
  );


  xnor
  g524
  (
    n473,
    n246,
    n256,
    n334,
    n309
  );


  xor
  g525
  (
    n381,
    n258,
    n287,
    n193,
    n219
  );


  or
  g526
  (
    n493,
    n293,
    n302,
    n183,
    n281
  );


  nand
  g527
  (
    n459,
    n288,
    n278,
    n332,
    n168
  );


  nand
  g528
  (
    n540,
    n309,
    n297,
    n189,
    n321
  );


  nor
  g529
  (
    n479,
    n206,
    n182,
    n190,
    n158
  );


  nand
  g530
  (
    n561,
    n308,
    n245,
    n235,
    n237
  );


  or
  g531
  (
    n359,
    n166,
    n231,
    n271,
    n79
  );


  xnor
  g532
  (
    n516,
    n78,
    n257,
    n275,
    n260
  );


  xnor
  g533
  (
    n394,
    n181,
    n170,
    n81,
    n85
  );


  nand
  g534
  (
    n519,
    n155,
    n291,
    n294,
    n313
  );


  xnor
  g535
  (
    n477,
    n144,
    n289,
    n266,
    n78
  );


  nand
  g536
  (
    n485,
    n240,
    n179,
    n248,
    n316
  );


  or
  g537
  (
    n445,
    n207,
    n214,
    n262,
    n300
  );


  buf
  g538
  (
    n576,
    n108
  );


  nand
  g539
  (
    n613,
    n375,
    n92,
    n100
  );


  or
  g540
  (
    n617,
    n341,
    n91,
    n112,
    n353
  );


  or
  g541
  (
    n594,
    n96,
    n110,
    n372,
    n375
  );


  or
  g542
  (
    n605,
    n370,
    n89,
    n86,
    n357
  );


  nand
  g543
  (
    n601,
    n88,
    n373,
    n103,
    n338
  );


  xor
  g544
  (
    n571,
    n373,
    n373,
    n344,
    n89
  );


  nor
  g545
  (
    n585,
    n372,
    n99,
    n363
  );


  nand
  g546
  (
    n583,
    n336,
    n93,
    n337,
    n374
  );


  nand
  g547
  (
    n603,
    n373,
    n109,
    n89,
    n349
  );


  nand
  g548
  (
    n574,
    n99,
    n103,
    n102,
    n100
  );


  or
  g549
  (
    n597,
    n92,
    n104,
    n98,
    n376
  );


  nand
  g550
  (
    n606,
    n90,
    n108,
    n92,
    n343
  );


  or
  g551
  (
    n579,
    n96,
    n374,
    n336,
    n106
  );


  and
  g552
  (
    n609,
    n336,
    n360,
    n372,
    n343
  );


  and
  g553
  (
    n611,
    n91,
    n375,
    n340,
    n104
  );


  xnor
  g554
  (
    n612,
    n102,
    n97,
    n93
  );


  nand
  g555
  (
    n584,
    n337,
    n99,
    n110,
    n348
  );


  nand
  g556
  (
    n581,
    n111,
    n91,
    n88,
    n100
  );


  xor
  g557
  (
    n610,
    n356,
    n101,
    n346,
    n105
  );


  and
  g558
  (
    n593,
    n94,
    n376,
    n335,
    n108
  );


  xor
  g559
  (
    n578,
    n358,
    n106,
    n101,
    n342
  );


  xor
  g560
  (
    n586,
    n337,
    n362,
    n95,
    n104
  );


  nand
  g561
  (
    n592,
    n368,
    n338,
    n341,
    n105
  );


  nor
  g562
  (
    n618,
    n110,
    n86,
    n361,
    n95
  );


  nor
  g563
  (
    n582,
    n375,
    n347,
    n339,
    n374
  );


  nor
  g564
  (
    n575,
    n336,
    n340,
    n342,
    n89
  );


  xnor
  g565
  (
    n608,
    n376,
    n90,
    n109,
    n365
  );


  or
  g566
  (
    n615,
    n94,
    n372,
    n345,
    n107
  );


  xor
  g567
  (
    n616,
    n91,
    n111,
    n107,
    n369
  );


  nor
  g568
  (
    n572,
    n112,
    n339,
    n352,
    n98
  );


  xnor
  g569
  (
    n589,
    n337,
    n341,
    n88,
    n103
  );


  nor
  g570
  (
    n591,
    n338,
    n90,
    n340,
    n95
  );


  and
  g571
  (
    n596,
    n87,
    n371,
    n101,
    n102
  );


  nand
  g572
  (
    n577,
    n339,
    n342,
    n374,
    n107
  );


  xor
  g573
  (
    n604,
    n111,
    n93,
    n376,
    n88
  );


  nor
  g574
  (
    n595,
    n100,
    n104,
    n339,
    n355
  );


  nand
  g575
  (
    n614,
    n105,
    n359,
    n350,
    n106
  );


  nand
  g576
  (
    n580,
    n87,
    n106,
    n335,
    n94
  );


  nand
  g577
  (
    n573,
    n93,
    n364,
    n98,
    n342
  );


  and
  g578
  (
    n599,
    n338,
    n97,
    n103,
    n108
  );


  nor
  g579
  (
    n598,
    n107,
    n95,
    n96,
    n92
  );


  nand
  g580
  (
    n590,
    n343,
    n96,
    n109,
    n97
  );


  nor
  g581
  (
    n602,
    n87,
    n367,
    n110,
    n354
  );


  nor
  g582
  (
    n607,
    n366,
    n105,
    n343,
    n94
  );


  xnor
  g583
  (
    n587,
    n340,
    n90,
    n112
  );


  nand
  g584
  (
    n600,
    n101,
    n351,
    n109,
    n111
  );


  xor
  g585
  (
    n588,
    n87,
    n98,
    n341,
    n102
  );


  and
  g586
  (
    KeyWire_0_30,
    n577,
    n409,
    n491
  );


  or
  g587
  (
    n681,
    n504,
    n415,
    n490,
    n602
  );


  xnor
  g588
  (
    n733,
    n452,
    n509,
    n595,
    n435
  );


  nand
  g589
  (
    n678,
    n519,
    n616,
    n456,
    n439
  );


  nand
  g590
  (
    KeyWire_0_1,
    n616,
    n497,
    n437,
    n435
  );


  or
  g591
  (
    n761,
    n489,
    n516,
    n519,
    n420
  );


  xor
  g592
  (
    n776,
    n401,
    n466,
    n405,
    n451
  );


  or
  g593
  (
    n757,
    n439,
    n440,
    n585,
    n378
  );


  and
  g594
  (
    n624,
    n396,
    n409,
    n492,
    n464
  );


  or
  g595
  (
    n747,
    n441,
    n599,
    n510,
    n488
  );


  xnor
  g596
  (
    n723,
    n464,
    n604,
    n395,
    n379
  );


  and
  g597
  (
    n638,
    n430,
    n470,
    n579,
    n397
  );


  and
  g598
  (
    n675,
    n575,
    n615,
    n428,
    n481
  );


  nand
  g599
  (
    n722,
    n498,
    n496,
    n470,
    n481
  );


  xnor
  g600
  (
    n720,
    n507,
    n506,
    n508,
    n468
  );


  and
  g601
  (
    n784,
    n589,
    n575,
    n488,
    n442
  );


  and
  g602
  (
    n657,
    n613,
    n472,
    n419,
    n583
  );


  xor
  g603
  (
    n654,
    n433,
    n494,
    n479,
    n498
  );


  xor
  g604
  (
    n752,
    n477,
    n601,
    n438,
    n511
  );


  or
  g605
  (
    n730,
    n475,
    n393,
    n605,
    n422
  );


  nand
  g606
  (
    n773,
    n408,
    n503,
    n592,
    n460
  );


  and
  g607
  (
    n808,
    n584,
    n425,
    n476,
    n388
  );


  or
  g608
  (
    n684,
    n592,
    n614,
    n451,
    n385
  );


  and
  g609
  (
    n651,
    n485,
    n579,
    n580,
    n406
  );


  nor
  g610
  (
    n754,
    n481,
    n445,
    n479,
    n505
  );


  xor
  g611
  (
    n689,
    n502,
    n476,
    n493,
    n397
  );


  or
  g612
  (
    n691,
    n379,
    n505,
    n611,
    n468
  );


  nand
  g613
  (
    KeyWire_0_3,
    n581,
    n380,
    n609,
    n510
  );


  xor
  g614
  (
    n628,
    n399,
    n385,
    n453,
    n482
  );


  nand
  g615
  (
    n688,
    n400,
    n470,
    n403,
    n612
  );


  nor
  g616
  (
    n724,
    n572,
    n424,
    n496,
    n463
  );


  xnor
  g617
  (
    n788,
    n406,
    n411,
    n394,
    n593
  );


  nand
  g618
  (
    n780,
    n420,
    n604,
    n453,
    n616
  );


  or
  g619
  (
    n745,
    n497,
    n441,
    n573,
    n449
  );


  nand
  g620
  (
    n759,
    n474,
    n386,
    n408,
    n513
  );


  xnor
  g621
  (
    n633,
    n401,
    n607,
    n489,
    n446
  );


  nor
  g622
  (
    n707,
    n580,
    n410,
    n511,
    n431
  );


  xor
  g623
  (
    n700,
    n418,
    n576,
    n518,
    n398
  );


  nor
  g624
  (
    n798,
    n441,
    n583,
    n438,
    n415
  );


  and
  g625
  (
    n726,
    n412,
    n394,
    n581,
    n517
  );


  xor
  g626
  (
    n644,
    n393,
    n587,
    n480,
    n513
  );


  and
  g627
  (
    n727,
    n378,
    n483,
    n447,
    n450
  );


  or
  g628
  (
    n721,
    n387,
    n458,
    n452,
    n520
  );


  or
  g629
  (
    n667,
    n380,
    n402,
    n436,
    n457
  );


  and
  g630
  (
    n658,
    n598,
    n382,
    n575,
    n396
  );


  nor
  g631
  (
    n660,
    n447,
    n472,
    n423,
    n383
  );


  nor
  g632
  (
    n706,
    n451,
    n394,
    n495,
    n587
  );


  nand
  g633
  (
    n765,
    n583,
    n586,
    n469,
    n496
  );


  nor
  g634
  (
    KeyWire_0_25,
    n595,
    n418,
    n473,
    n471
  );


  nand
  g635
  (
    n661,
    n490,
    n425,
    n433,
    n506
  );


  nand
  g636
  (
    n710,
    n615,
    n491,
    n508,
    n414
  );


  or
  g637
  (
    n630,
    n588,
    n590,
    n429,
    n389
  );


  xnor
  g638
  (
    n639,
    n458,
    n512,
    n460,
    n476
  );


  and
  g639
  (
    n637,
    n589,
    n511,
    n445,
    n579
  );


  or
  g640
  (
    KeyWire_0_5,
    n608,
    n428,
    n451,
    n469
  );


  nand
  g641
  (
    n717,
    n422,
    n500,
    n454,
    n418
  );


  nor
  g642
  (
    n627,
    n504,
    n516,
    n408,
    n606
  );


  or
  g643
  (
    n666,
    n472,
    n501,
    n407,
    n427
  );


  xor
  g644
  (
    n652,
    n441,
    n576,
    n399,
    n469
  );


  xor
  g645
  (
    n711,
    n385,
    n595,
    n389,
    n479
  );


  nand
  g646
  (
    n748,
    n476,
    n390,
    n613,
    n504
  );


  and
  g647
  (
    KeyWire_0_28,
    n582,
    n571,
    n607,
    n429
  );


  nand
  g648
  (
    n778,
    n609,
    n508,
    n510,
    n472
  );


  nand
  g649
  (
    n802,
    n413,
    n573,
    n506,
    n455
  );


  nor
  g650
  (
    n673,
    n573,
    n505,
    n383,
    n462
  );


  xnor
  g651
  (
    n622,
    n449,
    n475,
    n423,
    n386
  );


  nand
  g652
  (
    n664,
    n377,
    n377,
    n417,
    n384
  );


  nand
  g653
  (
    n737,
    n417,
    n484,
    n398,
    n584
  );


  xnor
  g654
  (
    n792,
    n610,
    n416,
    n512,
    n618
  );


  and
  g655
  (
    n782,
    n396,
    n485,
    n431,
    n421
  );


  xor
  g656
  (
    n696,
    n393,
    n605,
    n434,
    n391
  );


  xor
  g657
  (
    n695,
    n402,
    n444,
    n412,
    n600
  );


  and
  g658
  (
    n766,
    n512,
    n416,
    n617,
    n515
  );


  xor
  g659
  (
    n728,
    n502,
    n497,
    n465,
    n573
  );


  or
  g660
  (
    n671,
    n603,
    n612,
    n500,
    n436
  );


  and
  g661
  (
    n672,
    n594,
    n446,
    n413,
    n592
  );


  or
  g662
  (
    n648,
    n477,
    n483,
    n459,
    n576
  );


  nand
  g663
  (
    n665,
    n437,
    n606,
    n400,
    n419
  );


  nand
  g664
  (
    n685,
    n467,
    n503,
    n402,
    n431
  );


  or
  g665
  (
    n807,
    n404,
    n468,
    n450,
    n462
  );


  or
  g666
  (
    n682,
    n471,
    n377,
    n420,
    n602
  );


  nor
  g667
  (
    n756,
    n617,
    n518,
    n456,
    n453
  );


  or
  g668
  (
    n719,
    n483,
    n571,
    n435,
    n395
  );


  nand
  g669
  (
    n793,
    n446,
    n417,
    n518,
    n424
  );


  nor
  g670
  (
    n753,
    n578,
    n520,
    n460,
    n603
  );


  and
  g671
  (
    n626,
    n419,
    n484,
    n597,
    n416
  );


  nor
  g672
  (
    n740,
    n514,
    n616,
    n430,
    n432
  );


  xor
  g673
  (
    n749,
    n450,
    n495,
    n407,
    n517
  );


  nor
  g674
  (
    n805,
    n432,
    n607,
    n609,
    n467
  );


  xnor
  g675
  (
    n789,
    n461,
    n576,
    n397,
    n443
  );


  nor
  g676
  (
    n803,
    n473,
    n501,
    n405,
    n617
  );


  xnor
  g677
  (
    n683,
    n462,
    n505,
    n464,
    n488
  );


  xor
  g678
  (
    n646,
    n486,
    n431,
    n509,
    n577
  );


  xnor
  g679
  (
    KeyWire_0_27,
    n404,
    n480,
    n592,
    n400
  );


  and
  g680
  (
    n734,
    n427,
    n463,
    n426,
    n425
  );


  nand
  g681
  (
    n809,
    n410,
    n394,
    n435,
    n378
  );


  and
  g682
  (
    n714,
    n415,
    n438,
    n444,
    n482
  );


  nor
  g683
  (
    KeyWire_0_8,
    n454,
    n416,
    n404,
    n465
  );


  nand
  g684
  (
    n736,
    n519,
    n474,
    n488,
    n503
  );


  xnor
  g685
  (
    n697,
    n517,
    n610,
    n390,
    n590
  );


  nand
  g686
  (
    n647,
    n420,
    n399,
    n411,
    n422
  );


  or
  g687
  (
    n732,
    n614,
    n590,
    n577,
    n466
  );


  or
  g688
  (
    n738,
    n466,
    n459,
    n596,
    n477
  );


  xnor
  g689
  (
    n645,
    n583,
    n393,
    n390,
    n507
  );


  and
  g690
  (
    n643,
    n459,
    n406,
    n574,
    n601
  );


  xnor
  g691
  (
    n735,
    n392,
    n419,
    n411,
    n577
  );


  nor
  g692
  (
    n699,
    n586,
    n455,
    n572,
    n425
  );


  and
  g693
  (
    n701,
    n414,
    n613,
    n456,
    n499
  );


  nor
  g694
  (
    n758,
    n446,
    n407,
    n412,
    n496
  );


  xnor
  g695
  (
    n656,
    n611,
    n591,
    n596,
    n479
  );


  nor
  g696
  (
    n620,
    n590,
    n512,
    n440,
    n426
  );


  or
  g697
  (
    n783,
    n511,
    n614,
    n452,
    n515
  );


  nand
  g698
  (
    n744,
    n486,
    n387,
    n379,
    n430
  );


  xnor
  g699
  (
    n806,
    n397,
    n403,
    n571,
    n461
  );


  and
  g700
  (
    n642,
    n385,
    n502,
    n437,
    n414
  );


  xor
  g701
  (
    n662,
    n461,
    n378,
    n409,
    n464
  );


  xnor
  g702
  (
    n625,
    n388,
    n442,
    n432,
    n486
  );


  xor
  g703
  (
    n746,
    n482,
    n422,
    n387,
    n501
  );


  and
  g704
  (
    n669,
    n401,
    n434,
    n381,
    n405
  );


  and
  g705
  (
    n786,
    n491,
    n421,
    n609,
    n582
  );


  or
  g706
  (
    n768,
    n388,
    n581,
    n428,
    n603
  );


  or
  g707
  (
    n751,
    n392,
    n518,
    n465,
    n618
  );


  nor
  g708
  (
    n635,
    n445,
    n607,
    n589,
    n467
  );


  and
  g709
  (
    n715,
    n421,
    n509,
    n458,
    n485
  );


  xnor
  g710
  (
    n690,
    n587,
    n423,
    n443,
    n381
  );


  xor
  g711
  (
    n668,
    n465,
    n497,
    n601,
    n571
  );


  and
  g712
  (
    n770,
    n507,
    n482,
    n605,
    n480
  );


  xnor
  g713
  (
    n777,
    n391,
    n584,
    n478,
    n448
  );


  or
  g714
  (
    n709,
    n388,
    n380,
    n608
  );


  or
  g715
  (
    n698,
    n387,
    n606,
    n379,
    n448
  );


  or
  g716
  (
    n795,
    n389,
    n478,
    n513,
    n437
  );


  nand
  g717
  (
    n634,
    n439,
    n600,
    n447,
    n501
  );


  xor
  g718
  (
    n702,
    n581,
    n461,
    n613,
    n515
  );


  xor
  g719
  (
    n631,
    n593,
    n588,
    n618,
    n519
  );


  xnor
  g720
  (
    n797,
    n411,
    n407,
    n513,
    n587
  );


  nor
  g721
  (
    n621,
    n604,
    n598,
    n517,
    n384
  );


  xor
  g722
  (
    n679,
    n608,
    n598,
    n395,
    n584
  );


  xnor
  g723
  (
    n725,
    n586,
    n429,
    n575,
    n452
  );


  or
  g724
  (
    n787,
    n449,
    n383,
    n457,
    n474
  );


  xnor
  g725
  (
    n799,
    n490,
    n408,
    n484,
    n487
  );


  xnor
  g726
  (
    n674,
    n492,
    n484,
    n429,
    n588
  );


  xnor
  g727
  (
    n755,
    n478,
    n382,
    n608
  );


  or
  g728
  (
    KeyWire_0_20,
    n611,
    n582,
    n615,
    n428
  );


  and
  g729
  (
    n769,
    n591,
    n470,
    n426,
    n456
  );


  xor
  g730
  (
    n750,
    n392,
    n403,
    n596,
    n600
  );


  nand
  g731
  (
    n649,
    n398,
    n406,
    n399,
    n447
  );


  and
  g732
  (
    n796,
    n405,
    n457,
    n433,
    n612
  );


  and
  g733
  (
    n800,
    n448,
    n500,
    n604,
    n389
  );


  xnor
  g734
  (
    n653,
    n492,
    n574,
    n442,
    n423
  );


  and
  g735
  (
    n677,
    n618,
    n498,
    n585,
    n471
  );


  nand
  g736
  (
    n772,
    n489,
    n481,
    n591,
    n398
  );


  and
  g737
  (
    n705,
    n443,
    n386,
    n503,
    n466
  );


  xnor
  g738
  (
    n767,
    n597,
    n426,
    n510,
    n617
  );


  xnor
  g739
  (
    n810,
    n436,
    n414,
    n594,
    n415
  );


  nand
  g740
  (
    n694,
    n473,
    n504,
    n514,
    n508
  );


  or
  g741
  (
    n655,
    n469,
    n605,
    n580,
    n458
  );


  or
  g742
  (
    n670,
    n486,
    n460,
    n390,
    n396
  );


  xnor
  g743
  (
    n741,
    n520,
    n601,
    n453,
    n400
  );


  and
  g744
  (
    n693,
    n483,
    n480,
    n574,
    n404
  );


  or
  g745
  (
    n632,
    n391,
    n578,
    n595,
    n493
  );


  nand
  g746
  (
    n781,
    n507,
    n599,
    n442,
    n494
  );


  and
  g747
  (
    n629,
    n463,
    n448,
    n602,
    n494
  );


  or
  g748
  (
    n760,
    n430,
    n572,
    n610,
    n410
  );


  and
  g749
  (
    n703,
    n439,
    n612,
    n440,
    n392
  );


  xor
  g750
  (
    n659,
    n377,
    n440,
    n514,
    n487
  );


  nor
  g751
  (
    n716,
    n384,
    n427,
    n487,
    n591
  );


  and
  g752
  (
    n718,
    n475,
    n499,
    n445,
    n493
  );


  nand
  g753
  (
    n779,
    n599,
    n491,
    n432,
    n516
  );


  nand
  g754
  (
    n731,
    n489,
    n433,
    n574,
    n391
  );


  nor
  g755
  (
    n801,
    n597,
    n449,
    n603,
    n477
  );


  xor
  g756
  (
    n794,
    n487,
    n443,
    n478,
    n610
  );


  or
  g757
  (
    n641,
    n494,
    n471,
    n413,
    n438
  );


  xnor
  g758
  (
    n619,
    n382,
    n611,
    n413,
    n474
  );


  and
  g759
  (
    n636,
    n515,
    n599,
    n614,
    n602
  );


  and
  g760
  (
    n704,
    n450,
    n593,
    n578,
    n499
  );


  or
  g761
  (
    n712,
    n582,
    n401,
    n598,
    n600
  );


  or
  g762
  (
    n686,
    n572,
    n434,
    n412,
    n410
  );


  or
  g763
  (
    n742,
    n495,
    n502,
    n455,
    n615
  );


  or
  g764
  (
    n762,
    n444,
    n455,
    n421,
    n402
  );


  xor
  g765
  (
    n775,
    n381,
    n418,
    n514,
    n459
  );


  nor
  g766
  (
    n790,
    n468,
    n381,
    n516,
    n490
  );


  or
  g767
  (
    n623,
    n403,
    n454,
    n506,
    n588
  );


  and
  g768
  (
    n743,
    n593,
    n463,
    n500,
    n594
  );


  xor
  g769
  (
    n680,
    n498,
    n434,
    n395,
    n586
  );


  nor
  g770
  (
    n771,
    n454,
    n436,
    n485,
    n585
  );


  xor
  g771
  (
    n764,
    n462,
    n467,
    n457,
    n493
  );


  xnor
  g772
  (
    n676,
    n386,
    n417,
    n594,
    n606
  );


  and
  g773
  (
    n774,
    n424,
    n475,
    n579,
    n597
  );


  nor
  g774
  (
    n692,
    n580,
    n495,
    n384,
    n585
  );


  xor
  g775
  (
    n763,
    n473,
    n424,
    n427,
    n520
  );


  xor
  g776
  (
    n804,
    n509,
    n499,
    n492,
    n383
  );


  and
  g777
  (
    n739,
    n589,
    n444,
    n596,
    n578
  );


  buf
  g778
  (
    n814,
    n718
  );


  not
  g779
  (
    n919,
    n562
  );


  buf
  g780
  (
    n902,
    n560
  );


  not
  g781
  (
    n922,
    n661
  );


  buf
  g782
  (
    n812,
    n651
  );


  not
  g783
  (
    n824,
    n717
  );


  buf
  g784
  (
    n871,
    n561
  );


  not
  g785
  (
    n842,
    n756
  );


  xor
  g786
  (
    n836,
    n762,
    n747,
    n522,
    n732
  );


  xor
  g787
  (
    n848,
    n544,
    n731,
    n719,
    n648
  );


  nand
  g788
  (
    n823,
    n521,
    n723,
    n531,
    n764
  );


  xnor
  g789
  (
    n907,
    n623,
    n766,
    n568,
    n735
  );


  nor
  g790
  (
    n826,
    n528,
    n750,
    n732,
    n721
  );


  xor
  g791
  (
    n924,
    n522,
    n567,
    n546,
    n530
  );


  nand
  g792
  (
    n821,
    n563,
    n726,
    n765,
    n739
  );


  nand
  g793
  (
    KeyWire_0_11,
    n527,
    n760,
    n758,
    n754
  );


  nor
  g794
  (
    n940,
    n523,
    n535,
    n529,
    n545
  );


  xnor
  g795
  (
    n864,
    n751,
    n536,
    n667,
    n758
  );


  nor
  g796
  (
    n914,
    n541,
    n532,
    n570,
    n529
  );


  or
  g797
  (
    n927,
    n556,
    n707,
    n532,
    n756
  );


  xor
  g798
  (
    n820,
    n725,
    n552,
    n555,
    n738
  );


  nand
  g799
  (
    n854,
    n534,
    n759,
    n747,
    n741
  );


  and
  g800
  (
    n875,
    n541,
    n540,
    n682,
    n743
  );


  or
  g801
  (
    n831,
    n672,
    n538,
    n526,
    n710
  );


  nor
  g802
  (
    n938,
    n540,
    n713,
    n728,
    n521
  );


  or
  g803
  (
    n890,
    n742,
    n647,
    n727,
    n554
  );


  nor
  g804
  (
    n901,
    n696,
    n750,
    n738,
    n702
  );


  nor
  g805
  (
    n844,
    n717,
    n745,
    n529,
    n757
  );


  nand
  g806
  (
    n867,
    n736,
    n760,
    n664,
    n550
  );


  nor
  g807
  (
    n887,
    n742,
    n553,
    n748,
    n570
  );


  or
  g808
  (
    n846,
    n656,
    n749,
    n745,
    n558
  );


  nand
  g809
  (
    n866,
    n700,
    n552,
    n525,
    n692
  );


  xor
  g810
  (
    n896,
    n568,
    n558,
    n732,
    n756
  );


  and
  g811
  (
    n892,
    n737,
    n622,
    n666,
    n646
  );


  xor
  g812
  (
    n861,
    n668,
    n738,
    n524,
    n735
  );


  nand
  g813
  (
    n847,
    n552,
    n720,
    n636,
    n729
  );


  nor
  g814
  (
    n858,
    n643,
    n753,
    n746
  );


  or
  g815
  (
    n921,
    n556,
    n717,
    n534,
    n762
  );


  or
  g816
  (
    n937,
    n699,
    n719,
    n687,
    n525
  );


  or
  g817
  (
    n850,
    n663,
    n759,
    n533,
    n724
  );


  and
  g818
  (
    n884,
    n697,
    n543,
    n764,
    n675
  );


  or
  g819
  (
    n898,
    n529,
    n559,
    n759,
    n549
  );


  xnor
  g820
  (
    n834,
    n565,
    n681,
    n554,
    n734
  );


  xor
  g821
  (
    n888,
    n752,
    n709,
    n551,
    n721
  );


  or
  g822
  (
    n899,
    n740,
    n757,
    n539,
    n727
  );


  or
  g823
  (
    n935,
    n765,
    n521,
    n722,
    n726
  );


  nor
  g824
  (
    n839,
    n754,
    n752,
    n734,
    n522
  );


  or
  g825
  (
    n868,
    n550,
    n739,
    n543,
    n628
  );


  or
  g826
  (
    n828,
    n539,
    n557,
    n525,
    n536
  );


  xor
  g827
  (
    n853,
    n522,
    n743,
    n728,
    n538
  );


  xnor
  g828
  (
    n862,
    n650,
    n554,
    n548,
    n744
  );


  xnor
  g829
  (
    n873,
    n526,
    n569,
    n546,
    n632
  );


  xor
  g830
  (
    n897,
    n541,
    n670,
    n528,
    n757
  );


  or
  g831
  (
    n822,
    n743,
    n761,
    n723,
    n679
  );


  nand
  g832
  (
    n852,
    n759,
    n738,
    n674,
    n558
  );


  xor
  g833
  (
    n908,
    n686,
    n722,
    n564,
    n745
  );


  nor
  g834
  (
    n923,
    n760,
    n545,
    n557,
    n566
  );


  xor
  g835
  (
    n930,
    n523,
    n553,
    n530,
    n693
  );


  xor
  g836
  (
    n885,
    n753,
    n665,
    n763
  );


  or
  g837
  (
    n912,
    n560,
    n531,
    n737,
    n547
  );


  and
  g838
  (
    n833,
    n629,
    n718,
    n533,
    n569
  );


  and
  g839
  (
    n825,
    n727,
    n673,
    n748,
    n625
  );


  nor
  g840
  (
    n911,
    n705,
    n540,
    n530,
    n548
  );


  nor
  g841
  (
    n936,
    n721,
    n725,
    n730,
    n755
  );


  nand
  g842
  (
    n818,
    n750,
    n761,
    n723,
    n742
  );


  nor
  g843
  (
    n905,
    n547,
    n639,
    n569,
    n564
  );


  nand
  g844
  (
    n819,
    n566,
    n749,
    n565,
    n621
  );


  or
  g845
  (
    n904,
    n556,
    n640,
    n727,
    n542
  );


  xor
  g846
  (
    n856,
    n523,
    n534,
    n620,
    n676
  );


  or
  g847
  (
    n880,
    n695,
    n685,
    n561,
    n677
  );


  xor
  g848
  (
    n863,
    n535,
    n527,
    n757,
    n691
  );


  and
  g849
  (
    n838,
    n551,
    n657,
    n718,
    n546
  );


  xnor
  g850
  (
    n910,
    n523,
    n763,
    n530,
    n542
  );


  xor
  g851
  (
    n857,
    n524,
    n559,
    n566,
    n560
  );


  xnor
  g852
  (
    n913,
    n739,
    n566,
    n539,
    n729
  );


  xnor
  g853
  (
    KeyWire_0_31,
    n730,
    n543,
    n726,
    n536
  );


  and
  g854
  (
    n843,
    n562,
    n570,
    n540,
    n535
  );


  nand
  g855
  (
    n878,
    n655,
    n548,
    n538,
    n745
  );


  xor
  g856
  (
    n895,
    n555,
    n549,
    n550,
    n761
  );


  nand
  g857
  (
    n813,
    n750,
    n645,
    n706,
    n712
  );


  xor
  g858
  (
    n934,
    n626,
    n634,
    n723,
    n550
  );


  or
  g859
  (
    n939,
    n544,
    n720,
    n716,
    n658
  );


  nand
  g860
  (
    n916,
    n729,
    n546,
    n567,
    n641
  );


  xnor
  g861
  (
    n872,
    n537,
    n704,
    n562,
    n756
  );


  xnor
  g862
  (
    n889,
    n531,
    n736,
    n743,
    n549
  );


  xor
  g863
  (
    n929,
    n737,
    n749,
    n730,
    n744
  );


  nor
  g864
  (
    n915,
    n755,
    n538,
    n536,
    n724
  );


  nand
  g865
  (
    n882,
    n547,
    n558,
    n557,
    n741
  );


  nand
  g866
  (
    n865,
    n722,
    n764,
    n559,
    n624
  );


  or
  g867
  (
    n827,
    n725,
    n562,
    n703,
    n678
  );


  or
  g868
  (
    n851,
    n744,
    n531,
    n535,
    n728
  );


  nand
  g869
  (
    n816,
    n553,
    n542,
    n551,
    n557
  );


  or
  g870
  (
    n925,
    n690,
    n732,
    n542,
    n537
  );


  nand
  g871
  (
    n891,
    n718,
    n565,
    n537,
    n555
  );


  nor
  g872
  (
    n845,
    n737,
    n563,
    n548,
    n564
  );


  xnor
  g873
  (
    n855,
    n532,
    n551,
    n544,
    n527
  );


  nand
  g874
  (
    n876,
    n568,
    n635,
    n747,
    n627
  );


  or
  g875
  (
    n829,
    n720,
    n751,
    n554,
    n653
  );


  xor
  g876
  (
    n906,
    n739,
    n545,
    n733,
    n729
  );


  nand
  g877
  (
    n883,
    n740,
    n740,
    n735,
    n698
  );


  xor
  g878
  (
    n869,
    n747,
    n660,
    n556,
    n731
  );


  nand
  g879
  (
    n893,
    n720,
    n559,
    n526,
    n525
  );


  xor
  g880
  (
    n870,
    n528,
    n752,
    n755,
    n524
  );


  or
  g881
  (
    n815,
    n724,
    n711,
    n638,
    n521
  );


  nor
  g882
  (
    n928,
    n731,
    n537,
    n760,
    n733
  );


  xor
  g883
  (
    n859,
    n748,
    n736,
    n724,
    n547
  );


  nor
  g884
  (
    n903,
    n736,
    n659,
    n654,
    n543
  );


  and
  g885
  (
    n860,
    n532,
    n644,
    n751,
    n671
  );


  nand
  g886
  (
    n909,
    n721,
    n524,
    n733,
    n544
  );


  and
  g887
  (
    n894,
    n749,
    n725,
    n714,
    n528
  );


  or
  g888
  (
    n931,
    n734,
    n552,
    n719,
    n761
  );


  or
  g889
  (
    n920,
    n746,
    n541,
    n564,
    n569
  );


  nand
  g890
  (
    n837,
    n526,
    n533,
    n563,
    n731
  );


  xor
  g891
  (
    n918,
    n565,
    n560,
    n662,
    n684
  );


  or
  g892
  (
    n835,
    n766,
    n689,
    n534,
    n533
  );


  nand
  g893
  (
    n874,
    n741,
    n527,
    n758,
    n649
  );


  xnor
  g894
  (
    n832,
    n561,
    n568,
    n555,
    n753
  );


  xnor
  g895
  (
    KeyWire_0_17,
    n726,
    n637,
    n755,
    n744
  );


  xor
  g896
  (
    n933,
    n553,
    n765,
    n740,
    n722
  );


  nor
  g897
  (
    n840,
    n715,
    n728,
    n642,
    n758
  );


  xor
  g898
  (
    n817,
    n701,
    n765,
    n694,
    n751
  );


  nand
  g899
  (
    n841,
    n669,
    n735,
    n763,
    n680
  );


  nand
  g900
  (
    n900,
    n539,
    n746,
    n549,
    n748
  );


  or
  g901
  (
    KeyWire_0_21,
    n754,
    n730,
    n633,
    n630
  );


  and
  g902
  (
    n917,
    n652,
    n563,
    n734,
    n733
  );


  and
  g903
  (
    n886,
    n752,
    n754,
    n683,
    n688
  );


  nand
  g904
  (
    n830,
    n742,
    n619,
    n717,
    n719
  );


  xor
  g905
  (
    n926,
    n746,
    n762,
    n561,
    n708
  );


  nor
  g906
  (
    KeyWire_0_12,
    n631,
    n762,
    n567,
    n545
  );


  nand
  g907
  (
    KeyWire_0_2,
    n570,
    n764,
    n567,
    n741
  );


  nor
  g908
  (
    n964,
    n781,
    n795,
    n766,
    n777
  );


  or
  g909
  (
    n977,
    n780,
    n784,
    n795,
    n782
  );


  xor
  g910
  (
    n948,
    n788,
    n787,
    n785,
    n771
  );


  nand
  g911
  (
    n957,
    n794,
    n812,
    n790,
    n774
  );


  and
  g912
  (
    n950,
    n786,
    n774,
    n826,
    n780
  );


  nand
  g913
  (
    n953,
    n767,
    n822,
    n788,
    n837
  );


  and
  g914
  (
    KeyWire_0_0,
    n777,
    n818,
    n848,
    n794
  );


  xnor
  g915
  (
    n944,
    n832,
    n791,
    n792,
    n820
  );


  xnor
  g916
  (
    n946,
    n770,
    n785,
    n819,
    n844
  );


  xnor
  g917
  (
    n975,
    n793,
    n766,
    n771,
    n830
  );


  nor
  g918
  (
    n972,
    n782,
    n777,
    n767,
    n795
  );


  or
  g919
  (
    n942,
    n784,
    n786,
    n769,
    n773
  );


  and
  g920
  (
    n943,
    n831,
    n783,
    n842,
    n785
  );


  nor
  g921
  (
    n956,
    n767,
    n773,
    n796,
    n768
  );


  or
  g922
  (
    n966,
    n776,
    n777,
    n829,
    n792
  );


  or
  g923
  (
    n951,
    n814,
    n786,
    n778,
    n843
  );


  or
  g924
  (
    n947,
    n787,
    n784,
    n768,
    n811
  );


  xnor
  g925
  (
    n952,
    n834,
    n781,
    n776,
    n775
  );


  nor
  g926
  (
    n962,
    n779,
    n815,
    n769,
    n772
  );


  or
  g927
  (
    n961,
    n825,
    n791,
    n783,
    n790
  );


  xor
  g928
  (
    n967,
    n780,
    n778,
    n841,
    n788
  );


  xnor
  g929
  (
    n979,
    n769,
    n772,
    n840,
    n784
  );


  xnor
  g930
  (
    n969,
    n779,
    n770,
    n771,
    n772
  );


  xnor
  g931
  (
    n973,
    n767,
    n821,
    n836,
    n790
  );


  or
  g932
  (
    n971,
    n789,
    n791,
    n786,
    n823
  );


  nand
  g933
  (
    n963,
    n775,
    n770,
    n835,
    n828
  );


  xnor
  g934
  (
    n980,
    n787,
    n785,
    n776,
    n813
  );


  or
  g935
  (
    n958,
    n779,
    n793,
    n789,
    n791
  );


  nor
  g936
  (
    n968,
    n782,
    n792,
    n789,
    n775
  );


  xnor
  g937
  (
    n945,
    n850,
    n769,
    n783,
    n788
  );


  xnor
  g938
  (
    n949,
    n796,
    n846,
    n781,
    n770
  );


  xnor
  g939
  (
    n960,
    n847,
    n833,
    n792,
    n780
  );


  nor
  g940
  (
    n976,
    n774,
    n816,
    n771,
    n776
  );


  xor
  g941
  (
    n978,
    n839,
    n794,
    n779,
    n817
  );


  xor
  g942
  (
    n941,
    n787,
    n781,
    n845,
    n827
  );


  xor
  g943
  (
    n955,
    n790,
    n768,
    n778,
    n773
  );


  nor
  g944
  (
    n974,
    n783,
    n782,
    n774,
    n795
  );


  or
  g945
  (
    n959,
    n793,
    n838,
    n775,
    n778
  );


  nor
  g946
  (
    n970,
    n768,
    n789,
    n772,
    n849
  );


  xnor
  g947
  (
    n954,
    n794,
    n773,
    n793,
    n824
  );


  nor
  g948
  (
    n985,
    n943,
    n909,
    n874,
    n797
  );


  nor
  g949
  (
    n999,
    n893,
    n889,
    n936,
    n971
  );


  xor
  g950
  (
    n1006,
    n798,
    n927,
    n913,
    n901
  );


  nand
  g951
  (
    n997,
    n952,
    n959,
    n977,
    n911
  );


  or
  g952
  (
    n1000,
    n914,
    n968,
    n976,
    n879
  );


  xor
  g953
  (
    n1008,
    n966,
    n970,
    n975,
    n799
  );


  or
  g954
  (
    n990,
    n965,
    n941,
    n897,
    n929
  );


  xnor
  g955
  (
    n1007,
    n799,
    n866,
    n881,
    n932
  );


  nor
  g956
  (
    n1017,
    n886,
    n951,
    n851,
    n857
  );


  xor
  g957
  (
    n1016,
    n796,
    n947,
    n933,
    n870
  );


  or
  g958
  (
    n1010,
    n860,
    n872,
    n920,
    n796
  );


  xor
  g959
  (
    n998,
    n946,
    n892,
    n915,
    n853
  );


  and
  g960
  (
    n1002,
    n907,
    n926,
    n979,
    n938
  );


  nand
  g961
  (
    n996,
    n877,
    n880,
    n856,
    n905
  );


  nor
  g962
  (
    n1011,
    n859,
    n910,
    n935,
    n955
  );


  xor
  g963
  (
    n1004,
    n918,
    n930,
    n980,
    n800
  );


  and
  g964
  (
    n1015,
    n899,
    n876,
    n801,
    n948
  );


  nor
  g965
  (
    n993,
    n895,
    n937,
    n852,
    n928
  );


  xor
  g966
  (
    n995,
    n855,
    n882,
    n902,
    n896
  );


  nand
  g967
  (
    n1018,
    n888,
    n963,
    n904,
    n873
  );


  xnor
  g968
  (
    n983,
    n885,
    n878,
    n861,
    n868
  );


  xor
  g969
  (
    n987,
    n964,
    n922,
    n800,
    n801
  );


  nand
  g970
  (
    n1001,
    n798,
    n962,
    n950,
    n867
  );


  nand
  g971
  (
    n986,
    n883,
    n931,
    n957,
    n800
  );


  xor
  g972
  (
    n982,
    n799,
    n949,
    n969,
    n854
  );


  and
  g973
  (
    n1014,
    n798,
    n912,
    n801,
    n961
  );


  nand
  g974
  (
    n991,
    n973,
    n801,
    n884,
    n869
  );


  xor
  g975
  (
    n994,
    n958,
    n919,
    n925,
    n945
  );


  nand
  g976
  (
    n992,
    n799,
    n891,
    n894,
    n797
  );


  or
  g977
  (
    n1012,
    n898,
    n940,
    n972,
    n865
  );


  xnor
  g978
  (
    n988,
    n939,
    n944,
    n862,
    n978
  );


  xor
  g979
  (
    n981,
    n871,
    n916,
    n908,
    n797
  );


  nor
  g980
  (
    n1009,
    n890,
    n906,
    n974,
    n956
  );


  nand
  g981
  (
    n1005,
    n967,
    n953,
    n887,
    n921
  );


  nor
  g982
  (
    n984,
    n798,
    n903,
    n942,
    n858
  );


  or
  g983
  (
    n1013,
    n917,
    n864,
    n797,
    n900
  );


  nand
  g984
  (
    n1003,
    n960,
    n954,
    n800,
    n934
  );


  and
  g985
  (
    n989,
    n875,
    n924,
    n863,
    n923
  );


  nand
  g986
  (
    n1026,
    n1004,
    n1016,
    n807,
    n802
  );


  xor
  g987
  (
    n1019,
    n1013,
    n806,
    n1007,
    n1000
  );


  and
  g988
  (
    n1027,
    n802,
    n1008,
    n1017,
    n810
  );


  nand
  g989
  (
    n1028,
    n1001,
    n806,
    n805,
    n809
  );


  nor
  g990
  (
    n1022,
    n807,
    n1005,
    n1010,
    n805
  );


  nand
  g991
  (
    n1021,
    n803,
    n804,
    n808,
    n1002
  );


  xnor
  g992
  (
    n1031,
    n1009,
    n808,
    n999,
    n809
  );


  and
  g993
  (
    n1023,
    n1003,
    n810,
    n1018,
    n809
  );


  nand
  g994
  (
    n1030,
    n805,
    n804,
    n1015
  );


  xnor
  g995
  (
    n1032,
    n808,
    n803,
    n804
  );


  nor
  g996
  (
    n1024,
    n808,
    n809,
    n806,
    n802
  );


  nand
  g997
  (
    n1020,
    n806,
    n802,
    n810,
    n1012
  );


  xnor
  g998
  (
    n1025,
    n803,
    n1011,
    n807
  );


  nor
  g999
  (
    n1029,
    n1006,
    n1014,
    n805,
    n810
  );


  xor
  KeyGate_0_0
  (
    n965,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n708,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n932,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n729,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n525,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n713,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n78,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n192,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n663,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n186,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n219,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n877,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n879,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n260,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n258,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n84,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n467,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n811,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n155,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n169,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n640,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n881,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n451,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n527,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n337,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n785,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n376,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n650,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n687,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n225,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n791,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n849,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

