

module Stat_1418_20_7
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n1078,
  n1086,
  n1093,
  n1084,
  n1094,
  n1100,
  n1090,
  n1085,
  n1077,
  n1082,
  n1083,
  n1097,
  n1098,
  n1092,
  n1102,
  n1437,
  n1438,
  n1436,
  n1434,
  n1432,
  n1433,
  n1431,
  n1439,
  n1430,
  n1440,
  n1435,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1078;output n1086;output n1093;output n1084;output n1094;output n1100;output n1090;output n1085;output n1077;output n1082;output n1083;output n1097;output n1098;output n1092;output n1102;output n1437;output n1438;output n1436;output n1434;output n1432;output n1433;output n1431;output n1439;output n1430;output n1440;output n1435;
  wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1079;wire n1080;wire n1081;wire n1087;wire n1088;wire n1089;wire n1091;wire n1095;wire n1096;wire n1099;wire n1101;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  not
  g0
  (
    n108,
    n16
  );


  buf
  g1
  (
    n70,
    n22
  );


  buf
  g2
  (
    n45,
    n14
  );


  not
  g3
  (
    n105,
    n7
  );


  buf
  g4
  (
    n61,
    n13
  );


  buf
  g5
  (
    n39,
    n6
  );


  buf
  g6
  (
    n52,
    n13
  );


  buf
  g7
  (
    n42,
    n9
  );


  not
  g8
  (
    n91,
    n14
  );


  not
  g9
  (
    n76,
    n11
  );


  buf
  g10
  (
    n62,
    n21
  );


  not
  g11
  (
    n73,
    n2
  );


  not
  g12
  (
    n92,
    n1
  );


  not
  g13
  (
    n50,
    n18
  );


  buf
  g14
  (
    n85,
    n12
  );


  buf
  g15
  (
    n80,
    n13
  );


  buf
  g16
  (
    n43,
    n21
  );


  not
  g17
  (
    n98,
    n15
  );


  not
  g18
  (
    n109,
    n17
  );


  not
  g19
  (
    n82,
    n3
  );


  buf
  g20
  (
    n57,
    n7
  );


  buf
  g21
  (
    n44,
    n10
  );


  not
  g22
  (
    n32,
    n2
  );


  not
  g23
  (
    n65,
    n8
  );


  buf
  g24
  (
    KeyWire_0_24,
    n19
  );


  not
  g25
  (
    n75,
    n3
  );


  buf
  g26
  (
    n107,
    n14
  );


  buf
  g27
  (
    n31,
    n8
  );


  not
  g28
  (
    KeyWire_0_11,
    n17
  );


  buf
  g29
  (
    n100,
    n8
  );


  not
  g30
  (
    n63,
    n14
  );


  buf
  g31
  (
    n94,
    n11
  );


  not
  g32
  (
    n64,
    n10
  );


  buf
  g33
  (
    n104,
    n15
  );


  buf
  g34
  (
    n81,
    n19
  );


  not
  g35
  (
    n28,
    n11
  );


  not
  g36
  (
    KeyWire_0_14,
    n9
  );


  buf
  g37
  (
    n84,
    n20
  );


  buf
  g38
  (
    n25,
    n13
  );


  buf
  g39
  (
    n67,
    n2
  );


  not
  g40
  (
    n33,
    n20
  );


  not
  g41
  (
    n29,
    n17
  );


  buf
  g42
  (
    n38,
    n3
  );


  buf
  g43
  (
    n35,
    n22
  );


  buf
  g44
  (
    n97,
    n5
  );


  not
  g45
  (
    n78,
    n18
  );


  not
  g46
  (
    n27,
    n16
  );


  not
  g47
  (
    n54,
    n1
  );


  buf
  g48
  (
    n88,
    n4
  );


  buf
  g49
  (
    n77,
    n7
  );


  not
  g50
  (
    n110,
    n18
  );


  not
  g51
  (
    n46,
    n1
  );


  buf
  g52
  (
    n55,
    n10
  );


  buf
  g53
  (
    n51,
    n4
  );


  buf
  g54
  (
    n26,
    n8
  );


  buf
  g55
  (
    n106,
    n16
  );


  buf
  g56
  (
    n99,
    n3
  );


  buf
  g57
  (
    n53,
    n6
  );


  not
  g58
  (
    n30,
    n9
  );


  not
  g59
  (
    n59,
    n5
  );


  buf
  g60
  (
    n95,
    n5
  );


  not
  g61
  (
    n49,
    n18
  );


  buf
  g62
  (
    n60,
    n22
  );


  not
  g63
  (
    n23,
    n1
  );


  buf
  g64
  (
    n103,
    n19
  );


  buf
  g65
  (
    n66,
    n12
  );


  buf
  g66
  (
    n69,
    n9
  );


  not
  g67
  (
    n71,
    n6
  );


  buf
  g68
  (
    n47,
    n2
  );


  buf
  g69
  (
    n89,
    n12
  );


  buf
  g70
  (
    n79,
    n22
  );


  not
  g71
  (
    n24,
    n4
  );


  not
  g72
  (
    n58,
    n7
  );


  buf
  g73
  (
    n56,
    n12
  );


  not
  g74
  (
    n40,
    n19
  );


  buf
  g75
  (
    n37,
    n6
  );


  buf
  g76
  (
    n41,
    n17
  );


  not
  g77
  (
    n87,
    n11
  );


  buf
  g78
  (
    n90,
    n20
  );


  not
  g79
  (
    n102,
    n16
  );


  buf
  g80
  (
    n101,
    n20
  );


  buf
  g81
  (
    n48,
    n15
  );


  not
  g82
  (
    n72,
    n10
  );


  not
  g83
  (
    n93,
    n15
  );


  buf
  g84
  (
    n34,
    n4
  );


  not
  g85
  (
    n83,
    n21
  );


  buf
  g86
  (
    n86,
    n5
  );


  not
  g87
  (
    n68,
    n21
  );


  not
  g88
  (
    n260,
    n104
  );


  buf
  g89
  (
    n296,
    n35
  );


  buf
  g90
  (
    n428,
    n28
  );


  buf
  g91
  (
    n435,
    n88
  );


  buf
  g92
  (
    n249,
    n74
  );


  buf
  g93
  (
    n227,
    n102
  );


  not
  g94
  (
    n316,
    n36
  );


  buf
  g95
  (
    n379,
    n98
  );


  buf
  g96
  (
    n155,
    n71
  );


  not
  g97
  (
    n116,
    n41
  );


  buf
  g98
  (
    n186,
    n69
  );


  buf
  g99
  (
    n313,
    n59
  );


  buf
  g100
  (
    n262,
    n84
  );


  buf
  g101
  (
    n297,
    n29
  );


  not
  g102
  (
    n422,
    n47
  );


  buf
  g103
  (
    n354,
    n51
  );


  buf
  g104
  (
    n282,
    n29
  );


  not
  g105
  (
    n302,
    n91
  );


  not
  g106
  (
    n410,
    n73
  );


  buf
  g107
  (
    n138,
    n45
  );


  buf
  g108
  (
    n375,
    n25
  );


  buf
  g109
  (
    n277,
    n94
  );


  buf
  g110
  (
    n340,
    n28
  );


  buf
  g111
  (
    n373,
    n77
  );


  buf
  g112
  (
    n252,
    n85
  );


  not
  g113
  (
    n154,
    n108
  );


  buf
  g114
  (
    n188,
    n89
  );


  not
  g115
  (
    n216,
    n40
  );


  buf
  g116
  (
    n437,
    n71
  );


  buf
  g117
  (
    n221,
    n67
  );


  not
  g118
  (
    n180,
    n79
  );


  not
  g119
  (
    n268,
    n39
  );


  buf
  g120
  (
    KeyWire_0_29,
    n105
  );


  buf
  g121
  (
    n344,
    n62
  );


  not
  g122
  (
    n148,
    n60
  );


  not
  g123
  (
    n383,
    n107
  );


  not
  g124
  (
    n114,
    n94
  );


  not
  g125
  (
    n406,
    n48
  );


  buf
  g126
  (
    n125,
    n42
  );


  not
  g127
  (
    n184,
    n76
  );


  buf
  g128
  (
    n404,
    n89
  );


  buf
  g129
  (
    n234,
    n96
  );


  not
  g130
  (
    n285,
    n39
  );


  buf
  g131
  (
    n290,
    n85
  );


  not
  g132
  (
    n120,
    n78
  );


  buf
  g133
  (
    n195,
    n67
  );


  not
  g134
  (
    n300,
    n95
  );


  buf
  g135
  (
    n352,
    n98
  );


  buf
  g136
  (
    n309,
    n30
  );


  buf
  g137
  (
    n237,
    n86
  );


  not
  g138
  (
    n287,
    n49
  );


  buf
  g139
  (
    n112,
    n109
  );


  buf
  g140
  (
    n301,
    n103
  );


  not
  g141
  (
    n214,
    n70
  );


  not
  g142
  (
    n411,
    n61
  );


  not
  g143
  (
    n459,
    n27
  );


  not
  g144
  (
    n398,
    n81
  );


  not
  g145
  (
    n394,
    n88
  );


  not
  g146
  (
    n210,
    n27
  );


  not
  g147
  (
    n157,
    n92
  );


  buf
  g148
  (
    n205,
    n52
  );


  buf
  g149
  (
    n361,
    n92
  );


  not
  g150
  (
    n399,
    n65
  );


  buf
  g151
  (
    n130,
    n38
  );


  not
  g152
  (
    n265,
    n69
  );


  buf
  g153
  (
    n303,
    n104
  );


  not
  g154
  (
    n350,
    n31
  );


  buf
  g155
  (
    n259,
    n61
  );


  buf
  g156
  (
    n179,
    n109
  );


  buf
  g157
  (
    n289,
    n31
  );


  buf
  g158
  (
    n250,
    n50
  );


  buf
  g159
  (
    n450,
    n68
  );


  not
  g160
  (
    n161,
    n87
  );


  buf
  g161
  (
    n412,
    n32
  );


  buf
  g162
  (
    n246,
    n60
  );


  buf
  g163
  (
    n132,
    n44
  );


  not
  g164
  (
    n365,
    n100
  );


  buf
  g165
  (
    n390,
    n72
  );


  not
  g166
  (
    n315,
    n55
  );


  not
  g167
  (
    n229,
    n37
  );


  buf
  g168
  (
    n433,
    n45
  );


  not
  g169
  (
    n115,
    n83
  );


  buf
  g170
  (
    n167,
    n64
  );


  not
  g171
  (
    n121,
    n69
  );


  buf
  g172
  (
    n136,
    n25
  );


  buf
  g173
  (
    n454,
    n48
  );


  buf
  g174
  (
    n330,
    n90
  );


  buf
  g175
  (
    n335,
    n55
  );


  not
  g176
  (
    n141,
    n32
  );


  not
  g177
  (
    n322,
    n74
  );


  buf
  g178
  (
    n405,
    n79
  );


  buf
  g179
  (
    n152,
    n41
  );


  buf
  g180
  (
    n317,
    n42
  );


  not
  g181
  (
    n337,
    n37
  );


  buf
  g182
  (
    n181,
    n24
  );


  not
  g183
  (
    n407,
    n46
  );


  buf
  g184
  (
    n355,
    n63
  );


  not
  g185
  (
    n429,
    n95
  );


  buf
  g186
  (
    n182,
    n35
  );


  not
  g187
  (
    n423,
    n77
  );


  not
  g188
  (
    n360,
    n29
  );


  buf
  g189
  (
    n415,
    n38
  );


  buf
  g190
  (
    n147,
    n54
  );


  not
  g191
  (
    n291,
    n72
  );


  buf
  g192
  (
    n178,
    n23
  );


  not
  g193
  (
    n363,
    n89
  );


  not
  g194
  (
    n386,
    n61
  );


  buf
  g195
  (
    n253,
    n70
  );


  buf
  g196
  (
    KeyWire_0_18,
    n25
  );


  buf
  g197
  (
    n416,
    n110
  );


  buf
  g198
  (
    n206,
    n83
  );


  buf
  g199
  (
    n328,
    n56
  );


  buf
  g200
  (
    n408,
    n100
  );


  buf
  g201
  (
    KeyWire_0_23,
    n41
  );


  buf
  g202
  (
    n324,
    n99
  );


  buf
  g203
  (
    n164,
    n106
  );


  not
  g204
  (
    n308,
    n23
  );


  not
  g205
  (
    n175,
    n59
  );


  buf
  g206
  (
    n338,
    n57
  );


  buf
  g207
  (
    n424,
    n96
  );


  not
  g208
  (
    n312,
    n65
  );


  buf
  g209
  (
    n158,
    n78
  );


  not
  g210
  (
    KeyWire_0_25,
    n39
  );


  buf
  g211
  (
    n208,
    n26
  );


  not
  g212
  (
    n212,
    n82
  );


  not
  g213
  (
    n427,
    n79
  );


  buf
  g214
  (
    n370,
    n74
  );


  buf
  g215
  (
    n238,
    n97
  );


  not
  g216
  (
    n368,
    n75
  );


  not
  g217
  (
    n137,
    n57
  );


  buf
  g218
  (
    n134,
    n27
  );


  buf
  g219
  (
    n185,
    n48
  );


  not
  g220
  (
    n321,
    n99
  );


  not
  g221
  (
    n447,
    n45
  );


  buf
  g222
  (
    n430,
    n30
  );


  not
  g223
  (
    n357,
    n75
  );


  not
  g224
  (
    n451,
    n104
  );


  buf
  g225
  (
    n441,
    n26
  );


  not
  g226
  (
    n270,
    n47
  );


  buf
  g227
  (
    n209,
    n52
  );


  buf
  g228
  (
    n244,
    n33
  );


  buf
  g229
  (
    n233,
    n63
  );


  not
  g230
  (
    n353,
    n79
  );


  buf
  g231
  (
    n455,
    n84
  );


  not
  g232
  (
    n327,
    n53
  );


  not
  g233
  (
    n402,
    n44
  );


  not
  g234
  (
    n191,
    n100
  );


  buf
  g235
  (
    n444,
    n68
  );


  buf
  g236
  (
    n295,
    n49
  );


  buf
  g237
  (
    n286,
    n81
  );


  buf
  g238
  (
    n371,
    n48
  );


  not
  g239
  (
    n111,
    n95
  );


  buf
  g240
  (
    n333,
    n66
  );


  not
  g241
  (
    n162,
    n23
  );


  not
  g242
  (
    n393,
    n46
  );


  not
  g243
  (
    n272,
    n44
  );


  not
  g244
  (
    n425,
    n26
  );


  buf
  g245
  (
    KeyWire_0_16,
    n103
  );


  not
  g246
  (
    n248,
    n46
  );


  buf
  g247
  (
    n131,
    n69
  );


  buf
  g248
  (
    n264,
    n86
  );


  not
  g249
  (
    n204,
    n97
  );


  buf
  g250
  (
    n417,
    n96
  );


  not
  g251
  (
    n135,
    n93
  );


  buf
  g252
  (
    n160,
    n80
  );


  not
  g253
  (
    n426,
    n71
  );


  buf
  g254
  (
    n325,
    n83
  );


  not
  g255
  (
    n194,
    n107
  );


  buf
  g256
  (
    n456,
    n63
  );


  buf
  g257
  (
    n254,
    n40
  );


  buf
  g258
  (
    n156,
    n30
  );


  not
  g259
  (
    n163,
    n107
  );


  not
  g260
  (
    n359,
    n56
  );


  not
  g261
  (
    n172,
    n66
  );


  not
  g262
  (
    n224,
    n49
  );


  not
  g263
  (
    n391,
    n50
  );


  buf
  g264
  (
    n153,
    n86
  );


  not
  g265
  (
    n215,
    n51
  );


  buf
  g266
  (
    n228,
    n67
  );


  not
  g267
  (
    n366,
    n101
  );


  not
  g268
  (
    n192,
    n89
  );


  buf
  g269
  (
    n436,
    n88
  );


  not
  g270
  (
    n226,
    n97
  );


  not
  g271
  (
    n223,
    n53
  );


  not
  g272
  (
    n242,
    n59
  );


  buf
  g273
  (
    n241,
    n43
  );


  not
  g274
  (
    n124,
    n102
  );


  not
  g275
  (
    n122,
    n78
  );


  buf
  g276
  (
    n168,
    n95
  );


  buf
  g277
  (
    n171,
    n57
  );


  buf
  g278
  (
    n145,
    n49
  );


  buf
  g279
  (
    n293,
    n50
  );


  buf
  g280
  (
    n133,
    n58
  );


  buf
  g281
  (
    n142,
    n76
  );


  buf
  g282
  (
    n256,
    n45
  );


  not
  g283
  (
    n306,
    n90
  );


  buf
  g284
  (
    n385,
    n106
  );


  buf
  g285
  (
    n419,
    n55
  );


  not
  g286
  (
    n266,
    n97
  );


  not
  g287
  (
    n118,
    n26
  );


  not
  g288
  (
    n318,
    n39
  );


  buf
  g289
  (
    n140,
    n30
  );


  not
  g290
  (
    n183,
    n110
  );


  not
  g291
  (
    n358,
    n87
  );


  not
  g292
  (
    n255,
    n37
  );


  not
  g293
  (
    n413,
    n24
  );


  buf
  g294
  (
    n420,
    n28
  );


  not
  g295
  (
    n235,
    n82
  );


  not
  g296
  (
    n341,
    n33
  );


  not
  g297
  (
    n275,
    n40
  );


  not
  g298
  (
    n200,
    n23
  );


  buf
  g299
  (
    n173,
    n62
  );


  buf
  g300
  (
    n257,
    n64
  );


  buf
  g301
  (
    n174,
    n102
  );


  buf
  g302
  (
    n193,
    n81
  );


  not
  g303
  (
    n331,
    n43
  );


  not
  g304
  (
    n438,
    n107
  );


  not
  g305
  (
    n247,
    n93
  );


  not
  g306
  (
    n320,
    n29
  );


  buf
  g307
  (
    n431,
    n76
  );


  buf
  g308
  (
    n177,
    n77
  );


  buf
  g309
  (
    n263,
    n53
  );


  buf
  g310
  (
    n143,
    n31
  );


  buf
  g311
  (
    n284,
    n64
  );


  not
  g312
  (
    n146,
    n78
  );


  buf
  g313
  (
    n351,
    n58
  );


  buf
  g314
  (
    n139,
    n24
  );


  not
  g315
  (
    n288,
    n108
  );


  buf
  g316
  (
    n245,
    n35
  );


  not
  g317
  (
    n267,
    n75
  );


  not
  g318
  (
    n176,
    n72
  );


  not
  g319
  (
    n251,
    n72
  );


  buf
  g320
  (
    n240,
    n91
  );


  buf
  g321
  (
    n314,
    n27
  );


  buf
  g322
  (
    n243,
    n80
  );


  not
  g323
  (
    n332,
    n68
  );


  not
  g324
  (
    n144,
    n80
  );


  not
  g325
  (
    n149,
    n34
  );


  buf
  g326
  (
    n150,
    n62
  );


  buf
  g327
  (
    n117,
    n70
  );


  not
  g328
  (
    n461,
    n75
  );


  buf
  g329
  (
    n169,
    n42
  );


  buf
  g330
  (
    n273,
    n47
  );


  buf
  g331
  (
    n356,
    n33
  );


  not
  g332
  (
    n348,
    n105
  );


  buf
  g333
  (
    n392,
    n34
  );


  not
  g334
  (
    n281,
    n52
  );


  not
  g335
  (
    n376,
    n34
  );


  buf
  g336
  (
    n453,
    n62
  );


  not
  g337
  (
    n123,
    n54
  );


  buf
  g338
  (
    n190,
    n110
  );


  not
  g339
  (
    n443,
    n46
  );


  not
  g340
  (
    n346,
    n24
  );


  buf
  g341
  (
    n372,
    n56
  );


  buf
  g342
  (
    n377,
    n34
  );


  buf
  g343
  (
    n199,
    n94
  );


  not
  g344
  (
    n218,
    n93
  );


  not
  g345
  (
    n225,
    n33
  );


  not
  g346
  (
    n217,
    n32
  );


  not
  g347
  (
    n187,
    n84
  );


  not
  g348
  (
    n343,
    n108
  );


  not
  g349
  (
    n165,
    n61
  );


  not
  g350
  (
    n457,
    n82
  );


  buf
  g351
  (
    n445,
    n40
  );


  not
  g352
  (
    n271,
    n58
  );


  not
  g353
  (
    n311,
    n66
  );


  not
  g354
  (
    n403,
    n91
  );


  buf
  g355
  (
    n278,
    n44
  );


  buf
  g356
  (
    n369,
    n90
  );


  buf
  g357
  (
    n198,
    n38
  );


  buf
  g358
  (
    n170,
    n50
  );


  not
  g359
  (
    n239,
    n36
  );


  buf
  g360
  (
    n434,
    n42
  );


  buf
  g361
  (
    n397,
    n38
  );


  buf
  g362
  (
    n384,
    n68
  );


  not
  g363
  (
    n380,
    n54
  );


  not
  g364
  (
    n232,
    n106
  );


  buf
  g365
  (
    n400,
    n87
  );


  not
  g366
  (
    n283,
    n96
  );


  buf
  g367
  (
    n207,
    n82
  );


  buf
  g368
  (
    n261,
    n66
  );


  not
  g369
  (
    n258,
    n73
  );


  not
  g370
  (
    n448,
    n73
  );


  not
  g371
  (
    n307,
    n104
  );


  not
  g372
  (
    n294,
    n77
  );


  buf
  g373
  (
    n362,
    n101
  );


  buf
  g374
  (
    n202,
    n31
  );


  buf
  g375
  (
    n458,
    n109
  );


  buf
  g376
  (
    n166,
    n55
  );


  buf
  g377
  (
    n418,
    n100
  );


  not
  g378
  (
    n449,
    n28
  );


  not
  g379
  (
    n347,
    n59
  );


  buf
  g380
  (
    n128,
    n57
  );


  not
  g381
  (
    n439,
    n106
  );


  not
  g382
  (
    n339,
    n94
  );


  not
  g383
  (
    n336,
    n36
  );


  not
  g384
  (
    n440,
    n41
  );


  not
  g385
  (
    n421,
    n85
  );


  buf
  g386
  (
    n364,
    n60
  );


  buf
  g387
  (
    n279,
    n87
  );


  buf
  g388
  (
    n151,
    n51
  );


  buf
  g389
  (
    n329,
    n54
  );


  not
  g390
  (
    n276,
    n51
  );


  buf
  g391
  (
    n409,
    n37
  );


  buf
  g392
  (
    n432,
    n90
  );


  not
  g393
  (
    n345,
    n43
  );


  buf
  g394
  (
    n389,
    n74
  );


  not
  g395
  (
    n381,
    n67
  );


  not
  g396
  (
    n280,
    n80
  );


  not
  g397
  (
    n382,
    n98
  );


  not
  g398
  (
    n334,
    n101
  );


  not
  g399
  (
    n219,
    n105
  );


  not
  g400
  (
    n452,
    n103
  );


  not
  g401
  (
    n378,
    n99
  );


  buf
  g402
  (
    n396,
    n53
  );


  not
  g403
  (
    n213,
    n52
  );


  not
  g404
  (
    n310,
    n109
  );


  buf
  g405
  (
    n220,
    n88
  );


  not
  g406
  (
    n201,
    n93
  );


  not
  g407
  (
    n113,
    n91
  );


  buf
  g408
  (
    n203,
    n47
  );


  buf
  g409
  (
    n305,
    n99
  );


  buf
  g410
  (
    n401,
    n64
  );


  buf
  g411
  (
    n388,
    n92
  );


  buf
  g412
  (
    n374,
    n65
  );


  not
  g413
  (
    n236,
    n102
  );


  buf
  g414
  (
    n269,
    n84
  );


  not
  g415
  (
    n127,
    n60
  );


  buf
  g416
  (
    KeyWire_0_22,
    n86
  );


  buf
  g417
  (
    n189,
    n71
  );


  not
  g418
  (
    n460,
    n36
  );


  not
  g419
  (
    n323,
    n83
  );


  buf
  g420
  (
    n129,
    n85
  );


  not
  g421
  (
    n119,
    n76
  );


  not
  g422
  (
    n159,
    n25
  );


  not
  g423
  (
    n274,
    n43
  );


  buf
  g424
  (
    n319,
    n81
  );


  buf
  g425
  (
    n304,
    n73
  );


  buf
  g426
  (
    n230,
    n108
  );


  buf
  g427
  (
    n414,
    n56
  );


  not
  g428
  (
    n395,
    n32
  );


  buf
  g429
  (
    KeyWire_0_8,
    n35
  );


  not
  g430
  (
    n342,
    n63
  );


  not
  g431
  (
    n126,
    n58
  );


  not
  g432
  (
    n367,
    n70
  );


  not
  g433
  (
    n298,
    n105
  );


  buf
  g434
  (
    n231,
    n103
  );


  buf
  g435
  (
    n446,
    n98
  );


  buf
  g436
  (
    n387,
    n92
  );


  not
  g437
  (
    n442,
    n101
  );


  buf
  g438
  (
    n197,
    n65
  );


  not
  g439
  (
    n598,
    n266
  );


  buf
  g440
  (
    n679,
    n171
  );


  not
  g441
  (
    n652,
    n303
  );


  buf
  g442
  (
    n677,
    n305
  );


  not
  g443
  (
    n507,
    n273
  );


  not
  g444
  (
    n616,
    n309
  );


  buf
  g445
  (
    n551,
    n298
  );


  buf
  g446
  (
    n637,
    n239
  );


  not
  g447
  (
    n502,
    n116
  );


  not
  g448
  (
    n553,
    n121
  );


  not
  g449
  (
    n654,
    n179
  );


  not
  g450
  (
    n575,
    n304
  );


  not
  g451
  (
    n680,
    n259
  );


  buf
  g452
  (
    n512,
    n283
  );


  not
  g453
  (
    n538,
    n241
  );


  not
  g454
  (
    n481,
    n308
  );


  not
  g455
  (
    n664,
    n226
  );


  buf
  g456
  (
    n649,
    n172
  );


  not
  g457
  (
    n621,
    n210
  );


  buf
  g458
  (
    n479,
    n126
  );


  buf
  g459
  (
    n568,
    n305
  );


  not
  g460
  (
    n626,
    n189
  );


  not
  g461
  (
    n643,
    n304
  );


  not
  g462
  (
    n608,
    n134
  );


  buf
  g463
  (
    n625,
    n302
  );


  buf
  g464
  (
    n491,
    n136
  );


  buf
  g465
  (
    n501,
    n238
  );


  not
  g466
  (
    n676,
    n254
  );


  buf
  g467
  (
    KeyWire_0_0,
    n278
  );


  not
  g468
  (
    n647,
    n276
  );


  not
  g469
  (
    n498,
    n117
  );


  not
  g470
  (
    n511,
    n160
  );


  not
  g471
  (
    n651,
    n248
  );


  not
  g472
  (
    n504,
    n289
  );


  buf
  g473
  (
    n650,
    n234
  );


  not
  g474
  (
    n539,
    n308
  );


  not
  g475
  (
    n686,
    n143
  );


  not
  g476
  (
    n547,
    n240
  );


  buf
  g477
  (
    n544,
    n274
  );


  not
  g478
  (
    n674,
    n178
  );


  not
  g479
  (
    n632,
    n304
  );


  buf
  g480
  (
    n478,
    n242
  );


  not
  g481
  (
    n603,
    n146
  );


  not
  g482
  (
    n659,
    n300
  );


  buf
  g483
  (
    n573,
    n236
  );


  not
  g484
  (
    n618,
    n142
  );


  not
  g485
  (
    n584,
    n193
  );


  buf
  g486
  (
    n559,
    n137
  );


  buf
  g487
  (
    n462,
    n258
  );


  buf
  g488
  (
    n525,
    n295
  );


  not
  g489
  (
    n582,
    n293
  );


  not
  g490
  (
    n658,
    n145
  );


  not
  g491
  (
    n648,
    n263
  );


  buf
  g492
  (
    n609,
    n191
  );


  buf
  g493
  (
    n488,
    n199
  );


  not
  g494
  (
    n635,
    n112
  );


  not
  g495
  (
    n593,
    n118
  );


  not
  g496
  (
    n600,
    n224
  );


  buf
  g497
  (
    n683,
    n164
  );


  not
  g498
  (
    n569,
    n201
  );


  buf
  g499
  (
    n612,
    n214
  );


  not
  g500
  (
    n587,
    n306
  );


  buf
  g501
  (
    n503,
    n209
  );


  buf
  g502
  (
    n610,
    n268
  );


  buf
  g503
  (
    n644,
    n279
  );


  buf
  g504
  (
    n537,
    n129
  );


  buf
  g505
  (
    n601,
    n187
  );


  not
  g506
  (
    n566,
    n275
  );


  not
  g507
  (
    n510,
    n155
  );


  not
  g508
  (
    n556,
    n267
  );


  not
  g509
  (
    n528,
    n290
  );


  buf
  g510
  (
    n552,
    n183
  );


  not
  g511
  (
    n665,
    n288
  );


  buf
  g512
  (
    n662,
    n200
  );


  buf
  g513
  (
    n661,
    n271
  );


  buf
  g514
  (
    n567,
    n131
  );


  buf
  g515
  (
    n524,
    n249
  );


  not
  g516
  (
    n561,
    n303
  );


  not
  g517
  (
    n639,
    n303
  );


  not
  g518
  (
    n594,
    n272
  );


  buf
  g519
  (
    n536,
    n301
  );


  buf
  g520
  (
    n578,
    n153
  );


  buf
  g521
  (
    n619,
    n281
  );


  buf
  g522
  (
    KeyWire_0_10,
    n166
  );


  buf
  g523
  (
    n611,
    n237
  );


  buf
  g524
  (
    n638,
    n301
  );


  buf
  g525
  (
    n627,
    n306
  );


  not
  g526
  (
    n579,
    n150
  );


  not
  g527
  (
    n576,
    n173
  );


  not
  g528
  (
    n490,
    n306
  );


  buf
  g529
  (
    n673,
    n132
  );


  buf
  g530
  (
    n565,
    n264
  );


  not
  g531
  (
    n549,
    n211
  );


  buf
  g532
  (
    n470,
    n205
  );


  buf
  g533
  (
    n597,
    n308
  );


  not
  g534
  (
    n669,
    n207
  );


  buf
  g535
  (
    n520,
    n141
  );


  not
  g536
  (
    n666,
    n144
  );


  buf
  g537
  (
    n614,
    n303
  );


  not
  g538
  (
    n499,
    n128
  );


  buf
  g539
  (
    n489,
    n310
  );


  not
  g540
  (
    n533,
    n270
  );


  buf
  g541
  (
    n555,
    n218
  );


  not
  g542
  (
    n472,
    n251
  );


  buf
  g543
  (
    n596,
    n244
  );


  not
  g544
  (
    n592,
    n265
  );


  buf
  g545
  (
    n495,
    n232
  );


  not
  g546
  (
    n487,
    n161
  );


  buf
  g547
  (
    n623,
    n125
  );


  not
  g548
  (
    n494,
    n309
  );


  buf
  g549
  (
    n517,
    n188
  );


  not
  g550
  (
    n480,
    n194
  );


  buf
  g551
  (
    n467,
    n147
  );


  not
  g552
  (
    n475,
    n302
  );


  buf
  g553
  (
    n492,
    n149
  );


  buf
  g554
  (
    n497,
    n250
  );


  buf
  g555
  (
    n667,
    n185
  );


  buf
  g556
  (
    n585,
    n235
  );


  buf
  g557
  (
    n513,
    n306
  );


  buf
  g558
  (
    n469,
    n152
  );


  buf
  g559
  (
    n515,
    n287
  );


  buf
  g560
  (
    n531,
    n308
  );


  not
  g561
  (
    n684,
    n307
  );


  not
  g562
  (
    n506,
    n260
  );


  buf
  g563
  (
    n484,
    n158
  );


  not
  g564
  (
    n562,
    n301
  );


  buf
  g565
  (
    n532,
    n135
  );


  not
  g566
  (
    n671,
    n307
  );


  not
  g567
  (
    n570,
    n123
  );


  not
  g568
  (
    n595,
    n156
  );


  not
  g569
  (
    n586,
    n309
  );


  not
  g570
  (
    n633,
    n213
  );


  buf
  g571
  (
    n500,
    n177
  );


  not
  g572
  (
    n529,
    n124
  );


  not
  g573
  (
    n670,
    n122
  );


  not
  g574
  (
    n526,
    n269
  );


  not
  g575
  (
    n571,
    n151
  );


  buf
  g576
  (
    n485,
    n190
  );


  buf
  g577
  (
    n599,
    n277
  );


  not
  g578
  (
    n505,
    n162
  );


  buf
  g579
  (
    n523,
    n140
  );


  not
  g580
  (
    n477,
    n302
  );


  not
  g581
  (
    n535,
    n202
  );


  buf
  g582
  (
    n657,
    n222
  );


  not
  g583
  (
    n646,
    n133
  );


  buf
  g584
  (
    n534,
    n198
  );


  buf
  g585
  (
    n624,
    n299
  );


  not
  g586
  (
    n678,
    n216
  );


  buf
  g587
  (
    n486,
    n301
  );


  buf
  g588
  (
    n688,
    n294
  );


  buf
  g589
  (
    n493,
    n247
  );


  buf
  g590
  (
    n685,
    n223
  );


  buf
  g591
  (
    n605,
    n119
  );


  not
  g592
  (
    n617,
    n181
  );


  buf
  g593
  (
    n508,
    n252
  );


  not
  g594
  (
    n496,
    n196
  );


  not
  g595
  (
    n629,
    n163
  );


  not
  g596
  (
    n604,
    n286
  );


  buf
  g597
  (
    n518,
    n195
  );


  buf
  g598
  (
    n516,
    n233
  );


  not
  g599
  (
    n687,
    n253
  );


  not
  g600
  (
    n540,
    n212
  );


  buf
  g601
  (
    n548,
    n206
  );


  not
  g602
  (
    n542,
    n231
  );


  not
  g603
  (
    n473,
    n292
  );


  buf
  g604
  (
    n642,
    n115
  );


  not
  g605
  (
    n620,
    n245
  );


  not
  g606
  (
    n602,
    n217
  );


  buf
  g607
  (
    n466,
    n176
  );


  not
  g608
  (
    n591,
    n215
  );


  buf
  g609
  (
    n563,
    n175
  );


  buf
  g610
  (
    n580,
    n229
  );


  not
  g611
  (
    n645,
    n257
  );


  not
  g612
  (
    n519,
    n309
  );


  buf
  g613
  (
    n546,
    n227
  );


  not
  g614
  (
    n514,
    n221
  );


  not
  g615
  (
    n572,
    n307
  );


  buf
  g616
  (
    n672,
    n304
  );


  not
  g617
  (
    n636,
    n159
  );


  buf
  g618
  (
    n550,
    n282
  );


  buf
  g619
  (
    n588,
    n130
  );


  not
  g620
  (
    n465,
    n262
  );


  not
  g621
  (
    n630,
    n139
  );


  not
  g622
  (
    n606,
    n170
  );


  buf
  g623
  (
    n628,
    n280
  );


  buf
  g624
  (
    n583,
    n148
  );


  buf
  g625
  (
    n530,
    n208
  );


  not
  g626
  (
    n468,
    n261
  );


  buf
  g627
  (
    n681,
    n256
  );


  not
  g628
  (
    n541,
    n243
  );


  not
  g629
  (
    n545,
    n174
  );


  buf
  g630
  (
    n589,
    n220
  );


  not
  g631
  (
    n613,
    n228
  );


  buf
  g632
  (
    n682,
    n255
  );


  not
  g633
  (
    n675,
    n284
  );


  buf
  g634
  (
    n483,
    n169
  );


  buf
  g635
  (
    n476,
    n120
  );


  buf
  g636
  (
    n631,
    n285
  );


  buf
  g637
  (
    n464,
    n165
  );


  buf
  g638
  (
    n660,
    n305
  );


  buf
  g639
  (
    n554,
    n291
  );


  not
  g640
  (
    n474,
    n184
  );


  buf
  g641
  (
    n560,
    n230
  );


  not
  g642
  (
    n482,
    n114
  );


  not
  g643
  (
    n463,
    n186
  );


  not
  g644
  (
    n640,
    n168
  );


  buf
  g645
  (
    n527,
    n157
  );


  buf
  g646
  (
    n521,
    n182
  );


  not
  g647
  (
    n634,
    n138
  );


  not
  g648
  (
    n641,
    n127
  );


  buf
  g649
  (
    n622,
    n305
  );


  buf
  g650
  (
    n577,
    n307
  );


  not
  g651
  (
    n615,
    n219
  );


  buf
  g652
  (
    n656,
    n113
  );


  buf
  g653
  (
    n663,
    n180
  );


  not
  g654
  (
    n543,
    n297
  );


  buf
  g655
  (
    n509,
    n225
  );


  buf
  g656
  (
    n607,
    n192
  );


  not
  g657
  (
    n590,
    n111
  );


  buf
  g658
  (
    n581,
    n167
  );


  not
  g659
  (
    n653,
    n246
  );


  buf
  g660
  (
    n522,
    n302
  );


  buf
  g661
  (
    n557,
    n203
  );


  buf
  g662
  (
    n668,
    n204
  );


  buf
  g663
  (
    n558,
    n296
  );


  buf
  g664
  (
    n564,
    n154
  );


  buf
  g665
  (
    n574,
    n197
  );


  buf
  g666
  (
    n792,
    n326
  );


  not
  g667
  (
    n830,
    n351
  );


  buf
  g668
  (
    n711,
    n418
  );


  buf
  g669
  (
    n796,
    n537
  );


  not
  g670
  (
    n915,
    n398
  );


  buf
  g671
  (
    n811,
    n367
  );


  not
  g672
  (
    n759,
    n506
  );


  buf
  g673
  (
    n767,
    n312
  );


  buf
  g674
  (
    n754,
    n672
  );


  buf
  g675
  (
    n896,
    n441
  );


  buf
  g676
  (
    n746,
    n658
  );


  not
  g677
  (
    n847,
    n389
  );


  not
  g678
  (
    n698,
    n670
  );


  buf
  g679
  (
    n901,
    n667
  );


  not
  g680
  (
    n813,
    n353
  );


  not
  g681
  (
    n757,
    n376
  );


  not
  g682
  (
    n783,
    n374
  );


  buf
  g683
  (
    n713,
    n420
  );


  not
  g684
  (
    n881,
    n626
  );


  buf
  g685
  (
    n867,
    n431
  );


  buf
  g686
  (
    n753,
    n406
  );


  buf
  g687
  (
    n823,
    n379
  );


  not
  g688
  (
    n793,
    n591
  );


  not
  g689
  (
    n821,
    n392
  );


  buf
  g690
  (
    n787,
    n504
  );


  not
  g691
  (
    n727,
    n656
  );


  not
  g692
  (
    n869,
    n358
  );


  buf
  g693
  (
    n814,
    n328
  );


  xor
  g694
  (
    n911,
    n315,
    n542,
    n330,
    n454
  );


  and
  g695
  (
    n890,
    n675,
    n391,
    n530,
    n384
  );


  nor
  g696
  (
    n897,
    n434,
    n456,
    n440,
    n580
  );


  or
  g697
  (
    n872,
    n313,
    n435,
    n367,
    n453
  );


  xor
  g698
  (
    n837,
    n436,
    n374,
    n543,
    n437
  );


  nor
  g699
  (
    n702,
    n549,
    n337,
    n323,
    n356
  );


  xnor
  g700
  (
    n747,
    n635,
    n368,
    n401,
    n311
  );


  xnor
  g701
  (
    n817,
    n377,
    n638,
    n592,
    n349
  );


  or
  g702
  (
    n729,
    n510,
    n380,
    n342,
    n374
  );


  nand
  g703
  (
    n889,
    n450,
    n470,
    n383,
    n358
  );


  xnor
  g704
  (
    n871,
    n360,
    n419,
    n583,
    n413
  );


  nor
  g705
  (
    n894,
    n674,
    n401,
    n482,
    n567
  );


  or
  g706
  (
    n850,
    n643,
    n370,
    n476,
    n339
  );


  nand
  g707
  (
    n689,
    n333,
    n314,
    n324,
    n418
  );


  and
  g708
  (
    n775,
    n336,
    n405,
    n411,
    n483
  );


  nor
  g709
  (
    n806,
    n429,
    n312,
    n598,
    n632
  );


  or
  g710
  (
    n697,
    n317,
    n326,
    n528,
    n402
  );


  nand
  g711
  (
    n732,
    n351,
    n361,
    n341,
    n415
  );


  nand
  g712
  (
    n790,
    n376,
    n436,
    n664,
    n321
  );


  or
  g713
  (
    n726,
    n573,
    n399,
    n320,
    n343
  );


  and
  g714
  (
    n777,
    n392,
    n408,
    n641,
    n317
  );


  nor
  g715
  (
    n733,
    n408,
    n366,
    n686,
    n487
  );


  xor
  g716
  (
    n725,
    n331,
    n435,
    n557,
    n475
  );


  xor
  g717
  (
    n844,
    n366,
    n360,
    n443,
    n399
  );


  xor
  g718
  (
    n825,
    n352,
    n350,
    n415,
    n341
  );


  or
  g719
  (
    n887,
    n380,
    n509,
    n423,
    n644
  );


  and
  g720
  (
    n720,
    n391,
    n360,
    n439,
    n324
  );


  xnor
  g721
  (
    n780,
    n665,
    n428,
    n421,
    n616
  );


  xnor
  g722
  (
    n898,
    n605,
    n383,
    n458,
    n593
  );


  nand
  g723
  (
    n849,
    n347,
    n396,
    n516,
    n441
  );


  or
  g724
  (
    n841,
    n442,
    n467,
    n431,
    n333
  );


  or
  g725
  (
    n853,
    n417,
    n320,
    n325,
    n333
  );


  nand
  g726
  (
    n734,
    n427,
    n453,
    n400,
    n342
  );


  and
  g727
  (
    n838,
    n391,
    n522,
    n333,
    n400
  );


  xor
  g728
  (
    n724,
    n397,
    n365,
    n325,
    n421
  );


  xnor
  g729
  (
    n808,
    n451,
    n519,
    n579,
    n413
  );


  xnor
  g730
  (
    n828,
    n513,
    n428,
    n624,
    n455
  );


  nor
  g731
  (
    n905,
    n599,
    n421,
    n451,
    n463
  );


  or
  g732
  (
    n750,
    n415,
    n359,
    n340,
    n363
  );


  xnor
  g733
  (
    n886,
    n338,
    n640,
    n399,
    n477
  );


  nor
  g734
  (
    n778,
    n436,
    n369,
    n408,
    n327
  );


  nand
  g735
  (
    n851,
    n559,
    n410,
    n457,
    n326
  );


  nand
  g736
  (
    n876,
    n319,
    n582,
    n401,
    n322
  );


  xor
  g737
  (
    n818,
    n314,
    n442,
    n405,
    n359
  );


  xor
  g738
  (
    n820,
    n687,
    n390,
    n423,
    n468
  );


  nor
  g739
  (
    n760,
    n349,
    n316,
    n562,
    n437
  );


  xor
  g740
  (
    n840,
    n551,
    n393,
    n688,
    n439
  );


  xnor
  g741
  (
    n743,
    n310,
    n320,
    n404,
    n386
  );


  xor
  g742
  (
    n895,
    n359,
    n571,
    n452,
    n622
  );


  nand
  g743
  (
    n706,
    n311,
    n429,
    n419,
    n609
  );


  or
  g744
  (
    n888,
    n430,
    n338,
    n343,
    n404
  );


  nor
  g745
  (
    n832,
    n322,
    n405,
    n437,
    n382
  );


  or
  g746
  (
    n799,
    n630,
    n347,
    n446,
    n329
  );


  xnor
  g747
  (
    n755,
    n385,
    n402,
    n341,
    n382
  );


  nor
  g748
  (
    n913,
    n532,
    n427,
    n425,
    n454
  );


  nand
  g749
  (
    n701,
    n363,
    n435,
    n348,
    n422
  );


  xor
  g750
  (
    n858,
    n459,
    n438,
    n385,
    n362
  );


  nand
  g751
  (
    n776,
    n390,
    n350,
    n392,
    n485
  );


  and
  g752
  (
    n892,
    n651,
    n566,
    n451,
    n316
  );


  xnor
  g753
  (
    n865,
    n327,
    n448,
    n364,
    n393
  );


  nand
  g754
  (
    n846,
    n389,
    n355,
    n331,
    n455
  );


  nor
  g755
  (
    n914,
    n535,
    n449,
    n395,
    n390
  );


  or
  g756
  (
    n810,
    n472,
    n337,
    n494,
    n335
  );


  and
  g757
  (
    n705,
    n444,
    n621,
    n445,
    n488
  );


  or
  g758
  (
    n722,
    n634,
    n422,
    n354,
    n484
  );


  or
  g759
  (
    n904,
    n378,
    n331,
    n367,
    n332
  );


  xor
  g760
  (
    KeyWire_0_31,
    n409,
    n397,
    n661,
    n348
  );


  or
  g761
  (
    n795,
    n403,
    n443,
    n569,
    n427
  );


  and
  g762
  (
    n805,
    n335,
    n338,
    n330,
    n497
  );


  xnor
  g763
  (
    n740,
    n332,
    n360,
    n432,
    n318
  );


  or
  g764
  (
    n856,
    n449,
    n384,
    n353,
    n540
  );


  xor
  g765
  (
    KeyWire_0_1,
    n657,
    n427,
    n402,
    n453
  );


  nor
  g766
  (
    n848,
    n368,
    n413,
    n419,
    n439
  );


  xnor
  g767
  (
    n879,
    n429,
    n379,
    n412,
    n618
  );


  or
  g768
  (
    n883,
    n366,
    n346,
    n683,
    n432
  );


  nand
  g769
  (
    n715,
    n319,
    n575,
    n343,
    n310
  );


  nor
  g770
  (
    n824,
    n684,
    n348,
    n328,
    n386
  );


  xor
  g771
  (
    n692,
    n385,
    n404,
    n548,
    n681
  );


  nor
  g772
  (
    n700,
    n589,
    n363,
    n455,
    n620
  );


  or
  g773
  (
    n798,
    n404,
    n433,
    n357,
    n523
  );


  xnor
  g774
  (
    n762,
    n409,
    n492,
    n387,
    n346
  );


  xor
  g775
  (
    n903,
    n442,
    n420,
    n449,
    n388
  );


  and
  g776
  (
    n773,
    n321,
    n319,
    n560,
    n358
  );


  xor
  g777
  (
    n693,
    n402,
    n358,
    n682,
    n478
  );


  xor
  g778
  (
    n863,
    n405,
    n373,
    n323,
    n495
  );


  nand
  g779
  (
    n708,
    n446,
    n376,
    n334,
    n493
  );


  xnor
  g780
  (
    n696,
    n403,
    n508,
    n520,
    n426
  );


  or
  g781
  (
    n855,
    n446,
    n411,
    n365,
    n355
  );


  and
  g782
  (
    n721,
    n546,
    n371,
    n434,
    n329
  );


  and
  g783
  (
    n730,
    n444,
    n637,
    n671,
    n474
  );


  or
  g784
  (
    n906,
    n411,
    n652,
    n456,
    n349
  );


  nor
  g785
  (
    n728,
    n323,
    n454,
    n437,
    n505
  );


  xnor
  g786
  (
    n826,
    n525,
    n486,
    n357,
    n344
  );


  and
  g787
  (
    n745,
    n394,
    n576,
    n550,
    n568
  );


  or
  g788
  (
    n902,
    n314,
    n448,
    n668,
    n545
  );


  nand
  g789
  (
    n770,
    n660,
    n355,
    n447
  );


  and
  g790
  (
    n699,
    n443,
    n373,
    n361,
    n318
  );


  nor
  g791
  (
    n839,
    n396,
    n450,
    n327,
    n393
  );


  or
  g792
  (
    n822,
    n373,
    n450,
    n429,
    n334
  );


  xnor
  g793
  (
    n766,
    n320,
    n480,
    n453,
    n603
  );


  and
  g794
  (
    n694,
    n388,
    n334,
    n666,
    n353
  );


  and
  g795
  (
    n878,
    n447,
    n471,
    n459,
    n511
  );


  nand
  g796
  (
    n860,
    n597,
    n438,
    n655,
    n389
  );


  xnor
  g797
  (
    n816,
    n629,
    n538,
    n678,
    n627
  );


  nor
  g798
  (
    n809,
    n534,
    n636,
    n401,
    n362
  );


  xor
  g799
  (
    n854,
    n452,
    n313,
    n574,
    n418
  );


  nor
  g800
  (
    n739,
    n364,
    n444,
    n544,
    n585
  );


  and
  g801
  (
    n802,
    n398,
    n324,
    n369,
    n395
  );


  and
  g802
  (
    n714,
    n410,
    n679,
    n380,
    n312
  );


  or
  g803
  (
    n842,
    n558,
    n334,
    n440,
    n387
  );


  nor
  g804
  (
    n803,
    n426,
    n406,
    n445,
    n412
  );


  or
  g805
  (
    n800,
    n431,
    n369,
    n628
  );


  nand
  g806
  (
    n899,
    n378,
    n663,
    n372,
    n473
  );


  or
  g807
  (
    n752,
    n377,
    n531,
    n433,
    n399
  );


  nand
  g808
  (
    n771,
    n327,
    n385,
    n527,
    n348
  );


  nor
  g809
  (
    n829,
    n422,
    n336,
    n365,
    n368
  );


  xor
  g810
  (
    n703,
    n409,
    n337,
    n659,
    n368
  );


  or
  g811
  (
    n744,
    n447,
    n438,
    n642,
    n425
  );


  xnor
  g812
  (
    n831,
    n586,
    n349,
    n356,
    n411
  );


  nand
  g813
  (
    n884,
    n449,
    n373,
    n445,
    n396
  );


  nand
  g814
  (
    n815,
    n500,
    n418,
    n415,
    n324
  );


  or
  g815
  (
    n900,
    n514,
    n342,
    n353,
    n371
  );


  and
  g816
  (
    n742,
    n466,
    n469,
    n419,
    n326
  );


  and
  g817
  (
    n845,
    n345,
    n365,
    n340,
    n454
  );


  nor
  g818
  (
    n834,
    n413,
    n455,
    n361,
    n395
  );


  or
  g819
  (
    n882,
    n370,
    n452,
    n318,
    n328
  );


  nand
  g820
  (
    n710,
    n383,
    n412,
    n451,
    n491
  );


  and
  g821
  (
    n786,
    n332,
    n341,
    n403,
    n501
  );


  and
  g822
  (
    n748,
    n397,
    n388,
    n430,
    n371
  );


  or
  g823
  (
    n717,
    n645,
    n375,
    n613,
    n343
  );


  nor
  g824
  (
    n735,
    n370,
    n383,
    n595,
    n615
  );


  nand
  g825
  (
    n704,
    n336,
    n524,
    n315,
    n377
  );


  xor
  g826
  (
    n875,
    n489,
    n392,
    n515,
    n350
  );


  nor
  g827
  (
    n764,
    n417,
    n465,
    n600,
    n434
  );


  nand
  g828
  (
    n893,
    n394,
    n325,
    n444,
    n424
  );


  and
  g829
  (
    n794,
    n521,
    n650,
    n414,
    n379
  );


  nand
  g830
  (
    n835,
    n347,
    n325,
    n499,
    n407
  );


  nand
  g831
  (
    n857,
    n336,
    n364,
    n381,
    n445
  );


  nand
  g832
  (
    n709,
    n344,
    n347,
    n464,
    n371
  );


  or
  g833
  (
    n765,
    n356,
    n443,
    n502,
    n416
  );


  nand
  g834
  (
    n859,
    n315,
    n602,
    n625,
    n572
  );


  and
  g835
  (
    n772,
    n375,
    n408,
    n361,
    n457
  );


  or
  g836
  (
    n723,
    n407,
    n553,
    n352,
    n311
  );


  and
  g837
  (
    KeyWire_0_19,
    n381,
    n457,
    n581,
    n417
  );


  xor
  g838
  (
    n877,
    n354,
    n498,
    n555,
    n536
  );


  and
  g839
  (
    n738,
    n339,
    n565,
    n400,
    n496
  );


  xor
  g840
  (
    n789,
    n462,
    n346,
    n379,
    n344
  );


  xor
  g841
  (
    n862,
    n398,
    n458,
    n351,
    n321
  );


  and
  g842
  (
    KeyWire_0_20,
    n458,
    n518,
    n362,
    n601
  );


  and
  g843
  (
    n864,
    n676,
    n421,
    n623,
    n430
  );


  xor
  g844
  (
    n833,
    n319,
    n503,
    n375,
    n388
  );


  nand
  g845
  (
    n782,
    n362,
    n317,
    n619,
    n407
  );


  nor
  g846
  (
    n836,
    n434,
    n446,
    n669,
    n414
  );


  nand
  g847
  (
    n874,
    n617,
    n315,
    n612,
    n323
  );


  and
  g848
  (
    n804,
    n344,
    n570,
    n375,
    n337
  );


  xnor
  g849
  (
    n866,
    n438,
    n584,
    n386,
    n590
  );


  or
  g850
  (
    n763,
    n431,
    n578,
    n430,
    n512
  );


  and
  g851
  (
    n880,
    n387,
    n436,
    n539,
    n350
  );


  nor
  g852
  (
    n768,
    n352,
    n410,
    n456,
    n382
  );


  xor
  g853
  (
    n741,
    n440,
    n357,
    n312,
    n450
  );


  nand
  g854
  (
    n797,
    n420,
    n552,
    n554,
    n354
  );


  nand
  g855
  (
    n819,
    n441,
    n340,
    n414,
    n396
  );


  nand
  g856
  (
    n719,
    n377,
    n587,
    n614,
    n447
  );


  nor
  g857
  (
    n784,
    n416,
    n439,
    n406,
    n435
  );


  nand
  g858
  (
    n873,
    n677,
    n314,
    n342,
    n384
  );


  nand
  g859
  (
    n807,
    n577,
    n441,
    n529,
    n346
  );


  nor
  g860
  (
    n785,
    n378,
    n376,
    n328,
    n425
  );


  nor
  g861
  (
    n716,
    n490,
    n653,
    n372,
    n556
  );


  nor
  g862
  (
    n812,
    n685,
    n345,
    n400,
    n680
  );


  and
  g863
  (
    n791,
    n330,
    n426,
    n424,
    n367
  );


  and
  g864
  (
    n736,
    n384,
    n479,
    n426,
    n448
  );


  or
  g865
  (
    n827,
    n673,
    n452,
    n433,
    n422
  );


  xnor
  g866
  (
    n907,
    n372,
    n316,
    n359
  );


  xnor
  g867
  (
    n909,
    n394,
    n423,
    n313,
    n481
  );


  or
  g868
  (
    n910,
    n561,
    n338,
    n647,
    n432
  );


  nor
  g869
  (
    n868,
    n607,
    n395,
    n517,
    n335
  );


  xor
  g870
  (
    n718,
    n381,
    n352,
    n370,
    n389
  );


  xor
  g871
  (
    n769,
    n397,
    n594,
    n433,
    n564
  );


  nand
  g872
  (
    n756,
    n596,
    n608,
    n423,
    n380
  );


  and
  g873
  (
    n852,
    n381,
    n414,
    n507,
    n403
  );


  or
  g874
  (
    n749,
    n588,
    n331,
    n416,
    n339
  );


  xor
  g875
  (
    n712,
    n428,
    n364,
    n340,
    n322
  );


  nand
  g876
  (
    n801,
    n372,
    n412,
    n356,
    n526
  );


  or
  g877
  (
    n731,
    n391,
    n533,
    n424,
    n606
  );


  and
  g878
  (
    n788,
    n332,
    n410,
    n646,
    n633
  );


  and
  g879
  (
    n690,
    n351,
    n407,
    n424,
    n398
  );


  and
  g880
  (
    n761,
    n610,
    n335,
    n310,
    n648
  );


  nor
  g881
  (
    n861,
    n363,
    n457,
    n313,
    n639
  );


  and
  g882
  (
    n908,
    n631,
    n357,
    n382,
    n345
  );


  or
  g883
  (
    n912,
    n649,
    n440,
    n425,
    n322
  );


  xor
  g884
  (
    n870,
    n386,
    n420,
    n654,
    n378
  );


  or
  g885
  (
    KeyWire_0_26,
    n374,
    n458,
    n329,
    n321
  );


  and
  g886
  (
    n691,
    n366,
    n406,
    n611,
    n390
  );


  and
  g887
  (
    n779,
    n604,
    n456,
    n416,
    n387
  );


  nand
  g888
  (
    n781,
    n417,
    n428,
    n547,
    n339
  );


  and
  g889
  (
    n885,
    n318,
    n563,
    n432,
    n311
  );


  xor
  g890
  (
    n695,
    n317,
    n354,
    n394,
    n393
  );


  nor
  g891
  (
    n843,
    n409,
    n442,
    n329,
    n448
  );


  nor
  g892
  (
    n737,
    n662,
    n330,
    n541,
    n345
  );


  not
  g893
  (
    n926,
    n736
  );


  buf
  g894
  (
    n956,
    n717
  );


  buf
  g895
  (
    n955,
    n701
  );


  not
  g896
  (
    n934,
    n728
  );


  buf
  g897
  (
    n924,
    n713
  );


  not
  g898
  (
    n948,
    n711
  );


  not
  g899
  (
    n957,
    n729
  );


  buf
  g900
  (
    n932,
    n725
  );


  not
  g901
  (
    n949,
    n726
  );


  not
  g902
  (
    n921,
    n710
  );


  not
  g903
  (
    n927,
    n699
  );


  buf
  g904
  (
    n916,
    n706
  );


  buf
  g905
  (
    n963,
    n722
  );


  buf
  g906
  (
    KeyWire_0_13,
    n727
  );


  not
  g907
  (
    n958,
    n707
  );


  not
  g908
  (
    n945,
    n689
  );


  not
  g909
  (
    n935,
    n695
  );


  buf
  g910
  (
    n938,
    n698
  );


  buf
  g911
  (
    n961,
    n716
  );


  not
  g912
  (
    n918,
    n712
  );


  buf
  g913
  (
    n952,
    n721
  );


  buf
  g914
  (
    n937,
    n715
  );


  buf
  g915
  (
    n923,
    n708
  );


  buf
  g916
  (
    n939,
    n714
  );


  not
  g917
  (
    n936,
    n718
  );


  buf
  g918
  (
    n922,
    n700
  );


  buf
  g919
  (
    n942,
    n735
  );


  buf
  g920
  (
    n931,
    n692
  );


  buf
  g921
  (
    n925,
    n733
  );


  buf
  g922
  (
    n960,
    n734
  );


  not
  g923
  (
    n941,
    n719
  );


  buf
  g924
  (
    n947,
    n704
  );


  not
  g925
  (
    n940,
    n691
  );


  not
  g926
  (
    n943,
    n690
  );


  buf
  g927
  (
    n944,
    n724
  );


  buf
  g928
  (
    n920,
    n705
  );


  buf
  g929
  (
    n919,
    n732
  );


  not
  g930
  (
    n933,
    n731
  );


  buf
  g931
  (
    n953,
    n720
  );


  not
  g932
  (
    n951,
    n723
  );


  buf
  g933
  (
    n959,
    n702
  );


  buf
  g934
  (
    n962,
    n694
  );


  buf
  g935
  (
    n930,
    n730
  );


  not
  g936
  (
    n917,
    n703
  );


  not
  g937
  (
    KeyWire_0_28,
    n709
  );


  buf
  g938
  (
    n954,
    n693
  );


  buf
  g939
  (
    n928,
    n696
  );


  buf
  g940
  (
    n929,
    n697
  );


  xor
  g941
  (
    n987,
    n935,
    n815,
    n888,
    n937
  );


  xnor
  g942
  (
    n1011,
    n774,
    n921,
    n954,
    n956
  );


  xor
  g943
  (
    n1004,
    n782,
    n945,
    n738,
    n802
  );


  and
  g944
  (
    n976,
    n811,
    n862,
    n765,
    n885
  );


  nand
  g945
  (
    n1014,
    n833,
    n956,
    n742,
    n883
  );


  xor
  g946
  (
    n966,
    n805,
    n796,
    n804,
    n852
  );


  or
  g947
  (
    n1010,
    n841,
    n944,
    n939,
    n828
  );


  and
  g948
  (
    n981,
    n927,
    n770,
    n757,
    n956
  );


  nor
  g949
  (
    n965,
    n918,
    n885,
    n743,
    n949
  );


  and
  g950
  (
    n984,
    n791,
    n955,
    n838,
    n831
  );


  or
  g951
  (
    n975,
    n834,
    n764,
    n807,
    n888
  );


  xnor
  g952
  (
    n1001,
    n950,
    n957,
    n809,
    n775
  );


  xor
  g953
  (
    n986,
    n753,
    n865,
    n746,
    n823
  );


  or
  g954
  (
    n1016,
    n830,
    n957,
    n812,
    n760
  );


  and
  g955
  (
    n992,
    n886,
    n886,
    n759,
    n845
  );


  xor
  g956
  (
    n977,
    n886,
    n855,
    n744,
    n943
  );


  and
  g957
  (
    n967,
    n869,
    n763,
    n955,
    n924
  );


  nand
  g958
  (
    n998,
    n922,
    n884,
    n822,
    n938
  );


  xnor
  g959
  (
    n1013,
    n793,
    n837,
    n884,
    n936
  );


  nor
  g960
  (
    n1015,
    n767,
    n946,
    n850,
    n889
  );


  xor
  g961
  (
    n1007,
    n954,
    n952,
    n790,
    n955
  );


  xnor
  g962
  (
    n983,
    n788,
    n758,
    n947,
    n861
  );


  nor
  g963
  (
    n1021,
    n930,
    n826,
    n776,
    n777
  );


  or
  g964
  (
    n988,
    n801,
    n890,
    n747
  );


  xor
  g965
  (
    n1002,
    n925,
    n883,
    n794,
    n931
  );


  nand
  g966
  (
    n1022,
    n737,
    n885,
    n799,
    n958
  );


  xnor
  g967
  (
    n969,
    n878,
    n783,
    n940,
    n749
  );


  nand
  g968
  (
    n985,
    n929,
    n917,
    n870,
    n853
  );


  nor
  g969
  (
    n980,
    n785,
    n761,
    n919,
    n741
  );


  xor
  g970
  (
    n990,
    n820,
    n884,
    n882,
    n923
  );


  nand
  g971
  (
    n1008,
    n880,
    n818,
    n840,
    n886
  );


  and
  g972
  (
    n994,
    n768,
    n863,
    n795,
    n856
  );


  nand
  g973
  (
    n999,
    n867,
    n866,
    n854,
    n953
  );


  nand
  g974
  (
    n1006,
    n932,
    n772,
    n887,
    n958
  );


  and
  g975
  (
    n978,
    n808,
    n844,
    n800,
    n824
  );


  and
  g976
  (
    n1009,
    n848,
    n843,
    n885,
    n928
  );


  and
  g977
  (
    n1017,
    n819,
    n745,
    n916,
    n871
  );


  nor
  g978
  (
    n991,
    n889,
    n792,
    n881,
    n814
  );


  xor
  g979
  (
    n972,
    n882,
    n873,
    n836,
    n780
  );


  nand
  g980
  (
    n1023,
    n889,
    n784,
    n817,
    n920
  );


  xnor
  g981
  (
    n974,
    n951,
    n797,
    n948,
    n779
  );


  xor
  g982
  (
    n1020,
    n957,
    n857,
    n890,
    n874
  );


  nand
  g983
  (
    n1005,
    n887,
    n813,
    n953,
    n789
  );


  or
  g984
  (
    n1003,
    n882,
    n891,
    n750,
    n835
  );


  nor
  g985
  (
    n997,
    n879,
    n875,
    n756,
    n957
  );


  xor
  g986
  (
    n970,
    n762,
    n958,
    n887,
    n888
  );


  xor
  g987
  (
    n964,
    n890,
    n955,
    n851,
    n849
  );


  nand
  g988
  (
    n1024,
    n806,
    n810,
    n872,
    n883
  );


  and
  g989
  (
    n1012,
    n769,
    n821,
    n942,
    n787
  );


  nor
  g990
  (
    n982,
    n748,
    n781,
    n934,
    n755
  );


  or
  g991
  (
    n989,
    n827,
    n952,
    n887,
    n739
  );


  xnor
  g992
  (
    n1018,
    n846,
    n868,
    n839,
    n891
  );


  xor
  g993
  (
    n1000,
    n803,
    n754,
    n954,
    n859
  );


  xor
  g994
  (
    n979,
    n766,
    n926,
    n864,
    n959
  );


  nor
  g995
  (
    n973,
    n778,
    n740,
    n825,
    n954
  );


  nor
  g996
  (
    n971,
    n847,
    n798,
    n842,
    n786
  );


  nand
  g997
  (
    n968,
    n773,
    n882,
    n883,
    n771
  );


  nand
  g998
  (
    n993,
    n933,
    n889,
    n876,
    n752
  );


  xnor
  g999
  (
    n1019,
    n860,
    n884,
    n751,
    n958
  );


  or
  g1000
  (
    n996,
    n858,
    n888,
    n816,
    n956
  );


  nand
  g1001
  (
    n995,
    n829,
    n832,
    n941,
    n877
  );


  not
  g1002
  (
    n1047,
    n998
  );


  not
  g1003
  (
    n1041,
    n1000
  );


  not
  g1004
  (
    n1068,
    n976
  );


  not
  g1005
  (
    KeyWire_0_2,
    n989
  );


  not
  g1006
  (
    n1066,
    n1002
  );


  not
  g1007
  (
    n1051,
    n996
  );


  buf
  g1008
  (
    n1030,
    n973
  );


  not
  g1009
  (
    n1045,
    n1004
  );


  buf
  g1010
  (
    n1059,
    n1009
  );


  not
  g1011
  (
    n1054,
    n970
  );


  not
  g1012
  (
    n1040,
    n977
  );


  not
  g1013
  (
    n1050,
    n995
  );


  not
  g1014
  (
    n1056,
    n994
  );


  buf
  g1015
  (
    n1026,
    n981
  );


  buf
  g1016
  (
    n1067,
    n1001
  );


  buf
  g1017
  (
    n1058,
    n991
  );


  buf
  g1018
  (
    n1029,
    n986
  );


  buf
  g1019
  (
    n1069,
    n980
  );


  not
  g1020
  (
    n1027,
    n982
  );


  not
  g1021
  (
    n1064,
    n984
  );


  not
  g1022
  (
    n1034,
    n967
  );


  buf
  g1023
  (
    n1046,
    n972
  );


  buf
  g1024
  (
    n1033,
    n979
  );


  not
  g1025
  (
    n1031,
    n964
  );


  not
  g1026
  (
    n1049,
    n987
  );


  buf
  g1027
  (
    n1025,
    n983
  );


  buf
  g1028
  (
    n1055,
    n965
  );


  buf
  g1029
  (
    n1032,
    n1007
  );


  buf
  g1030
  (
    n1043,
    n974
  );


  buf
  g1031
  (
    n1048,
    n969
  );


  not
  g1032
  (
    n1060,
    n1003
  );


  buf
  g1033
  (
    n1070,
    n971
  );


  not
  g1034
  (
    KeyWire_0_4,
    n988
  );


  not
  g1035
  (
    n1063,
    n1006
  );


  buf
  g1036
  (
    n1061,
    n999
  );


  buf
  g1037
  (
    n1035,
    n993
  );


  not
  g1038
  (
    n1044,
    n975
  );


  not
  g1039
  (
    n1057,
    n990
  );


  buf
  g1040
  (
    n1038,
    n1008
  );


  buf
  g1041
  (
    n1037,
    n1005
  );


  buf
  g1042
  (
    n1042,
    n997
  );


  buf
  g1043
  (
    n1036,
    n985
  );


  not
  g1044
  (
    n1065,
    n992
  );


  not
  g1045
  (
    n1062,
    n966
  );


  not
  g1046
  (
    n1028,
    n968
  );


  buf
  g1047
  (
    n1039,
    n978
  );


  xor
  g1048
  (
    n1090,
    n1056,
    n1024,
    n1057,
    n899
  );


  xor
  g1049
  (
    n1073,
    n1030,
    n896,
    n1020,
    n1043
  );


  and
  g1050
  (
    n1083,
    n1023,
    n1054,
    n1015,
    n1039
  );


  nor
  g1051
  (
    n1080,
    n897,
    n895,
    n893,
    n1055
  );


  or
  g1052
  (
    n1099,
    n897,
    n1052,
    n892,
    n895
  );


  xnor
  g1053
  (
    n1077,
    n1047,
    n1056,
    n893,
    n1032
  );


  or
  g1054
  (
    n1092,
    n900,
    n902,
    n893,
    n894
  );


  nor
  g1055
  (
    n1100,
    n893,
    n1012,
    n896,
    n1055
  );


  xnor
  g1056
  (
    n1097,
    n898,
    n1057,
    n1010,
    n905
  );


  nand
  g1057
  (
    n1095,
    n901,
    n904,
    n1021,
    n1049
  );


  and
  g1058
  (
    n1087,
    n1055,
    n902,
    n904
  );


  and
  g1059
  (
    n1076,
    n904,
    n900,
    n1048,
    n905
  );


  and
  g1060
  (
    n1098,
    n1056,
    n899,
    n1044,
    n898
  );


  nor
  g1061
  (
    n1082,
    n1054,
    n1054,
    n894,
    n896
  );


  and
  g1062
  (
    n1096,
    n1050,
    n1057,
    n1033,
    n897
  );


  or
  g1063
  (
    n1086,
    n1038,
    n1041,
    n1026,
    n903
  );


  xnor
  g1064
  (
    n1071,
    n900,
    n900,
    n1042,
    n894
  );


  nor
  g1065
  (
    n1088,
    n897,
    n892,
    n901,
    n1057
  );


  xor
  g1066
  (
    n1091,
    n1017,
    n1025,
    n1056,
    n891
  );


  xnor
  g1067
  (
    n1081,
    n903,
    n1011,
    n1013,
    n895
  );


  xnor
  g1068
  (
    n1084,
    n1022,
    n1019,
    n906,
    n1045
  );


  xor
  g1069
  (
    n1089,
    n891,
    n902,
    n904,
    n1054
  );


  and
  g1070
  (
    n1094,
    n905,
    n895,
    n1036,
    n1040
  );


  xnor
  g1071
  (
    n1072,
    n903,
    n1016,
    n905,
    n1034
  );


  and
  g1072
  (
    n1093,
    n892,
    n1035,
    n1031,
    n1037
  );


  xor
  g1073
  (
    n1075,
    n892,
    n901,
    n899,
    n898
  );


  nor
  g1074
  (
    n1079,
    n1028,
    n899,
    n1051,
    n898
  );


  nor
  g1075
  (
    n1078,
    n1029,
    n896,
    n1053
  );


  xnor
  g1076
  (
    n1085,
    n1055,
    n903,
    n901,
    n1014
  );


  or
  g1077
  (
    n1074,
    n1018,
    n894,
    n1027,
    n1046
  );


  buf
  g1078
  (
    n1102,
    n1088
  );


  buf
  g1079
  (
    n1104,
    n1087
  );


  buf
  g1080
  (
    n1101,
    n1086
  );


  not
  g1081
  (
    n1103,
    n1085
  );


  and
  g1082
  (
    n1106,
    n1104,
    n1059
  );


  nor
  g1083
  (
    n1105,
    n1059,
    n1058,
    n1102
  );


  or
  g1084
  (
    n1107,
    n1060,
    n1103,
    n1058
  );


  buf
  g1085
  (
    n1119,
    n1107
  );


  buf
  g1086
  (
    n1109,
    n1107
  );


  not
  g1087
  (
    n1113,
    n1105
  );


  not
  g1088
  (
    n1118,
    n1106
  );


  not
  g1089
  (
    n1111,
    n1107
  );


  buf
  g1090
  (
    n1108,
    n1107
  );


  not
  g1091
  (
    n1112,
    n1106
  );


  buf
  g1092
  (
    n1114,
    n1105
  );


  buf
  g1093
  (
    n1117,
    n1106
  );


  buf
  g1094
  (
    n1110,
    n1105
  );


  not
  g1095
  (
    n1115,
    n1105
  );


  not
  g1096
  (
    n1116,
    n1106
  );


  not
  g1097
  (
    n1146,
    n960
  );


  not
  g1098
  (
    n1153,
    n1119
  );


  not
  g1099
  (
    n1134,
    n908
  );


  not
  g1100
  (
    n1162,
    n910
  );


  not
  g1101
  (
    n1136,
    n960
  );


  not
  g1102
  (
    n1138,
    n909
  );


  buf
  g1103
  (
    n1148,
    n959
  );


  buf
  g1104
  (
    n1130,
    n1089
  );


  not
  g1105
  (
    n1147,
    n459
  );


  not
  g1106
  (
    n1143,
    n1100
  );


  buf
  g1107
  (
    n1127,
    n910
  );


  buf
  g1108
  (
    KeyWire_0_5,
    n1114
  );


  buf
  g1109
  (
    n1126,
    n906
  );


  buf
  g1110
  (
    n1137,
    n962
  );


  not
  g1111
  (
    n1150,
    n961
  );


  buf
  g1112
  (
    n1140,
    n1117
  );


  buf
  g1113
  (
    n1128,
    n963
  );


  buf
  g1114
  (
    n1167,
    n1108
  );


  not
  g1115
  (
    n1166,
    n1115
  );


  not
  g1116
  (
    n1149,
    n1111
  );


  buf
  g1117
  (
    n1129,
    n959
  );


  buf
  g1118
  (
    n1156,
    n1090
  );


  buf
  g1119
  (
    n1142,
    n962
  );


  buf
  g1120
  (
    n1159,
    n907
  );


  not
  g1121
  (
    n1155,
    n910
  );


  not
  g1122
  (
    n1122,
    n1112
  );


  not
  g1123
  (
    n1152,
    n1108
  );


  not
  g1124
  (
    n1139,
    n1060
  );


  and
  g1125
  (
    n1135,
    n1099,
    n1119,
    n1112,
    n908
  );


  and
  g1126
  (
    n1163,
    n1097,
    n906,
    n1114,
    n1118
  );


  xnor
  g1127
  (
    n1157,
    n1117,
    n1098,
    n908
  );


  nand
  g1128
  (
    n1141,
    n959,
    n1116,
    n963,
    n1109
  );


  and
  g1129
  (
    n1121,
    n1061,
    n909,
    n1118,
    n1108
  );


  xnor
  g1130
  (
    n1124,
    n1117,
    n907,
    n962,
    n1115
  );


  xnor
  g1131
  (
    n1120,
    n1113,
    n1115,
    n1112,
    n1118
  );


  xnor
  g1132
  (
    n1144,
    n1113,
    n1108,
    n910,
    n960
  );


  or
  g1133
  (
    n1158,
    n1094,
    n907,
    n961,
    n962
  );


  and
  g1134
  (
    n1154,
    n1092,
    n1110,
    n1119,
    n1061
  );


  or
  g1135
  (
    n1131,
    n1110,
    n907,
    n1116,
    n963
  );


  or
  g1136
  (
    n1165,
    n1093,
    n1114,
    n960,
    n1061
  );


  or
  g1137
  (
    n1145,
    n1116,
    n1109,
    n1060,
    n909
  );


  or
  g1138
  (
    n1132,
    n911,
    n1110,
    n963
  );


  and
  g1139
  (
    n1151,
    n1115,
    n1111,
    n1117,
    n1060
  );


  and
  g1140
  (
    n1161,
    n1095,
    n961,
    n1061,
    n1109
  );


  nand
  g1141
  (
    n1164,
    n1118,
    n1109,
    n1112,
    n1114
  );


  and
  g1142
  (
    n1160,
    n1111,
    n961,
    n1113,
    n906
  );


  xnor
  g1143
  (
    n1133,
    n1096,
    n1111,
    n1116,
    n1119
  );


  or
  g1144
  (
    n1123,
    n1113,
    n909,
    n1091,
    n1062
  );


  not
  g1145
  (
    n1203,
    n1130
  );


  buf
  g1146
  (
    n1177,
    n1137
  );


  buf
  g1147
  (
    n1199,
    n1128
  );


  not
  g1148
  (
    n1196,
    n1126
  );


  buf
  g1149
  (
    n1198,
    n1135
  );


  buf
  g1150
  (
    n1179,
    n1133
  );


  buf
  g1151
  (
    n1180,
    n1124
  );


  not
  g1152
  (
    n1168,
    n1131
  );


  not
  g1153
  (
    n1184,
    n1136
  );


  buf
  g1154
  (
    n1175,
    n1124
  );


  buf
  g1155
  (
    n1204,
    n1132
  );


  buf
  g1156
  (
    n1185,
    n1139
  );


  buf
  g1157
  (
    n1189,
    n1137
  );


  not
  g1158
  (
    n1169,
    n1130
  );


  not
  g1159
  (
    n1172,
    n1134
  );


  not
  g1160
  (
    n1192,
    n1138
  );


  not
  g1161
  (
    n1170,
    n1122
  );


  buf
  g1162
  (
    n1183,
    n1125
  );


  buf
  g1163
  (
    n1182,
    n1123
  );


  not
  g1164
  (
    n1202,
    n1120
  );


  buf
  g1165
  (
    n1187,
    n1139
  );


  buf
  g1166
  (
    n1171,
    n1122
  );


  buf
  g1167
  (
    n1195,
    n1133
  );


  not
  g1168
  (
    n1201,
    n1121
  );


  buf
  g1169
  (
    n1174,
    n1125
  );


  not
  g1170
  (
    n1205,
    n1136
  );


  not
  g1171
  (
    n1173,
    n1129
  );


  not
  g1172
  (
    n1176,
    n1120
  );


  not
  g1173
  (
    n1197,
    n1132
  );


  not
  g1174
  (
    n1193,
    n1128
  );


  not
  g1175
  (
    n1181,
    n1126
  );


  not
  g1176
  (
    n1190,
    n1134
  );


  not
  g1177
  (
    n1191,
    n1131
  );


  buf
  g1178
  (
    n1207,
    n1127
  );


  buf
  g1179
  (
    n1186,
    n1135
  );


  buf
  g1180
  (
    n1206,
    n1129
  );


  buf
  g1181
  (
    n1194,
    n1121
  );


  not
  g1182
  (
    n1188,
    n1123
  );


  buf
  g1183
  (
    n1178,
    n1127
  );


  not
  g1184
  (
    n1200,
    n1138
  );


  buf
  g1185
  (
    n1220,
    n1201
  );


  buf
  g1186
  (
    n1213,
    n1195
  );


  buf
  g1187
  (
    n1284,
    n1062
  );


  buf
  g1188
  (
    n1242,
    n1198
  );


  buf
  g1189
  (
    n1250,
    n1199
  );


  not
  g1190
  (
    n1239,
    n1189
  );


  not
  g1191
  (
    n1280,
    n1141
  );


  buf
  g1192
  (
    n1278,
    n1195
  );


  buf
  g1193
  (
    n1266,
    n1198
  );


  buf
  g1194
  (
    n1238,
    n1194
  );


  buf
  g1195
  (
    n1210,
    n1170
  );


  buf
  g1196
  (
    n1215,
    n1193
  );


  buf
  g1197
  (
    n1232,
    n1143
  );


  buf
  g1198
  (
    n1246,
    n1062
  );


  not
  g1199
  (
    n1268,
    n1200
  );


  buf
  g1200
  (
    n1241,
    n1197
  );


  buf
  g1201
  (
    n1245,
    n1187
  );


  not
  g1202
  (
    n1271,
    n1185
  );


  not
  g1203
  (
    n1287,
    n1145
  );


  not
  g1204
  (
    n1282,
    n1207
  );


  not
  g1205
  (
    n1216,
    n1178
  );


  not
  g1206
  (
    n1249,
    n1141
  );


  buf
  g1207
  (
    n1217,
    n1199
  );


  buf
  g1208
  (
    n1262,
    n1188
  );


  not
  g1209
  (
    n1222,
    n1199
  );


  not
  g1210
  (
    n1214,
    n1196
  );


  not
  g1211
  (
    n1209,
    n1144
  );


  not
  g1212
  (
    n1251,
    n1179
  );


  buf
  g1213
  (
    n1256,
    n1203
  );


  not
  g1214
  (
    n1265,
    n1207
  );


  buf
  g1215
  (
    n1261,
    n1196
  );


  not
  g1216
  (
    n1258,
    n1205
  );


  not
  g1217
  (
    n1229,
    n1206
  );


  not
  g1218
  (
    n1237,
    n1190
  );


  not
  g1219
  (
    n1263,
    n1147
  );


  not
  g1220
  (
    n1286,
    n1203
  );


  not
  g1221
  (
    n1235,
    n1063
  );


  buf
  g1222
  (
    n1219,
    n1197
  );


  not
  g1223
  (
    n1226,
    n1196
  );


  buf
  g1224
  (
    n1281,
    n1181
  );


  buf
  g1225
  (
    n1211,
    n1201
  );


  buf
  g1226
  (
    n1255,
    n1146
  );


  buf
  g1227
  (
    n1269,
    n1182
  );


  not
  g1228
  (
    n1236,
    n1194
  );


  buf
  g1229
  (
    n1274,
    n1204
  );


  not
  g1230
  (
    n1253,
    n1140
  );


  buf
  g1231
  (
    n1252,
    n1062
  );


  not
  g1232
  (
    n1264,
    n1196
  );


  buf
  g1233
  (
    n1277,
    n1207
  );


  buf
  g1234
  (
    n1254,
    n1173
  );


  buf
  g1235
  (
    n1260,
    n1204
  );


  not
  g1236
  (
    n1234,
    n1186
  );


  not
  g1237
  (
    n1212,
    n1204
  );


  not
  g1238
  (
    n1224,
    n1198
  );


  not
  g1239
  (
    n1218,
    n1204
  );


  buf
  g1240
  (
    n1270,
    n1202
  );


  buf
  g1241
  (
    n1227,
    n1147
  );


  not
  g1242
  (
    n1208,
    n1142
  );


  not
  g1243
  (
    n1240,
    n1140
  );


  not
  g1244
  (
    n1273,
    n1202
  );


  not
  g1245
  (
    n1285,
    n1191
  );


  not
  g1246
  (
    n1233,
    n1168
  );


  not
  g1247
  (
    n1221,
    n1148
  );


  not
  g1248
  (
    n1257,
    n1201
  );


  not
  g1249
  (
    n1267,
    n1195
  );


  buf
  g1250
  (
    n1275,
    n1143
  );


  buf
  g1251
  (
    n1244,
    n1144
  );


  not
  g1252
  (
    n1276,
    n1180
  );


  buf
  g1253
  (
    n1279,
    n1197
  );


  xnor
  g1254
  (
    n1228,
    n1174,
    n1169,
    n1146
  );


  xnor
  g1255
  (
    n1230,
    n1203,
    n1206,
    n1195
  );


  and
  g1256
  (
    n1272,
    n1197,
    n1206,
    n1205
  );


  and
  g1257
  (
    n1247,
    n1205,
    n1200
  );


  or
  g1258
  (
    n1283,
    n1148,
    n1142,
    n1206
  );


  xor
  g1259
  (
    n1259,
    n1192,
    n1199,
    n1176
  );


  nand
  g1260
  (
    n1248,
    n1203,
    n1201,
    n1202
  );


  nand
  g1261
  (
    KeyWire_0_27,
    n1145,
    n1207,
    n1171
  );


  nor
  g1262
  (
    n1243,
    n1177,
    n1172,
    n1175
  );


  xnor
  g1263
  (
    n1223,
    n1200,
    n1184,
    n1183
  );


  and
  g1264
  (
    n1231,
    n1205,
    n1198,
    n1202
  );


  not
  g1265
  (
    n1317,
    n1151
  );


  buf
  g1266
  (
    n1308,
    n460
  );


  buf
  g1267
  (
    n1319,
    n1154
  );


  not
  g1268
  (
    n1290,
    n461
  );


  buf
  g1269
  (
    n1309,
    n1157
  );


  buf
  g1270
  (
    n1310,
    n1212
  );


  not
  g1271
  (
    n1320,
    n1222
  );


  buf
  g1272
  (
    n1323,
    n1221
  );


  not
  g1273
  (
    n1307,
    n461
  );


  buf
  g1274
  (
    n1322,
    n1156
  );


  buf
  g1275
  (
    n1306,
    n1226
  );


  buf
  g1276
  (
    n1295,
    n1223
  );


  buf
  g1277
  (
    n1291,
    n1238
  );


  buf
  g1278
  (
    n1299,
    n1219
  );


  not
  g1279
  (
    n1298,
    n1153
  );


  buf
  g1280
  (
    n1300,
    n1240
  );


  buf
  g1281
  (
    n1315,
    n1218
  );


  buf
  g1282
  (
    n1297,
    n1244
  );


  buf
  g1283
  (
    n1293,
    n1217
  );


  not
  g1284
  (
    n1305,
    n1227
  );


  not
  g1285
  (
    n1303,
    n1233
  );


  not
  g1286
  (
    n1301,
    n1156
  );


  not
  g1287
  (
    n1294,
    n1243
  );


  buf
  g1288
  (
    n1316,
    n1209
  );


  not
  g1289
  (
    n1288,
    n460
  );


  not
  g1290
  (
    KeyWire_0_17,
    n1242
  );


  buf
  g1291
  (
    n1302,
    n461
  );


  not
  g1292
  (
    KeyWire_0_7,
    n1150
  );


  xor
  g1293
  (
    n1292,
    n1224,
    n1155,
    n459,
    n1236
  );


  and
  g1294
  (
    n1296,
    n1228,
    n1232,
    n1154,
    n1241
  );


  xnor
  g1295
  (
    n1304,
    n1225,
    n1208,
    n1149,
    n1155
  );


  and
  g1296
  (
    n1324,
    n1149,
    n1230,
    n1152
  );


  and
  g1297
  (
    n1313,
    n1150,
    n1214,
    n1151,
    n1210
  );


  xor
  g1298
  (
    n1312,
    n1153,
    n461,
    n1239,
    n1237
  );


  xor
  g1299
  (
    n1321,
    n1220,
    n460,
    n1229,
    n1213
  );


  xor
  g1300
  (
    n1314,
    n1234,
    n1215,
    n460,
    n1231
  );


  nor
  g1301
  (
    n1318,
    n1216,
    n1157,
    n1211,
    n1235
  );


  not
  g1302
  (
    n1337,
    n1285
  );


  not
  g1303
  (
    n1361,
    n1292
  );


  buf
  g1304
  (
    n1362,
    n1324
  );


  not
  g1305
  (
    n1330,
    n1272
  );


  not
  g1306
  (
    n1334,
    n1253
  );


  not
  g1307
  (
    n1350,
    n1255
  );


  buf
  g1308
  (
    n1332,
    n1314
  );


  buf
  g1309
  (
    n1352,
    n1278
  );


  not
  g1310
  (
    n1329,
    n1310
  );


  not
  g1311
  (
    n1358,
    n1271
  );


  not
  g1312
  (
    n1342,
    n1300
  );


  not
  g1313
  (
    n1343,
    n1066
  );


  buf
  g1314
  (
    n1360,
    n1267
  );


  buf
  g1315
  (
    n1344,
    n1259
  );


  buf
  g1316
  (
    KeyWire_0_9,
    n1251
  );


  buf
  g1317
  (
    n1356,
    n1276
  );


  buf
  g1318
  (
    KeyWire_0_30,
    n1063
  );


  nand
  g1319
  (
    n1348,
    n1067,
    n1067,
    n1295,
    n1268
  );


  and
  g1320
  (
    n1339,
    n1293,
    n1282,
    n1321,
    n1068
  );


  and
  g1321
  (
    n1359,
    n1065,
    n1317,
    n1064
  );


  xnor
  g1322
  (
    KeyWire_0_15,
    n1280,
    n1065,
    n1290,
    n1298
  );


  xor
  g1323
  (
    n1345,
    n1262,
    n1065,
    n1312,
    n1301
  );


  nand
  g1324
  (
    n1355,
    n1319,
    n1297,
    n1281,
    n1273
  );


  or
  g1325
  (
    n1338,
    n1286,
    n1279,
    n1302,
    n1263
  );


  or
  g1326
  (
    KeyWire_0_6,
    n1320,
    n1266,
    n1260,
    n1274
  );


  nand
  g1327
  (
    n1349,
    n1064,
    n1063,
    n1287,
    n1066
  );


  nor
  g1328
  (
    n1354,
    n1275,
    n1323,
    n1289,
    n1256
  );


  xnor
  g1329
  (
    n1353,
    n1258,
    n1306,
    n1318,
    n1309
  );


  nor
  g1330
  (
    n1328,
    n1247,
    n1063,
    n1265,
    n1249
  );


  nand
  g1331
  (
    n1357,
    n1252,
    n1303,
    n1313,
    n1264
  );


  nand
  g1332
  (
    n1335,
    n1299,
    n1322,
    n1245,
    n1316
  );


  and
  g1333
  (
    n1340,
    n1311,
    n1284,
    n1248,
    n1277
  );


  and
  g1334
  (
    n1326,
    n1254,
    n1250,
    n1294,
    n1066
  );


  xor
  g1335
  (
    n1341,
    n1257,
    n1304,
    n1246,
    n1324
  );


  or
  g1336
  (
    KeyWire_0_21,
    n1305,
    n1270,
    n1288,
    n1269
  );


  and
  g1337
  (
    n1331,
    n1261,
    n1308,
    n1283,
    n1067
  );


  nor
  g1338
  (
    n1336,
    n1067,
    n1291,
    n1066,
    n1315
  );


  nand
  g1339
  (
    KeyWire_0_3,
    n1296,
    n1065,
    n1064,
    n1307
  );


  buf
  g1340
  (
    n1367,
    n1328
  );


  not
  g1341
  (
    n1363,
    n1328
  );


  not
  g1342
  (
    n1364,
    n1327
  );


  not
  g1343
  (
    n1368,
    n1325
  );


  not
  g1344
  (
    n1366,
    n1329
  );


  buf
  g1345
  (
    n1365,
    n1326
  );


  buf
  g1346
  (
    n1371,
    n1338
  );


  buf
  g1347
  (
    n1382,
    n913
  );


  nor
  g1348
  (
    n1377,
    n913,
    n1068
  );


  nand
  g1349
  (
    n1375,
    n1367,
    n1337,
    n1333,
    n914
  );


  nand
  g1350
  (
    n1373,
    n1368,
    n1331,
    n1329,
    n911
  );


  or
  g1351
  (
    n1372,
    n1338,
    n1339,
    n1365,
    n1336
  );


  or
  g1352
  (
    n1384,
    n1367,
    n915,
    n912
  );


  nand
  g1353
  (
    n1376,
    n911,
    n911,
    n1368,
    n1366
  );


  nand
  g1354
  (
    n1369,
    n1365,
    n1336,
    n1363,
    n1332
  );


  and
  g1355
  (
    n1378,
    n1331,
    n1332,
    n1334,
    n1335
  );


  nor
  g1356
  (
    n1383,
    n1337,
    n1068,
    n912,
    n1341
  );


  or
  g1357
  (
    n1380,
    n913,
    n1364,
    n1366
  );


  and
  g1358
  (
    n1374,
    n914,
    n1330,
    n1367
  );


  xnor
  g1359
  (
    n1379,
    n1339,
    n912,
    n1340,
    n1334
  );


  nor
  g1360
  (
    n1385,
    n1368,
    n1333,
    n1366,
    n1364
  );


  nand
  g1361
  (
    n1381,
    n914,
    n913,
    n1341,
    n1340
  );


  or
  g1362
  (
    n1370,
    n1335,
    n1367,
    n914,
    n1368
  );


  not
  g1363
  (
    n1400,
    n1359
  );


  nor
  g1364
  (
    n1426,
    n1375,
    n1378
  );


  xnor
  g1365
  (
    n1395,
    n1360,
    n1158
  );


  nor
  g1366
  (
    n1410,
    n1377,
    n110
  );


  nor
  g1367
  (
    n1406,
    n1159,
    n1068
  );


  nor
  g1368
  (
    n1409,
    n1369,
    n1351
  );


  or
  g1369
  (
    n1411,
    n1362,
    n1382
  );


  or
  g1370
  (
    n1407,
    n1355,
    n1349
  );


  nand
  g1371
  (
    n1415,
    n915,
    n1348
  );


  xnor
  g1372
  (
    n1405,
    n1347,
    n1354
  );


  nand
  g1373
  (
    n1408,
    n1070,
    n1355
  );


  nor
  g1374
  (
    n1393,
    n1161,
    n1380
  );


  nor
  g1375
  (
    n1425,
    n1160,
    n1357,
    n1356,
    n1377
  );


  xnor
  g1376
  (
    n1399,
    n1358,
    n1380,
    n1353,
    n1343
  );


  nor
  g1377
  (
    n1401,
    n1379,
    n1162,
    n1361,
    n1069
  );


  and
  g1378
  (
    n1387,
    n1360,
    n1350,
    n1361,
    n1378
  );


  nor
  g1379
  (
    n1392,
    n1344,
    n1344,
    n1372,
    n1349
  );


  or
  g1380
  (
    n1402,
    n1385,
    n1381,
    n1348,
    n1350
  );


  and
  g1381
  (
    n1403,
    n1357,
    n1358,
    n1164,
    n1343
  );


  xor
  g1382
  (
    n1398,
    n915,
    n1353,
    n1351,
    n1362
  );


  or
  g1383
  (
    n1413,
    n1346,
    n1381,
    n1350,
    n1069
  );


  xnor
  g1384
  (
    n1389,
    n1342,
    n1383,
    n1161
  );


  xnor
  g1385
  (
    n1420,
    n1160,
    n1070,
    n1382,
    n1347
  );


  xor
  g1386
  (
    n1423,
    n1351,
    n1163,
    n1355,
    n1166
  );


  or
  g1387
  (
    n1416,
    n1165,
    n1384,
    n1359,
    n1356
  );


  xor
  g1388
  (
    n1396,
    n1069,
    n915,
    n1362,
    n1358
  );


  or
  g1389
  (
    n1421,
    n1164,
    n1357,
    n1379,
    n1355
  );


  nand
  g1390
  (
    n1427,
    n1377,
    n1383,
    n1347,
    n1382
  );


  xor
  g1391
  (
    n1414,
    n1352,
    n1352,
    n1162,
    n1350
  );


  xnor
  g1392
  (
    n1391,
    n1351,
    n1354,
    n1361,
    n1384
  );


  or
  g1393
  (
    n1386,
    n1362,
    n1352,
    n1346,
    n1374
  );


  nand
  g1394
  (
    n1422,
    n1349,
    n1373,
    n1070,
    n1371
  );


  and
  g1395
  (
    n1404,
    n1376,
    n1165,
    n1342,
    n1070
  );


  nand
  g1396
  (
    n1388,
    n1379,
    n1353,
    n1163,
    n1380
  );


  nand
  g1397
  (
    n1424,
    n1360,
    n1381,
    n1345
  );


  nor
  g1398
  (
    n1412,
    n1348,
    n1385,
    n1384
  );


  and
  g1399
  (
    n1417,
    n1347,
    n1383,
    n1353,
    n1167
  );


  and
  g1400
  (
    n1394,
    n1349,
    n1361,
    n1380,
    n1359
  );


  and
  g1401
  (
    n1418,
    n1159,
    n1378,
    n1384,
    n1379
  );


  xor
  g1402
  (
    n1390,
    n1385,
    n1370,
    n1377,
    n1354
  );


  and
  g1403
  (
    n1419,
    n1158,
    n1357,
    n1356,
    n1358
  );


  nor
  g1404
  (
    n1397,
    n1354,
    n1378,
    n1069,
    n1382
  );


  or
  g1405
  (
    n1429,
    n1352,
    n1359,
    n1360,
    n1345
  );


  and
  g1406
  (
    KeyWire_0_12,
    n1356,
    n1166,
    n1167,
    n1348
  );


  and
  g1407
  (
    n1440,
    n1423,
    n1424,
    n1419,
    n1397
  );


  xor
  g1408
  (
    n1432,
    n1421,
    n1388,
    n1429,
    n1400
  );


  nor
  g1409
  (
    n1437,
    n1422,
    n1415,
    n1427,
    n1412
  );


  xor
  g1410
  (
    n1438,
    n1398,
    n1390,
    n1414,
    n1428
  );


  xnor
  g1411
  (
    n1436,
    n1408,
    n1426,
    n1420,
    n1410
  );


  nand
  g1412
  (
    n1434,
    n1391,
    n1418,
    n1416,
    n1395
  );


  xor
  g1413
  (
    n1431,
    n1403,
    n1406,
    n1407,
    n1417
  );


  xnor
  g1414
  (
    n1435,
    n1399,
    n1392,
    n1386,
    n1389
  );


  nand
  g1415
  (
    n1439,
    n1409,
    n1387,
    n1402,
    n1411
  );


  or
  g1416
  (
    n1430,
    n1404,
    n1405,
    n1413,
    n1425
  );


  and
  g1417
  (
    n1433,
    n1394,
    n1393,
    n1401,
    n1396
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n471,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n891,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1053,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1327,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n1052,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1125,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1333,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1311,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n292,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1325,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n655,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n74,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n1428,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n946,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n36,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1346,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n349,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1289,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n211,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n758,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n707,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1347,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n326,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n196,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n96,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n222,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n751,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1225,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n950,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n299,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1351,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n774,
    KeyNOTWire_0_31
  );


endmodule

