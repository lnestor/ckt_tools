

module Stat_3107_39_9
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n2232,
  n2229,
  n2226,
  n2249,
  n2298,
  n2307,
  n2300,
  n2297,
  n2290,
  n2308,
  n2303,
  n2292,
  n3116,
  n3127,
  n3111,
  n3117,
  n3120,
  n3108,
  n3123,
  n3107,
  n3106,
  n3121,
  n3105,
  n3113,
  n3118,
  n3131,
  n3126,
  n3125,
  n3112,
  n3122,
  n3115,
  n3129,
  n3128,
  n3109,
  n3119,
  n3110,
  n3124,
  n3114,
  n3130,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n2232;
  output n2229;
  output n2226;
  output n2249;
  output n2298;
  output n2307;
  output n2300;
  output n2297;
  output n2290;
  output n2308;
  output n2303;
  output n2292;
  output n3116;
  output n3127;
  output n3111;
  output n3117;
  output n3120;
  output n3108;
  output n3123;
  output n3107;
  output n3106;
  output n3121;
  output n3105;
  output n3113;
  output n3118;
  output n3131;
  output n3126;
  output n3125;
  output n3112;
  output n3122;
  output n3115;
  output n3129;
  output n3128;
  output n3109;
  output n3119;
  output n3110;
  output n3124;
  output n3114;
  output n3130;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2227;
  wire n2228;
  wire n2230;
  wire n2231;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2291;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2299;
  wire n2301;
  wire n2302;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire n3030;
  wire n3031;
  wire n3032;
  wire n3033;
  wire n3034;
  wire n3035;
  wire n3036;
  wire n3037;
  wire n3038;
  wire n3039;
  wire n3040;
  wire n3041;
  wire n3042;
  wire n3043;
  wire n3044;
  wire n3045;
  wire n3046;
  wire n3047;
  wire n3048;
  wire n3049;
  wire n3050;
  wire n3051;
  wire n3052;
  wire n3053;
  wire n3054;
  wire n3055;
  wire n3056;
  wire n3057;
  wire n3058;
  wire n3059;
  wire n3060;
  wire n3061;
  wire n3062;
  wire n3063;
  wire n3064;
  wire n3065;
  wire n3066;
  wire n3067;
  wire n3068;
  wire n3069;
  wire n3070;
  wire n3071;
  wire n3072;
  wire n3073;
  wire n3074;
  wire n3075;
  wire n3076;
  wire n3077;
  wire n3078;
  wire n3079;
  wire n3080;
  wire n3081;
  wire n3082;
  wire n3083;
  wire n3084;
  wire n3085;
  wire n3086;
  wire n3087;
  wire n3088;
  wire n3089;
  wire n3090;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire n3095;
  wire n3096;
  wire n3097;
  wire n3098;
  wire n3099;
  wire n3100;
  wire n3101;
  wire n3102;
  wire n3103;
  wire n3104;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n97,
    n1
  );


  not
  g1
  (
    n27,
    n20
  );


  not
  g2
  (
    n51,
    n18
  );


  buf
  g3
  (
    n108,
    n18
  );


  not
  g4
  (
    n88,
    n8
  );


  not
  g5
  (
    n70,
    n18
  );


  not
  g6
  (
    n58,
    n3
  );


  buf
  g7
  (
    n72,
    n3
  );


  buf
  g8
  (
    n95,
    n9
  );


  buf
  g9
  (
    n48,
    n5
  );


  not
  g10
  (
    n81,
    n15
  );


  not
  g11
  (
    n54,
    n14
  );


  buf
  g12
  (
    n115,
    n21
  );


  not
  g13
  (
    n38,
    n14
  );


  buf
  g14
  (
    n92,
    n23
  );


  buf
  g15
  (
    n101,
    n10
  );


  buf
  g16
  (
    n91,
    n5
  );


  buf
  g17
  (
    n33,
    n19
  );


  not
  g18
  (
    n100,
    n10
  );


  not
  g19
  (
    n30,
    n16
  );


  not
  g20
  (
    n107,
    n16
  );


  not
  g21
  (
    n36,
    n24
  );


  buf
  g22
  (
    n74,
    n23
  );


  not
  g23
  (
    n49,
    n18
  );


  buf
  g24
  (
    n68,
    n17
  );


  not
  g25
  (
    n39,
    n24
  );


  not
  g26
  (
    n102,
    n8
  );


  buf
  g27
  (
    n80,
    n6
  );


  buf
  g28
  (
    n34,
    n7
  );


  not
  g29
  (
    n65,
    n14
  );


  buf
  g30
  (
    n110,
    n8
  );


  buf
  g31
  (
    n28,
    n12
  );


  not
  g32
  (
    n116,
    n12
  );


  not
  g33
  (
    n55,
    n4
  );


  not
  g34
  (
    n73,
    n2
  );


  not
  g35
  (
    n41,
    n21
  );


  buf
  g36
  (
    n113,
    n7
  );


  buf
  g37
  (
    n114,
    n13
  );


  not
  g38
  (
    n90,
    n10
  );


  buf
  g39
  (
    n75,
    n2
  );


  buf
  g40
  (
    n98,
    n9
  );


  not
  g41
  (
    n50,
    n7
  );


  buf
  g42
  (
    n86,
    n16
  );


  not
  g43
  (
    n111,
    n9
  );


  buf
  g44
  (
    n119,
    n20
  );


  not
  g45
  (
    n106,
    n19
  );


  not
  g46
  (
    n40,
    n24
  );


  buf
  g47
  (
    n52,
    n13
  );


  not
  g48
  (
    n56,
    n3
  );


  buf
  g49
  (
    n62,
    n3
  );


  buf
  g50
  (
    n32,
    n11
  );


  buf
  g51
  (
    n25,
    n23
  );


  buf
  g52
  (
    n29,
    n15
  );


  buf
  g53
  (
    n87,
    n6
  );


  buf
  g54
  (
    n60,
    n22
  );


  not
  g55
  (
    n45,
    n2
  );


  buf
  g56
  (
    n103,
    n17
  );


  buf
  g57
  (
    n112,
    n2
  );


  buf
  g58
  (
    n44,
    n4
  );


  not
  g59
  (
    n93,
    n6
  );


  buf
  g60
  (
    n71,
    n15
  );


  buf
  g61
  (
    n84,
    n1
  );


  not
  g62
  (
    n89,
    n9
  );


  buf
  g63
  (
    n35,
    n5
  );


  not
  g64
  (
    n57,
    n13
  );


  buf
  g65
  (
    n59,
    n12
  );


  not
  g66
  (
    n104,
    n20
  );


  not
  g67
  (
    n63,
    n4
  );


  not
  g68
  (
    n99,
    n13
  );


  not
  g69
  (
    n120,
    n16
  );


  not
  g70
  (
    n69,
    n4
  );


  not
  g71
  (
    n105,
    n17
  );


  buf
  g72
  (
    n96,
    n11
  );


  not
  g73
  (
    n118,
    n15
  );


  buf
  g74
  (
    n26,
    n11
  );


  not
  g75
  (
    n61,
    n22
  );


  buf
  g76
  (
    n83,
    n22
  );


  not
  g77
  (
    n109,
    n6
  );


  not
  g78
  (
    n42,
    n21
  );


  not
  g79
  (
    n85,
    n11
  );


  buf
  g80
  (
    n79,
    n21
  );


  buf
  g81
  (
    n78,
    n19
  );


  not
  g82
  (
    n66,
    n17
  );


  buf
  g83
  (
    n46,
    n1
  );


  not
  g84
  (
    n67,
    n7
  );


  buf
  g85
  (
    n43,
    n1
  );


  buf
  g86
  (
    n117,
    n22
  );


  not
  g87
  (
    n47,
    n5
  );


  buf
  g88
  (
    n76,
    n24
  );


  buf
  g89
  (
    n77,
    n19
  );


  buf
  g90
  (
    n37,
    n10
  );


  not
  g91
  (
    n94,
    n12
  );


  buf
  g92
  (
    n64,
    n8
  );


  buf
  g93
  (
    n82,
    n20
  );


  not
  g94
  (
    n31,
    n23
  );


  buf
  g95
  (
    n53,
    n14
  );


  not
  g96
  (
    n305,
    n84
  );


  not
  g97
  (
    n183,
    n113
  );


  not
  g98
  (
    n231,
    n88
  );


  not
  g99
  (
    n388,
    n42
  );


  buf
  g100
  (
    n262,
    n45
  );


  not
  g101
  (
    n352,
    n99
  );


  buf
  g102
  (
    n167,
    n46
  );


  buf
  g103
  (
    n164,
    n102
  );


  buf
  g104
  (
    n481,
    n94
  );


  not
  g105
  (
    n479,
    n86
  );


  buf
  g106
  (
    n446,
    n92
  );


  buf
  g107
  (
    n220,
    n45
  );


  buf
  g108
  (
    n138,
    n89
  );


  not
  g109
  (
    n132,
    n96
  );


  buf
  g110
  (
    n139,
    n99
  );


  not
  g111
  (
    n314,
    n110
  );


  not
  g112
  (
    n154,
    n37
  );


  not
  g113
  (
    n144,
    n110
  );


  not
  g114
  (
    n405,
    n29
  );


  not
  g115
  (
    n238,
    n81
  );


  not
  g116
  (
    n470,
    n116
  );


  not
  g117
  (
    n413,
    n55
  );


  not
  g118
  (
    n488,
    n100
  );


  buf
  g119
  (
    n222,
    n52
  );


  not
  g120
  (
    n445,
    n109
  );


  buf
  g121
  (
    n131,
    n69
  );


  buf
  g122
  (
    n122,
    n78
  );


  not
  g123
  (
    n324,
    n73
  );


  not
  g124
  (
    n353,
    n50
  );


  buf
  g125
  (
    n386,
    n116
  );


  not
  g126
  (
    n333,
    n92
  );


  not
  g127
  (
    n423,
    n28
  );


  not
  g128
  (
    n253,
    n112
  );


  not
  g129
  (
    n412,
    n72
  );


  not
  g130
  (
    n190,
    n42
  );


  not
  g131
  (
    n419,
    n68
  );


  buf
  g132
  (
    n365,
    n66
  );


  buf
  g133
  (
    n442,
    n41
  );


  not
  g134
  (
    n434,
    n51
  );


  buf
  g135
  (
    n438,
    n40
  );


  buf
  g136
  (
    n245,
    n115
  );


  not
  g137
  (
    n258,
    n108
  );


  not
  g138
  (
    n462,
    n56
  );


  buf
  g139
  (
    n483,
    n107
  );


  not
  g140
  (
    n206,
    n32
  );


  not
  g141
  (
    n387,
    n39
  );


  not
  g142
  (
    n177,
    n42
  );


  buf
  g143
  (
    n246,
    n85
  );


  not
  g144
  (
    n148,
    n77
  );


  buf
  g145
  (
    n156,
    n108
  );


  buf
  g146
  (
    n227,
    n31
  );


  not
  g147
  (
    n179,
    n89
  );


  buf
  g148
  (
    n151,
    n105
  );


  buf
  g149
  (
    n406,
    n65
  );


  not
  g150
  (
    n150,
    n53
  );


  buf
  g151
  (
    n340,
    n83
  );


  buf
  g152
  (
    n436,
    n35
  );


  not
  g153
  (
    n255,
    n75
  );


  not
  g154
  (
    n494,
    n34
  );


  buf
  g155
  (
    n303,
    n101
  );


  buf
  g156
  (
    n391,
    n92
  );


  not
  g157
  (
    n424,
    n111
  );


  not
  g158
  (
    n230,
    n52
  );


  buf
  g159
  (
    n301,
    n64
  );


  buf
  g160
  (
    n404,
    n78
  );


  not
  g161
  (
    n444,
    n74
  );


  buf
  g162
  (
    n399,
    n79
  );


  not
  g163
  (
    n256,
    n59
  );


  buf
  g164
  (
    n384,
    n63
  );


  buf
  g165
  (
    n322,
    n64
  );


  not
  g166
  (
    n130,
    n45
  );


  not
  g167
  (
    n326,
    n107
  );


  not
  g168
  (
    n234,
    n78
  );


  buf
  g169
  (
    n425,
    n82
  );


  not
  g170
  (
    n276,
    n55
  );


  not
  g171
  (
    n327,
    n27
  );


  buf
  g172
  (
    n395,
    n49
  );


  buf
  g173
  (
    n466,
    n30
  );


  buf
  g174
  (
    n473,
    n75
  );


  not
  g175
  (
    n250,
    n67
  );


  buf
  g176
  (
    n221,
    n57
  );


  not
  g177
  (
    n485,
    n60
  );


  not
  g178
  (
    n441,
    n83
  );


  not
  g179
  (
    n199,
    n93
  );


  buf
  g180
  (
    n398,
    n54
  );


  not
  g181
  (
    n459,
    n37
  );


  not
  g182
  (
    n341,
    n76
  );


  buf
  g183
  (
    n338,
    n44
  );


  buf
  g184
  (
    n282,
    n87
  );


  not
  g185
  (
    n373,
    n52
  );


  buf
  g186
  (
    n123,
    n97
  );


  buf
  g187
  (
    n382,
    n55
  );


  buf
  g188
  (
    n414,
    n27
  );


  not
  g189
  (
    n225,
    n57
  );


  buf
  g190
  (
    n235,
    n62
  );


  buf
  g191
  (
    n178,
    n62
  );


  buf
  g192
  (
    n328,
    n114
  );


  buf
  g193
  (
    n216,
    n56
  );


  buf
  g194
  (
    n366,
    n49
  );


  not
  g195
  (
    n394,
    n28
  );


  not
  g196
  (
    n455,
    n82
  );


  not
  g197
  (
    n280,
    n91
  );


  buf
  g198
  (
    n430,
    n113
  );


  buf
  g199
  (
    n347,
    n58
  );


  buf
  g200
  (
    n292,
    n69
  );


  not
  g201
  (
    n370,
    n90
  );


  buf
  g202
  (
    n209,
    n119
  );


  buf
  g203
  (
    n482,
    n110
  );


  not
  g204
  (
    n486,
    n103
  );


  buf
  g205
  (
    n126,
    n105
  );


  buf
  g206
  (
    n415,
    n26
  );


  not
  g207
  (
    n196,
    n44
  );


  buf
  g208
  (
    n332,
    n43
  );


  not
  g209
  (
    n267,
    n68
  );


  not
  g210
  (
    n233,
    n30
  );


  buf
  g211
  (
    n166,
    n61
  );


  not
  g212
  (
    n173,
    n75
  );


  not
  g213
  (
    n224,
    n33
  );


  buf
  g214
  (
    n359,
    n112
  );


  not
  g215
  (
    n211,
    n94
  );


  not
  g216
  (
    n428,
    n43
  );


  buf
  g217
  (
    n411,
    n29
  );


  buf
  g218
  (
    n153,
    n47
  );


  buf
  g219
  (
    n329,
    n50
  );


  buf
  g220
  (
    n458,
    n114
  );


  buf
  g221
  (
    n187,
    n84
  );


  buf
  g222
  (
    n193,
    n103
  );


  not
  g223
  (
    n294,
    n60
  );


  buf
  g224
  (
    n439,
    n104
  );


  buf
  g225
  (
    n315,
    n82
  );


  not
  g226
  (
    n279,
    n53
  );


  not
  g227
  (
    n283,
    n118
  );


  not
  g228
  (
    n121,
    n86
  );


  buf
  g229
  (
    n307,
    n87
  );


  not
  g230
  (
    n496,
    n88
  );


  buf
  g231
  (
    n480,
    n76
  );


  not
  g232
  (
    n313,
    n49
  );


  not
  g233
  (
    n429,
    n105
  );


  buf
  g234
  (
    n135,
    n86
  );


  not
  g235
  (
    n277,
    n59
  );


  not
  g236
  (
    n192,
    n113
  );


  not
  g237
  (
    n499,
    n35
  );


  not
  g238
  (
    n378,
    n40
  );


  not
  g239
  (
    n460,
    n119
  );


  buf
  g240
  (
    n318,
    n84
  );


  buf
  g241
  (
    n133,
    n57
  );


  buf
  g242
  (
    n448,
    n85
  );


  not
  g243
  (
    n364,
    n86
  );


  buf
  g244
  (
    n194,
    n95
  );


  not
  g245
  (
    n208,
    n118
  );


  buf
  g246
  (
    n437,
    n66
  );


  buf
  g247
  (
    KeyWire_0_0,
    n111
  );


  not
  g248
  (
    n357,
    n38
  );


  buf
  g249
  (
    n330,
    n76
  );


  not
  g250
  (
    n207,
    n63
  );


  buf
  g251
  (
    n240,
    n99
  );


  not
  g252
  (
    n360,
    n60
  );


  buf
  g253
  (
    n270,
    n67
  );


  buf
  g254
  (
    n375,
    n51
  );


  not
  g255
  (
    n200,
    n119
  );


  not
  g256
  (
    n219,
    n53
  );


  buf
  g257
  (
    n478,
    n54
  );


  not
  g258
  (
    n477,
    n65
  );


  buf
  g259
  (
    n427,
    n56
  );


  buf
  g260
  (
    n214,
    n31
  );


  buf
  g261
  (
    n204,
    n48
  );


  not
  g262
  (
    n181,
    n77
  );


  buf
  g263
  (
    n497,
    n28
  );


  not
  g264
  (
    n409,
    n107
  );


  buf
  g265
  (
    n475,
    n53
  );


  buf
  g266
  (
    n312,
    n64
  );


  buf
  g267
  (
    n464,
    n57
  );


  not
  g268
  (
    n308,
    n43
  );


  buf
  g269
  (
    n146,
    n65
  );


  not
  g270
  (
    n127,
    n73
  );


  not
  g271
  (
    n161,
    n76
  );


  not
  g272
  (
    n362,
    n26
  );


  buf
  g273
  (
    n182,
    n46
  );


  buf
  g274
  (
    n321,
    n62
  );


  buf
  g275
  (
    n472,
    n91
  );


  buf
  g276
  (
    n431,
    n31
  );


  not
  g277
  (
    n356,
    n98
  );


  buf
  g278
  (
    n371,
    n116
  );


  buf
  g279
  (
    n215,
    n83
  );


  not
  g280
  (
    n311,
    n83
  );


  not
  g281
  (
    n463,
    n117
  );


  buf
  g282
  (
    n418,
    n119
  );


  not
  g283
  (
    n316,
    n118
  );


  buf
  g284
  (
    n249,
    n51
  );


  buf
  g285
  (
    n197,
    n40
  );


  not
  g286
  (
    n205,
    n37
  );


  not
  g287
  (
    n269,
    n70
  );


  not
  g288
  (
    n420,
    n89
  );


  not
  g289
  (
    n383,
    n37
  );


  buf
  g290
  (
    n278,
    n46
  );


  buf
  g291
  (
    n241,
    n49
  );


  not
  g292
  (
    n291,
    n29
  );


  not
  g293
  (
    n218,
    n40
  );


  buf
  g294
  (
    n342,
    n79
  );


  buf
  g295
  (
    n201,
    n97
  );


  buf
  g296
  (
    n296,
    n72
  );


  not
  g297
  (
    n259,
    n36
  );


  buf
  g298
  (
    n467,
    n61
  );


  buf
  g299
  (
    n495,
    n70
  );


  buf
  g300
  (
    n223,
    n74
  );


  not
  g301
  (
    n152,
    n54
  );


  buf
  g302
  (
    n410,
    n75
  );


  not
  g303
  (
    n440,
    n117
  );


  buf
  g304
  (
    n374,
    n44
  );


  buf
  g305
  (
    n176,
    n32
  );


  not
  g306
  (
    n210,
    n69
  );


  not
  g307
  (
    n325,
    n73
  );


  not
  g308
  (
    n376,
    n94
  );


  buf
  g309
  (
    n407,
    n96
  );


  not
  g310
  (
    n355,
    n74
  );


  buf
  g311
  (
    n377,
    n112
  );


  buf
  g312
  (
    n162,
    n50
  );


  not
  g313
  (
    n229,
    n33
  );


  not
  g314
  (
    n487,
    n70
  );


  buf
  g315
  (
    n396,
    n93
  );


  not
  g316
  (
    KeyWire_0_12,
    n110
  );


  not
  g317
  (
    n454,
    n41
  );


  not
  g318
  (
    n421,
    n58
  );


  not
  g319
  (
    n174,
    n106
  );


  not
  g320
  (
    n381,
    n109
  );


  buf
  g321
  (
    n149,
    n63
  );


  not
  g322
  (
    n195,
    n71
  );


  buf
  g323
  (
    n336,
    n79
  );


  buf
  g324
  (
    n287,
    n38
  );


  not
  g325
  (
    n389,
    n80
  );


  buf
  g326
  (
    n157,
    n34
  );


  not
  g327
  (
    n251,
    n87
  );


  not
  g328
  (
    n186,
    n115
  );


  not
  g329
  (
    n266,
    n32
  );


  not
  g330
  (
    n129,
    n48
  );


  not
  g331
  (
    n275,
    n95
  );


  buf
  g332
  (
    n498,
    n100
  );


  not
  g333
  (
    n317,
    n101
  );


  buf
  g334
  (
    n416,
    n104
  );


  not
  g335
  (
    n476,
    n74
  );


  buf
  g336
  (
    n203,
    n108
  );


  buf
  g337
  (
    n299,
    n39
  );


  buf
  g338
  (
    n319,
    n62
  );


  not
  g339
  (
    n271,
    n25
  );


  not
  g340
  (
    n247,
    n36
  );


  not
  g341
  (
    n335,
    n88
  );


  not
  g342
  (
    n172,
    n81
  );


  not
  g343
  (
    n358,
    n61
  );


  buf
  g344
  (
    n289,
    n93
  );


  buf
  g345
  (
    n422,
    n41
  );


  buf
  g346
  (
    n169,
    n106
  );


  buf
  g347
  (
    n500,
    n72
  );


  not
  g348
  (
    n300,
    n78
  );


  buf
  g349
  (
    n397,
    n47
  );


  not
  g350
  (
    n293,
    n111
  );


  buf
  g351
  (
    n302,
    n81
  );


  buf
  g352
  (
    n239,
    n61
  );


  not
  g353
  (
    n254,
    n25
  );


  buf
  g354
  (
    n492,
    n27
  );


  not
  g355
  (
    n217,
    n107
  );


  buf
  g356
  (
    n142,
    n97
  );


  buf
  g357
  (
    n408,
    n97
  );


  buf
  g358
  (
    n331,
    n102
  );


  not
  g359
  (
    n165,
    n54
  );


  buf
  g360
  (
    KeyWire_0_7,
    n80
  );


  not
  g361
  (
    n484,
    n64
  );


  not
  g362
  (
    n237,
    n56
  );


  buf
  g363
  (
    n184,
    n115
  );


  buf
  g364
  (
    n125,
    n115
  );


  buf
  g365
  (
    KeyWire_0_13,
    n80
  );


  not
  g366
  (
    n264,
    n80
  );


  buf
  g367
  (
    n160,
    n73
  );


  not
  g368
  (
    n426,
    n39
  );


  not
  g369
  (
    n143,
    n77
  );


  buf
  g370
  (
    n469,
    n66
  );


  not
  g371
  (
    n385,
    n103
  );


  buf
  g372
  (
    n159,
    n59
  );


  buf
  g373
  (
    n134,
    n90
  );


  buf
  g374
  (
    n349,
    n98
  );


  buf
  g375
  (
    n344,
    n116
  );


  not
  g376
  (
    n297,
    n59
  );


  buf
  g377
  (
    n145,
    n67
  );


  not
  g378
  (
    n304,
    n26
  );


  not
  g379
  (
    n402,
    n32
  );


  not
  g380
  (
    n465,
    n44
  );


  buf
  g381
  (
    n306,
    n38
  );


  not
  g382
  (
    n273,
    n34
  );


  buf
  g383
  (
    n274,
    n65
  );


  buf
  g384
  (
    n369,
    n38
  );


  buf
  g385
  (
    n433,
    n67
  );


  buf
  g386
  (
    n202,
    n118
  );


  not
  g387
  (
    n449,
    n41
  );


  buf
  g388
  (
    KeyWire_0_26,
    n101
  );


  not
  g389
  (
    n260,
    n34
  );


  buf
  g390
  (
    n168,
    n60
  );


  buf
  g391
  (
    n450,
    n35
  );


  not
  g392
  (
    n191,
    n96
  );


  not
  g393
  (
    n451,
    n71
  );


  not
  g394
  (
    n501,
    n85
  );


  buf
  g395
  (
    n443,
    n92
  );


  not
  g396
  (
    n393,
    n89
  );


  not
  g397
  (
    n128,
    n58
  );


  not
  g398
  (
    n309,
    n95
  );


  buf
  g399
  (
    n212,
    n99
  );


  not
  g400
  (
    n489,
    n95
  );


  not
  g401
  (
    n252,
    n30
  );


  not
  g402
  (
    n348,
    n52
  );


  not
  g403
  (
    n367,
    n100
  );


  buf
  g404
  (
    n379,
    n90
  );


  buf
  g405
  (
    n261,
    n28
  );


  not
  g406
  (
    n372,
    n48
  );


  buf
  g407
  (
    n163,
    n106
  );


  not
  g408
  (
    n350,
    n26
  );


  buf
  g409
  (
    n137,
    n30
  );


  not
  g410
  (
    n298,
    n82
  );


  not
  g411
  (
    n345,
    n109
  );


  buf
  g412
  (
    n310,
    n91
  );


  not
  g413
  (
    n268,
    n77
  );


  not
  g414
  (
    n198,
    n102
  );


  buf
  g415
  (
    n354,
    n88
  );


  not
  g416
  (
    n170,
    n42
  );


  buf
  g417
  (
    n363,
    n98
  );


  not
  g418
  (
    n368,
    n104
  );


  not
  g419
  (
    n474,
    n81
  );


  buf
  g420
  (
    n403,
    n72
  );


  buf
  g421
  (
    n147,
    n106
  );


  not
  g422
  (
    n124,
    n111
  );


  buf
  g423
  (
    n189,
    n55
  );


  buf
  g424
  (
    n285,
    n69
  );


  buf
  g425
  (
    n337,
    n104
  );


  not
  g426
  (
    n213,
    n47
  );


  not
  g427
  (
    n244,
    n33
  );


  buf
  g428
  (
    n334,
    n98
  );


  not
  g429
  (
    n380,
    n31
  );


  buf
  g430
  (
    n232,
    n109
  );


  not
  g431
  (
    n188,
    n71
  );


  not
  g432
  (
    n281,
    n29
  );


  not
  g433
  (
    n432,
    n25
  );


  not
  g434
  (
    n392,
    n91
  );


  buf
  g435
  (
    n320,
    n68
  );


  buf
  g436
  (
    n457,
    n66
  );


  buf
  g437
  (
    n361,
    n47
  );


  buf
  g438
  (
    n461,
    n79
  );


  not
  g439
  (
    n468,
    n114
  );


  not
  g440
  (
    n290,
    n114
  );


  not
  g441
  (
    n185,
    n71
  );


  buf
  g442
  (
    n456,
    n90
  );


  buf
  g443
  (
    n284,
    n117
  );


  not
  g444
  (
    n417,
    n101
  );


  buf
  g445
  (
    n295,
    n70
  );


  not
  g446
  (
    n228,
    n120
  );


  buf
  g447
  (
    n263,
    n39
  );


  not
  g448
  (
    n158,
    n112
  );


  buf
  g449
  (
    n171,
    n100
  );


  not
  g450
  (
    n400,
    n102
  );


  buf
  g451
  (
    n323,
    n35
  );


  not
  g452
  (
    n272,
    n25
  );


  buf
  g453
  (
    n343,
    n117
  );


  not
  g454
  (
    n493,
    n48
  );


  buf
  g455
  (
    n175,
    n45
  );


  buf
  g456
  (
    n155,
    n68
  );


  buf
  g457
  (
    n286,
    n63
  );


  buf
  g458
  (
    n471,
    n113
  );


  not
  g459
  (
    n226,
    n51
  );


  buf
  g460
  (
    n346,
    n103
  );


  buf
  g461
  (
    n243,
    n84
  );


  not
  g462
  (
    n435,
    n87
  );


  not
  g463
  (
    n141,
    n36
  );


  not
  g464
  (
    n140,
    n108
  );


  not
  g465
  (
    n401,
    n46
  );


  not
  g466
  (
    n242,
    n85
  );


  buf
  g467
  (
    n351,
    n105
  );


  buf
  g468
  (
    n452,
    n94
  );


  buf
  g469
  (
    n453,
    n50
  );


  buf
  g470
  (
    n339,
    n27
  );


  not
  g471
  (
    n491,
    n96
  );


  not
  g472
  (
    n248,
    n36
  );


  buf
  g473
  (
    n136,
    n93
  );


  buf
  g474
  (
    n265,
    n43
  );


  buf
  g475
  (
    n288,
    n58
  );


  buf
  g476
  (
    n180,
    n33
  );


  not
  g477
  (
    n792,
    n143
  );


  buf
  g478
  (
    n1230,
    n324
  );


  not
  g479
  (
    n1029,
    n321
  );


  buf
  g480
  (
    KeyWire_0_15,
    n184
  );


  not
  g481
  (
    n653,
    n388
  );


  buf
  g482
  (
    n1354,
    n175
  );


  buf
  g483
  (
    n565,
    n159
  );


  not
  g484
  (
    n768,
    n371
  );


  buf
  g485
  (
    n505,
    n169
  );


  not
  g486
  (
    n1044,
    n311
  );


  not
  g487
  (
    n1385,
    n292
  );


  buf
  g488
  (
    n678,
    n260
  );


  not
  g489
  (
    n1439,
    n367
  );


  buf
  g490
  (
    n1315,
    n175
  );


  buf
  g491
  (
    n1259,
    n361
  );


  buf
  g492
  (
    n677,
    n304
  );


  not
  g493
  (
    n1189,
    n157
  );


  not
  g494
  (
    n727,
    n343
  );


  buf
  g495
  (
    n735,
    n306
  );


  buf
  g496
  (
    n1160,
    n222
  );


  not
  g497
  (
    n912,
    n354
  );


  buf
  g498
  (
    n1061,
    n261
  );


  buf
  g499
  (
    n1172,
    n277
  );


  not
  g500
  (
    n902,
    n260
  );


  buf
  g501
  (
    n502,
    n190
  );


  not
  g502
  (
    n1426,
    n259
  );


  buf
  g503
  (
    n1124,
    n211
  );


  buf
  g504
  (
    n1241,
    n128
  );


  buf
  g505
  (
    n1398,
    n357
  );


  buf
  g506
  (
    n1470,
    n206
  );


  not
  g507
  (
    n843,
    n314
  );


  not
  g508
  (
    n1456,
    n337
  );


  buf
  g509
  (
    n692,
    n239
  );


  not
  g510
  (
    n1348,
    n267
  );


  not
  g511
  (
    n863,
    n131
  );


  buf
  g512
  (
    n625,
    n223
  );


  buf
  g513
  (
    n1097,
    n128
  );


  buf
  g514
  (
    n1482,
    n343
  );


  not
  g515
  (
    n594,
    n209
  );


  not
  g516
  (
    n1043,
    n204
  );


  not
  g517
  (
    n1091,
    n268
  );


  buf
  g518
  (
    n503,
    n158
  );


  not
  g519
  (
    n1009,
    n142
  );


  buf
  g520
  (
    n1473,
    n208
  );


  buf
  g521
  (
    n577,
    n299
  );


  not
  g522
  (
    n872,
    n223
  );


  not
  g523
  (
    n1074,
    n244
  );


  buf
  g524
  (
    n1353,
    n322
  );


  not
  g525
  (
    n1051,
    n249
  );


  not
  g526
  (
    n1069,
    n311
  );


  not
  g527
  (
    n1250,
    n122
  );


  buf
  g528
  (
    n518,
    n144
  );


  buf
  g529
  (
    n786,
    n174
  );


  not
  g530
  (
    n1316,
    n321
  );


  buf
  g531
  (
    n1382,
    n198
  );


  not
  g532
  (
    n751,
    n167
  );


  buf
  g533
  (
    n970,
    n125
  );


  buf
  g534
  (
    n812,
    n314
  );


  buf
  g535
  (
    n1056,
    n204
  );


  not
  g536
  (
    n941,
    n300
  );


  not
  g537
  (
    n811,
    n134
  );


  not
  g538
  (
    n1296,
    n145
  );


  buf
  g539
  (
    n628,
    n331
  );


  not
  g540
  (
    n973,
    n132
  );


  buf
  g541
  (
    n743,
    n275
  );


  not
  g542
  (
    n1286,
    n209
  );


  not
  g543
  (
    n659,
    n216
  );


  not
  g544
  (
    n1361,
    n369
  );


  not
  g545
  (
    n724,
    n276
  );


  not
  g546
  (
    n916,
    n299
  );


  buf
  g547
  (
    n509,
    n295
  );


  not
  g548
  (
    n747,
    n264
  );


  buf
  g549
  (
    n635,
    n276
  );


  not
  g550
  (
    n574,
    n126
  );


  buf
  g551
  (
    n757,
    n339
  );


  not
  g552
  (
    n1168,
    n276
  );


  not
  g553
  (
    n510,
    n226
  );


  buf
  g554
  (
    n1035,
    n195
  );


  buf
  g555
  (
    n774,
    n196
  );


  buf
  g556
  (
    n763,
    n183
  );


  buf
  g557
  (
    n830,
    n178
  );


  buf
  g558
  (
    n1132,
    n263
  );


  not
  g559
  (
    n1411,
    n325
  );


  not
  g560
  (
    n880,
    n233
  );


  not
  g561
  (
    n1063,
    n306
  );


  buf
  g562
  (
    n1360,
    n279
  );


  not
  g563
  (
    n674,
    n279
  );


  not
  g564
  (
    n834,
    n170
  );


  not
  g565
  (
    n1210,
    n366
  );


  not
  g566
  (
    n562,
    n258
  );


  buf
  g567
  (
    n1220,
    n241
  );


  not
  g568
  (
    n1330,
    n387
  );


  not
  g569
  (
    KeyWire_0_9,
    n129
  );


  not
  g570
  (
    n546,
    n152
  );


  not
  g571
  (
    n1182,
    n180
  );


  buf
  g572
  (
    n672,
    n335
  );


  buf
  g573
  (
    n1487,
    n315
  );


  buf
  g574
  (
    n1016,
    n147
  );


  buf
  g575
  (
    n938,
    n225
  );


  not
  g576
  (
    n1046,
    n254
  );


  not
  g577
  (
    n890,
    n334
  );


  not
  g578
  (
    n942,
    n227
  );


  not
  g579
  (
    n1404,
    n345
  );


  buf
  g580
  (
    n1239,
    n134
  );


  buf
  g581
  (
    n922,
    n286
  );


  not
  g582
  (
    n1012,
    n352
  );


  buf
  g583
  (
    n1170,
    n289
  );


  buf
  g584
  (
    n1090,
    n174
  );


  buf
  g585
  (
    KeyWire_0_8,
    n212
  );


  buf
  g586
  (
    n564,
    n208
  );


  buf
  g587
  (
    n764,
    n143
  );


  not
  g588
  (
    n985,
    n224
  );


  buf
  g589
  (
    n818,
    n367
  );


  not
  g590
  (
    n1326,
    n234
  );


  buf
  g591
  (
    n1409,
    n320
  );


  not
  g592
  (
    n1447,
    n184
  );


  buf
  g593
  (
    n1134,
    n383
  );


  buf
  g594
  (
    n1373,
    n257
  );


  buf
  g595
  (
    n867,
    n363
  );


  buf
  g596
  (
    n645,
    n378
  );


  buf
  g597
  (
    n1460,
    n139
  );


  not
  g598
  (
    n707,
    n255
  );


  buf
  g599
  (
    n1011,
    n311
  );


  not
  g600
  (
    n865,
    n182
  );


  not
  g601
  (
    n640,
    n136
  );


  not
  g602
  (
    n1464,
    n293
  );


  not
  g603
  (
    n1190,
    n207
  );


  buf
  g604
  (
    n1082,
    n250
  );


  not
  g605
  (
    n819,
    n304
  );


  buf
  g606
  (
    n905,
    n350
  );


  buf
  g607
  (
    n1384,
    n210
  );


  not
  g608
  (
    n1071,
    n222
  );


  not
  g609
  (
    n643,
    n121
  );


  buf
  g610
  (
    n946,
    n228
  );


  not
  g611
  (
    n1085,
    n135
  );


  buf
  g612
  (
    n874,
    n340
  );


  buf
  g613
  (
    n1308,
    n139
  );


  buf
  g614
  (
    n1185,
    n244
  );


  buf
  g615
  (
    n803,
    n216
  );


  not
  g616
  (
    n900,
    n294
  );


  not
  g617
  (
    n759,
    n275
  );


  not
  g618
  (
    n513,
    n342
  );


  not
  g619
  (
    n1100,
    n132
  );


  not
  g620
  (
    n627,
    n176
  );


  buf
  g621
  (
    n709,
    n350
  );


  not
  g622
  (
    n1167,
    n263
  );


  buf
  g623
  (
    n1175,
    n216
  );


  buf
  g624
  (
    n1480,
    n329
  );


  not
  g625
  (
    n1471,
    n242
  );


  not
  g626
  (
    n630,
    n362
  );


  buf
  g627
  (
    n1476,
    n296
  );


  buf
  g628
  (
    n539,
    n344
  );


  buf
  g629
  (
    n1040,
    n375
  );


  buf
  g630
  (
    n669,
    n183
  );


  not
  g631
  (
    n895,
    n346
  );


  buf
  g632
  (
    n808,
    n168
  );


  not
  g633
  (
    n875,
    n133
  );


  not
  g634
  (
    n711,
    n203
  );


  not
  g635
  (
    n1135,
    n295
  );


  not
  g636
  (
    n532,
    n243
  );


  not
  g637
  (
    n1045,
    n258
  );


  not
  g638
  (
    n675,
    n318
  );


  not
  g639
  (
    n858,
    n355
  );


  buf
  g640
  (
    n1058,
    n164
  );


  not
  g641
  (
    n1033,
    n274
  );


  buf
  g642
  (
    n1021,
    n173
  );


  not
  g643
  (
    n1025,
    n159
  );


  not
  g644
  (
    n815,
    n133
  );


  buf
  g645
  (
    n1481,
    n266
  );


  buf
  g646
  (
    n1352,
    n245
  );


  buf
  g647
  (
    n1400,
    n262
  );


  buf
  g648
  (
    n554,
    n167
  );


  not
  g649
  (
    n1219,
    n304
  );


  buf
  g650
  (
    n572,
    n176
  );


  not
  g651
  (
    n986,
    n278
  );


  not
  g652
  (
    n1010,
    n226
  );


  buf
  g653
  (
    n689,
    n320
  );


  buf
  g654
  (
    n655,
    n183
  );


  buf
  g655
  (
    n561,
    n230
  );


  not
  g656
  (
    n903,
    n242
  );


  not
  g657
  (
    n1014,
    n282
  );


  not
  g658
  (
    n1386,
    n387
  );


  buf
  g659
  (
    n1419,
    n182
  );


  buf
  g660
  (
    n1064,
    n199
  );


  not
  g661
  (
    n1133,
    n250
  );


  buf
  g662
  (
    n1054,
    n364
  );


  buf
  g663
  (
    n1454,
    n256
  );


  not
  g664
  (
    n1248,
    n290
  );


  buf
  g665
  (
    n1295,
    n287
  );


  buf
  g666
  (
    n847,
    n234
  );


  not
  g667
  (
    n1150,
    n287
  );


  not
  g668
  (
    n1217,
    n379
  );


  not
  g669
  (
    n883,
    n185
  );


  not
  g670
  (
    n1146,
    n176
  );


  buf
  g671
  (
    n1371,
    n267
  );


  buf
  g672
  (
    n708,
    n227
  );


  buf
  g673
  (
    n878,
    n179
  );


  buf
  g674
  (
    n681,
    n174
  );


  buf
  g675
  (
    n899,
    n320
  );


  buf
  g676
  (
    n1003,
    n386
  );


  buf
  g677
  (
    n713,
    n163
  );


  buf
  g678
  (
    n636,
    n221
  );


  buf
  g679
  (
    n1483,
    n171
  );


  buf
  g680
  (
    n740,
    n204
  );


  not
  g681
  (
    n1293,
    n353
  );


  buf
  g682
  (
    n1027,
    n215
  );


  buf
  g683
  (
    n791,
    n355
  );


  buf
  g684
  (
    n1320,
    n240
  );


  not
  g685
  (
    n1433,
    n328
  );


  buf
  g686
  (
    n1203,
    n363
  );


  not
  g687
  (
    n1484,
    n224
  );


  buf
  g688
  (
    n714,
    n147
  );


  not
  g689
  (
    n1343,
    n290
  );


  not
  g690
  (
    n1281,
    n296
  );


  buf
  g691
  (
    n620,
    n199
  );


  buf
  g692
  (
    n950,
    n344
  );


  buf
  g693
  (
    n1077,
    n294
  );


  buf
  g694
  (
    n846,
    n266
  );


  buf
  g695
  (
    n813,
    n232
  );


  buf
  g696
  (
    n789,
    n136
  );


  buf
  g697
  (
    n1425,
    n212
  );


  buf
  g698
  (
    n1455,
    n346
  );


  buf
  g699
  (
    n918,
    n143
  );


  buf
  g700
  (
    n1365,
    n314
  );


  not
  g701
  (
    n806,
    n386
  );


  not
  g702
  (
    n790,
    n385
  );


  buf
  g703
  (
    n1268,
    n203
  );


  buf
  g704
  (
    n825,
    n251
  );


  buf
  g705
  (
    n1479,
    n359
  );


  not
  g706
  (
    n571,
    n178
  );


  not
  g707
  (
    KeyWire_0_31,
    n247
  );


  buf
  g708
  (
    n1391,
    n128
  );


  buf
  g709
  (
    n773,
    n269
  );


  buf
  g710
  (
    n1107,
    n373
  );


  not
  g711
  (
    n1084,
    n170
  );


  not
  g712
  (
    n524,
    n224
  );


  buf
  g713
  (
    n515,
    n190
  );


  buf
  g714
  (
    n1313,
    n211
  );


  buf
  g715
  (
    n1262,
    n240
  );


  buf
  g716
  (
    n927,
    n379
  );


  buf
  g717
  (
    n1466,
    n342
  );


  not
  g718
  (
    n1192,
    n203
  );


  not
  g719
  (
    n1363,
    n185
  );


  buf
  g720
  (
    n1468,
    n209
  );


  not
  g721
  (
    n1118,
    n152
  );


  buf
  g722
  (
    n798,
    n152
  );


  buf
  g723
  (
    n619,
    n146
  );


  buf
  g724
  (
    n1050,
    n255
  );


  buf
  g725
  (
    n887,
    n279
  );


  buf
  g726
  (
    n736,
    n268
  );


  not
  g727
  (
    n598,
    n264
  );


  not
  g728
  (
    n1137,
    n366
  );


  buf
  g729
  (
    n644,
    n260
  );


  not
  g730
  (
    n1402,
    n202
  );


  buf
  g731
  (
    n584,
    n218
  );


  buf
  g732
  (
    n976,
    n340
  );


  buf
  g733
  (
    n576,
    n160
  );


  buf
  g734
  (
    n1272,
    n194
  );


  buf
  g735
  (
    n964,
    n272
  );


  not
  g736
  (
    n1463,
    n232
  );


  not
  g737
  (
    n1161,
    n303
  );


  buf
  g738
  (
    n971,
    n301
  );


  not
  g739
  (
    n1323,
    n269
  );


  buf
  g740
  (
    n991,
    n163
  );


  not
  g741
  (
    n1086,
    n163
  );


  not
  g742
  (
    n1188,
    n219
  );


  buf
  g743
  (
    n1350,
    n169
  );


  not
  g744
  (
    n647,
    n124
  );


  not
  g745
  (
    n1006,
    n137
  );


  not
  g746
  (
    n664,
    n191
  );


  buf
  g747
  (
    n873,
    n291
  );


  not
  g748
  (
    n519,
    n205
  );


  not
  g749
  (
    n1186,
    n173
  );


  buf
  g750
  (
    n1156,
    n153
  );


  not
  g751
  (
    n881,
    n261
  );


  buf
  g752
  (
    n1452,
    n156
  );


  not
  g753
  (
    n698,
    n348
  );


  not
  g754
  (
    KeyWire_0_29,
    n320
  );


  buf
  g755
  (
    n1184,
    n380
  );


  buf
  g756
  (
    n1112,
    n192
  );


  not
  g757
  (
    n587,
    n247
  );


  not
  g758
  (
    n646,
    n306
  );


  buf
  g759
  (
    n869,
    n369
  );


  not
  g760
  (
    n1453,
    n272
  );


  buf
  g761
  (
    n1042,
    n133
  );


  not
  g762
  (
    n650,
    n250
  );


  not
  g763
  (
    n844,
    n217
  );


  not
  g764
  (
    n1225,
    n353
  );


  buf
  g765
  (
    n1098,
    n365
  );


  not
  g766
  (
    n1148,
    n357
  );


  not
  g767
  (
    n1216,
    n330
  );


  not
  g768
  (
    n746,
    n295
  );


  not
  g769
  (
    n1206,
    n331
  );


  not
  g770
  (
    n679,
    n197
  );


  buf
  g771
  (
    n921,
    n189
  );


  buf
  g772
  (
    n1449,
    n239
  );


  buf
  g773
  (
    n1235,
    n252
  );


  buf
  g774
  (
    n531,
    n200
  );


  buf
  g775
  (
    n893,
    n180
  );


  not
  g776
  (
    n1234,
    n161
  );


  buf
  g777
  (
    n1153,
    n298
  );


  not
  g778
  (
    n580,
    n376
  );


  not
  g779
  (
    n1087,
    n167
  );


  buf
  g780
  (
    n1446,
    n291
  );


  not
  g781
  (
    n1459,
    n221
  );


  not
  g782
  (
    n972,
    n313
  );


  buf
  g783
  (
    n1207,
    n210
  );


  buf
  g784
  (
    n1242,
    n378
  );


  buf
  g785
  (
    n1194,
    n194
  );


  not
  g786
  (
    n667,
    n121
  );


  not
  g787
  (
    n1076,
    n386
  );


  buf
  g788
  (
    n1443,
    n193
  );


  buf
  g789
  (
    n859,
    n259
  );


  not
  g790
  (
    n632,
    n170
  );


  buf
  g791
  (
    n857,
    n133
  );


  not
  g792
  (
    n660,
    n282
  );


  buf
  g793
  (
    n862,
    n192
  );


  not
  g794
  (
    n1261,
    n360
  );


  not
  g795
  (
    n1004,
    n346
  );


  buf
  g796
  (
    n1013,
    n150
  );


  not
  g797
  (
    n1240,
    n121
  );


  buf
  g798
  (
    n1157,
    n222
  );


  buf
  g799
  (
    n777,
    n385
  );


  not
  g800
  (
    n871,
    n151
  );


  buf
  g801
  (
    n831,
    n288
  );


  buf
  g802
  (
    n780,
    n363
  );


  buf
  g803
  (
    n1123,
    n244
  );


  not
  g804
  (
    n526,
    n349
  );


  buf
  g805
  (
    n596,
    n237
  );


  not
  g806
  (
    n1428,
    n374
  );


  not
  g807
  (
    n886,
    n228
  );


  buf
  g808
  (
    n782,
    n197
  );


  buf
  g809
  (
    n823,
    n292
  );


  buf
  g810
  (
    n686,
    n145
  );


  buf
  g811
  (
    n533,
    n219
  );


  not
  g812
  (
    n1290,
    n281
  );


  buf
  g813
  (
    n1034,
    n232
  );


  not
  g814
  (
    n1039,
    n311
  );


  buf
  g815
  (
    n604,
    n338
  );


  not
  g816
  (
    n1109,
    n252
  );


  buf
  g817
  (
    n548,
    n294
  );


  not
  g818
  (
    n1269,
    n151
  );


  buf
  g819
  (
    n1031,
    n315
  );


  not
  g820
  (
    n1304,
    n367
  );


  buf
  g821
  (
    n586,
    n217
  );


  buf
  g822
  (
    n1231,
    n147
  );


  not
  g823
  (
    n563,
    n245
  );


  buf
  g824
  (
    n719,
    n280
  );


  buf
  g825
  (
    n877,
    n345
  );


  buf
  g826
  (
    n1356,
    n348
  );


  not
  g827
  (
    n855,
    n214
  );


  not
  g828
  (
    n1396,
    n229
  );


  not
  g829
  (
    n974,
    n388
  );


  not
  g830
  (
    n975,
    n172
  );


  not
  g831
  (
    n1047,
    n192
  );


  buf
  g832
  (
    n1114,
    n169
  );


  buf
  g833
  (
    n936,
    n253
  );


  buf
  g834
  (
    n593,
    n376
  );


  not
  g835
  (
    n860,
    n343
  );


  buf
  g836
  (
    n1162,
    n306
  );


  buf
  g837
  (
    n605,
    n269
  );


  not
  g838
  (
    n1164,
    n127
  );


  not
  g839
  (
    n892,
    n300
  );


  not
  g840
  (
    n528,
    n329
  );


  buf
  g841
  (
    n573,
    n283
  );


  buf
  g842
  (
    n1368,
    n156
  );


  not
  g843
  (
    n897,
    n342
  );


  buf
  g844
  (
    n608,
    n299
  );


  not
  g845
  (
    n1445,
    n160
  );


  buf
  g846
  (
    n793,
    n150
  );


  buf
  g847
  (
    n1342,
    n213
  );


  buf
  g848
  (
    n1325,
    n193
  );


  not
  g849
  (
    n845,
    n359
  );


  not
  g850
  (
    n1407,
    n175
  );


  buf
  g851
  (
    n1437,
    n319
  );


  not
  g852
  (
    n810,
    n341
  );


  not
  g853
  (
    n779,
    n147
  );


  not
  g854
  (
    n1126,
    n335
  );


  buf
  g855
  (
    n861,
    n160
  );


  buf
  g856
  (
    n882,
    n327
  );


  not
  g857
  (
    n1332,
    n166
  );


  not
  g858
  (
    n1279,
    n228
  );


  buf
  g859
  (
    n1440,
    n360
  );


  buf
  g860
  (
    n1275,
    n126
  );


  not
  g861
  (
    n1270,
    n161
  );


  buf
  g862
  (
    n1362,
    n235
  );


  buf
  g863
  (
    n1357,
    n256
  );


  buf
  g864
  (
    n568,
    n356
  );


  not
  g865
  (
    n919,
    n368
  );


  buf
  g866
  (
    n1211,
    n257
  );


  buf
  g867
  (
    n696,
    n379
  );


  not
  g868
  (
    n582,
    n142
  );


  not
  g869
  (
    n1486,
    n233
  );


  buf
  g870
  (
    n555,
    n259
  );


  buf
  g871
  (
    n1285,
    n332
  );


  buf
  g872
  (
    n992,
    n161
  );


  not
  g873
  (
    n799,
    n172
  );


  buf
  g874
  (
    n700,
    n157
  );


  buf
  g875
  (
    n1331,
    n191
  );


  buf
  g876
  (
    n1128,
    n389
  );


  buf
  g877
  (
    n1193,
    n351
  );


  not
  g878
  (
    n1438,
    n130
  );


  buf
  g879
  (
    n690,
    n371
  );


  not
  g880
  (
    n1244,
    n301
  );


  buf
  g881
  (
    n984,
    n156
  );


  buf
  g882
  (
    n1236,
    n295
  );


  not
  g883
  (
    n896,
    n214
  );


  buf
  g884
  (
    n1258,
    n354
  );


  buf
  g885
  (
    n1020,
    n339
  );


  buf
  g886
  (
    n704,
    n290
  );


  not
  g887
  (
    n626,
    n229
  );


  not
  g888
  (
    n1410,
    n281
  );


  not
  g889
  (
    n618,
    n267
  );


  buf
  g890
  (
    n1345,
    n286
  );


  buf
  g891
  (
    n765,
    n149
  );


  buf
  g892
  (
    n1317,
    n358
  );


  buf
  g893
  (
    n745,
    n121
  );


  buf
  g894
  (
    n787,
    n327
  );


  not
  g895
  (
    n1403,
    n184
  );


  not
  g896
  (
    n800,
    n219
  );


  not
  g897
  (
    n884,
    n376
  );


  buf
  g898
  (
    n739,
    n262
  );


  not
  g899
  (
    n1370,
    n353
  );


  buf
  g900
  (
    n671,
    n271
  );


  buf
  g901
  (
    n754,
    n385
  );


  buf
  g902
  (
    n722,
    n292
  );


  buf
  g903
  (
    n521,
    n248
  );


  buf
  g904
  (
    n926,
    n323
  );


  buf
  g905
  (
    n603,
    n240
  );


  not
  g906
  (
    n1106,
    n140
  );


  buf
  g907
  (
    n506,
    n388
  );


  not
  g908
  (
    n701,
    n272
  );


  not
  g909
  (
    n1399,
    n129
  );


  buf
  g910
  (
    n940,
    n123
  );


  not
  g911
  (
    n1298,
    n282
  );


  buf
  g912
  (
    n1117,
    n161
  );


  not
  g913
  (
    n726,
    n176
  );


  not
  g914
  (
    n1142,
    n188
  );


  buf
  g915
  (
    n1380,
    n281
  );


  not
  g916
  (
    n538,
    n333
  );


  not
  g917
  (
    n981,
    n172
  );


  not
  g918
  (
    n1367,
    n285
  );


  not
  g919
  (
    n1254,
    n262
  );


  not
  g920
  (
    n959,
    n250
  );


  buf
  g921
  (
    n954,
    n352
  );


  not
  g922
  (
    n738,
    n293
  );


  not
  g923
  (
    n1197,
    n380
  );


  not
  g924
  (
    n1257,
    n303
  );


  not
  g925
  (
    n1227,
    n144
  );


  buf
  g926
  (
    n1078,
    n313
  );


  buf
  g927
  (
    n924,
    n224
  );


  buf
  g928
  (
    n889,
    n186
  );


  not
  g929
  (
    n550,
    n283
  );


  not
  g930
  (
    n1310,
    n165
  );


  not
  g931
  (
    n1263,
    n140
  );


  not
  g932
  (
    n989,
    n183
  );


  buf
  g933
  (
    n988,
    n181
  );


  buf
  g934
  (
    n993,
    n158
  );


  buf
  g935
  (
    n931,
    n369
  );


  not
  g936
  (
    n552,
    n139
  );


  buf
  g937
  (
    n1319,
    n370
  );


  buf
  g938
  (
    n1416,
    n225
  );


  buf
  g939
  (
    n1237,
    n170
  );


  not
  g940
  (
    n527,
    n275
  );


  not
  g941
  (
    n589,
    n271
  );


  buf
  g942
  (
    n688,
    n325
  );


  buf
  g943
  (
    n828,
    n177
  );


  not
  g944
  (
    n1388,
    n203
  );


  not
  g945
  (
    n575,
    n218
  );


  not
  g946
  (
    n994,
    n168
  );


  buf
  g947
  (
    n534,
    n336
  );


  buf
  g948
  (
    n1376,
    n205
  );


  not
  g949
  (
    n559,
    n149
  );


  not
  g950
  (
    n609,
    n376
  );


  not
  g951
  (
    n761,
    n194
  );


  buf
  g952
  (
    n657,
    n152
  );


  not
  g953
  (
    n540,
    n327
  );


  not
  g954
  (
    n569,
    n289
  );


  buf
  g955
  (
    n516,
    n146
  );


  buf
  g956
  (
    n1472,
    n142
  );


  buf
  g957
  (
    n1120,
    n283
  );


  not
  g958
  (
    n631,
    n372
  );


  not
  g959
  (
    n1378,
    n301
  );


  not
  g960
  (
    n1346,
    n249
  );


  buf
  g961
  (
    n662,
    n164
  );


  buf
  g962
  (
    n842,
    n310
  );


  buf
  g963
  (
    n1450,
    n138
  );


  buf
  g964
  (
    n1347,
    n351
  );


  buf
  g965
  (
    n535,
    n342
  );


  not
  g966
  (
    n1022,
    n282
  );


  not
  g967
  (
    n1019,
    n327
  );


  buf
  g968
  (
    n1374,
    n333
  );


  buf
  g969
  (
    n553,
    n345
  );


  buf
  g970
  (
    n1334,
    n291
  );


  not
  g971
  (
    n599,
    n350
  );


  not
  g972
  (
    n566,
    n225
  );


  not
  g973
  (
    n511,
    n307
  );


  not
  g974
  (
    n1300,
    n273
  );


  buf
  g975
  (
    n1375,
    n384
  );


  not
  g976
  (
    n687,
    n348
  );


  buf
  g977
  (
    n1277,
    n302
  );


  not
  g978
  (
    n1333,
    n216
  );


  not
  g979
  (
    n1273,
    n248
  );


  not
  g980
  (
    n829,
    n365
  );


  buf
  g981
  (
    n1066,
    n375
  );


  not
  g982
  (
    n1271,
    n337
  );


  buf
  g983
  (
    n545,
    n193
  );


  not
  g984
  (
    n1251,
    n384
  );


  not
  g985
  (
    n1017,
    n150
  );


  not
  g986
  (
    n851,
    n215
  );


  buf
  g987
  (
    n956,
    n300
  );


  buf
  g988
  (
    n904,
    n362
  );


  buf
  g989
  (
    n1477,
    n257
  );


  not
  g990
  (
    n1475,
    n188
  );


  buf
  g991
  (
    n1284,
    n273
  );


  buf
  g992
  (
    n983,
    n318
  );


  buf
  g993
  (
    n685,
    n226
  );


  not
  g994
  (
    n1129,
    n227
  );


  not
  g995
  (
    n838,
    n309
  );


  not
  g996
  (
    n654,
    n249
  );


  not
  g997
  (
    n1420,
    n338
  );


  buf
  g998
  (
    n1155,
    n293
  );


  buf
  g999
  (
    n1249,
    n350
  );


  buf
  g1000
  (
    n1282,
    n352
  );


  not
  g1001
  (
    n1392,
    n324
  );


  buf
  g1002
  (
    n1366,
    n254
  );


  buf
  g1003
  (
    n703,
    n289
  );


  not
  g1004
  (
    n1457,
    n245
  );


  not
  g1005
  (
    n969,
    n195
  );


  buf
  g1006
  (
    n1204,
    n344
  );


  buf
  g1007
  (
    n537,
    n365
  );


  not
  g1008
  (
    n621,
    n179
  );


  not
  g1009
  (
    n1393,
    n303
  );


  buf
  g1010
  (
    n1113,
    n127
  );


  not
  g1011
  (
    n1306,
    n169
  );


  buf
  g1012
  (
    n1288,
    n180
  );


  buf
  g1013
  (
    n1289,
    n159
  );


  not
  g1014
  (
    n1149,
    n313
  );


  not
  g1015
  (
    n1072,
    n302
  );


  not
  g1016
  (
    n641,
    n326
  );


  not
  g1017
  (
    n1144,
    n288
  );


  not
  g1018
  (
    n770,
    n127
  );


  not
  g1019
  (
    n542,
    n181
  );


  buf
  g1020
  (
    n1324,
    n371
  );


  buf
  g1021
  (
    n1212,
    n208
  );


  not
  g1022
  (
    n910,
    n331
  );


  buf
  g1023
  (
    n822,
    n198
  );


  buf
  g1024
  (
    n1057,
    n383
  );


  buf
  g1025
  (
    n522,
    n230
  );


  buf
  g1026
  (
    n588,
    n187
  );


  buf
  g1027
  (
    n721,
    n385
  );


  not
  g1028
  (
    n1461,
    n196
  );


  not
  g1029
  (
    n652,
    n171
  );


  buf
  g1030
  (
    n1213,
    n186
  );


  buf
  g1031
  (
    n957,
    n197
  );


  not
  g1032
  (
    n1215,
    n362
  );


  not
  g1033
  (
    n1015,
    n125
  );


  buf
  g1034
  (
    n925,
    n220
  );


  not
  g1035
  (
    n1138,
    n326
  );


  not
  g1036
  (
    n952,
    n213
  );


  not
  g1037
  (
    n876,
    n246
  );


  buf
  g1038
  (
    n784,
    n387
  );


  not
  g1039
  (
    n507,
    n242
  );


  not
  g1040
  (
    n514,
    n340
  );


  buf
  g1041
  (
    n1173,
    n239
  );


  buf
  g1042
  (
    n682,
    n238
  );


  buf
  g1043
  (
    n804,
    n255
  );


  buf
  g1044
  (
    n642,
    n181
  );


  buf
  g1045
  (
    n908,
    n155
  );


  not
  g1046
  (
    n1312,
    n188
  );


  not
  g1047
  (
    n1297,
    n373
  );


  not
  g1048
  (
    n1052,
    n240
  );


  not
  g1049
  (
    n1089,
    n206
  );


  buf
  g1050
  (
    n1094,
    n252
  );


  not
  g1051
  (
    n1264,
    n211
  );


  not
  g1052
  (
    n1119,
    n239
  );


  buf
  g1053
  (
    n1383,
    n132
  );


  buf
  g1054
  (
    n833,
    n175
  );


  buf
  g1055
  (
    n1278,
    n349
  );


  buf
  g1056
  (
    n639,
    n333
  );


  buf
  g1057
  (
    n944,
    n347
  );


  not
  g1058
  (
    n1053,
    n122
  );


  not
  g1059
  (
    n597,
    n172
  );


  not
  g1060
  (
    n595,
    n337
  );


  not
  g1061
  (
    n723,
    n196
  );


  not
  g1062
  (
    n1181,
    n182
  );


  not
  g1063
  (
    n517,
    n164
  );


  not
  g1064
  (
    n1023,
    n188
  );


  buf
  g1065
  (
    n1202,
    n312
  );


  not
  g1066
  (
    n1414,
    n357
  );


  not
  g1067
  (
    n1122,
    n138
  );


  buf
  g1068
  (
    n1314,
    n276
  );


  not
  g1069
  (
    n615,
    n388
  );


  not
  g1070
  (
    n788,
    n254
  );


  buf
  g1071
  (
    n821,
    n273
  );


  not
  g1072
  (
    n856,
    n220
  );


  not
  g1073
  (
    n1205,
    n287
  );


  buf
  g1074
  (
    n1377,
    n126
  );


  not
  g1075
  (
    n1423,
    n220
  );


  not
  g1076
  (
    n909,
    n138
  );


  buf
  g1077
  (
    n737,
    n125
  );


  not
  g1078
  (
    n1406,
    n234
  );


  buf
  g1079
  (
    n888,
    n191
  );


  not
  g1080
  (
    n879,
    n232
  );


  buf
  g1081
  (
    n715,
    n382
  );


  buf
  g1082
  (
    n996,
    n197
  );


  not
  g1083
  (
    n616,
    n144
  );


  not
  g1084
  (
    n906,
    n372
  );


  buf
  g1085
  (
    n1283,
    n204
  );


  not
  g1086
  (
    n1145,
    n316
  );


  not
  g1087
  (
    n866,
    n237
  );


  not
  g1088
  (
    n1395,
    n262
  );


  buf
  g1089
  (
    n915,
    n230
  );


  buf
  g1090
  (
    n1093,
    n141
  );


  buf
  g1091
  (
    n1096,
    n288
  );


  not
  g1092
  (
    n1340,
    n315
  );


  buf
  g1093
  (
    n1274,
    n246
  );


  not
  g1094
  (
    n928,
    n265
  );


  not
  g1095
  (
    n1435,
    n336
  );


  not
  g1096
  (
    n835,
    n341
  );


  not
  g1097
  (
    n1018,
    n341
  );


  buf
  g1098
  (
    n995,
    n191
  );


  not
  g1099
  (
    n820,
    n130
  );


  not
  g1100
  (
    n1305,
    n238
  );


  buf
  g1101
  (
    n634,
    n281
  );


  buf
  g1102
  (
    n1469,
    n221
  );


  buf
  g1103
  (
    n1232,
    n186
  );


  not
  g1104
  (
    n1478,
    n217
  );


  buf
  g1105
  (
    n1488,
    n189
  );


  not
  g1106
  (
    n1299,
    n151
  );


  buf
  g1107
  (
    n1372,
    n241
  );


  not
  g1108
  (
    n1121,
    n318
  );


  not
  g1109
  (
    n781,
    n231
  );


  buf
  g1110
  (
    n1099,
    n178
  );


  not
  g1111
  (
    n623,
    n277
  );


  not
  g1112
  (
    n826,
    n361
  );


  buf
  g1113
  (
    n1302,
    n242
  );


  buf
  g1114
  (
    n1311,
    n235
  );


  not
  g1115
  (
    n693,
    n148
  );


  buf
  g1116
  (
    n1037,
    n332
  );


  buf
  g1117
  (
    n1442,
    n379
  );


  not
  g1118
  (
    n1265,
    n308
  );


  buf
  g1119
  (
    n613,
    n153
  );


  not
  g1120
  (
    n1228,
    n261
  );


  buf
  g1121
  (
    n663,
    n205
  );


  not
  g1122
  (
    n523,
    n368
  );


  not
  g1123
  (
    n797,
    n374
  );


  buf
  g1124
  (
    n633,
    n254
  );


  not
  g1125
  (
    n748,
    n319
  );


  not
  g1126
  (
    n673,
    n336
  );


  not
  g1127
  (
    n1048,
    n265
  );


  not
  g1128
  (
    n1080,
    n284
  );


  not
  g1129
  (
    n1246,
    n150
  );


  buf
  g1130
  (
    n610,
    n243
  );


  not
  g1131
  (
    n741,
    n238
  );


  not
  g1132
  (
    n1434,
    n212
  );


  buf
  g1133
  (
    n961,
    n200
  );


  buf
  g1134
  (
    n758,
    n382
  );


  buf
  g1135
  (
    n601,
    n305
  );


  buf
  g1136
  (
    n607,
    n310
  );


  not
  g1137
  (
    n849,
    n155
  );


  not
  g1138
  (
    n1335,
    n339
  );


  buf
  g1139
  (
    n684,
    n335
  );


  buf
  g1140
  (
    n1200,
    n347
  );


  buf
  g1141
  (
    n836,
    n136
  );


  buf
  g1142
  (
    n801,
    n377
  );


  buf
  g1143
  (
    n547,
    n154
  );


  buf
  g1144
  (
    n590,
    n377
  );


  not
  g1145
  (
    n840,
    n297
  );


  buf
  g1146
  (
    n1049,
    n283
  );


  buf
  g1147
  (
    n794,
    n387
  );


  not
  g1148
  (
    n749,
    n185
  );


  not
  g1149
  (
    n930,
    n174
  );


  buf
  g1150
  (
    n578,
    n303
  );


  not
  g1151
  (
    n1055,
    n148
  );


  buf
  g1152
  (
    n1130,
    n322
  );


  buf
  g1153
  (
    n1424,
    n141
  );


  not
  g1154
  (
    n1028,
    n255
  );


  buf
  g1155
  (
    n1038,
    n241
  );


  not
  g1156
  (
    n960,
    n305
  );


  not
  g1157
  (
    n1467,
    n338
  );


  not
  g1158
  (
    n1412,
    n227
  );


  not
  g1159
  (
    n756,
    n277
  );


  not
  g1160
  (
    n1387,
    n199
  );


  buf
  g1161
  (
    n1159,
    n264
  );


  buf
  g1162
  (
    n1245,
    n171
  );


  not
  g1163
  (
    n1158,
    n373
  );


  not
  g1164
  (
    n1218,
    n381
  );


  not
  g1165
  (
    n953,
    n213
  );


  not
  g1166
  (
    n1151,
    n368
  );


  buf
  g1167
  (
    n907,
    n233
  );


  buf
  g1168
  (
    n898,
    n140
  );


  buf
  g1169
  (
    n817,
    n335
  );


  buf
  g1170
  (
    n1081,
    n345
  );


  not
  g1171
  (
    n1379,
    n334
  );


  not
  g1172
  (
    n730,
    n122
  );


  buf
  g1173
  (
    n1344,
    n138
  );


  buf
  g1174
  (
    n581,
    n372
  );


  not
  g1175
  (
    n894,
    n251
  );


  buf
  g1176
  (
    n1405,
    n237
  );


  buf
  g1177
  (
    n752,
    n270
  );


  buf
  g1178
  (
    n891,
    n123
  );


  not
  g1179
  (
    n1256,
    n193
  );


  not
  g1180
  (
    n718,
    n217
  );


  not
  g1181
  (
    n1171,
    n247
  );


  buf
  g1182
  (
    n1292,
    n153
  );


  not
  g1183
  (
    n1199,
    n316
  );


  not
  g1184
  (
    n549,
    n358
  );


  not
  g1185
  (
    n753,
    n330
  );


  buf
  g1186
  (
    n837,
    n135
  );


  buf
  g1187
  (
    n778,
    n351
  );


  buf
  g1188
  (
    n525,
    n358
  );


  not
  g1189
  (
    n1195,
    n149
  );


  buf
  g1190
  (
    n1127,
    n389
  );


  buf
  g1191
  (
    n920,
    n340
  );


  buf
  g1192
  (
    n520,
    n253
  );


  not
  g1193
  (
    n864,
    n131
  );


  not
  g1194
  (
    n1007,
    n187
  );


  not
  g1195
  (
    n661,
    n307
  );


  buf
  g1196
  (
    KeyWire_0_21,
    n317
  );


  buf
  g1197
  (
    n760,
    n324
  );


  buf
  g1198
  (
    n611,
    n166
  );


  not
  g1199
  (
    n1485,
    n166
  );


  not
  g1200
  (
    n504,
    n356
  );


  buf
  g1201
  (
    n744,
    n210
  );


  buf
  g1202
  (
    n1222,
    n378
  );


  buf
  g1203
  (
    n1065,
    n202
  );


  not
  g1204
  (
    n958,
    n344
  );


  not
  g1205
  (
    n1209,
    n248
  );


  not
  g1206
  (
    n680,
    n234
  );


  buf
  g1207
  (
    n816,
    n259
  );


  not
  g1208
  (
    n702,
    n375
  );


  buf
  g1209
  (
    n1329,
    n270
  );


  buf
  g1210
  (
    n853,
    n266
  );


  buf
  g1211
  (
    n1421,
    n195
  );


  buf
  g1212
  (
    n775,
    n154
  );


  buf
  g1213
  (
    n1444,
    n207
  );


  buf
  g1214
  (
    n1026,
    n361
  );


  not
  g1215
  (
    n917,
    n359
  );


  not
  g1216
  (
    n1083,
    n356
  );


  buf
  g1217
  (
    n1238,
    n263
  );


  not
  g1218
  (
    n769,
    n280
  );


  not
  g1219
  (
    n651,
    n141
  );


  buf
  g1220
  (
    n841,
    n271
  );


  buf
  g1221
  (
    n999,
    n195
  );


  not
  g1222
  (
    n977,
    n267
  );


  buf
  g1223
  (
    n1364,
    n285
  );


  not
  g1224
  (
    n583,
    n156
  );


  buf
  g1225
  (
    n1000,
    n277
  );


  buf
  g1226
  (
    n814,
    n330
  );


  buf
  g1227
  (
    n1102,
    n300
  );


  not
  g1228
  (
    n544,
    n139
  );


  buf
  g1229
  (
    n949,
    n178
  );


  not
  g1230
  (
    n1110,
    n165
  );


  buf
  g1231
  (
    n766,
    n235
  );


  not
  g1232
  (
    n668,
    n251
  );


  not
  g1233
  (
    n1252,
    n366
  );


  buf
  g1234
  (
    n1221,
    n362
  );


  buf
  g1235
  (
    n1116,
    n309
  );


  buf
  g1236
  (
    n762,
    n288
  );


  buf
  g1237
  (
    n934,
    n317
  );


  not
  g1238
  (
    n706,
    n297
  );


  not
  g1239
  (
    n666,
    n351
  );


  not
  g1240
  (
    n1321,
    n337
  );


  buf
  g1241
  (
    n1451,
    n192
  );


  buf
  g1242
  (
    n1294,
    n334
  );


  buf
  g1243
  (
    n1163,
    n199
  );


  buf
  g1244
  (
    n911,
    n353
  );


  buf
  g1245
  (
    n658,
    n279
  );


  not
  g1246
  (
    n1280,
    n366
  );


  buf
  g1247
  (
    n1427,
    n229
  );


  not
  g1248
  (
    n832,
    n278
  );


  not
  g1249
  (
    n1147,
    n179
  );


  buf
  g1250
  (
    n979,
    n371
  );


  buf
  g1251
  (
    n1417,
    n349
  );


  buf
  g1252
  (
    n997,
    n384
  );


  not
  g1253
  (
    n945,
    n302
  );


  buf
  g1254
  (
    n1338,
    n309
  );


  buf
  g1255
  (
    n1059,
    n358
  );


  buf
  g1256
  (
    n695,
    n381
  );


  not
  g1257
  (
    n1092,
    n140
  );


  buf
  g1258
  (
    n1291,
    n177
  );


  buf
  g1259
  (
    n962,
    n220
  );


  buf
  g1260
  (
    n1267,
    n236
  );


  buf
  g1261
  (
    n1243,
    n159
  );


  buf
  g1262
  (
    n1095,
    n157
  );


  not
  g1263
  (
    n716,
    n270
  );


  buf
  g1264
  (
    n614,
    n189
  );


  not
  g1265
  (
    n617,
    n299
  );


  buf
  g1266
  (
    n1260,
    n298
  );


  buf
  g1267
  (
    n612,
    n231
  );


  not
  g1268
  (
    n1322,
    n355
  );


  buf
  g1269
  (
    n1328,
    n205
  );


  not
  g1270
  (
    n1458,
    n208
  );


  not
  g1271
  (
    n870,
    n148
  );


  not
  g1272
  (
    n1073,
    n321
  );


  not
  g1273
  (
    n1339,
    n215
  );


  not
  g1274
  (
    n1408,
    n179
  );


  buf
  g1275
  (
    KeyWire_0_24,
    n321
  );


  not
  g1276
  (
    n694,
    n166
  );


  not
  g1277
  (
    n868,
    n122
  );


  not
  g1278
  (
    n965,
    n200
  );


  not
  g1279
  (
    n670,
    n381
  );


  not
  g1280
  (
    n1154,
    n301
  );


  not
  g1281
  (
    n1341,
    n328
  );


  buf
  g1282
  (
    n809,
    n372
  );


  buf
  g1283
  (
    n1183,
    n257
  );


  buf
  g1284
  (
    n560,
    n370
  );


  buf
  g1285
  (
    n1005,
    n355
  );


  not
  g1286
  (
    n839,
    n364
  );


  buf
  g1287
  (
    n1125,
    n343
  );


  buf
  g1288
  (
    n1136,
    n187
  );


  not
  g1289
  (
    n1131,
    n123
  );


  not
  g1290
  (
    n771,
    n198
  );


  buf
  g1291
  (
    n592,
    n218
  );


  buf
  g1292
  (
    n602,
    n207
  );


  buf
  g1293
  (
    n854,
    n230
  );


  buf
  g1294
  (
    n1432,
    n164
  );


  not
  g1295
  (
    n558,
    n307
  );


  not
  g1296
  (
    n1369,
    n210
  );


  not
  g1297
  (
    n1178,
    n374
  );


  buf
  g1298
  (
    n802,
    n322
  );


  not
  g1299
  (
    n1430,
    n162
  );


  not
  g1300
  (
    n1276,
    n206
  );


  not
  g1301
  (
    n1008,
    n352
  );


  not
  g1302
  (
    n1327,
    n145
  );


  not
  g1303
  (
    n720,
    n286
  );


  buf
  g1304
  (
    n734,
    n329
  );


  buf
  g1305
  (
    n827,
    n233
  );


  not
  g1306
  (
    n1030,
    n357
  );


  buf
  g1307
  (
    n1307,
    n275
  );


  not
  g1308
  (
    n1062,
    n312
  );


  buf
  g1309
  (
    n933,
    n382
  );


  buf
  g1310
  (
    n1465,
    n236
  );


  buf
  g1311
  (
    n600,
    n364
  );


  buf
  g1312
  (
    n648,
    n236
  );


  not
  g1313
  (
    n1115,
    n222
  );


  not
  g1314
  (
    n1351,
    n271
  );


  not
  g1315
  (
    n929,
    n171
  );


  not
  g1316
  (
    n1143,
    n225
  );


  not
  g1317
  (
    n728,
    n145
  );


  not
  g1318
  (
    n967,
    n356
  );


  buf
  g1319
  (
    n1187,
    n130
  );


  not
  g1320
  (
    n1140,
    n190
  );


  not
  g1321
  (
    n543,
    n315
  );


  buf
  g1322
  (
    n665,
    n238
  );


  not
  g1323
  (
    n824,
    n231
  );


  not
  g1324
  (
    n556,
    n130
  );


  not
  g1325
  (
    n1390,
    n190
  );


  buf
  g1326
  (
    n1105,
    n308
  );


  not
  g1327
  (
    n914,
    n339
  );


  buf
  g1328
  (
    n1174,
    n162
  );


  not
  g1329
  (
    n807,
    n332
  );


  buf
  g1330
  (
    n1229,
    n312
  );


  buf
  g1331
  (
    n637,
    n246
  );


  buf
  g1332
  (
    n901,
    n323
  );


  buf
  g1333
  (
    n1075,
    n314
  );


  not
  g1334
  (
    n1349,
    n185
  );


  not
  g1335
  (
    n699,
    n200
  );


  not
  g1336
  (
    n1429,
    n363
  );


  buf
  g1337
  (
    n1024,
    n146
  );


  not
  g1338
  (
    n705,
    n324
  );


  buf
  g1339
  (
    n885,
    n132
  );


  buf
  g1340
  (
    n1152,
    n280
  );


  buf
  g1341
  (
    n1318,
    n278
  );


  not
  g1342
  (
    n935,
    n218
  );


  not
  g1343
  (
    n785,
    n219
  );


  buf
  g1344
  (
    n729,
    n168
  );


  not
  g1345
  (
    n1223,
    n304
  );


  buf
  g1346
  (
    n1413,
    n157
  );


  buf
  g1347
  (
    n1139,
    n163
  );


  buf
  g1348
  (
    n848,
    n310
  );


  not
  g1349
  (
    n1108,
    n158
  );


  buf
  g1350
  (
    n1226,
    n243
  );


  not
  g1351
  (
    n551,
    n305
  );


  buf
  g1352
  (
    n1422,
    n260
  );


  buf
  g1353
  (
    n567,
    n127
  );


  not
  g1354
  (
    n1474,
    n383
  );


  not
  g1355
  (
    n1180,
    n151
  );


  buf
  g1356
  (
    n1394,
    n162
  );


  not
  g1357
  (
    n1431,
    n134
  );


  not
  g1358
  (
    n796,
    n223
  );


  buf
  g1359
  (
    n1191,
    n215
  );


  not
  g1360
  (
    n783,
    n265
  );


  buf
  g1361
  (
    n570,
    n237
  );


  not
  g1362
  (
    n579,
    n158
  );


  not
  g1363
  (
    n1358,
    n349
  );


  not
  g1364
  (
    n541,
    n293
  );


  buf
  g1365
  (
    n557,
    n361
  );


  buf
  g1366
  (
    n1111,
    n313
  );


  not
  g1367
  (
    n1165,
    n202
  );


  not
  g1368
  (
    n1355,
    n258
  );


  not
  g1369
  (
    n1067,
    n134
  );


  buf
  g1370
  (
    n932,
    n380
  );


  not
  g1371
  (
    n1224,
    n386
  );


  not
  g1372
  (
    n1104,
    n316
  );


  not
  g1373
  (
    n1103,
    n360
  );


  not
  g1374
  (
    n1176,
    n319
  );


  buf
  g1375
  (
    n697,
    n317
  );


  buf
  g1376
  (
    n591,
    n377
  );


  and
  g1377
  (
    n1359,
    n338,
    n196
  );


  and
  g1378
  (
    n1041,
    n285,
    n297
  );


  xnor
  g1379
  (
    n732,
    n375,
    n146
  );


  and
  g1380
  (
    n717,
    n290,
    n268
  );


  xor
  g1381
  (
    n767,
    n334,
    n201
  );


  xor
  g1382
  (
    n710,
    n251,
    n383
  );


  and
  g1383
  (
    n733,
    n211,
    n284
  );


  xor
  g1384
  (
    n980,
    n384,
    n184
  );


  xor
  g1385
  (
    n1166,
    n246,
    n221
  );


  or
  g1386
  (
    n963,
    n206,
    n173
  );


  xnor
  g1387
  (
    n913,
    n153,
    n201
  );


  nand
  g1388
  (
    n512,
    n245,
    n269
  );


  xnor
  g1389
  (
    KeyWire_0_10,
    n274,
    n378
  );


  nor
  g1390
  (
    n1401,
    n284,
    n187
  );


  nand
  g1391
  (
    n978,
    n333,
    n326
  );


  and
  g1392
  (
    n585,
    n336,
    n322
  );


  nor
  g1393
  (
    n638,
    n226,
    n256
  );


  and
  g1394
  (
    n755,
    n186,
    n148
  );


  and
  g1395
  (
    n606,
    n155,
    n249
  );


  nand
  g1396
  (
    n1179,
    n135,
    n268
  );


  xor
  g1397
  (
    n947,
    n258,
    n318
  );


  and
  g1398
  (
    n1088,
    n273,
    n332
  );


  xnor
  g1399
  (
    n1208,
    n266,
    n253
  );


  or
  g1400
  (
    n1418,
    n235,
    n341
  );


  or
  g1401
  (
    n948,
    n354,
    n167
  );


  nor
  g1402
  (
    n1441,
    n142,
    n317
  );


  and
  g1403
  (
    KeyWire_0_27,
    n137,
    n165
  );


  xor
  g1404
  (
    n966,
    n228,
    n177
  );


  xor
  g1405
  (
    n1036,
    n247,
    n129
  );


  nand
  g1406
  (
    n1301,
    n328,
    n198
  );


  nor
  g1407
  (
    n1381,
    n272,
    n229
  );


  and
  g1408
  (
    n982,
    n209,
    n181
  );


  or
  g1409
  (
    n1415,
    n370,
    n124
  );


  xnor
  g1410
  (
    n536,
    n325,
    n173
  );


  xnor
  g1411
  (
    n1002,
    n346,
    n310
  );


  nand
  g1412
  (
    n629,
    n287,
    n154
  );


  nor
  g1413
  (
    n852,
    n316,
    n286
  );


  nand
  g1414
  (
    n923,
    n177,
    n261
  );


  nand
  g1415
  (
    n683,
    n330,
    n354
  );


  nor
  g1416
  (
    n1198,
    n201,
    n264
  );


  and
  g1417
  (
    n1169,
    n253,
    n308
  );


  nor
  g1418
  (
    n622,
    n292,
    n182
  );


  nor
  g1419
  (
    n955,
    n326,
    n291
  );


  nor
  g1420
  (
    n1068,
    n307,
    n274
  );


  nor
  g1421
  (
    n1448,
    n278,
    n294
  );


  xor
  g1422
  (
    n968,
    n248,
    n168
  );


  nor
  g1423
  (
    n1266,
    n131,
    n124
  );


  and
  g1424
  (
    n776,
    n213,
    n270
  );


  nand
  g1425
  (
    n712,
    n207,
    n296
  );


  xor
  g1426
  (
    n1177,
    n319,
    n129
  );


  or
  g1427
  (
    n508,
    n212,
    n285
  );


  and
  g1428
  (
    n1101,
    n309,
    n323
  );


  nor
  g1429
  (
    n1247,
    n141,
    n160
  );


  xor
  g1430
  (
    n649,
    n223,
    n263
  );


  xor
  g1431
  (
    n742,
    n373,
    n180
  );


  nand
  g1432
  (
    n1233,
    n214,
    n289
  );


  xnor
  g1433
  (
    n725,
    n323,
    n365
  );


  and
  g1434
  (
    n987,
    n256,
    n194
  );


  nand
  g1435
  (
    n624,
    n126,
    n252
  );


  nand
  g1436
  (
    n1060,
    n137,
    n284
  );


  nor
  g1437
  (
    n731,
    n370,
    n305
  );


  nand
  g1438
  (
    n1079,
    n137,
    n202
  );


  nor
  g1439
  (
    n691,
    n243,
    n374
  );


  nand
  g1440
  (
    n1141,
    n201,
    n124
  );


  or
  g1441
  (
    n1196,
    n125,
    n265
  );


  nand
  g1442
  (
    n1462,
    n128,
    n154
  );


  nand
  g1443
  (
    n937,
    n231,
    n312
  );


  or
  g1444
  (
    n795,
    n241,
    n123
  );


  xor
  g1445
  (
    n1214,
    n328,
    n380
  );


  or
  g1446
  (
    n1303,
    n280,
    n165
  );


  xnor
  g1447
  (
    n1070,
    n143,
    n368
  );


  or
  g1448
  (
    n1287,
    n381,
    n367
  );


  and
  g1449
  (
    n1337,
    n244,
    n347
  );


  xnor
  g1450
  (
    n1436,
    n214,
    n359
  );


  nor
  g1451
  (
    n1397,
    n308,
    n348
  );


  nand
  g1452
  (
    n530,
    n325,
    n135
  );


  xor
  g1453
  (
    n805,
    n298,
    n131
  );


  or
  g1454
  (
    n1309,
    n274,
    n298
  );


  and
  g1455
  (
    n990,
    n329,
    n377
  );


  nand
  g1456
  (
    n1032,
    n149,
    n155
  );


  xnor
  g1457
  (
    n750,
    n144,
    n360
  );


  nor
  g1458
  (
    n939,
    n369,
    n347
  );


  xnor
  g1459
  (
    n1255,
    n331,
    n136
  );


  xor
  g1460
  (
    n656,
    n382,
    n297
  );


  or
  g1461
  (
    n943,
    n236,
    n364
  );


  and
  g1462
  (
    n772,
    n302,
    n162
  );


  nor
  g1463
  (
    n951,
    n296,
    n189
  );


  not
  g1464
  (
    n1498,
    n514
  );


  buf
  g1465
  (
    n1496,
    n524
  );


  buf
  g1466
  (
    n1492,
    n509
  );


  not
  g1467
  (
    n1504,
    n523
  );


  buf
  g1468
  (
    n1499,
    n504
  );


  not
  g1469
  (
    n1489,
    n515
  );


  buf
  g1470
  (
    n1502,
    n527
  );


  not
  g1471
  (
    n1501,
    n518
  );


  buf
  g1472
  (
    n1495,
    n507
  );


  buf
  g1473
  (
    n1497,
    n502
  );


  not
  g1474
  (
    n1494,
    n516
  );


  buf
  g1475
  (
    n1490,
    n510
  );


  xor
  g1476
  (
    n1491,
    n521,
    n512,
    n520,
    n513
  );


  xnor
  g1477
  (
    n1493,
    n506,
    n503,
    n522,
    n508
  );


  xnor
  g1478
  (
    n1503,
    n528,
    n517,
    n505,
    n511
  );


  xnor
  g1479
  (
    n1500,
    n525,
    n526,
    n519,
    n529
  );


  not
  g1480
  (
    n1527,
    n1498
  );


  not
  g1481
  (
    n1518,
    n1501
  );


  not
  g1482
  (
    n1534,
    n1491
  );


  buf
  g1483
  (
    n1508,
    n1489
  );


  buf
  g1484
  (
    n1528,
    n1499
  );


  buf
  g1485
  (
    n1533,
    n1502
  );


  not
  g1486
  (
    n1532,
    n1501
  );


  not
  g1487
  (
    n1523,
    n1503
  );


  buf
  g1488
  (
    n1505,
    n1499
  );


  not
  g1489
  (
    n1529,
    n1498
  );


  not
  g1490
  (
    n1522,
    n1498
  );


  not
  g1491
  (
    n1520,
    n1495
  );


  not
  g1492
  (
    n1514,
    n1499
  );


  not
  g1493
  (
    n1517,
    n1501
  );


  not
  g1494
  (
    n1509,
    n1498
  );


  not
  g1495
  (
    n1510,
    n1500
  );


  not
  g1496
  (
    n1512,
    n1499
  );


  not
  g1497
  (
    n1526,
    n1493
  );


  buf
  g1498
  (
    n1525,
    n1494
  );


  not
  g1499
  (
    n1513,
    n1502
  );


  buf
  g1500
  (
    n1521,
    n1500
  );


  not
  g1501
  (
    n1530,
    n1496
  );


  buf
  g1502
  (
    n1515,
    n1502
  );


  not
  g1503
  (
    n1511,
    n1500
  );


  not
  g1504
  (
    n1531,
    n1501
  );


  not
  g1505
  (
    n1524,
    n1497
  );


  buf
  g1506
  (
    n1506,
    n1492
  );


  not
  g1507
  (
    n1507,
    n1490
  );


  not
  g1508
  (
    n1516,
    n1502
  );


  buf
  g1509
  (
    n1519,
    n1500
  );


  buf
  g1510
  (
    n1565,
    n1532
  );


  not
  g1511
  (
    n1552,
    n1528
  );


  buf
  g1512
  (
    n1607,
    n1522
  );


  buf
  g1513
  (
    n1557,
    n1508
  );


  not
  g1514
  (
    n1586,
    n1519
  );


  buf
  g1515
  (
    n1560,
    n1531
  );


  not
  g1516
  (
    n1548,
    n1518
  );


  buf
  g1517
  (
    n1641,
    n1508
  );


  not
  g1518
  (
    n1577,
    n1510
  );


  not
  g1519
  (
    n1640,
    n1534
  );


  not
  g1520
  (
    n1626,
    n1507
  );


  not
  g1521
  (
    n1608,
    n1527
  );


  buf
  g1522
  (
    n1570,
    n1516
  );


  not
  g1523
  (
    n1553,
    n1514
  );


  buf
  g1524
  (
    n1591,
    n1504
  );


  buf
  g1525
  (
    n1623,
    n1519
  );


  buf
  g1526
  (
    n1631,
    n1522
  );


  buf
  g1527
  (
    n1582,
    n1524
  );


  not
  g1528
  (
    n1619,
    n1530
  );


  not
  g1529
  (
    n1618,
    n1511
  );


  not
  g1530
  (
    n1601,
    n1515
  );


  not
  g1531
  (
    n1537,
    n1530
  );


  not
  g1532
  (
    n1599,
    n1517
  );


  not
  g1533
  (
    n1540,
    n1519
  );


  not
  g1534
  (
    n1651,
    n1524
  );


  buf
  g1535
  (
    n1654,
    n1529
  );


  not
  g1536
  (
    n1544,
    n1508
  );


  buf
  g1537
  (
    n1632,
    n1507
  );


  buf
  g1538
  (
    n1612,
    n1509
  );


  not
  g1539
  (
    n1593,
    n1517
  );


  buf
  g1540
  (
    n1606,
    n1523
  );


  buf
  g1541
  (
    n1539,
    n1523
  );


  buf
  g1542
  (
    n1638,
    n1508
  );


  buf
  g1543
  (
    n1590,
    n1513
  );


  buf
  g1544
  (
    n1580,
    n1530
  );


  buf
  g1545
  (
    n1653,
    n1529
  );


  not
  g1546
  (
    n1614,
    n1519
  );


  not
  g1547
  (
    n1652,
    n1515
  );


  not
  g1548
  (
    n1541,
    n1523
  );


  not
  g1549
  (
    n1643,
    n1531
  );


  buf
  g1550
  (
    n1551,
    n1526
  );


  buf
  g1551
  (
    n1648,
    n1516
  );


  buf
  g1552
  (
    n1579,
    n1518
  );


  not
  g1553
  (
    n1639,
    n1518
  );


  not
  g1554
  (
    n1636,
    n1504
  );


  buf
  g1555
  (
    n1535,
    n1528
  );


  buf
  g1556
  (
    n1566,
    n1525
  );


  not
  g1557
  (
    n1545,
    n1526
  );


  not
  g1558
  (
    n1562,
    n1524
  );


  buf
  g1559
  (
    n1635,
    n1503
  );


  buf
  g1560
  (
    n1620,
    n1514
  );


  buf
  g1561
  (
    n1568,
    n1504
  );


  not
  g1562
  (
    n1574,
    n1533
  );


  buf
  g1563
  (
    n1611,
    n1528
  );


  not
  g1564
  (
    n1613,
    n1512
  );


  not
  g1565
  (
    n1609,
    n1532
  );


  not
  g1566
  (
    n1555,
    n1507
  );


  not
  g1567
  (
    n1584,
    n1517
  );


  buf
  g1568
  (
    n1538,
    n1514
  );


  not
  g1569
  (
    n1646,
    n1505
  );


  not
  g1570
  (
    n1558,
    n1533
  );


  not
  g1571
  (
    n1616,
    n1506
  );


  not
  g1572
  (
    n1576,
    n1523
  );


  not
  g1573
  (
    n1628,
    n1512
  );


  not
  g1574
  (
    n1634,
    n1532
  );


  buf
  g1575
  (
    n1645,
    n1529
  );


  buf
  g1576
  (
    n1542,
    n1514
  );


  not
  g1577
  (
    n1603,
    n1516
  );


  buf
  g1578
  (
    n1595,
    n1513
  );


  buf
  g1579
  (
    KeyWire_0_25,
    n1520
  );


  not
  g1580
  (
    n1561,
    n1529
  );


  buf
  g1581
  (
    n1602,
    n1506
  );


  buf
  g1582
  (
    n1617,
    n1522
  );


  buf
  g1583
  (
    n1642,
    n1510
  );


  not
  g1584
  (
    n1647,
    n1512
  );


  not
  g1585
  (
    n1546,
    n1506
  );


  not
  g1586
  (
    n1564,
    n1531
  );


  buf
  g1587
  (
    n1581,
    n1513
  );


  buf
  g1588
  (
    n1594,
    n1505
  );


  buf
  g1589
  (
    n1571,
    n1521
  );


  buf
  g1590
  (
    n1536,
    n1520
  );


  not
  g1591
  (
    n1588,
    n1526
  );


  buf
  g1592
  (
    n1650,
    n1527
  );


  buf
  g1593
  (
    n1621,
    n1532
  );


  not
  g1594
  (
    n1630,
    n1533
  );


  not
  g1595
  (
    n1592,
    n1520
  );


  not
  g1596
  (
    n1567,
    n1505
  );


  buf
  g1597
  (
    n1610,
    n1525
  );


  buf
  g1598
  (
    n1598,
    n1507
  );


  not
  g1599
  (
    n1543,
    n1525
  );


  buf
  g1600
  (
    n1587,
    n1521
  );


  buf
  g1601
  (
    n1649,
    n1512
  );


  buf
  g1602
  (
    n1622,
    n1505
  );


  not
  g1603
  (
    n1583,
    n1517
  );


  buf
  g1604
  (
    n1633,
    n1534
  );


  buf
  g1605
  (
    n1604,
    n1509
  );


  not
  g1606
  (
    n1575,
    n1534
  );


  buf
  g1607
  (
    n1547,
    n1525
  );


  buf
  g1608
  (
    n1585,
    n1511
  );


  buf
  g1609
  (
    n1600,
    n1509
  );


  not
  g1610
  (
    n1550,
    n1511
  );


  buf
  g1611
  (
    n1549,
    n1521
  );


  not
  g1612
  (
    n1625,
    n1530
  );


  buf
  g1613
  (
    n1572,
    n1503
  );


  not
  g1614
  (
    n1569,
    n1518
  );


  buf
  g1615
  (
    n1627,
    n1513
  );


  not
  g1616
  (
    n1563,
    n1533
  );


  buf
  g1617
  (
    n1589,
    n1524
  );


  buf
  g1618
  (
    n1644,
    n1527
  );


  buf
  g1619
  (
    n1578,
    n1506
  );


  not
  g1620
  (
    n1596,
    n1527
  );


  buf
  g1621
  (
    n1573,
    n1531
  );


  not
  g1622
  (
    n1624,
    n1503
  );


  nand
  g1623
  (
    n1554,
    n1521,
    n1516
  );


  and
  g1624
  (
    n1559,
    n1510,
    n1504
  );


  nor
  g1625
  (
    n1556,
    n1520,
    n1515
  );


  and
  g1626
  (
    n1637,
    n1528,
    n1511
  );


  nor
  g1627
  (
    n1597,
    n1509,
    n1522
  );


  xnor
  g1628
  (
    n1605,
    n1534,
    n1510
  );


  and
  g1629
  (
    n1615,
    n1515,
    n1526
  );


  buf
  g1630
  (
    n1863,
    n1606
  );


  buf
  g1631
  (
    n1967,
    n1647
  );


  not
  g1632
  (
    n2062,
    n1602
  );


  buf
  g1633
  (
    n1873,
    n1614
  );


  not
  g1634
  (
    n1879,
    n1632
  );


  not
  g1635
  (
    n2009,
    n1582
  );


  not
  g1636
  (
    n2128,
    n1614
  );


  buf
  g1637
  (
    n1936,
    n1641
  );


  not
  g1638
  (
    n1991,
    n1623
  );


  buf
  g1639
  (
    n2122,
    n1645
  );


  not
  g1640
  (
    n1862,
    n1589
  );


  not
  g1641
  (
    n1881,
    n1627
  );


  buf
  g1642
  (
    n2080,
    n1544
  );


  not
  g1643
  (
    n1833,
    n1559
  );


  not
  g1644
  (
    n1885,
    n1586
  );


  buf
  g1645
  (
    n1770,
    n1599
  );


  not
  g1646
  (
    n1753,
    n1604
  );


  buf
  g1647
  (
    n1840,
    n1600
  );


  not
  g1648
  (
    n1791,
    n1565
  );


  buf
  g1649
  (
    n2048,
    n1628
  );


  buf
  g1650
  (
    n2005,
    n1571
  );


  not
  g1651
  (
    n1888,
    n1645
  );


  not
  g1652
  (
    n1670,
    n1571
  );


  not
  g1653
  (
    n2041,
    n1564
  );


  not
  g1654
  (
    n2001,
    n1541
  );


  buf
  g1655
  (
    n1868,
    n1613
  );


  not
  g1656
  (
    n1695,
    n1570
  );


  not
  g1657
  (
    n2015,
    n1552
  );


  not
  g1658
  (
    n1864,
    n1645
  );


  buf
  g1659
  (
    n1766,
    n1651
  );


  buf
  g1660
  (
    n1929,
    n1626
  );


  not
  g1661
  (
    n1758,
    n1571
  );


  not
  g1662
  (
    n1886,
    n1589
  );


  not
  g1663
  (
    n2091,
    n1600
  );


  not
  g1664
  (
    n1764,
    n1616
  );


  buf
  g1665
  (
    n1836,
    n1574
  );


  not
  g1666
  (
    n2099,
    n1643
  );


  not
  g1667
  (
    n1801,
    n1588
  );


  buf
  g1668
  (
    n1997,
    n1585
  );


  buf
  g1669
  (
    n1725,
    n1609
  );


  buf
  g1670
  (
    n1665,
    n1565
  );


  buf
  g1671
  (
    n2056,
    n1622
  );


  not
  g1672
  (
    n1706,
    n1627
  );


  buf
  g1673
  (
    n2025,
    n1629
  );


  not
  g1674
  (
    n2011,
    n1651
  );


  not
  g1675
  (
    n1760,
    n1638
  );


  not
  g1676
  (
    n1702,
    n1652
  );


  buf
  g1677
  (
    KeyWire_0_22,
    n1644
  );


  not
  g1678
  (
    n1923,
    n1624
  );


  buf
  g1679
  (
    n1950,
    n1619
  );


  not
  g1680
  (
    n1955,
    n1640
  );


  not
  g1681
  (
    n1690,
    n1568
  );


  not
  g1682
  (
    n1907,
    n1589
  );


  not
  g1683
  (
    n1804,
    n1567
  );


  buf
  g1684
  (
    n1975,
    n1553
  );


  buf
  g1685
  (
    n1932,
    n1554
  );


  buf
  g1686
  (
    n1747,
    n1550
  );


  buf
  g1687
  (
    n1931,
    n1611
  );


  not
  g1688
  (
    n2109,
    n1611
  );


  not
  g1689
  (
    n1782,
    n1643
  );


  buf
  g1690
  (
    n1847,
    n1593
  );


  buf
  g1691
  (
    n2077,
    n1632
  );


  buf
  g1692
  (
    n1814,
    n1601
  );


  not
  g1693
  (
    n1780,
    n1587
  );


  not
  g1694
  (
    n1977,
    n1572
  );


  not
  g1695
  (
    n2112,
    n1581
  );


  buf
  g1696
  (
    n2007,
    n1646
  );


  buf
  g1697
  (
    n2035,
    n1551
  );


  buf
  g1698
  (
    n1812,
    n1635
  );


  not
  g1699
  (
    n1943,
    n1639
  );


  buf
  g1700
  (
    n1984,
    n1575
  );


  not
  g1701
  (
    n1948,
    n1561
  );


  buf
  g1702
  (
    n1867,
    n1577
  );


  not
  g1703
  (
    n1820,
    n1617
  );


  buf
  g1704
  (
    n2093,
    n1605
  );


  not
  g1705
  (
    n1857,
    n1580
  );


  buf
  g1706
  (
    n1785,
    n1577
  );


  buf
  g1707
  (
    n1743,
    n1641
  );


  not
  g1708
  (
    n2117,
    n1604
  );


  buf
  g1709
  (
    n2051,
    n1553
  );


  buf
  g1710
  (
    n1774,
    n1622
  );


  buf
  g1711
  (
    n1754,
    n1550
  );


  buf
  g1712
  (
    n1667,
    n1562
  );


  buf
  g1713
  (
    n1998,
    n1605
  );


  not
  g1714
  (
    n1749,
    n1639
  );


  buf
  g1715
  (
    n2076,
    n1583
  );


  buf
  g1716
  (
    n1876,
    n1567
  );


  not
  g1717
  (
    n1808,
    n1573
  );


  not
  g1718
  (
    KeyWire_0_4,
    n1604
  );


  buf
  g1719
  (
    n2075,
    n1557
  );


  buf
  g1720
  (
    n2124,
    n1614
  );


  buf
  g1721
  (
    n1687,
    n1580
  );


  not
  g1722
  (
    n1976,
    n1556
  );


  not
  g1723
  (
    n1821,
    n1601
  );


  not
  g1724
  (
    n2132,
    n1594
  );


  buf
  g1725
  (
    n2002,
    n1593
  );


  buf
  g1726
  (
    n2029,
    n1566
  );


  not
  g1727
  (
    n2102,
    n1637
  );


  buf
  g1728
  (
    n1918,
    n1650
  );


  not
  g1729
  (
    n1884,
    n1581
  );


  buf
  g1730
  (
    KeyWire_0_16,
    n1546
  );


  buf
  g1731
  (
    n1996,
    n1603
  );


  not
  g1732
  (
    n1656,
    n1541
  );


  not
  g1733
  (
    n1830,
    n1591
  );


  not
  g1734
  (
    n1894,
    n1578
  );


  not
  g1735
  (
    n1737,
    n1549
  );


  buf
  g1736
  (
    n1703,
    n1572
  );


  buf
  g1737
  (
    n1970,
    n1646
  );


  not
  g1738
  (
    n1889,
    n1554
  );


  not
  g1739
  (
    n1896,
    n1617
  );


  not
  g1740
  (
    n2022,
    n1543
  );


  buf
  g1741
  (
    n1824,
    n1603
  );


  not
  g1742
  (
    n1949,
    n1560
  );


  buf
  g1743
  (
    n1883,
    n1654
  );


  not
  g1744
  (
    n2018,
    n1642
  );


  buf
  g1745
  (
    n1837,
    n1620
  );


  buf
  g1746
  (
    n1783,
    n1583
  );


  buf
  g1747
  (
    n1941,
    n1572
  );


  not
  g1748
  (
    n2068,
    n1561
  );


  not
  g1749
  (
    n1979,
    n1648
  );


  not
  g1750
  (
    n1819,
    n1569
  );


  not
  g1751
  (
    n2131,
    n1555
  );


  buf
  g1752
  (
    n1887,
    n1622
  );


  buf
  g1753
  (
    n1815,
    n1536
  );


  not
  g1754
  (
    n1709,
    n1597
  );


  not
  g1755
  (
    n1963,
    n1581
  );


  not
  g1756
  (
    n1700,
    n1609
  );


  buf
  g1757
  (
    n1712,
    n1652
  );


  buf
  g1758
  (
    n1757,
    n1596
  );


  not
  g1759
  (
    n1657,
    n1556
  );


  not
  g1760
  (
    n1726,
    n1560
  );


  not
  g1761
  (
    n2033,
    n1602
  );


  not
  g1762
  (
    n1685,
    n1543
  );


  not
  g1763
  (
    n1683,
    n1590
  );


  not
  g1764
  (
    n1663,
    n1580
  );


  buf
  g1765
  (
    n1677,
    n1631
  );


  not
  g1766
  (
    n1912,
    n1553
  );


  not
  g1767
  (
    n1715,
    n1575
  );


  buf
  g1768
  (
    n1895,
    n1535
  );


  not
  g1769
  (
    n1908,
    n1542
  );


  not
  g1770
  (
    n2090,
    n1586
  );


  buf
  g1771
  (
    n1927,
    n1597
  );


  not
  g1772
  (
    n1773,
    n1565
  );


  buf
  g1773
  (
    n1865,
    n1537
  );


  not
  g1774
  (
    n1718,
    n1562
  );


  not
  g1775
  (
    n2046,
    n1633
  );


  buf
  g1776
  (
    n2012,
    n1558
  );


  not
  g1777
  (
    n1680,
    n1615
  );


  not
  g1778
  (
    n1675,
    n1633
  );


  not
  g1779
  (
    n2134,
    n1620
  );


  buf
  g1780
  (
    n1745,
    n1565
  );


  buf
  g1781
  (
    n1767,
    n1580
  );


  not
  g1782
  (
    n1696,
    n1653
  );


  not
  g1783
  (
    n2053,
    n1586
  );


  buf
  g1784
  (
    n2108,
    n1594
  );


  not
  g1785
  (
    n1826,
    n1645
  );


  not
  g1786
  (
    n1985,
    n1539
  );


  not
  g1787
  (
    n2073,
    n1605
  );


  not
  g1788
  (
    n1916,
    n1646
  );


  not
  g1789
  (
    n1871,
    n1548
  );


  not
  g1790
  (
    n1662,
    n1537
  );


  buf
  g1791
  (
    n2106,
    n1617
  );


  not
  g1792
  (
    n2127,
    n1584
  );


  not
  g1793
  (
    n1678,
    n1548
  );


  buf
  g1794
  (
    n1980,
    n1545
  );


  buf
  g1795
  (
    KeyWire_0_14,
    n1574
  );


  buf
  g1796
  (
    n1947,
    n1642
  );


  buf
  g1797
  (
    n1739,
    n1582
  );


  not
  g1798
  (
    n1856,
    n1605
  );


  buf
  g1799
  (
    n1779,
    n1628
  );


  not
  g1800
  (
    n2069,
    n1541
  );


  buf
  g1801
  (
    n1786,
    n1635
  );


  buf
  g1802
  (
    n1850,
    n1653
  );


  buf
  g1803
  (
    n1959,
    n1632
  );


  not
  g1804
  (
    n1992,
    n1614
  );


  buf
  g1805
  (
    n1874,
    n1618
  );


  buf
  g1806
  (
    n1756,
    n1649
  );


  buf
  g1807
  (
    n2032,
    n1644
  );


  buf
  g1808
  (
    n1838,
    n1609
  );


  not
  g1809
  (
    n2043,
    n1563
  );


  buf
  g1810
  (
    n2027,
    n1551
  );


  not
  g1811
  (
    n1746,
    n1570
  );


  buf
  g1812
  (
    n1831,
    n1549
  );


  not
  g1813
  (
    n1834,
    n1636
  );


  buf
  g1814
  (
    n1822,
    n1552
  );


  not
  g1815
  (
    n1939,
    n1621
  );


  buf
  g1816
  (
    n2024,
    n1547
  );


  not
  g1817
  (
    n2008,
    n1615
  );


  buf
  g1818
  (
    n2037,
    n1585
  );


  not
  g1819
  (
    n1858,
    n1589
  );


  not
  g1820
  (
    n1684,
    n1593
  );


  not
  g1821
  (
    n1828,
    n1606
  );


  not
  g1822
  (
    n1763,
    n1539
  );


  not
  g1823
  (
    n1733,
    n1616
  );


  not
  g1824
  (
    n1778,
    n1643
  );


  buf
  g1825
  (
    n2003,
    n1548
  );


  buf
  g1826
  (
    n2114,
    n1615
  );


  buf
  g1827
  (
    n1999,
    n1560
  );


  buf
  g1828
  (
    n1818,
    n1654
  );


  not
  g1829
  (
    n2105,
    n1574
  );


  not
  g1830
  (
    n1717,
    n1636
  );


  buf
  g1831
  (
    n1842,
    n1598
  );


  not
  g1832
  (
    n2071,
    n1537
  );


  buf
  g1833
  (
    n1742,
    n1642
  );


  buf
  g1834
  (
    n1915,
    n1599
  );


  not
  g1835
  (
    n2092,
    n1652
  );


  buf
  g1836
  (
    n1698,
    n1552
  );


  buf
  g1837
  (
    n1859,
    n1650
  );


  buf
  g1838
  (
    n1988,
    n1596
  );


  buf
  g1839
  (
    n1800,
    n1542
  );


  not
  g1840
  (
    n1710,
    n1555
  );


  buf
  g1841
  (
    n1679,
    n1647
  );


  not
  g1842
  (
    n1954,
    n1587
  );


  not
  g1843
  (
    n1671,
    n1612
  );


  not
  g1844
  (
    n1892,
    n1634
  );


  not
  g1845
  (
    n1669,
    n1535
  );


  not
  g1846
  (
    n1744,
    n1650
  );


  not
  g1847
  (
    n2101,
    n1634
  );


  buf
  g1848
  (
    n2126,
    n1621
  );


  buf
  g1849
  (
    n1891,
    n1575
  );


  not
  g1850
  (
    n1962,
    n1650
  );


  not
  g1851
  (
    n1655,
    n1598
  );


  buf
  g1852
  (
    n1741,
    n1637
  );


  buf
  g1853
  (
    n2030,
    n1535
  );


  not
  g1854
  (
    n1707,
    n1613
  );


  not
  g1855
  (
    n2006,
    n1606
  );


  not
  g1856
  (
    n1704,
    n1625
  );


  not
  g1857
  (
    n1969,
    n1545
  );


  not
  g1858
  (
    n1978,
    n1575
  );


  buf
  g1859
  (
    n1816,
    n1629
  );


  buf
  g1860
  (
    n1776,
    n1638
  );


  not
  g1861
  (
    n2039,
    n1616
  );


  buf
  g1862
  (
    n1901,
    n1615
  );


  not
  g1863
  (
    n2023,
    n1573
  );


  buf
  g1864
  (
    n1990,
    n1546
  );


  buf
  g1865
  (
    n1781,
    n1607
  );


  buf
  g1866
  (
    n1719,
    n1629
  );


  not
  g1867
  (
    n1953,
    n1559
  );


  not
  g1868
  (
    n1930,
    n1646
  );


  buf
  g1869
  (
    n1694,
    n1595
  );


  not
  g1870
  (
    n2067,
    n1557
  );


  buf
  g1871
  (
    n2079,
    n1637
  );


  not
  g1872
  (
    n2036,
    n1576
  );


  not
  g1873
  (
    n2017,
    n1638
  );


  not
  g1874
  (
    n1810,
    n1601
  );


  not
  g1875
  (
    n1771,
    n1573
  );


  buf
  g1876
  (
    n1900,
    n1628
  );


  not
  g1877
  (
    n2049,
    n1536
  );


  buf
  g1878
  (
    n1839,
    n1627
  );


  buf
  g1879
  (
    n2129,
    n1573
  );


  not
  g1880
  (
    n1761,
    n1630
  );


  not
  g1881
  (
    n2047,
    n1560
  );


  buf
  g1882
  (
    n1914,
    n1609
  );


  not
  g1883
  (
    n2088,
    n1607
  );


  not
  g1884
  (
    n2083,
    n1619
  );


  buf
  g1885
  (
    n1825,
    n1635
  );


  buf
  g1886
  (
    n2085,
    n1576
  );


  buf
  g1887
  (
    n1937,
    n1595
  );


  buf
  g1888
  (
    n1674,
    n1590
  );


  not
  g1889
  (
    n1995,
    n1581
  );


  not
  g1890
  (
    n1807,
    n1618
  );


  not
  g1891
  (
    n1853,
    n1612
  );


  not
  g1892
  (
    n1869,
    n1608
  );


  buf
  g1893
  (
    n1809,
    n1641
  );


  buf
  g1894
  (
    n1933,
    n1653
  );


  not
  g1895
  (
    n1668,
    n1596
  );


  not
  g1896
  (
    n2013,
    n1564
  );


  buf
  g1897
  (
    n1994,
    n1578
  );


  not
  g1898
  (
    n1806,
    n1643
  );


  buf
  g1899
  (
    n1983,
    n1547
  );


  not
  g1900
  (
    n1875,
    n1625
  );


  buf
  g1901
  (
    n1993,
    n1567
  );


  buf
  g1902
  (
    n1860,
    n1619
  );


  not
  g1903
  (
    n2087,
    n1576
  );


  not
  g1904
  (
    n2057,
    n1640
  );


  not
  g1905
  (
    n1934,
    n1593
  );


  buf
  g1906
  (
    n1788,
    n1648
  );


  buf
  g1907
  (
    n1676,
    n1566
  );


  buf
  g1908
  (
    n1795,
    n1616
  );


  buf
  g1909
  (
    n1942,
    n1537
  );


  not
  g1910
  (
    n1799,
    n1594
  );


  not
  g1911
  (
    n1673,
    n1576
  );


  buf
  g1912
  (
    n2045,
    n1651
  );


  not
  g1913
  (
    n1817,
    n1579
  );


  not
  g1914
  (
    n2054,
    n1611
  );


  not
  g1915
  (
    n1952,
    n1542
  );


  not
  g1916
  (
    n1823,
    n1587
  );


  not
  g1917
  (
    n2097,
    n1548
  );


  not
  g1918
  (
    n1987,
    n1591
  );


  buf
  g1919
  (
    n2111,
    n1600
  );


  buf
  g1920
  (
    n1713,
    n1538
  );


  buf
  g1921
  (
    n1855,
    n1599
  );


  buf
  g1922
  (
    n2123,
    n1568
  );


  not
  g1923
  (
    n2084,
    n1603
  );


  buf
  g1924
  (
    n1843,
    n1569
  );


  not
  g1925
  (
    n1692,
    n1536
  );


  buf
  g1926
  (
    n1762,
    n1617
  );


  not
  g1927
  (
    n1861,
    n1553
  );


  buf
  g1928
  (
    n1922,
    n1610
  );


  buf
  g1929
  (
    n1905,
    n1635
  );


  buf
  g1930
  (
    n1724,
    n1592
  );


  not
  g1931
  (
    n1917,
    n1618
  );


  not
  g1932
  (
    n2130,
    n1558
  );


  not
  g1933
  (
    n2089,
    n1582
  );


  buf
  g1934
  (
    n2016,
    n1584
  );


  buf
  g1935
  (
    n1708,
    n1550
  );


  not
  g1936
  (
    n1972,
    n1546
  );


  not
  g1937
  (
    n1796,
    n1597
  );


  buf
  g1938
  (
    n1666,
    n1596
  );


  not
  g1939
  (
    n2086,
    n1603
  );


  not
  g1940
  (
    n1752,
    n1546
  );


  not
  g1941
  (
    n2119,
    n1594
  );


  buf
  g1942
  (
    n1877,
    n1608
  );


  not
  g1943
  (
    n1732,
    n1606
  );


  buf
  g1944
  (
    n1841,
    n1624
  );


  not
  g1945
  (
    n1909,
    n1569
  );


  buf
  g1946
  (
    n1897,
    n1653
  );


  buf
  g1947
  (
    n1910,
    n1564
  );


  not
  g1948
  (
    n1974,
    n1639
  );


  buf
  g1949
  (
    n2082,
    n1625
  );


  not
  g1950
  (
    n2044,
    n1597
  );


  not
  g1951
  (
    n1723,
    n1566
  );


  buf
  g1952
  (
    n2010,
    n1540
  );


  buf
  g1953
  (
    n1705,
    n1549
  );


  buf
  g1954
  (
    n1924,
    n1542
  );


  not
  g1955
  (
    n2113,
    n1536
  );


  buf
  g1956
  (
    n2107,
    n1558
  );


  not
  g1957
  (
    n2133,
    n1577
  );


  buf
  g1958
  (
    n1835,
    n1578
  );


  buf
  g1959
  (
    n1716,
    n1551
  );


  not
  g1960
  (
    n2052,
    n1654
  );


  not
  g1961
  (
    n2038,
    n1637
  );


  buf
  g1962
  (
    n1787,
    n1631
  );


  buf
  g1963
  (
    n1971,
    n1535
  );


  buf
  g1964
  (
    n1701,
    n1584
  );


  buf
  g1965
  (
    n1851,
    n1622
  );


  buf
  g1966
  (
    n1768,
    n1652
  );


  buf
  g1967
  (
    n1944,
    n1578
  );


  buf
  g1968
  (
    n2081,
    n1588
  );


  buf
  g1969
  (
    n2061,
    n1568
  );


  buf
  g1970
  (
    n1870,
    n1604
  );


  not
  g1971
  (
    n1920,
    n1583
  );


  buf
  g1972
  (
    n1951,
    n1640
  );


  buf
  g1973
  (
    n1945,
    n1539
  );


  not
  g1974
  (
    n1973,
    n1638
  );


  buf
  g1975
  (
    n1769,
    n1649
  );


  not
  g1976
  (
    n1921,
    n1654
  );


  buf
  g1977
  (
    n1803,
    n1623
  );


  buf
  g1978
  (
    n1982,
    n1547
  );


  buf
  g1979
  (
    n2098,
    n1627
  );


  not
  g1980
  (
    n1890,
    n1624
  );


  buf
  g1981
  (
    n2050,
    n1538
  );


  buf
  g1982
  (
    n1872,
    n1538
  );


  buf
  g1983
  (
    n2019,
    n1570
  );


  buf
  g1984
  (
    n2014,
    n1610
  );


  buf
  g1985
  (
    n2094,
    n1624
  );


  buf
  g1986
  (
    n1904,
    n1607
  );


  not
  g1987
  (
    n1880,
    n1568
  );


  not
  g1988
  (
    n1738,
    n1567
  );


  buf
  g1989
  (
    n1956,
    n1543
  );


  not
  g1990
  (
    n1811,
    n1612
  );


  not
  g1991
  (
    n2070,
    n1572
  );


  buf
  g1992
  (
    n1813,
    n1540
  );


  buf
  g1993
  (
    n1755,
    n1649
  );


  buf
  g1994
  (
    n2060,
    n1647
  );


  buf
  g1995
  (
    n1852,
    n1554
  );


  not
  g1996
  (
    n1734,
    n1590
  );


  not
  g1997
  (
    n1965,
    n1602
  );


  buf
  g1998
  (
    n2026,
    n1579
  );


  not
  g1999
  (
    n1893,
    n1551
  );


  not
  g2000
  (
    n1693,
    n1630
  );


  buf
  g2001
  (
    n1845,
    n1538
  );


  buf
  g2002
  (
    n1784,
    n1556
  );


  not
  g2003
  (
    n2042,
    n1559
  );


  buf
  g2004
  (
    n2040,
    n1590
  );


  not
  g2005
  (
    n1829,
    n1588
  );


  not
  g2006
  (
    n1659,
    n1544
  );


  buf
  g2007
  (
    n1898,
    n1595
  );


  buf
  g2008
  (
    n2095,
    n1585
  );


  not
  g2009
  (
    n1899,
    n1591
  );


  not
  g2010
  (
    n2034,
    n1610
  );


  buf
  g2011
  (
    KeyWire_0_17,
    n1649
  );


  buf
  g2012
  (
    n1735,
    n1554
  );


  not
  g2013
  (
    n2120,
    n1561
  );


  buf
  g2014
  (
    n2031,
    n1586
  );


  not
  g2015
  (
    n1958,
    n1563
  );


  not
  g2016
  (
    n1986,
    n1544
  );


  not
  g2017
  (
    n1794,
    n1555
  );


  buf
  g2018
  (
    n1848,
    n1561
  );


  not
  g2019
  (
    n1688,
    n1651
  );


  not
  g2020
  (
    n2104,
    n1582
  );


  not
  g2021
  (
    n1938,
    n1556
  );


  not
  g2022
  (
    n2000,
    n1647
  );


  buf
  g2023
  (
    n1866,
    n1557
  );


  buf
  g2024
  (
    n2118,
    n1626
  );


  not
  g2025
  (
    n2078,
    n1636
  );


  not
  g2026
  (
    n1957,
    n1539
  );


  buf
  g2027
  (
    n1798,
    n1636
  );


  buf
  g2028
  (
    n1792,
    n1626
  );


  not
  g2029
  (
    n1699,
    n1598
  );


  not
  g2030
  (
    n1849,
    n1600
  );


  buf
  g2031
  (
    n1731,
    n1623
  );


  not
  g2032
  (
    n1805,
    n1644
  );


  buf
  g2033
  (
    n1964,
    n1583
  );


  not
  g2034
  (
    n1727,
    n1621
  );


  buf
  g2035
  (
    n1919,
    n1564
  );


  not
  g2036
  (
    n1748,
    n1620
  );


  not
  g2037
  (
    n2066,
    n1566
  );


  buf
  g2038
  (
    n1926,
    n1595
  );


  buf
  g2039
  (
    n2055,
    n1629
  );


  not
  g2040
  (
    n1660,
    n1620
  );


  not
  g2041
  (
    n1844,
    n1587
  );


  buf
  g2042
  (
    n1802,
    n1547
  );


  not
  g2043
  (
    n1681,
    n1623
  );


  not
  g2044
  (
    n1961,
    n1640
  );


  buf
  g2045
  (
    n1832,
    n1557
  );


  not
  g2046
  (
    n1772,
    n1630
  );


  buf
  g2047
  (
    n1775,
    n1571
  );


  buf
  g2048
  (
    n1751,
    n1608
  );


  not
  g2049
  (
    KeyWire_0_2,
    n1574
  );


  not
  g2050
  (
    n1960,
    n1619
  );


  buf
  g2051
  (
    n1740,
    n1543
  );


  not
  g2052
  (
    n2121,
    n1641
  );


  not
  g2053
  (
    n1711,
    n1563
  );


  not
  g2054
  (
    n2096,
    n1611
  );


  buf
  g2055
  (
    n1928,
    n1621
  );


  not
  g2056
  (
    n2059,
    n1648
  );


  not
  g2057
  (
    n2103,
    n1577
  );


  not
  g2058
  (
    n1846,
    n1588
  );


  not
  g2059
  (
    n1911,
    n1610
  );


  not
  g2060
  (
    n2110,
    n1601
  );


  buf
  g2061
  (
    n1827,
    n1544
  );


  buf
  g2062
  (
    n1689,
    n1632
  );


  not
  g2063
  (
    n1697,
    n1598
  );


  not
  g2064
  (
    n1682,
    n1648
  );


  not
  g2065
  (
    n1728,
    n1608
  );


  not
  g2066
  (
    n2021,
    n1634
  );


  not
  g2067
  (
    n1906,
    n1552
  );


  buf
  g2068
  (
    n1902,
    n1628
  );


  not
  g2069
  (
    n2074,
    n1613
  );


  buf
  g2070
  (
    n1729,
    n1585
  );


  not
  g2071
  (
    n1722,
    n1555
  );


  not
  g2072
  (
    n1789,
    n1569
  );


  buf
  g2073
  (
    n1878,
    n1579
  );


  not
  g2074
  (
    n2028,
    n1545
  );


  buf
  g2075
  (
    n1714,
    n1591
  );


  buf
  g2076
  (
    n1968,
    n1570
  );


  buf
  g2077
  (
    n1935,
    n1602
  );


  not
  g2078
  (
    n2004,
    n1562
  );


  not
  g2079
  (
    n2125,
    n1540
  );


  not
  g2080
  (
    n1854,
    n1626
  );


  not
  g2081
  (
    n1981,
    n1625
  );


  buf
  g2082
  (
    n2058,
    n1562
  );


  buf
  g2083
  (
    n1720,
    n1558
  );


  buf
  g2084
  (
    n2020,
    n1642
  );


  not
  g2085
  (
    n2064,
    n1607
  );


  not
  g2086
  (
    n1790,
    n1540
  );


  buf
  g2087
  (
    n1793,
    n1545
  );


  not
  g2088
  (
    n2115,
    n1549
  );


  not
  g2089
  (
    n1913,
    n1633
  );


  not
  g2090
  (
    n1940,
    n1579
  );


  buf
  g2091
  (
    n1882,
    n1644
  );


  not
  g2092
  (
    n1658,
    n1613
  );


  not
  g2093
  (
    n1966,
    n1631
  );


  not
  g2094
  (
    n1664,
    n1633
  );


  not
  g2095
  (
    n1661,
    n1541
  );


  not
  g2096
  (
    n1730,
    n1599
  );


  not
  g2097
  (
    n1903,
    n1630
  );


  buf
  g2098
  (
    n1797,
    n1559
  );


  buf
  g2099
  (
    n1750,
    n1634
  );


  not
  g2100
  (
    n1686,
    n1592
  );


  buf
  g2101
  (
    n2063,
    n1631
  );


  buf
  g2102
  (
    n1777,
    n1584
  );


  buf
  g2103
  (
    n1759,
    n1618
  );


  not
  g2104
  (
    n2100,
    n1592
  );


  not
  g2105
  (
    n1721,
    n1550
  );


  not
  g2106
  (
    n1925,
    n1612
  );


  not
  g2107
  (
    n1691,
    n1592
  );


  buf
  g2108
  (
    n1765,
    n1563
  );


  buf
  g2109
  (
    n1989,
    n1639
  );


  buf
  g2110
  (
    n2145,
    n1673
  );


  not
  g2111
  (
    n2188,
    n1705
  );


  not
  g2112
  (
    n2136,
    n1696
  );


  not
  g2113
  (
    n2182,
    n1693
  );


  not
  g2114
  (
    n2149,
    n1689
  );


  buf
  g2115
  (
    n2138,
    n1677
  );


  buf
  g2116
  (
    n2161,
    n1700
  );


  buf
  g2117
  (
    n2146,
    n1662
  );


  not
  g2118
  (
    n2190,
    n1667
  );


  buf
  g2119
  (
    n2152,
    n1685
  );


  buf
  g2120
  (
    n2189,
    n1710
  );


  buf
  g2121
  (
    n2155,
    n1656
  );


  not
  g2122
  (
    n2186,
    n1671
  );


  buf
  g2123
  (
    n2147,
    n1682
  );


  buf
  g2124
  (
    n2174,
    n1704
  );


  buf
  g2125
  (
    n2176,
    n1666
  );


  buf
  g2126
  (
    n2162,
    n1707
  );


  not
  g2127
  (
    n2151,
    n1698
  );


  buf
  g2128
  (
    n2185,
    n1690
  );


  not
  g2129
  (
    n2173,
    n1664
  );


  not
  g2130
  (
    n2148,
    n1706
  );


  not
  g2131
  (
    n2180,
    n1679
  );


  not
  g2132
  (
    n2165,
    n1683
  );


  buf
  g2133
  (
    n2153,
    n1669
  );


  buf
  g2134
  (
    n2170,
    n1709
  );


  not
  g2135
  (
    n2156,
    n1686
  );


  not
  g2136
  (
    n2177,
    n1660
  );


  not
  g2137
  (
    n2172,
    n1657
  );


  buf
  g2138
  (
    n2167,
    n1702
  );


  buf
  g2139
  (
    n2158,
    n1663
  );


  not
  g2140
  (
    n2140,
    n1674
  );


  not
  g2141
  (
    n2160,
    n1697
  );


  not
  g2142
  (
    n2144,
    n1678
  );


  not
  g2143
  (
    n2157,
    n1680
  );


  not
  g2144
  (
    n2164,
    n1688
  );


  not
  g2145
  (
    n2142,
    n1658
  );


  not
  g2146
  (
    n2178,
    n1675
  );


  buf
  g2147
  (
    n2169,
    n1681
  );


  buf
  g2148
  (
    n2187,
    n1655
  );


  buf
  g2149
  (
    KeyWire_0_30,
    n1670
  );


  buf
  g2150
  (
    n2159,
    n1691
  );


  not
  g2151
  (
    n2181,
    n1695
  );


  buf
  g2152
  (
    n2150,
    n1672
  );


  not
  g2153
  (
    n2171,
    n1668
  );


  not
  g2154
  (
    n2135,
    n1661
  );


  not
  g2155
  (
    n2179,
    n1703
  );


  not
  g2156
  (
    n2141,
    n1692
  );


  buf
  g2157
  (
    n2166,
    n1699
  );


  not
  g2158
  (
    n2143,
    n1687
  );


  not
  g2159
  (
    n2163,
    n1676
  );


  buf
  g2160
  (
    n2137,
    n1694
  );


  not
  g2161
  (
    n2168,
    n1665
  );


  not
  g2162
  (
    n2183,
    n1659
  );


  not
  g2163
  (
    n2184,
    n1684
  );


  not
  g2164
  (
    n2154,
    n1701
  );


  buf
  g2165
  (
    n2139,
    n1708
  );


  buf
  g2166
  (
    n2192,
    n2135
  );


  buf
  g2167
  (
    n2193,
    n2135
  );


  not
  g2168
  (
    n2191,
    n2135
  );


  buf
  g2169
  (
    n2194,
    n2135
  );


  or
  g2170
  (
    n2202,
    n2193,
    n2140,
    n2137,
    n2139
  );


  nand
  g2171
  (
    n2207,
    n2194,
    n2146,
    n2139,
    n2192
  );


  or
  g2172
  (
    n2209,
    n2192,
    n2192,
    n2144,
    n2147
  );


  or
  g2173
  (
    n2203,
    n2140,
    n2136,
    n2137,
    n2138
  );


  or
  g2174
  (
    n2204,
    n2141,
    n2146,
    n2136
  );


  and
  g2175
  (
    n2200,
    n2192,
    n2138,
    n2139
  );


  nor
  g2176
  (
    n2199,
    n2193,
    n2144,
    n2145,
    n2138
  );


  xnor
  g2177
  (
    n2198,
    n2146,
    n2136,
    n2137,
    n2141
  );


  xnor
  g2178
  (
    KeyWire_0_11,
    n2144,
    n2191,
    n2136,
    n2140
  );


  nor
  g2179
  (
    n2201,
    n2191,
    n2142,
    n2193,
    n2137
  );


  or
  g2180
  (
    n2195,
    n2139,
    n2142,
    n2144,
    n2141
  );


  nand
  g2181
  (
    n2206,
    n2191,
    n2142,
    n2141
  );


  nand
  g2182
  (
    n2197,
    n2191,
    n2194,
    n2140,
    n2143
  );


  nand
  g2183
  (
    n2196,
    n2193,
    n2143
  );


  xnor
  g2184
  (
    n2208,
    n2194,
    n2145
  );


  or
  g2185
  (
    n2211,
    n396,
    n399,
    n2199,
    n398
  );


  or
  g2186
  (
    n2214,
    n400,
    n2200,
    n390
  );


  xor
  g2187
  (
    n2219,
    n2201,
    n390,
    n2198
  );


  xnor
  g2188
  (
    n2221,
    n395,
    n395,
    n2202,
    n530
  );


  and
  g2189
  (
    n2210,
    n2200,
    n394,
    n391,
    n397
  );


  xor
  g2190
  (
    n2225,
    n399,
    n2196,
    n392
  );


  or
  g2191
  (
    n2224,
    n394,
    n399,
    n391,
    n2201
  );


  xor
  g2192
  (
    n2220,
    n389,
    n397,
    n391,
    n2197
  );


  nor
  g2193
  (
    n2213,
    n396,
    n392,
    n395,
    n394
  );


  xor
  g2194
  (
    n2216,
    n399,
    n2195,
    n396,
    n395
  );


  nand
  g2195
  (
    n2218,
    n2201,
    n2202,
    n396
  );


  xnor
  g2196
  (
    n2215,
    n531,
    n2201,
    n393
  );


  and
  g2197
  (
    n2217,
    n397,
    n392,
    n398,
    n400
  );


  and
  g2198
  (
    n2222,
    n390,
    n393,
    n389
  );


  nor
  g2199
  (
    n2212,
    n400,
    n394,
    n398
  );


  xnor
  g2200
  (
    n2223,
    n391,
    n397,
    n400,
    n2200
  );


  nor
  g2201
  (
    n2227,
    n2217,
    n553,
    n534,
    n548
  );


  nor
  g2202
  (
    n2230,
    n2212,
    n540,
    n539,
    n538
  );


  xnor
  g2203
  (
    n2226,
    n543,
    n542,
    n559,
    n558
  );


  xor
  g2204
  (
    n2235,
    n2215,
    n550,
    n536,
    n537
  );


  nor
  g2205
  (
    n2231,
    n557,
    n561,
    n533,
    n560
  );


  nand
  g2206
  (
    n2228,
    n552,
    n2211,
    n532,
    n2214
  );


  and
  g2207
  (
    n2232,
    n546,
    n544,
    n549,
    n2210
  );


  nor
  g2208
  (
    n2234,
    n545,
    n541,
    n2218,
    n2216
  );


  nor
  g2209
  (
    n2233,
    n2213,
    n554,
    n535,
    n547
  );


  and
  g2210
  (
    n2229,
    n2219,
    n551,
    n555,
    n556
  );


  buf
  g2211
  (
    n2236,
    n2235
  );


  not
  g2212
  (
    n2242,
    n2231
  );


  buf
  g2213
  (
    n2241,
    n2229
  );


  not
  g2214
  (
    n2238,
    n2232
  );


  buf
  g2215
  (
    n2237,
    n2234
  );


  buf
  g2216
  (
    n2240,
    n2233
  );


  not
  g2217
  (
    n2239,
    n2230
  );


  buf
  g2218
  (
    n2243,
    n2237
  );


  buf
  g2219
  (
    n2246,
    n2236
  );


  buf
  g2220
  (
    n2245,
    n2238
  );


  and
  g2221
  (
    n2244,
    n2237,
    n2236,
    n2239
  );


  and
  g2222
  (
    n2247,
    n2238,
    n2236,
    n2237
  );


  nand
  g2223
  (
    n2251,
    n1712,
    n401,
    n1716
  );


  xor
  g2224
  (
    n2250,
    n1713,
    n2245,
    n401,
    n402
  );


  xnor
  g2225
  (
    n2249,
    n2244,
    n1711,
    n401,
    n402
  );


  nand
  g2226
  (
    n2248,
    n1714,
    n1715,
    n2246,
    n2243
  );


  buf
  g2227
  (
    n2253,
    n1717
  );


  not
  g2228
  (
    n2252,
    n2251
  );


  or
  g2229
  (
    n2254,
    n1719,
    n2250,
    n1718,
    n2249
  );


  xor
  g2230
  (
    n2256,
    n2254,
    n566,
    n569,
    n562
  );


  or
  g2231
  (
    n2257,
    n571,
    n570,
    n565,
    n563
  );


  or
  g2232
  (
    n2255,
    n567,
    n572,
    n2252,
    n2254
  );


  or
  g2233
  (
    n2258,
    n568,
    n573,
    n2253,
    n564
  );


  not
  g2234
  (
    n2271,
    n2256
  );


  not
  g2235
  (
    n2264,
    n2258
  );


  buf
  g2236
  (
    n2267,
    n2257
  );


  not
  g2237
  (
    n2269,
    n2256
  );


  buf
  g2238
  (
    n2262,
    n120
  );


  buf
  g2239
  (
    n2270,
    n2255
  );


  not
  g2240
  (
    n2263,
    n2257
  );


  not
  g2241
  (
    n2268,
    n2256
  );


  not
  g2242
  (
    n2265,
    n2255
  );


  not
  g2243
  (
    n2259,
    n2255
  );


  not
  g2244
  (
    n2266,
    n2257
  );


  buf
  g2245
  (
    n2260,
    n120
  );


  nor
  g2246
  (
    n2261,
    n2256,
    n2257,
    n120,
    n2255
  );


  nand
  g2247
  (
    n2284,
    n402,
    n403,
    n411,
    n410
  );


  or
  g2248
  (
    n2274,
    n411,
    n410,
    n409
  );


  or
  g2249
  (
    n2283,
    n2268,
    n2259,
    n406,
    n403
  );


  xnor
  g2250
  (
    n2277,
    n404,
    n411,
    n405,
    n407
  );


  and
  g2251
  (
    n2272,
    n2270,
    n407,
    n404,
    n2265
  );


  nand
  g2252
  (
    n2276,
    n411,
    n405,
    n402
  );


  xor
  g2253
  (
    n2279,
    n408,
    n2271,
    n407,
    n403
  );


  or
  g2254
  (
    n2275,
    n410,
    n407,
    n408,
    n409
  );


  nand
  g2255
  (
    n2273,
    n2264,
    n406,
    n2262,
    n404
  );


  nand
  g2256
  (
    n2280,
    n406,
    n2260,
    n2267,
    n408
  );


  and
  g2257
  (
    n2282,
    n406,
    n405,
    n412,
    n404
  );


  nand
  g2258
  (
    n2281,
    n410,
    n2269,
    n408,
    n2261
  );


  nand
  g2259
  (
    n2278,
    n2263,
    n409,
    n403,
    n2266
  );


  or
  g2260
  (
    n2288,
    n576,
    n584
  );


  xor
  g2261
  (
    n2286,
    n574,
    n583
  );


  nand
  g2262
  (
    KeyWire_0_20,
    n2273,
    n577,
    n2274,
    n582
  );


  and
  g2263
  (
    n2287,
    n2274,
    n581,
    n575,
    n580
  );


  xnor
  g2264
  (
    n2289,
    n2275,
    n578,
    n579,
    n2272
  );


  xnor
  g2265
  (
    n2307,
    n2286,
    n2287,
    n613,
    n2288
  );


  nand
  g2266
  (
    n2300,
    n588,
    n600,
    n639,
    n585
  );


  and
  g2267
  (
    n2299,
    n590,
    n621,
    n591,
    n619
  );


  xor
  g2268
  (
    n2308,
    n2287,
    n629,
    n2285,
    n607
  );


  xor
  g2269
  (
    n2302,
    n641,
    n2285,
    n586,
    n597
  );


  or
  g2270
  (
    n2309,
    n632,
    n610,
    n592,
    n635
  );


  xnor
  g2271
  (
    n2291,
    n609,
    n2287,
    n2288,
    n623
  );


  xor
  g2272
  (
    n2301,
    n2285,
    n2288,
    n596
  );


  and
  g2273
  (
    n2306,
    n587,
    n599,
    n601,
    n620
  );


  nand
  g2274
  (
    n2292,
    n2285,
    n612,
    n626,
    n2289
  );


  nor
  g2275
  (
    n2294,
    n606,
    n595,
    n622,
    n608
  );


  and
  g2276
  (
    n2296,
    n2289,
    n605,
    n2286,
    n594
  );


  nor
  g2277
  (
    n2298,
    n627,
    n625,
    n638,
    n615
  );


  xor
  g2278
  (
    n2295,
    n589,
    n616,
    n644,
    n643
  );


  or
  g2279
  (
    n2293,
    n617,
    n593,
    n630,
    n634
  );


  xnor
  g2280
  (
    n2305,
    n633,
    n603,
    n2286,
    n614
  );


  or
  g2281
  (
    n2304,
    n598,
    n631,
    n2286,
    n2287
  );


  nor
  g2282
  (
    n2303,
    n636,
    n618,
    n628,
    n640
  );


  nand
  g2283
  (
    n2297,
    n637,
    n611,
    n642,
    n602
  );


  or
  g2284
  (
    n2290,
    n624,
    n604,
    n2289
  );


  nor
  g2285
  (
    n2310,
    n2305,
    n413,
    n2147,
    n2240
  );


  xnor
  g2286
  (
    n2314,
    n661,
    n647,
    n652,
    n412
  );


  nor
  g2287
  (
    n2319,
    n656,
    n654,
    n2309,
    n2302
  );


  and
  g2288
  (
    n2313,
    n413,
    n2301,
    n2298,
    n658
  );


  or
  g2289
  (
    n2312,
    n2240,
    n2239,
    n2299,
    n645
  );


  xnor
  g2290
  (
    n2321,
    n2147,
    n651,
    n646,
    n413
  );


  and
  g2291
  (
    n2311,
    n414,
    n660,
    n2239,
    n2307
  );


  and
  g2292
  (
    n2315,
    n2240,
    n649,
    n653,
    n2300
  );


  xnor
  g2293
  (
    n2317,
    n2241,
    n412,
    n657,
    n2303
  );


  nor
  g2294
  (
    n2316,
    n2304,
    n648,
    n2240,
    n655
  );


  or
  g2295
  (
    n2320,
    n2241,
    n659,
    n412,
    n2308
  );


  xnor
  g2296
  (
    n2318,
    n413,
    n650,
    n2239,
    n2306
  );


  buf
  g2297
  (
    n2322,
    n2310
  );


  buf
  g2298
  (
    n2323,
    n2311
  );


  nor
  g2299
  (
    n2324,
    n1720,
    n2322
  );


  or
  g2300
  (
    n2328,
    n2149,
    n2149,
    n2148,
    n2324
  );


  xor
  g2301
  (
    n2327,
    n2148,
    n2147,
    n2150,
    n2324
  );


  xor
  g2302
  (
    n2326,
    n2324,
    n2324,
    n662,
    n2149
  );


  and
  g2303
  (
    n2325,
    n2149,
    n2148,
    n2150
  );


  and
  g2304
  (
    n2337,
    n2327,
    n669,
    n692,
    n681
  );


  xor
  g2305
  (
    KeyWire_0_19,
    n667,
    n2327,
    n664,
    n684
  );


  or
  g2306
  (
    n2333,
    n679,
    n2325,
    n2327,
    n680
  );


  nand
  g2307
  (
    n2331,
    n668,
    n2328,
    n674,
    n686
  );


  and
  g2308
  (
    n2329,
    n2327,
    n678,
    n2328,
    n691
  );


  xnor
  g2309
  (
    n2338,
    n665,
    n672,
    n685,
    n687
  );


  or
  g2310
  (
    n2330,
    n666,
    n673,
    n663,
    n675
  );


  xor
  g2311
  (
    n2332,
    n671,
    n688,
    n690,
    n670
  );


  and
  g2312
  (
    n2334,
    n2326,
    n677,
    n2328,
    n676
  );


  nor
  g2313
  (
    n2336,
    n682,
    n2328,
    n683,
    n689
  );


  buf
  g2314
  (
    n2339,
    n2330
  );


  buf
  g2315
  (
    n2340,
    n2329
  );


  and
  g2316
  (
    n2346,
    n2332,
    n2331,
    n2340
  );


  and
  g2317
  (
    n2341,
    n2334,
    n2333
  );


  nor
  g2318
  (
    n2345,
    n2331,
    n2340,
    n2330
  );


  or
  g2319
  (
    n2343,
    n2330,
    n2332,
    n2334
  );


  nor
  g2320
  (
    n2342,
    n2331,
    n2330,
    n2332
  );


  nor
  g2321
  (
    n2344,
    n2333,
    n2339,
    n2331
  );


  nor
  g2322
  (
    n2347,
    n712,
    n2343,
    n696,
    n2346
  );


  nor
  g2323
  (
    KeyWire_0_1,
    n699,
    n2341,
    n714,
    n705
  );


  nor
  g2324
  (
    n2353,
    n713,
    n706,
    n709,
    n710
  );


  nor
  g2325
  (
    n2352,
    n698,
    n711,
    n701,
    n708
  );


  nor
  g2326
  (
    n2354,
    n707,
    n2346,
    n704,
    n702
  );


  or
  g2327
  (
    n2348,
    n2342,
    n716,
    n718,
    n2345
  );


  xor
  g2328
  (
    n2355,
    n715,
    n697,
    n2346,
    n694
  );


  xnor
  g2329
  (
    n2349,
    n700,
    n717,
    n2346,
    n693
  );


  or
  g2330
  (
    n2351,
    n719,
    n703,
    n695,
    n2344
  );


  or
  g2331
  (
    n2376,
    n1741,
    n1729,
    n720,
    n2353
  );


  or
  g2332
  (
    n2359,
    n2353,
    n724,
    n738,
    n1780
  );


  nor
  g2333
  (
    n2388,
    n2348,
    n1789,
    n1772,
    n729
  );


  nor
  g2334
  (
    n2370,
    n1781,
    n1787,
    n736,
    n1759
  );


  nand
  g2335
  (
    n2356,
    n1766,
    n1757,
    n1769,
    n1779
  );


  xor
  g2336
  (
    n2377,
    n2350,
    n728,
    n2242,
    n2347
  );


  and
  g2337
  (
    n2383,
    n1753,
    n2355,
    n733,
    n1751
  );


  xnor
  g2338
  (
    n2357,
    n1754,
    n2354,
    n1723,
    n1740
  );


  xnor
  g2339
  (
    n2362,
    n1762,
    n1786,
    n2352,
    n734
  );


  and
  g2340
  (
    n2389,
    n1790,
    n2352,
    n2354,
    n1767
  );


  nand
  g2341
  (
    n2364,
    n725,
    n2351,
    n1737,
    n2352
  );


  nand
  g2342
  (
    n2367,
    n1770,
    n1777,
    n1746,
    n2350
  );


  or
  g2343
  (
    n2382,
    n737,
    n2241,
    n748,
    n732
  );


  and
  g2344
  (
    n2360,
    n730,
    n1727,
    n2354,
    n2347
  );


  nor
  g2345
  (
    n2379,
    n1756,
    n1776,
    n2349,
    n1725
  );


  nor
  g2346
  (
    n2369,
    n1749,
    n2350,
    n1761,
    n743
  );


  or
  g2347
  (
    n2373,
    n2351,
    n2355,
    n1733,
    n1739
  );


  xnor
  g2348
  (
    n2390,
    n2348,
    n2241,
    n1726,
    n1747
  );


  xnor
  g2349
  (
    n2361,
    n746,
    n2353,
    n1722,
    n1721
  );


  xor
  g2350
  (
    n2371,
    n2354,
    n1764,
    n723,
    n1765
  );


  or
  g2351
  (
    n2385,
    n2355,
    n1744,
    n1750,
    n1791
  );


  and
  g2352
  (
    n2386,
    n2242,
    n1742,
    n739,
    n2348
  );


  xnor
  g2353
  (
    n2365,
    n1774,
    n2349,
    n1785,
    n1743
  );


  and
  g2354
  (
    n2391,
    n1732,
    n1736,
    n1730,
    n1734
  );


  and
  g2355
  (
    n2358,
    n1731,
    n1775,
    n2349,
    n1768
  );


  xor
  g2356
  (
    n2384,
    n1782,
    n1735,
    n1778,
    n2351
  );


  xor
  g2357
  (
    n2366,
    n1760,
    n2351,
    n1748,
    n2242
  );


  nor
  g2358
  (
    n2363,
    n2355,
    n1771,
    n727,
    n2350
  );


  or
  g2359
  (
    n2378,
    n741,
    n2348,
    n2353,
    n747
  );


  and
  g2360
  (
    n2381,
    n2347,
    n735,
    n1788,
    n2349
  );


  xnor
  g2361
  (
    n2372,
    n1724,
    n1758,
    n1745,
    n2242
  );


  xnor
  g2362
  (
    n2374,
    n1773,
    n1738,
    n726,
    n2352
  );


  nor
  g2363
  (
    n2380,
    n745,
    n1793,
    n1755,
    n1763
  );


  nor
  g2364
  (
    n2375,
    n1783,
    n744,
    n740,
    n721
  );


  xor
  g2365
  (
    n2387,
    n1792,
    n1752,
    n722,
    n2347
  );


  nor
  g2366
  (
    n2368,
    n1728,
    n1784,
    n731,
    n742
  );


  nand
  g2367
  (
    n2444,
    n2387,
    n1052,
    n1137,
    n937
  );


  or
  g2368
  (
    n2522,
    n876,
    n990,
    n2372,
    n2379
  );


  nor
  g2369
  (
    n2394,
    n885,
    n981,
    n947,
    n2359
  );


  xor
  g2370
  (
    n2462,
    n2386,
    n2376,
    n2389,
    n1124
  );


  nand
  g2371
  (
    n2427,
    n763,
    n843,
    n2383,
    n925
  );


  or
  g2372
  (
    n2524,
    n934,
    n2319,
    n2391,
    n1161
  );


  xnor
  g2373
  (
    n2528,
    n2367,
    n2365,
    n1144,
    n906
  );


  and
  g2374
  (
    n2441,
    n770,
    n2383,
    n2385,
    n1105
  );


  xnor
  g2375
  (
    n2509,
    n2379,
    n886,
    n2377
  );


  and
  g2376
  (
    n2454,
    n815,
    n2375,
    n1093,
    n2383
  );


  and
  g2377
  (
    n2472,
    n984,
    n973,
    n846,
    n2363
  );


  xnor
  g2378
  (
    n2520,
    n1113,
    n1067,
    n2379,
    n1162
  );


  or
  g2379
  (
    n2464,
    n1062,
    n1123,
    n2375,
    n2357
  );


  xor
  g2380
  (
    n2434,
    n980,
    n936,
    n1007,
    n1058
  );


  and
  g2381
  (
    n2455,
    n793,
    n870,
    n804,
    n1077
  );


  nand
  g2382
  (
    n2478,
    n789,
    n1023,
    n884,
    n1072
  );


  nand
  g2383
  (
    n2413,
    n2363,
    n1033,
    n1156,
    n942
  );


  and
  g2384
  (
    n2430,
    n1010,
    n780,
    n2382,
    n941
  );


  nor
  g2385
  (
    n2503,
    n1014,
    n2314,
    n919,
    n2372
  );


  nor
  g2386
  (
    n2480,
    n2356,
    n2359,
    n898,
    n760
  );


  nor
  g2387
  (
    n2510,
    n2370,
    n841,
    n1063,
    n828
  );


  and
  g2388
  (
    n2450,
    n950,
    n2379,
    n2320,
    n1003
  );


  nor
  g2389
  (
    n2496,
    n894,
    n2389,
    n813,
    n773
  );


  xor
  g2390
  (
    n2461,
    n878,
    n2360,
    n764,
    n2361
  );


  xor
  g2391
  (
    n2517,
    n949,
    n851,
    n749,
    n2360
  );


  xnor
  g2392
  (
    n2392,
    n871,
    n970,
    n899,
    n2382
  );


  nand
  g2393
  (
    n2443,
    n924,
    n2319,
    n1017,
    n1026
  );


  nor
  g2394
  (
    n2471,
    n1122,
    n869,
    n963,
    n818
  );


  xor
  g2395
  (
    n2421,
    n756,
    n1142,
    n1108,
    n1114
  );


  xnor
  g2396
  (
    n2438,
    n2371,
    n2371,
    n801,
    n1005
  );


  nor
  g2397
  (
    n2417,
    n777,
    n986,
    n959,
    n1000
  );


  and
  g2398
  (
    n2446,
    n1061,
    n938,
    n1024,
    n1021
  );


  nor
  g2399
  (
    n2416,
    n850,
    n2387,
    n2372,
    n914
  );


  xor
  g2400
  (
    n2516,
    n859,
    n953,
    n1112,
    n1069
  );


  nor
  g2401
  (
    n2426,
    n944,
    n993,
    n2391,
    n1111
  );


  or
  g2402
  (
    n2400,
    n882,
    n765,
    n893,
    n1106
  );


  xor
  g2403
  (
    n2484,
    n857,
    n930,
    n922,
    n1071
  );


  or
  g2404
  (
    n2457,
    n852,
    n1102,
    n2384,
    n1053
  );


  or
  g2405
  (
    n2415,
    n1046,
    n2361,
    n909,
    n1147
  );


  xor
  g2406
  (
    n2435,
    n781,
    n978,
    n1029,
    n2368
  );


  and
  g2407
  (
    n2475,
    n844,
    n2381,
    n1031,
    n915
  );


  xor
  g2408
  (
    n2399,
    n921,
    n800,
    n1015,
    n809
  );


  xor
  g2409
  (
    n2420,
    n2390,
    n796,
    n957,
    n982
  );


  xnor
  g2410
  (
    n2397,
    n794,
    n790,
    n1059,
    n2390
  );


  and
  g2411
  (
    n2476,
    n912,
    n2313,
    n964,
    n933
  );


  and
  g2412
  (
    n2532,
    n1076,
    n1022,
    n814,
    n824
  );


  nand
  g2413
  (
    n2519,
    n798,
    n2391,
    n926,
    n868
  );


  xor
  g2414
  (
    n2429,
    n863,
    n1151,
    n1060,
    n1100
  );


  or
  g2415
  (
    n2447,
    n2312,
    n792,
    n2358
  );


  and
  g2416
  (
    n2470,
    n2381,
    n1070,
    n811,
    n1089
  );


  nand
  g2417
  (
    n2490,
    n839,
    n1164,
    n2374,
    n994
  );


  and
  g2418
  (
    n2456,
    n2386,
    n2387,
    n889,
    n860
  );


  xnor
  g2419
  (
    n2493,
    n943,
    n2359,
    n920,
    n2373
  );


  nand
  g2420
  (
    n2498,
    n1157,
    n833,
    n1098,
    n1118
  );


  xor
  g2421
  (
    n2501,
    n1032,
    n791,
    n1136,
    n782
  );


  and
  g2422
  (
    n2526,
    n2381,
    n2320,
    n864,
    n1073
  );


  and
  g2423
  (
    n2500,
    n837,
    n2363,
    n865,
    n1129
  );


  and
  g2424
  (
    n2491,
    n2367,
    n879,
    n2369,
    n2366
  );


  nand
  g2425
  (
    n2393,
    n965,
    n2376,
    n1115,
    n975
  );


  nor
  g2426
  (
    n2433,
    n795,
    n891,
    n951,
    n1131
  );


  nor
  g2427
  (
    n2432,
    n2378,
    n783,
    n913,
    n1041
  );


  nand
  g2428
  (
    n2486,
    n887,
    n989,
    n2364,
    n1016
  );


  and
  g2429
  (
    n2409,
    n2358,
    n969,
    n2388,
    n872
  );


  nand
  g2430
  (
    n2489,
    n1056,
    n1078,
    n935,
    n916
  );


  xnor
  g2431
  (
    n2405,
    n1009,
    n988,
    n1152,
    n955
  );


  and
  g2432
  (
    n2398,
    n1038,
    n888,
    n1092,
    n1163
  );


  or
  g2433
  (
    n2530,
    n1080,
    n2389,
    n1008,
    n976
  );


  nand
  g2434
  (
    n2408,
    n2390,
    n2364,
    n2385
  );


  xnor
  g2435
  (
    n2418,
    n1050,
    n769,
    n1154,
    n855
  );


  xor
  g2436
  (
    n2507,
    n758,
    n753,
    n2362,
    n803
  );


  or
  g2437
  (
    n2497,
    n2382,
    n840,
    n849,
    n1121
  );


  nand
  g2438
  (
    n2459,
    n2319,
    n967,
    n1051,
    n1018
  );


  or
  g2439
  (
    n2411,
    n752,
    n1039,
    n1040,
    n767
  );


  and
  g2440
  (
    n2463,
    n2357,
    n1047,
    n2370,
    n2317
  );


  xor
  g2441
  (
    n2495,
    n805,
    n873,
    n827,
    n2362
  );


  nor
  g2442
  (
    n2439,
    n2359,
    n1084,
    n1045,
    n917
  );


  xnor
  g2443
  (
    n2404,
    n2369,
    n1107,
    n821,
    n806
  );


  xnor
  g2444
  (
    n2488,
    n779,
    n858,
    n1138,
    n838
  );


  xor
  g2445
  (
    n2402,
    n940,
    n2378,
    n778,
    n2380
  );


  xor
  g2446
  (
    n2440,
    n991,
    n2367,
    n883,
    n761
  );


  and
  g2447
  (
    n2479,
    n1074,
    n1117,
    n2384,
    n2377
  );


  nand
  g2448
  (
    n2487,
    n2361,
    n787,
    n856,
    n2362
  );


  xor
  g2449
  (
    n2437,
    n786,
    n1160,
    n822,
    n825
  );


  xnor
  g2450
  (
    n2502,
    n983,
    n996,
    n1150,
    n896
  );


  xnor
  g2451
  (
    n2512,
    n2380,
    n2376,
    n2362,
    n1068
  );


  nand
  g2452
  (
    n2465,
    n892,
    n995,
    n1110,
    n2386
  );


  xor
  g2453
  (
    n2453,
    n768,
    n961,
    n866,
    n2388
  );


  xor
  g2454
  (
    n2410,
    n771,
    n2387,
    n759,
    n830
  );


  nor
  g2455
  (
    n2451,
    n831,
    n890,
    n1109,
    n992
  );


  or
  g2456
  (
    n2445,
    n877,
    n2384,
    n946,
    n819
  );


  or
  g2457
  (
    n2514,
    n907,
    n1116,
    n1049,
    n807
  );


  nor
  g2458
  (
    n2436,
    n1153,
    n2386,
    n1139,
    n956
  );


  and
  g2459
  (
    n2492,
    n931,
    n2385,
    n842,
    n968
  );


  xor
  g2460
  (
    n2428,
    n784,
    n1091,
    n2368,
    n1042
  );


  nor
  g2461
  (
    n2499,
    n901,
    n848,
    n832,
    n2382
  );


  xor
  g2462
  (
    n2460,
    n1011,
    n1133,
    n802,
    n757
  );


  xor
  g2463
  (
    n2424,
    n750,
    n1006,
    n2375,
    n1035
  );


  nor
  g2464
  (
    n2452,
    n826,
    n1159,
    n1034,
    n1141
  );


  nor
  g2465
  (
    n2431,
    n1012,
    n2371,
    n903,
    n910
  );


  xnor
  g2466
  (
    n2423,
    n2374,
    n2388,
    n2383,
    n2371
  );


  or
  g2467
  (
    n2531,
    n862,
    n875,
    n2381,
    n2372
  );


  xnor
  g2468
  (
    n2403,
    n1043,
    n2364,
    n2374,
    n897
  );


  or
  g2469
  (
    n2506,
    n1130,
    n1004,
    n772,
    n911
  );


  nand
  g2470
  (
    n2458,
    n881,
    n2363,
    n2366,
    n1037
  );


  xor
  g2471
  (
    n2466,
    n788,
    n2365,
    n835,
    n1082
  );


  nor
  g2472
  (
    n2469,
    n2356,
    n979,
    n918,
    n766
  );


  nand
  g2473
  (
    n2468,
    n755,
    n1065,
    n960,
    n776
  );


  xnor
  g2474
  (
    n2534,
    n1132,
    n1088,
    n1025,
    n785
  );


  xnor
  g2475
  (
    n2448,
    n2368,
    n2315,
    n1145,
    n2367
  );


  xor
  g2476
  (
    n2419,
    n2380,
    n1085,
    n2378,
    n1094
  );


  xnor
  g2477
  (
    n2396,
    n1001,
    n1165,
    n880,
    n2375
  );


  and
  g2478
  (
    n2529,
    n923,
    n927,
    n1054,
    n999
  );


  nor
  g2479
  (
    n2515,
    n2378,
    n2356,
    n939
  );


  nor
  g2480
  (
    n2485,
    n2318,
    n817,
    n2373,
    n2366
  );


  xnor
  g2481
  (
    n2406,
    n2365,
    n812,
    n2360,
    n823
  );


  nor
  g2482
  (
    n2483,
    n1075,
    n900,
    n1125,
    n2357
  );


  xnor
  g2483
  (
    n2505,
    n1158,
    n1019,
    n2373,
    n1048
  );


  xor
  g2484
  (
    n2533,
    n954,
    n1020,
    n2391,
    n1083
  );


  or
  g2485
  (
    n2467,
    n1120,
    n1002,
    n1134,
    n2384
  );


  and
  g2486
  (
    n2518,
    n1119,
    n2380,
    n1057,
    n1149
  );


  and
  g2487
  (
    n2508,
    n2360,
    n1027,
    n2366,
    n847
  );


  xnor
  g2488
  (
    n2504,
    n1099,
    n2389,
    n854,
    n977
  );


  or
  g2489
  (
    n2481,
    n2357,
    n799,
    n962,
    n1096
  );


  xnor
  g2490
  (
    n2412,
    n867,
    n1148,
    n861,
    n797
  );


  nor
  g2491
  (
    n2474,
    n820,
    n1155,
    n974,
    n2376
  );


  and
  g2492
  (
    n2523,
    n1090,
    n958,
    n1103,
    n908
  );


  nand
  g2493
  (
    n2511,
    n1036,
    n774,
    n905,
    n762
  );


  nand
  g2494
  (
    n2407,
    n2365,
    n972,
    n1064,
    n1128
  );


  xnor
  g2495
  (
    n2513,
    n2368,
    n952,
    n1079,
    n751
  );


  xor
  g2496
  (
    n2449,
    n928,
    n1044,
    n874,
    n1101
  );


  or
  g2497
  (
    n2535,
    n1028,
    n836,
    n1104,
    n1013
  );


  nand
  g2498
  (
    n2527,
    n754,
    n929,
    n987,
    n816
  );


  nor
  g2499
  (
    n2401,
    n932,
    n902,
    n948,
    n845
  );


  nand
  g2500
  (
    n2414,
    n2320,
    n1087,
    n2361,
    n2390
  );


  xnor
  g2501
  (
    n2442,
    n2370,
    n1066,
    n2247,
    n2316
  );


  xor
  g2502
  (
    n2477,
    n829,
    n810,
    n1146,
    n2385
  );


  nand
  g2503
  (
    n2494,
    n1055,
    n2358,
    n1081,
    n985
  );


  nor
  g2504
  (
    n2395,
    n1127,
    n1086,
    n1140,
    n2369
  );


  or
  g2505
  (
    n2521,
    n1143,
    n971,
    n2370,
    n2377
  );


  or
  g2506
  (
    n2482,
    n998,
    n834,
    n1135,
    n1095
  );


  nor
  g2507
  (
    n2422,
    n808,
    n1126,
    n2369,
    n853
  );


  xor
  g2508
  (
    n2425,
    n2388,
    n1097,
    n945,
    n1030
  );


  and
  g2509
  (
    n2473,
    n966,
    n775,
    n2373,
    n2319
  );


  and
  g2510
  (
    n2525,
    n997,
    n2374,
    n895,
    n904
  );


  xnor
  g2511
  (
    n2708,
    n2124,
    n471,
    n474,
    n464
  );


  xor
  g2512
  (
    n2593,
    n416,
    n2023,
    n2446,
    n425
  );


  or
  g2513
  (
    n2758,
    n1936,
    n2126,
    n2194,
    n2507
  );


  xor
  g2514
  (
    n2667,
    n2115,
    n1969,
    n1986,
    n1839
  );


  xor
  g2515
  (
    n2662,
    n429,
    n2125,
    n483,
    n2510
  );


  xor
  g2516
  (
    n2701,
    n2402,
    n2153,
    n481,
    n2075
  );


  xnor
  g2517
  (
    n2730,
    n1884,
    n1965,
    n2110,
    n1909
  );


  nand
  g2518
  (
    n2562,
    n2442,
    n469,
    n468,
    n2066
  );


  xor
  g2519
  (
    n2588,
    n1836,
    n2500,
    n467,
    n2395
  );


  nand
  g2520
  (
    n2555,
    n460,
    n2517,
    n418,
    n2054
  );


  or
  g2521
  (
    n2601,
    n1819,
    n420,
    n1912,
    n2534
  );


  and
  g2522
  (
    n2564,
    n416,
    n430,
    n1947,
    n488
  );


  or
  g2523
  (
    n2729,
    n2514,
    n499,
    n1924,
    n2464
  );


  nor
  g2524
  (
    n2631,
    n2203,
    n1985,
    n2151,
    n1923
  );


  xor
  g2525
  (
    n2704,
    n446,
    n455,
    n480,
    n2503
  );


  or
  g2526
  (
    n2561,
    n2503,
    n2486,
    n463,
    n2031
  );


  xor
  g2527
  (
    n2579,
    n1821,
    n1966,
    n445,
    n1892
  );


  nor
  g2528
  (
    n2795,
    n2120,
    n1859,
    n1991,
    n2117
  );


  nand
  g2529
  (
    n2589,
    n2419,
    n495,
    n2117,
    n2505
  );


  xor
  g2530
  (
    n2682,
    n473,
    n2497,
    n2403,
    n1857
  );


  or
  g2531
  (
    n2717,
    n429,
    n488,
    n2516,
    n1917
  );


  xnor
  g2532
  (
    n2609,
    n2520,
    n2494,
    n424,
    n2065
  );


  xnor
  g2533
  (
    n2663,
    n2466,
    n444,
    n2512,
    n2012
  );


  and
  g2534
  (
    n2539,
    n1855,
    n1838,
    n428,
    n1914
  );


  and
  g2535
  (
    n2775,
    n499,
    n2127,
    n2492,
    n2133
  );


  nand
  g2536
  (
    n2627,
    n2535,
    n2408,
    n1860,
    n480
  );


  xnor
  g2537
  (
    n2574,
    n1990,
    n2028,
    n475,
    n2469
  );


  and
  g2538
  (
    n2632,
    n474,
    n2111,
    n2513,
    n2027
  );


  and
  g2539
  (
    n2797,
    n419,
    n1815,
    n1953,
    n495
  );


  xor
  g2540
  (
    n2678,
    n2526,
    n450,
    n1825,
    n1968
  );


  nor
  g2541
  (
    n2731,
    n2500,
    n2524,
    n437,
    n2501
  );


  xor
  g2542
  (
    n2573,
    n438,
    n2050,
    n422,
    n2443
  );


  nand
  g2543
  (
    n2711,
    n1946,
    n2089,
    n2493,
    n1899
  );


  nand
  g2544
  (
    n2592,
    n2528,
    n1898,
    n1960,
    n493
  );


  nand
  g2545
  (
    n2571,
    n2504,
    n487,
    n2040,
    n2117
  );


  and
  g2546
  (
    n2638,
    n451,
    n2428,
    n2532,
    n2115
  );


  nand
  g2547
  (
    n2789,
    n452,
    n2113,
    n421,
    n2516
  );


  xor
  g2548
  (
    n2728,
    n481,
    n1944,
    n2527,
    n2522
  );


  nand
  g2549
  (
    n2559,
    n466,
    n2515,
    n471,
    n1867
  );


  xnor
  g2550
  (
    n2751,
    n452,
    n2467,
    n2113,
    n437
  );


  nand
  g2551
  (
    n2560,
    n1951,
    n478,
    n418,
    n2496
  );


  xor
  g2552
  (
    n2706,
    n2523,
    n2451,
    n463,
    n2131
  );


  or
  g2553
  (
    n2748,
    n472,
    n432,
    n2430,
    n1988
  );


  xor
  g2554
  (
    n2674,
    n449,
    n2501,
    n1844,
    n2002
  );


  xnor
  g2555
  (
    n2725,
    n1942,
    n2534,
    n2530,
    n2059
  );


  xor
  g2556
  (
    n2642,
    n1943,
    n432,
    n2132,
    n1875
  );


  and
  g2557
  (
    n2726,
    n2515,
    n2501,
    n1170,
    n2527
  );


  xnor
  g2558
  (
    n2607,
    n2529,
    n2055,
    n414,
    n2102
  );


  xnor
  g2559
  (
    n2693,
    n2447,
    n2478,
    n2049,
    n2481
  );


  or
  g2560
  (
    n2787,
    n2035,
    n2150,
    n1903,
    n2007
  );


  xor
  g2561
  (
    n2733,
    n2514,
    n493,
    n471,
    n2154
  );


  nor
  g2562
  (
    n2695,
    n2152,
    n2513,
    n465,
    n2520
  );


  xnor
  g2563
  (
    n2750,
    n1906,
    n1981,
    n1846,
    n2151
  );


  xnor
  g2564
  (
    n2702,
    n1896,
    n2399,
    n476,
    n2522
  );


  xnor
  g2565
  (
    n2616,
    n2506,
    n2115,
    n1907,
    n478
  );


  nand
  g2566
  (
    n2645,
    n2525,
    n463,
    n1935,
    n492
  );


  nand
  g2567
  (
    n2790,
    n460,
    n2498,
    n1804,
    n494
  );


  nor
  g2568
  (
    n2699,
    n459,
    n461,
    n2392,
    n2415
  );


  and
  g2569
  (
    n2603,
    n415,
    n2452,
    n1938,
    n2426
  );


  or
  g2570
  (
    n2595,
    n484,
    n2004,
    n2459,
    n2449
  );


  or
  g2571
  (
    n2630,
    n2525,
    n1806,
    n2116,
    n2123
  );


  nand
  g2572
  (
    n2615,
    n1169,
    n2510,
    n1956,
    n1994
  );


  nor
  g2573
  (
    n2581,
    n1890,
    n421,
    n2397,
    n462
  );


  or
  g2574
  (
    n2781,
    n500,
    n489,
    n451,
    n2503
  );


  xor
  g2575
  (
    n2689,
    n2506,
    n479,
    n1957,
    n451
  );


  and
  g2576
  (
    n2732,
    n1893,
    n1967,
    n1824,
    n2122
  );


  nor
  g2577
  (
    n2779,
    n2129,
    n443,
    n492,
    n479
  );


  nor
  g2578
  (
    n2685,
    n2523,
    n2154,
    n474,
    n453
  );


  xnor
  g2579
  (
    n2657,
    n2508,
    n2116,
    n2071,
    n485
  );


  nand
  g2580
  (
    n2544,
    n1879,
    n2131,
    n1989,
    n2530
  );


  or
  g2581
  (
    n2620,
    n2108,
    n2106,
    n2116,
    n2512
  );


  nor
  g2582
  (
    n2577,
    n2037,
    n493,
    n486,
    n2522
  );


  xor
  g2583
  (
    KeyWire_0_28,
    n1814,
    n457,
    n451,
    n483
  );


  and
  g2584
  (
    n2742,
    n424,
    n2505,
    n1877,
    n2123
  );


  or
  g2585
  (
    n2796,
    n2203,
    n2134,
    n456,
    n496
  );


  xnor
  g2586
  (
    n2600,
    n491,
    n2116,
    n2150,
    n2500
  );


  nor
  g2587
  (
    n2683,
    n492,
    n481,
    n483,
    n2413
  );


  xnor
  g2588
  (
    n2692,
    n1984,
    n2057,
    n2103,
    n448
  );


  nand
  g2589
  (
    n2672,
    n1818,
    n1928,
    n2153,
    n425
  );


  nor
  g2590
  (
    n2697,
    n2514,
    n2036,
    n458,
    n2041
  );


  nand
  g2591
  (
    n2703,
    n1843,
    n2501,
    n1992,
    n2082
  );


  xor
  g2592
  (
    n2651,
    n2323,
    n1871,
    n1897,
    n1832
  );


  nor
  g2593
  (
    n2715,
    n1811,
    n439,
    n460,
    n2056
  );


  or
  g2594
  (
    n2550,
    n1929,
    n2508,
    n2130,
    n1886
  );


  xor
  g2595
  (
    n2759,
    n445,
    n2533,
    n2506,
    n2484
  );


  nand
  g2596
  (
    n2794,
    n2414,
    n2072,
    n455,
    n2468
  );


  nand
  g2597
  (
    n2635,
    n2152,
    n2530,
    n465,
    n2091
  );


  xnor
  g2598
  (
    n2700,
    n2437,
    n2502,
    n1998,
    n2491
  );


  xnor
  g2599
  (
    n2656,
    n2471,
    n2118,
    n2453,
    n1872
  );


  xor
  g2600
  (
    KeyWire_0_6,
    n2323,
    n2128,
    n476,
    n1885
  );


  xnor
  g2601
  (
    n2576,
    n1168,
    n425,
    n1987,
    n2519
  );


  nor
  g2602
  (
    n2598,
    n434,
    n2112,
    n2422,
    n2456
  );


  xor
  g2603
  (
    n2636,
    n2033,
    n1904,
    n429,
    n422
  );


  and
  g2604
  (
    n2778,
    n475,
    n426,
    n1167,
    n2462
  );


  xnor
  g2605
  (
    n2621,
    n470,
    n2047,
    n419,
    n1808
  );


  nor
  g2606
  (
    n2643,
    n462,
    n1807,
    n1841,
    n1940
  );


  or
  g2607
  (
    n2769,
    n2017,
    n457,
    n430,
    n1889
  );


  xnor
  g2608
  (
    n2661,
    n2432,
    n2123,
    n2130,
    n2431
  );


  xnor
  g2609
  (
    n2719,
    n1830,
    n2533,
    n1800,
    n2516
  );


  xnor
  g2610
  (
    n2666,
    n2460,
    n2511,
    n2405,
    n2498
  );


  and
  g2611
  (
    n2671,
    n496,
    n2125,
    n2113,
    n488
  );


  nor
  g2612
  (
    n2712,
    n2506,
    n459,
    n2436,
    n2134
  );


  nand
  g2613
  (
    n2557,
    n2495,
    n2153,
    n416,
    n2128
  );


  nand
  g2614
  (
    n2792,
    n1854,
    n439,
    n2043,
    n1961
  );


  nor
  g2615
  (
    n2694,
    n1995,
    n2532,
    n1919,
    n2404
  );


  xor
  g2616
  (
    n2659,
    n2505,
    n439,
    n423,
    n497
  );


  xor
  g2617
  (
    n2743,
    n2433,
    n1977,
    n448,
    n2507
  );


  and
  g2618
  (
    n2768,
    n1801,
    n1997,
    n2435,
    n2058
  );


  nor
  g2619
  (
    n2780,
    n1973,
    n2122,
    n1932,
    n484
  );


  xor
  g2620
  (
    n2640,
    n2097,
    n415,
    n495,
    n2153
  );


  xor
  g2621
  (
    n2707,
    n2128,
    n433,
    n1902,
    n1794
  );


  nand
  g2622
  (
    n2687,
    n2396,
    n475,
    n435,
    n454
  );


  nor
  g2623
  (
    n2543,
    n468,
    n2513,
    n1795,
    n2016
  );


  nand
  g2624
  (
    n2629,
    n482,
    n455,
    n436,
    n1816
  );


  nor
  g2625
  (
    n2676,
    n1948,
    n2202,
    n2104,
    n1980
  );


  or
  g2626
  (
    n2583,
    n423,
    n1970,
    n1862,
    n2019
  );


  and
  g2627
  (
    n2658,
    n2120,
    n467,
    n1933,
    n1894
  );


  xor
  g2628
  (
    n2605,
    n2476,
    n2044,
    n1972,
    n453
  );


  xor
  g2629
  (
    n2757,
    n2034,
    n2440,
    n1858,
    n501
  );


  xor
  g2630
  (
    n2580,
    n465,
    n1950,
    n2450,
    n2132
  );


  nand
  g2631
  (
    n2542,
    n2401,
    n2502,
    n435,
    n2127
  );


  nor
  g2632
  (
    n2772,
    n2081,
    n501,
    n1869,
    n2006
  );


  nand
  g2633
  (
    n2720,
    n2532,
    n2482,
    n2011,
    n2509
  );


  xor
  g2634
  (
    n2608,
    n464,
    n2499,
    n428,
    n1817
  );


  or
  g2635
  (
    n2716,
    n447,
    n1842,
    n2528,
    n420
  );


  nand
  g2636
  (
    n2756,
    n467,
    n473,
    n1979,
    n1829
  );


  xnor
  g2637
  (
    n2553,
    n2126,
    n499,
    n440,
    n421
  );


  and
  g2638
  (
    n2738,
    n2000,
    n446,
    n2497,
    n2463
  );


  and
  g2639
  (
    n2723,
    n2105,
    n2118,
    n2052,
    n421
  );


  nor
  g2640
  (
    n2558,
    n466,
    n2107,
    n2499,
    n2409
  );


  xnor
  g2641
  (
    n2718,
    n434,
    n2479,
    n1835,
    n2092
  );


  nor
  g2642
  (
    n2765,
    n2124,
    n440,
    n2508,
    n2086
  );


  xnor
  g2643
  (
    n2799,
    n449,
    n2014,
    n1874,
    n1812
  );


  nand
  g2644
  (
    n2785,
    n1822,
    n2005,
    n2083,
    n2514
  );


  nor
  g2645
  (
    n2679,
    n2026,
    n466,
    n1810,
    n2444
  );


  xor
  g2646
  (
    n2617,
    n2095,
    n477,
    n2076,
    n473
  );


  or
  g2647
  (
    n2753,
    n423,
    n487,
    n448,
    n498
  );


  nand
  g2648
  (
    n2641,
    n2531,
    n437,
    n2517,
    n477
  );


  xor
  g2649
  (
    n2541,
    n2457,
    n2513,
    n1913,
    n491
  );


  or
  g2650
  (
    n2547,
    n428,
    n2121,
    n1945,
    n2474
  );


  nor
  g2651
  (
    n2538,
    n2487,
    n2526,
    n500,
    n469
  );


  xnor
  g2652
  (
    n2548,
    n496,
    n431,
    n2512,
    n1982
  );


  nor
  g2653
  (
    n2664,
    n2407,
    n2134,
    n438,
    n1922
  );


  nor
  g2654
  (
    n2686,
    n2121,
    n2520,
    n497,
    n472
  );


  or
  g2655
  (
    n2625,
    n2504,
    n2131,
    n1918,
    n417
  );


  xnor
  g2656
  (
    n2572,
    n2393,
    n2220,
    n2087,
    n432
  );


  xor
  g2657
  (
    n2554,
    n1823,
    n2015,
    n2114,
    n2499
  );


  nor
  g2658
  (
    n2545,
    n416,
    n489,
    n454,
    n2496
  );


  nor
  g2659
  (
    n2612,
    n443,
    n476,
    n446,
    n442
  );


  nor
  g2660
  (
    n2665,
    n1911,
    n477,
    n469,
    n449
  );


  xnor
  g2661
  (
    n2654,
    n2517,
    n2531,
    n478,
    n2003
  );


  and
  g2662
  (
    n2734,
    n488,
    n445,
    n1999,
    n2425
  );


  xor
  g2663
  (
    n2614,
    n472,
    n1976,
    n2470,
    n427
  );


  nand
  g2664
  (
    n2565,
    n501,
    n468,
    n489,
    n454
  );


  or
  g2665
  (
    n2760,
    n2203,
    n449,
    n1916,
    n490
  );


  nor
  g2666
  (
    n2634,
    n2121,
    n2521,
    n2461,
    n2125
  );


  nor
  g2667
  (
    n2546,
    n2130,
    n2117,
    n1954,
    n420
  );


  nand
  g2668
  (
    n2633,
    n450,
    n2531,
    n2067,
    n1955
  );


  xor
  g2669
  (
    n2713,
    n1826,
    n2060,
    n2062,
    n2441
  );


  xnor
  g2670
  (
    n2746,
    n433,
    n492,
    n432,
    n2113
  );


  xnor
  g2671
  (
    n2798,
    n2009,
    n2424,
    n1803,
    n417
  );


  nand
  g2672
  (
    n2552,
    n2524,
    n2008,
    n1937,
    n2421
  );


  nor
  g2673
  (
    n2721,
    n1963,
    n2322,
    n2507,
    n2045
  );


  or
  g2674
  (
    n2637,
    n2529,
    n2473,
    n1895,
    n490
  );


  xor
  g2675
  (
    n2652,
    n2420,
    n1865,
    n490,
    n2510
  );


  and
  g2676
  (
    n2604,
    n2024,
    n2524,
    n472,
    n430
  );


  xnor
  g2677
  (
    KeyWire_0_5,
    n2525,
    n2518,
    n1934,
    n2132
  );


  xnor
  g2678
  (
    n2761,
    n475,
    n2509,
    n500,
    n417
  );


  nor
  g2679
  (
    n2587,
    n2100,
    n2131,
    n456,
    n418
  );


  or
  g2680
  (
    n2696,
    n438,
    n2517,
    n1883,
    n1971
  );


  xnor
  g2681
  (
    n2764,
    n1962,
    n474,
    n2120,
    n2533
  );


  xor
  g2682
  (
    n2690,
    n498,
    n2151,
    n2127,
    n2531
  );


  xor
  g2683
  (
    n2578,
    n486,
    n2323,
    n1881,
    n481
  );


  and
  g2684
  (
    n2747,
    n2132,
    n463,
    n2128,
    n2101
  );


  or
  g2685
  (
    n2569,
    n414,
    n436,
    n2439,
    n2021
  );


  xor
  g2686
  (
    n2594,
    n2511,
    n2013,
    n427
  );


  xor
  g2687
  (
    n2575,
    n1901,
    n434,
    n491,
    n431
  );


  or
  g2688
  (
    n2597,
    n456,
    n1941,
    n1847,
    n1796
  );


  and
  g2689
  (
    n2777,
    n2509,
    n1834,
    n2124,
    n2527
  );


  xnor
  g2690
  (
    n2639,
    n2394,
    n441,
    n424,
    n2122
  );


  or
  g2691
  (
    n2776,
    n1958,
    n2411,
    n438,
    n2472
  );


  or
  g2692
  (
    n2788,
    n2523,
    n458,
    n2412,
    n2529
  );


  or
  g2693
  (
    n2655,
    n2125,
    n2483,
    n431,
    n447
  );


  nor
  g2694
  (
    n2739,
    n2521,
    n2084,
    n2133,
    n2516
  );


  and
  g2695
  (
    n2774,
    n477,
    n484,
    n2133,
    n2497
  );


  nor
  g2696
  (
    n2762,
    n2528,
    n2511,
    n2118,
    n419
  );


  nand
  g2697
  (
    n2740,
    n436,
    n441,
    n452,
    n494
  );


  xor
  g2698
  (
    n2567,
    n1798,
    n1833,
    n2020,
    n2498
  );


  xor
  g2699
  (
    n2688,
    n445,
    n2120,
    n466,
    n2114
  );


  and
  g2700
  (
    n2766,
    n497,
    n1166,
    n2048,
    n2416
  );


  xnor
  g2701
  (
    n2646,
    n1848,
    n2465,
    n2508,
    n467
  );


  xor
  g2702
  (
    n2653,
    n453,
    n2502,
    n418,
    n499
  );


  nand
  g2703
  (
    n2584,
    n2073,
    n448,
    n422,
    n425
  );


  or
  g2704
  (
    n2714,
    n441,
    n1863,
    n501,
    n426
  );


  xor
  g2705
  (
    n2784,
    n1820,
    n1827,
    n470,
    n2119
  );


  xnor
  g2706
  (
    n2537,
    n2535,
    n2119,
    n1851,
    n2152
  );


  xor
  g2707
  (
    n2624,
    n480,
    n464,
    n484,
    n2512
  );


  or
  g2708
  (
    n2752,
    n2398,
    n2046,
    n1959,
    n444
  );


  and
  g2709
  (
    n2684,
    n2410,
    n2129,
    n415,
    n2519
  );


  nand
  g2710
  (
    n2549,
    n2119,
    n480,
    n469,
    n1870
  );


  nor
  g2711
  (
    n2770,
    n1915,
    n1983,
    n2534,
    n1850
  );


  xnor
  g2712
  (
    n2613,
    n1880,
    n431,
    n2042,
    n2130
  );


  and
  g2713
  (
    n2786,
    n1866,
    n2496,
    n458,
    n2429
  );


  or
  g2714
  (
    n2606,
    n2030,
    n2454,
    n2529,
    n2068
  );


  or
  g2715
  (
    n2705,
    n1837,
    n457,
    n2051,
    n2445
  );


  nand
  g2716
  (
    n2618,
    n1802,
    n2510,
    n486,
    n2427
  );


  xor
  g2717
  (
    n2591,
    n427,
    n2522,
    n1876,
    n485
  );


  or
  g2718
  (
    n2648,
    n1868,
    n2001,
    n2126,
    n2518
  );


  and
  g2719
  (
    n2745,
    n1856,
    n1799,
    n455,
    n2322
  );


  or
  g2720
  (
    n2590,
    n2521,
    n2129,
    n2519,
    n2080
  );


  and
  g2721
  (
    n2563,
    n476,
    n2500,
    n1996,
    n1845
  );


  xnor
  g2722
  (
    n2623,
    n1900,
    n2521,
    n1949,
    n440
  );


  xor
  g2723
  (
    n2610,
    n459,
    n482,
    n461,
    n1925
  );


  xnor
  g2724
  (
    n2668,
    n2489,
    n2438,
    n454,
    n2070
  );


  or
  g2725
  (
    n2536,
    n2032,
    n2509,
    n417,
    n428
  );


  nand
  g2726
  (
    n2570,
    n2079,
    n452,
    n2123,
    n442
  );


  and
  g2727
  (
    n2767,
    n1974,
    n460,
    n1952,
    n2490
  );


  nor
  g2728
  (
    n2566,
    n419,
    n2505,
    n414,
    n2423
  );


  or
  g2729
  (
    n2681,
    n422,
    n1926,
    n1852,
    n2520
  );


  and
  g2730
  (
    n2709,
    n2010,
    n2114,
    n1964,
    n2458
  );


  nand
  g2731
  (
    n2622,
    n462,
    n2534,
    n487,
    n486
  );


  nor
  g2732
  (
    n2551,
    n2488,
    n2480,
    n2022,
    n2064
  );


  xnor
  g2733
  (
    n2741,
    n482,
    n450,
    n457,
    n2096
  );


  nor
  g2734
  (
    n2670,
    n2502,
    n2133,
    n429,
    n2115
  );


  xnor
  g2735
  (
    n2727,
    n1882,
    n2535,
    n468,
    n420
  );


  xor
  g2736
  (
    n2650,
    n458,
    n2417,
    n2498,
    n459
  );


  and
  g2737
  (
    n2602,
    n2134,
    n2053,
    n426,
    n462
  );


  xor
  g2738
  (
    n2782,
    n497,
    n2400,
    n2528,
    n1849
  );


  xnor
  g2739
  (
    n2556,
    n498,
    n2533,
    n2518,
    n430
  );


  xor
  g2740
  (
    n2744,
    n436,
    n2515,
    n1920,
    n2126
  );


  xor
  g2741
  (
    n2673,
    n495,
    n1891,
    n2507,
    n426
  );


  xnor
  g2742
  (
    n2677,
    n485,
    n1805,
    n2025,
    n1853
  );


  nand
  g2743
  (
    n2755,
    n435,
    n2523,
    n1978,
    n415
  );


  or
  g2744
  (
    n2540,
    n461,
    n1831,
    n447,
    n2455
  );


  or
  g2745
  (
    n2586,
    n443,
    n1878,
    n2122,
    n494
  );


  nand
  g2746
  (
    n2754,
    n442,
    n1905,
    n1887,
    n2526
  );


  xor
  g2747
  (
    n2626,
    n435,
    n2129,
    n2127,
    n2038
  );


  xnor
  g2748
  (
    n2691,
    n1975,
    n443,
    n465,
    n456
  );


  xnor
  g2749
  (
    n2596,
    n2098,
    n2099,
    n433,
    n1828
  );


  and
  g2750
  (
    n2599,
    n473,
    n2119,
    n2061,
    n1930
  );


  nor
  g2751
  (
    n2735,
    n1813,
    n2152,
    n470,
    n2530
  );


  xnor
  g2752
  (
    n2773,
    n2088,
    n1993,
    n487,
    n450
  );


  or
  g2753
  (
    n2611,
    n493,
    n479,
    n453,
    n461
  );


  xor
  g2754
  (
    n2710,
    n2063,
    n2477,
    n439,
    n2525
  );


  nor
  g2755
  (
    n2619,
    n489,
    n2526,
    n2118,
    n2322
  );


  xnor
  g2756
  (
    n2736,
    n1809,
    n2074,
    n478,
    n2069
  );


  nor
  g2757
  (
    n2582,
    n1861,
    n1908,
    n2018,
    n482
  );


  nor
  g2758
  (
    n2771,
    n2093,
    n1864,
    n2518,
    n2121
  );


  nor
  g2759
  (
    n2749,
    n433,
    n2078,
    n2527,
    n500
  );


  xnor
  g2760
  (
    n2644,
    n1910,
    n2029,
    n2511,
    n2515
  );


  or
  g2761
  (
    n2793,
    n2434,
    n2151,
    n2519,
    n1931
  );


  or
  g2762
  (
    n2724,
    n2524,
    n491,
    n485,
    n1921
  );


  or
  g2763
  (
    n2675,
    n1840,
    n479,
    n2504,
    n496
  );


  xnor
  g2764
  (
    n2568,
    n2124,
    n2090,
    n483,
    n2114
  );


  nand
  g2765
  (
    n2763,
    n444,
    n2535,
    n2499,
    n1939
  );


  nand
  g2766
  (
    n2783,
    n442,
    n2504,
    n2448,
    n2094
  );


  xor
  g2767
  (
    n2585,
    n1927,
    n2475,
    n444,
    n471
  );


  xnor
  g2768
  (
    n2722,
    n446,
    n2406,
    n440,
    n447
  );


  xnor
  g2769
  (
    n2698,
    n2485,
    n1873,
    n1888,
    n437
  );


  nand
  g2770
  (
    n2669,
    n2532,
    n2109,
    n498,
    n441
  );


  nor
  g2771
  (
    n2649,
    n2323,
    n2039,
    n2085,
    n490
  );


  or
  g2772
  (
    n2791,
    n2077,
    n424,
    n2503,
    n470
  );


  nor
  g2773
  (
    n2680,
    n494,
    n434,
    n1797,
    n2496
  );


  or
  g2774
  (
    n2737,
    n423,
    n464,
    n2418,
    n2497
  );


  or
  g2775
  (
    n2808,
    n2786,
    n2777,
    n2696,
    n2621
  );


  xor
  g2776
  (
    n2853,
    n2563,
    n2596,
    n2739,
    n2742
  );


  nor
  g2777
  (
    n2817,
    n2650,
    n2691,
    n2655,
    n2736
  );


  nand
  g2778
  (
    n2815,
    n2746,
    n2597,
    n2758,
    n2616
  );


  xnor
  g2779
  (
    n2820,
    n2669,
    n2683,
    n2545,
    n2725
  );


  nor
  g2780
  (
    n2824,
    n2711,
    n2724,
    n2658,
    n2600
  );


  xor
  g2781
  (
    n2852,
    n2783,
    n2636,
    n2769,
    n2744
  );


  nor
  g2782
  (
    n2813,
    n2543,
    n2751,
    n2699,
    n2720
  );


  and
  g2783
  (
    n2807,
    n2601,
    n2768,
    n2712,
    n2569
  );


  or
  g2784
  (
    n2839,
    n2635,
    n2793,
    n2555,
    n2646
  );


  and
  g2785
  (
    n2819,
    n2564,
    n2755,
    n2790,
    n2659
  );


  and
  g2786
  (
    n2860,
    n2704,
    n2747,
    n2714,
    n2542
  );


  xor
  g2787
  (
    n2803,
    n2690,
    n2578,
    n2750,
    n2678
  );


  or
  g2788
  (
    n2856,
    n2689,
    n2548,
    n2759,
    n2716
  );


  xnor
  g2789
  (
    n2802,
    n2792,
    n2589,
    n2776,
    n2722
  );


  nor
  g2790
  (
    n2864,
    n2730,
    n2713,
    n2587,
    n2681
  );


  xor
  g2791
  (
    n2814,
    n2671,
    n2640,
    n2607,
    n2677
  );


  and
  g2792
  (
    n2809,
    n2623,
    n2595,
    n2694,
    n2546
  );


  xor
  g2793
  (
    n2822,
    n2585,
    n2552,
    n2610,
    n2743
  );


  or
  g2794
  (
    n2812,
    n2710,
    n2784,
    n2727,
    n2664
  );


  nor
  g2795
  (
    n2854,
    n2559,
    n2615,
    n2705,
    n2565
  );


  and
  g2796
  (
    n2831,
    n2673,
    n2741,
    n2684,
    n2656
  );


  nand
  g2797
  (
    n2842,
    n2612,
    n2791,
    n2603,
    n2574
  );


  nor
  g2798
  (
    n2846,
    n2654,
    n2645,
    n2674,
    n2719
  );


  nand
  g2799
  (
    n2828,
    n2707,
    n2773,
    n2576,
    n2570
  );


  and
  g2800
  (
    n2858,
    n2581,
    n2772,
    n2651,
    n2660
  );


  nand
  g2801
  (
    n2806,
    n2794,
    n2631,
    n2622,
    n2785
  );


  nor
  g2802
  (
    n2826,
    n2676,
    n2735,
    n2708,
    n2561
  );


  and
  g2803
  (
    n2836,
    n2787,
    n2675,
    n2605,
    n2731
  );


  xnor
  g2804
  (
    n2804,
    n2551,
    n2630,
    n2609,
    n2706
  );


  nor
  g2805
  (
    n2844,
    n2611,
    n2560,
    n2598,
    n2756
  );


  and
  g2806
  (
    n2861,
    n2703,
    n2771,
    n2682,
    n2637
  );


  or
  g2807
  (
    n2863,
    n2639,
    n2618,
    n2764,
    n2753
  );


  or
  g2808
  (
    n2840,
    n2737,
    n2738,
    n2579,
    n2634
  );


  or
  g2809
  (
    n2855,
    n2663,
    n2586,
    n2672,
    n2572
  );


  nand
  g2810
  (
    n2805,
    n2553,
    n2754,
    n2728,
    n2593
  );


  xnor
  g2811
  (
    n2849,
    n2698,
    n2575,
    n2679,
    n2604
  );


  xnor
  g2812
  (
    n2848,
    n2558,
    n2619,
    n2729,
    n2740
  );


  xor
  g2813
  (
    n2801,
    n2766,
    n2624,
    n2638,
    n2592
  );


  nand
  g2814
  (
    n2832,
    n2680,
    n2748,
    n2625,
    n2617
  );


  nor
  g2815
  (
    n2857,
    n2762,
    n2721,
    n2541,
    n2643
  );


  xor
  g2816
  (
    n2833,
    n2668,
    n2757,
    n2778,
    n2661
  );


  xnor
  g2817
  (
    n2821,
    n2632,
    n2760,
    n2577,
    n2620
  );


  nor
  g2818
  (
    n2862,
    n2539,
    n2795,
    n2780,
    n2614
  );


  xnor
  g2819
  (
    n2829,
    n2775,
    n2688,
    n2538,
    n2599
  );


  and
  g2820
  (
    n2838,
    n2573,
    n2657,
    n2745,
    n2540
  );


  nand
  g2821
  (
    n2834,
    n2591,
    n2765,
    n2761,
    n2692
  );


  nand
  g2822
  (
    n2810,
    n2644,
    n2590,
    n2702,
    n2717
  );


  nor
  g2823
  (
    n2850,
    n2568,
    n2608,
    n2562,
    n2782
  );


  xor
  g2824
  (
    n2845,
    n2613,
    n2781,
    n2549,
    n2709
  );


  and
  g2825
  (
    n2830,
    n2571,
    n2547,
    n2697,
    n2774
  );


  nand
  g2826
  (
    n2818,
    n2715,
    n2718,
    n2554,
    n2536
  );


  or
  g2827
  (
    n2816,
    n2767,
    n2752,
    n2594,
    n2580
  );


  xnor
  g2828
  (
    n2800,
    n2789,
    n2652,
    n2582,
    n2670
  );


  xnor
  g2829
  (
    n2841,
    n2763,
    n2733,
    n2641,
    n2788
  );


  or
  g2830
  (
    n2859,
    n2648,
    n2685,
    n2665,
    n2537
  );


  xnor
  g2831
  (
    n2847,
    n2588,
    n2726,
    n2700,
    n2628
  );


  xor
  g2832
  (
    n2827,
    n2686,
    n2662,
    n2749,
    n2734
  );


  or
  g2833
  (
    n2837,
    n2602,
    n2693,
    n2642,
    n2653
  );


  or
  g2834
  (
    n2843,
    n2629,
    n2550,
    n2557,
    n2732
  );


  and
  g2835
  (
    n2823,
    n2667,
    n2544,
    n2701,
    n2779
  );


  and
  g2836
  (
    n2835,
    n2626,
    n2770,
    n2666,
    n2583
  );


  and
  g2837
  (
    n2811,
    n2695,
    n2566,
    n2687,
    n2556
  );


  nor
  g2838
  (
    n2851,
    n2584,
    n2627,
    n2647,
    n2606
  );


  xor
  g2839
  (
    n2825,
    n2723,
    n2633,
    n2649,
    n2567
  );


  buf
  g2840
  (
    n2867,
    n2806
  );


  buf
  g2841
  (
    n2872,
    n2811
  );


  buf
  g2842
  (
    n2876,
    n2804
  );


  buf
  g2843
  (
    n2865,
    n2809
  );


  buf
  g2844
  (
    n2866,
    n2802
  );


  not
  g2845
  (
    n2874,
    n2813
  );


  not
  g2846
  (
    n2873,
    n2807
  );


  buf
  g2847
  (
    n2878,
    n2801
  );


  not
  g2848
  (
    n2868,
    n2812
  );


  not
  g2849
  (
    n2875,
    n2805
  );


  buf
  g2850
  (
    n2870,
    n2808
  );


  buf
  g2851
  (
    n2871,
    n2803
  );


  buf
  g2852
  (
    n2877,
    n2810
  );


  buf
  g2853
  (
    n2869,
    n2800
  );


  not
  g2854
  (
    n2881,
    n2868
  );


  buf
  g2855
  (
    n2885,
    n2867
  );


  buf
  g2856
  (
    n2884,
    n2868
  );


  buf
  g2857
  (
    n2882,
    n2868
  );


  not
  g2858
  (
    n2880,
    n2866
  );


  not
  g2859
  (
    n2879,
    n2868
  );


  not
  g2860
  (
    n2883,
    n2865
  );


  or
  g2861
  (
    n2893,
    n1171,
    n2875,
    n2279,
    n2336
  );


  and
  g2862
  (
    n2886,
    n2874,
    n2880,
    n2819,
    n2882
  );


  nor
  g2863
  (
    n2903,
    n2883,
    n2871,
    n2885,
    n2878
  );


  nand
  g2864
  (
    n2892,
    n2871,
    n2883,
    n2873,
    n2279
  );


  xnor
  g2865
  (
    n2898,
    n2875,
    n2826,
    n2869,
    n2335
  );


  nor
  g2866
  (
    n2908,
    n2882,
    n2335,
    n2277,
    n2885
  );


  xnor
  g2867
  (
    n2897,
    n2870,
    n2818,
    n2821,
    n2881
  );


  xnor
  g2868
  (
    n2906,
    n2881,
    n2815,
    n2825,
    n2279
  );


  xor
  g2869
  (
    n2889,
    n2816,
    n2878,
    n2276
  );


  or
  g2870
  (
    n2905,
    n2871,
    n2869,
    n2877
  );


  or
  g2871
  (
    n2896,
    n2276,
    n2870,
    n2879,
    n2827
  );


  nand
  g2872
  (
    n2890,
    n2877,
    n2881,
    n2879,
    n2872
  );


  and
  g2873
  (
    n2909,
    n2882,
    n2880,
    n2280,
    n2277
  );


  nand
  g2874
  (
    n2899,
    n2884,
    n2884,
    n2878,
    n2276
  );


  xnor
  g2875
  (
    n2900,
    n2336,
    n2872,
    n2882,
    n2279
  );


  nand
  g2876
  (
    n2888,
    n2822,
    n2883,
    n2881,
    n2873
  );


  nand
  g2877
  (
    n2910,
    n2873,
    n2278,
    n2883,
    n2877
  );


  xor
  g2878
  (
    n2907,
    n2879,
    n2277,
    n2824,
    n2874
  );


  xnor
  g2879
  (
    n2911,
    n2884,
    n2817,
    n2876,
    n2276
  );


  or
  g2880
  (
    n2902,
    n2879,
    n2275,
    n2876,
    n2334
  );


  xor
  g2881
  (
    n2895,
    n2876,
    n2874,
    n2823,
    n2877
  );


  nand
  g2882
  (
    n2887,
    n2880,
    n2278,
    n2870,
    n2875
  );


  nand
  g2883
  (
    n2894,
    n2880,
    n2875,
    n2876,
    n2278
  );


  xor
  g2884
  (
    n2904,
    n2874,
    n2335,
    n2885,
    n2870
  );


  nand
  g2885
  (
    n2913,
    n2872,
    n2820,
    n2280,
    n2814
  );


  xnor
  g2886
  (
    n2891,
    n2873,
    n2884,
    n2277,
    n2869
  );


  nor
  g2887
  (
    n2901,
    n2275,
    n2275,
    n2872,
    n2336
  );


  xor
  g2888
  (
    n2912,
    n2278,
    n2871,
    n2885,
    n2335
  );


  xnor
  g2889
  (
    n3019,
    n2904,
    n1268,
    n1476,
    n1186
  );


  and
  g2890
  (
    n3012,
    n1263,
    n2904,
    n1310,
    n1449
  );


  and
  g2891
  (
    n2946,
    n1406,
    n2897,
    n1326,
    n1413
  );


  nand
  g2892
  (
    n2958,
    n1371,
    n1482,
    n1261,
    n2889
  );


  xor
  g2893
  (
    n2950,
    n1303,
    n2912,
    n1396,
    n1321
  );


  and
  g2894
  (
    n2967,
    n1392,
    n1260,
    n2828,
    n1391
  );


  nor
  g2895
  (
    n3005,
    n1430,
    n1424,
    n1421,
    n2886
  );


  xor
  g2896
  (
    n2932,
    n2900,
    n1372,
    n1225,
    n1337
  );


  xor
  g2897
  (
    n2930,
    n2905,
    n1187,
    n2912,
    n1381
  );


  or
  g2898
  (
    n2947,
    n1264,
    n1368,
    n1477,
    n1415
  );


  or
  g2899
  (
    n2970,
    n1286,
    n2887,
    n1458,
    n1447
  );


  or
  g2900
  (
    n2926,
    n1172,
    n2909,
    n2284,
    n1182
  );


  nor
  g2901
  (
    n2995,
    n1300,
    n1294,
    n1238,
    n1213
  );


  nand
  g2902
  (
    n2933,
    n1332,
    n2282,
    n1357,
    n1444
  );


  nand
  g2903
  (
    n2959,
    n1190,
    n1347,
    n2911,
    n2899
  );


  or
  g2904
  (
    n3007,
    n1464,
    n2913,
    n1414,
    n1317
  );


  nor
  g2905
  (
    n2921,
    n1237,
    n2906,
    n1295,
    n1288
  );


  and
  g2906
  (
    n2939,
    n1226,
    n1240,
    n1282,
    n1446
  );


  nand
  g2907
  (
    n2919,
    n1486,
    n2897,
    n1233,
    n2893
  );


  nand
  g2908
  (
    n2915,
    n2911,
    n1252,
    n1191,
    n2902
  );


  and
  g2909
  (
    n2987,
    n1276,
    n1407,
    n1232,
    n2281
  );


  xor
  g2910
  (
    n2957,
    n1196,
    n1433,
    n1390,
    n1229
  );


  or
  g2911
  (
    n2928,
    n1253,
    n1367,
    n1230,
    n1203
  );


  xnor
  g2912
  (
    n3022,
    n1179,
    n2888,
    n1445
  );


  xor
  g2913
  (
    n2997,
    n1360,
    n1275,
    n1206,
    n1409
  );


  xnor
  g2914
  (
    n2991,
    n1320,
    n2902,
    n1331,
    n1296
  );


  xor
  g2915
  (
    n2934,
    n2909,
    n2892,
    n1370,
    n1345
  );


  and
  g2916
  (
    n3020,
    n2908,
    n1198,
    n2888,
    n2905
  );


  nor
  g2917
  (
    n2948,
    n1395,
    n1343,
    n1218,
    n1329
  );


  nand
  g2918
  (
    n2960,
    n1224,
    n1359,
    n1488,
    n2280
  );


  or
  g2919
  (
    n3010,
    n1420,
    n1327,
    n1346,
    n1183
  );


  or
  g2920
  (
    n2977,
    n1463,
    n1195,
    n1350,
    n1279
  );


  or
  g2921
  (
    n3021,
    n1308,
    n1278,
    n1416,
    n2901
  );


  xnor
  g2922
  (
    n2966,
    n1451,
    n2912,
    n1349,
    n2904
  );


  nand
  g2923
  (
    n2982,
    n1313,
    n1324,
    n1478,
    n2892
  );


  nor
  g2924
  (
    n2993,
    n1319,
    n1456,
    n1184,
    n1304
  );


  or
  g2925
  (
    n2974,
    n1484,
    n1358,
    n1335,
    n2902
  );


  nor
  g2926
  (
    n3002,
    n1242,
    n2886,
    n1292,
    n1334
  );


  or
  g2927
  (
    n2918,
    n1417,
    n1418,
    n2896,
    n2913
  );


  xor
  g2928
  (
    n2992,
    n2284,
    n1199,
    n1475,
    n1425
  );


  xor
  g2929
  (
    n3023,
    n2896,
    n2890,
    n2906,
    n2899
  );


  nor
  g2930
  (
    n2917,
    n1379,
    n2283,
    n2912,
    n1411
  );


  or
  g2931
  (
    n2961,
    n1364,
    n1221,
    n1204,
    n2891
  );


  xor
  g2932
  (
    n3013,
    n1384,
    n1442,
    n1339,
    n2909
  );


  or
  g2933
  (
    n2938,
    n2906,
    n1215,
    n2896,
    n2908
  );


  or
  g2934
  (
    n2956,
    n1272,
    n2282,
    n1454,
    n2899
  );


  xnor
  g2935
  (
    n2923,
    n2892,
    n2889,
    n1312,
    n1353
  );


  xor
  g2936
  (
    n2954,
    n2891,
    n2900,
    n2280,
    n1375
  );


  or
  g2937
  (
    n2994,
    n1254,
    n1479,
    n1440,
    n1257
  );


  xor
  g2938
  (
    n2914,
    n2898,
    n1205,
    n1373,
    n1231
  );


  nand
  g2939
  (
    n2978,
    n1267,
    n1382,
    n2908,
    n1438
  );


  xnor
  g2940
  (
    n2931,
    n1471,
    n2891,
    n1265,
    n2899
  );


  xor
  g2941
  (
    n2935,
    n1462,
    n1262,
    n1466,
    n2283
  );


  or
  g2942
  (
    n2924,
    n1419,
    n1251,
    n1448,
    n2887
  );


  xnor
  g2943
  (
    n3015,
    n1287,
    n1378,
    n1428,
    n1338
  );


  and
  g2944
  (
    n3014,
    n1173,
    n2281,
    n1220,
    n2901
  );


  nor
  g2945
  (
    n3003,
    n1325,
    n1361,
    n1427,
    n1185
  );


  or
  g2946
  (
    n2951,
    n1468,
    n1309,
    n2903,
    n1188
  );


  or
  g2947
  (
    n2996,
    n1298,
    n1209,
    n2896,
    n2907
  );


  xnor
  g2948
  (
    n2981,
    n1250,
    n1328,
    n2282,
    n1452
  );


  nand
  g2949
  (
    n2979,
    n1178,
    n1470,
    n2905,
    n2283
  );


  or
  g2950
  (
    KeyWire_0_23,
    n1344,
    n2894,
    n1259,
    n1469
  );


  and
  g2951
  (
    n2942,
    n2891,
    n1394,
    n1403,
    n1437
  );


  or
  g2952
  (
    n3009,
    n2893,
    n2886,
    n1284,
    n2905
  );


  and
  g2953
  (
    n2952,
    n1431,
    n2897,
    n1236,
    n1239
  );


  or
  g2954
  (
    n2944,
    n1366,
    n1393,
    n2907,
    n1228
  );


  nand
  g2955
  (
    n2969,
    n1227,
    n1351,
    n2890,
    n1336
  );


  and
  g2956
  (
    n3017,
    n1241,
    n1374,
    n1429,
    n2898
  );


  xnor
  g2957
  (
    n2929,
    n1271,
    n1376,
    n1333,
    n1404
  );


  xnor
  g2958
  (
    n2925,
    n1245,
    n1302,
    n1352,
    n2281
  );


  and
  g2959
  (
    n2920,
    n1299,
    n1387,
    n1210,
    n1340
  );


  or
  g2960
  (
    n2936,
    n2895,
    n1247,
    n2910,
    n1175
  );


  nor
  g2961
  (
    n2973,
    n1219,
    n1255,
    n2895,
    n1244
  );


  xor
  g2962
  (
    n3018,
    n1256,
    n1342,
    n1483,
    n1281
  );


  and
  g2963
  (
    n2963,
    n2900,
    n2900,
    n2903,
    n2895
  );


  nor
  g2964
  (
    n2945,
    n1269,
    n1305,
    n1480,
    n2903
  );


  and
  g2965
  (
    n2943,
    n1297,
    n1461,
    n1274,
    n1356
  );


  xor
  g2966
  (
    n2989,
    n2887,
    n1283,
    n1405,
    n2889
  );


  and
  g2967
  (
    n2972,
    n2913,
    n1412,
    n1362,
    n1365
  );


  nand
  g2968
  (
    n2990,
    n1441,
    n2895,
    n1280,
    n1485
  );


  xnor
  g2969
  (
    n2949,
    n2890,
    n1398,
    n1216,
    n2908
  );


  nand
  g2970
  (
    n2988,
    n1306,
    n1181,
    n2889,
    n1348
  );


  and
  g2971
  (
    n2968,
    n1243,
    n1214,
    n1249,
    n1180
  );


  nand
  g2972
  (
    n2916,
    n1467,
    n1318,
    n1323,
    n1439
  );


  and
  g2973
  (
    KeyWire_0_18,
    n1194,
    n1289,
    n1246,
    n1273
  );


  nor
  g2974
  (
    n2999,
    n1234,
    n1487,
    n1201,
    n1341
  );


  xor
  g2975
  (
    n2940,
    n2913,
    n2910,
    n1457,
    n1266
  );


  nor
  g2976
  (
    n2962,
    n1277,
    n1363,
    n2897,
    n1453
  );


  or
  g2977
  (
    n3001,
    n1389,
    n2910,
    n1174,
    n1223
  );


  xnor
  g2978
  (
    n2941,
    n1402,
    n1397,
    n1385,
    n1436
  );


  nand
  g2979
  (
    n2927,
    n1193,
    n1465,
    n2887,
    n1330
  );


  nand
  g2980
  (
    n2984,
    n1426,
    n2284,
    n1177,
    n1212
  );


  nand
  g2981
  (
    n2955,
    n1197,
    n1200,
    n2894,
    n1474
  );


  xnor
  g2982
  (
    n3008,
    n2893,
    n2910,
    n2903,
    n1401
  );


  or
  g2983
  (
    n2976,
    n1450,
    n1176,
    n1316,
    n1432
  );


  or
  g2984
  (
    n2922,
    n2284,
    n2281,
    n1434,
    n1443
  );


  and
  g2985
  (
    n2983,
    n1380,
    n1290,
    n1293,
    n2888
  );


  nand
  g2986
  (
    n3025,
    n1248,
    n2894,
    n1258
  );


  and
  g2987
  (
    n3016,
    n2911,
    n2904,
    n1459,
    n1388
  );


  nor
  g2988
  (
    n2965,
    n2907,
    n1423,
    n1472,
    n1410
  );


  nand
  g2989
  (
    n2971,
    n1314,
    n2282,
    n2909,
    n2901
  );


  or
  g2990
  (
    n2964,
    n1235,
    n2898,
    n2906,
    n1315
  );


  and
  g2991
  (
    n2985,
    n1399,
    n2898,
    n1285,
    n1386
  );


  xor
  g2992
  (
    n3024,
    n2283,
    n1208,
    n2901,
    n1377
  );


  nand
  g2993
  (
    n3006,
    n2902,
    n1435,
    n1270,
    n1192
  );


  and
  g2994
  (
    n2980,
    n1322,
    n1222,
    n1291,
    n1217
  );


  nand
  g2995
  (
    n3004,
    n1211,
    n1400,
    n1383,
    n1355
  );


  xnor
  g2996
  (
    n2986,
    n1202,
    n2890,
    n1369,
    n1481
  );


  or
  g2997
  (
    n2953,
    n1422,
    n1307,
    n1301,
    n2886
  );


  xor
  g2998
  (
    n3000,
    n1354,
    n1311,
    n1460,
    n2907
  );


  xnor
  g2999
  (
    n2998,
    n1207,
    n1473,
    n1408,
    n1189
  );


  nand
  g3000
  (
    n2937,
    n2893,
    n2892,
    n1455,
    n2911
  );


  xor
  g3001
  (
    n3047,
    n2951,
    n2160,
    n2166,
    n2162
  );


  or
  g3002
  (
    n3063,
    n2169,
    n2224,
    n2845,
    n2969
  );


  or
  g3003
  (
    n3087,
    n2955,
    n2161,
    n2184,
    n2917
  );


  nand
  g3004
  (
    n3028,
    n2184,
    n2169,
    n2221,
    n3013
  );


  and
  g3005
  (
    n3048,
    n2165,
    n2915,
    n2182,
    n2841
  );


  xor
  g3006
  (
    n3081,
    n2171,
    n2156,
    n3000,
    n2829
  );


  and
  g3007
  (
    n3043,
    n2178,
    n2982,
    n2993,
    n2992
  );


  xor
  g3008
  (
    n3040,
    n2926,
    n2181,
    n2921,
    n2164
  );


  nand
  g3009
  (
    n3082,
    n3018,
    n2972,
    n2183,
    n2930
  );


  or
  g3010
  (
    n3026,
    n2157,
    n2975,
    n2932,
    n2209
  );


  nand
  g3011
  (
    KeyWire_0_3,
    n2183,
    n2188,
    n2842,
    n2167
  );


  nand
  g3012
  (
    n3027,
    n2946,
    n2162,
    n2158,
    n2207
  );


  nand
  g3013
  (
    n3033,
    n2156,
    n2173,
    n2321,
    n2175
  );


  and
  g3014
  (
    n3080,
    n2916,
    n2172,
    n2956,
    n2173
  );


  xnor
  g3015
  (
    n3074,
    n2966,
    n2172,
    n2156,
    n2170
  );


  and
  g3016
  (
    n3062,
    n2187,
    n2994,
    n2206,
    n2174
  );


  nand
  g3017
  (
    n3031,
    n2164,
    n2225,
    n3023,
    n2258
  );


  nand
  g3018
  (
    n3038,
    n2208,
    n2925,
    n2177,
    n2160
  );


  and
  g3019
  (
    n3029,
    n2180,
    n2205,
    n2964,
    n2168
  );


  xnor
  g3020
  (
    n3092,
    n2171,
    n2173,
    n2203,
    n3006
  );


  nor
  g3021
  (
    n3057,
    n2160,
    n2952,
    n2178,
    n2166
  );


  nand
  g3022
  (
    n3069,
    n2185,
    n2844,
    n2959,
    n3010
  );


  and
  g3023
  (
    n3058,
    n2963,
    n2974,
    n2209,
    n2984
  );


  and
  g3024
  (
    n3077,
    n3005,
    n2189,
    n2176,
    n3003
  );


  nand
  g3025
  (
    n3061,
    n2179,
    n2163,
    n2838,
    n2207
  );


  nor
  g3026
  (
    n3037,
    n2190,
    n2175,
    n2976,
    n2184
  );


  xor
  g3027
  (
    n3055,
    n2205,
    n2181,
    n2999,
    n2182
  );


  nor
  g3028
  (
    n3068,
    n2168,
    n2206,
    n2185,
    n2165
  );


  xnor
  g3029
  (
    n3091,
    n2185,
    n2934,
    n2169,
    n2168
  );


  xor
  g3030
  (
    n3042,
    n2950,
    n2169,
    n2167,
    n2161
  );


  nand
  g3031
  (
    n3099,
    n2258,
    n2190,
    n2188,
    n2939
  );


  or
  g3032
  (
    n3071,
    n2961,
    n2987,
    n2998,
    n2920
  );


  or
  g3033
  (
    n3097,
    n2948,
    n2180,
    n2942,
    n2155
  );


  and
  g3034
  (
    n3089,
    n2178,
    n2208,
    n2161,
    n2164
  );


  xor
  g3035
  (
    n3053,
    n2936,
    n2941,
    n2208,
    n2923
  );


  nor
  g3036
  (
    n3085,
    n2973,
    n2321,
    n2155,
    n2931
  );


  and
  g3037
  (
    n3030,
    n2160,
    n2837,
    n2174,
    n2163
  );


  xor
  g3038
  (
    n3052,
    n2991,
    n2937,
    n2177,
    n2163
  );


  xor
  g3039
  (
    n3096,
    n2846,
    n2321,
    n2940,
    n2172
  );


  xor
  g3040
  (
    n3104,
    n2848,
    n3012,
    n2843,
    n2258
  );


  or
  g3041
  (
    n3102,
    n2204,
    n2207,
    n2175,
    n2187
  );


  and
  g3042
  (
    n3049,
    n2164,
    n2166,
    n2186,
    n2830
  );


  nor
  g3043
  (
    n3065,
    n2205,
    n2177,
    n2180,
    n2938
  );


  xor
  g3044
  (
    n3094,
    n3014,
    n2176,
    n2835,
    n2159
  );


  nand
  g3045
  (
    n3078,
    n2836,
    n2173,
    n3020,
    n2181
  );


  nand
  g3046
  (
    n3070,
    n2176,
    n2177,
    n2183,
    n2943
  );


  or
  g3047
  (
    n3056,
    n3021,
    n2949,
    n2161,
    n3011
  );


  xnor
  g3048
  (
    n3083,
    n2914,
    n3019,
    n3007,
    n2163
  );


  or
  g3049
  (
    n3090,
    n3017,
    n2981,
    n2154,
    n2958
  );


  nor
  g3050
  (
    n3050,
    n2176,
    n2204,
    n2209,
    n3002
  );


  or
  g3051
  (
    n3075,
    n3015,
    n2178,
    n2922,
    n2971
  );


  xnor
  g3052
  (
    n3098,
    n2935,
    n2967,
    n3001,
    n2978
  );


  or
  g3053
  (
    n3044,
    n2175,
    n2209,
    n2159,
    n2832
  );


  and
  g3054
  (
    n3079,
    n2995,
    n2933,
    n2957,
    n2182
  );


  and
  g3055
  (
    n3046,
    n2186,
    n2206,
    n3009,
    n2179
  );


  xor
  g3056
  (
    n3066,
    n2167,
    n2172,
    n2174,
    n2321
  );


  xor
  g3057
  (
    n3064,
    n2928,
    n2189,
    n2320,
    n2162
  );


  xnor
  g3058
  (
    n3072,
    n2154,
    n2831,
    n2186,
    n2179
  );


  and
  g3059
  (
    n3060,
    n2208,
    n2187,
    n2223,
    n2186
  );


  or
  g3060
  (
    n3101,
    n2187,
    n2158,
    n2954,
    n2944
  );


  nand
  g3061
  (
    n3032,
    n2927,
    n2989,
    n2165,
    n2159
  );


  nor
  g3062
  (
    n3067,
    n2833,
    n2988,
    n2181,
    n2970
  );


  nand
  g3063
  (
    n3034,
    n2204,
    n2183,
    n2986,
    n2924
  );


  xor
  g3064
  (
    n3093,
    n2184,
    n2180,
    n2207,
    n2962
  );


  or
  g3065
  (
    n3054,
    n2996,
    n2188,
    n2945,
    n2190
  );


  and
  g3066
  (
    n3103,
    n2171,
    n2919,
    n2155,
    n3025
  );


  xnor
  g3067
  (
    n3084,
    n2174,
    n2847,
    n2997,
    n2162
  );


  and
  g3068
  (
    n3039,
    n2977,
    n2947,
    n2190,
    n2980
  );


  or
  g3069
  (
    n3059,
    n3004,
    n2166,
    n2188,
    n2167
  );


  nand
  g3070
  (
    n3036,
    n3016,
    n2189,
    n2159,
    n2157
  );


  nor
  g3071
  (
    n3045,
    n2918,
    n3008,
    n2206,
    n2985
  );


  and
  g3072
  (
    n3073,
    n2179,
    n3024,
    n3022,
    n2839
  );


  or
  g3073
  (
    n3035,
    n2170,
    n2990,
    n2979,
    n2157
  );


  xnor
  g3074
  (
    n3086,
    n2222,
    n2170,
    n2171,
    n2960
  );


  and
  g3075
  (
    n3100,
    n2158,
    n2157,
    n2168,
    n2189
  );


  nor
  g3076
  (
    n3041,
    n2965,
    n2204,
    n2929,
    n2840
  );


  or
  g3077
  (
    n3095,
    n2983,
    n2170,
    n2156,
    n2185
  );


  xnor
  g3078
  (
    n3076,
    n2155,
    n2182,
    n2165,
    n2205
  );


  or
  g3079
  (
    n3088,
    n2834,
    n2968,
    n2953,
    n2158
  );


  nand
  g3080
  (
    n3119,
    n3051,
    n3080,
    n3039,
    n3059
  );


  xor
  g3081
  (
    n3108,
    n3072,
    n2859,
    n3054,
    n3087
  );


  nor
  g3082
  (
    n3116,
    n3050,
    n3101,
    n2864,
    n3055
  );


  xor
  g3083
  (
    n3113,
    n3098,
    n2338,
    n3060,
    n2851
  );


  nand
  g3084
  (
    n3118,
    n3041,
    n2861,
    n3095,
    n2857
  );


  xnor
  g3085
  (
    n3117,
    n2855,
    n3104,
    n3096,
    n3053
  );


  xor
  g3086
  (
    n3122,
    n3100,
    n2860,
    n3084,
    n3036
  );


  xor
  g3087
  (
    n3115,
    n3089,
    n3074,
    n2338,
    n3048
  );


  nand
  g3088
  (
    n3123,
    n2798,
    n3057,
    n3027,
    n2850
  );


  or
  g3089
  (
    n3126,
    n3032,
    n3042,
    n2338,
    n3077
  );


  nand
  g3090
  (
    n3120,
    n3097,
    n3035,
    n3056,
    n3086
  );


  or
  g3091
  (
    n3106,
    n3065,
    n3043,
    n3070,
    n3090
  );


  nor
  g3092
  (
    n3131,
    n2337,
    n3085,
    n3064,
    n2849
  );


  or
  g3093
  (
    n3111,
    n2863,
    n3066,
    n3063,
    n2852
  );


  and
  g3094
  (
    n3130,
    n3026,
    n3079,
    n3028,
    n3069
  );


  xor
  g3095
  (
    n3125,
    n3031,
    n2338,
    n2799,
    n2797
  );


  or
  g3096
  (
    n3114,
    n2337,
    n3049,
    n3093,
    n3092
  );


  and
  g3097
  (
    n3105,
    n3062,
    n3040,
    n3045,
    n3081
  );


  nand
  g3098
  (
    n3109,
    n3034,
    n3061,
    n3091,
    n3046
  );


  or
  g3099
  (
    n3110,
    n3067,
    n3071,
    n3102,
    n2337
  );


  and
  g3100
  (
    n3128,
    n3068,
    n3078,
    n2796,
    n2862
  );


  or
  g3101
  (
    n3129,
    n3099,
    n3058,
    n3094,
    n3076
  );


  or
  g3102
  (
    n3127,
    n3073,
    n3082,
    n2336,
    n3083
  );


  nor
  g3103
  (
    n3107,
    n3103,
    n3052,
    n3029,
    n2853
  );


  nand
  g3104
  (
    n3112,
    n3047,
    n2858,
    n3030,
    n3075
  );


  xnor
  g3105
  (
    n3121,
    n3037,
    n2337,
    n3038,
    n3088
  );


  nor
  g3106
  (
    n3124,
    n3033,
    n2856,
    n2854,
    n3044
  );


  xor
  KeyGate_0_0
  (
    n390,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n2350,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n2072,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n3051,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1946,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n2660,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n2628,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n490,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n529,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1253,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n850,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n2205,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n236,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n257,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1672,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1001,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1736,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n2116,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n2975,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n2335,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n2285,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1201,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n2065,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n3011,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1336,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1629,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n447,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n676,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n2647,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1389,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n2175,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n998,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

