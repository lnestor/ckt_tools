

module Stat_1940_64_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n165,
  n347,
  n350,
  n588,
  n584,
  n587,
  n581,
  n582,
  n904,
  n910,
  n1958,
  n1959,
  n1954,
  n1965,
  n1960,
  n1964,
  n1950,
  n1955,
  n1962,
  n1957,
  n1948,
  n1952,
  n1963,
  n1966,
  n1951,
  n1961,
  n1956,
  n1949,
  n1953
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n165;output n347;output n350;output n588;output n584;output n587;output n581;output n582;output n904;output n910;output n1958;output n1959;output n1954;output n1965;output n1960;output n1964;output n1950;output n1955;output n1962;output n1957;output n1948;output n1952;output n1963;output n1966;output n1951;output n1961;output n1956;output n1949;output n1953;
  wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n348;wire n349;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n583;wire n585;wire n586;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n905;wire n906;wire n907;wire n908;wire n909;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n28,
    n1
  );


  buf
  g1
  (
    n27,
    n2
  );


  not
  g2
  (
    n30,
    n1
  );


  not
  g3
  (
    n31,
    n1
  );


  buf
  g4
  (
    n29,
    n1
  );


  buf
  g5
  (
    n49,
    n27
  );


  buf
  g6
  (
    n38,
    n28
  );


  not
  g7
  (
    KeyWire_0_9,
    n27
  );


  not
  g8
  (
    n48,
    n29
  );


  not
  g9
  (
    n40,
    n30
  );


  not
  g10
  (
    n42,
    n28
  );


  buf
  g11
  (
    n47,
    n27
  );


  buf
  g12
  (
    n45,
    n30
  );


  buf
  g13
  (
    n43,
    n30
  );


  buf
  g14
  (
    n44,
    n30
  );


  not
  g15
  (
    n32,
    n28
  );


  buf
  g16
  (
    n41,
    n29
  );


  not
  g17
  (
    n33,
    n29
  );


  buf
  g18
  (
    n35,
    n28
  );


  buf
  g19
  (
    n37,
    n27
  );


  not
  g20
  (
    n39,
    n29
  );


  not
  g21
  (
    n34,
    n31
  );


  buf
  g22
  (
    n46,
    n31
  );


  not
  g23
  (
    n96,
    n43
  );


  buf
  g24
  (
    n111,
    n42
  );


  not
  g25
  (
    n60,
    n46
  );


  buf
  g26
  (
    n77,
    n36
  );


  not
  g27
  (
    n110,
    n42
  );


  buf
  g28
  (
    n75,
    n43
  );


  buf
  g29
  (
    n105,
    n36
  );


  buf
  g30
  (
    n89,
    n41
  );


  buf
  g31
  (
    n101,
    n35
  );


  not
  g32
  (
    n92,
    n46
  );


  not
  g33
  (
    n86,
    n36
  );


  not
  g34
  (
    n91,
    n42
  );


  buf
  g35
  (
    n70,
    n35
  );


  buf
  g36
  (
    n95,
    n45
  );


  buf
  g37
  (
    n118,
    n49
  );


  not
  g38
  (
    n107,
    n38
  );


  buf
  g39
  (
    n106,
    n36
  );


  not
  g40
  (
    n83,
    n46
  );


  not
  g41
  (
    n69,
    n33
  );


  buf
  g42
  (
    n66,
    n32
  );


  buf
  g43
  (
    n99,
    n35
  );


  buf
  g44
  (
    n50,
    n41
  );


  not
  g45
  (
    n56,
    n33
  );


  buf
  g46
  (
    n102,
    n46
  );


  buf
  g47
  (
    n74,
    n40
  );


  buf
  g48
  (
    n82,
    n42
  );


  buf
  g49
  (
    n78,
    n38
  );


  not
  g50
  (
    n112,
    n40
  );


  not
  g51
  (
    n87,
    n37
  );


  buf
  g52
  (
    n55,
    n48
  );


  buf
  g53
  (
    n98,
    n32
  );


  not
  g54
  (
    n72,
    n32
  );


  buf
  g55
  (
    n71,
    n33
  );


  buf
  g56
  (
    n97,
    n40
  );


  buf
  g57
  (
    n93,
    n44
  );


  buf
  g58
  (
    n114,
    n39
  );


  not
  g59
  (
    n52,
    n34
  );


  buf
  g60
  (
    n68,
    n44
  );


  buf
  g61
  (
    n73,
    n39
  );


  not
  g62
  (
    n117,
    n48
  );


  not
  g63
  (
    n104,
    n32
  );


  buf
  g64
  (
    n109,
    n45
  );


  not
  g65
  (
    n85,
    n33
  );


  not
  g66
  (
    n51,
    n47
  );


  not
  g67
  (
    n108,
    n40
  );


  not
  g68
  (
    n81,
    n44
  );


  buf
  g69
  (
    n67,
    n48
  );


  not
  g70
  (
    n90,
    n47
  );


  not
  g71
  (
    n63,
    n38
  );


  not
  g72
  (
    n88,
    n48
  );


  not
  g73
  (
    n80,
    n47
  );


  not
  g74
  (
    n94,
    n44
  );


  buf
  g75
  (
    n62,
    n34
  );


  buf
  g76
  (
    KeyWire_0_26,
    n35
  );


  not
  g77
  (
    n64,
    n37
  );


  not
  g78
  (
    n115,
    n47
  );


  buf
  g79
  (
    n58,
    n45
  );


  not
  g80
  (
    n84,
    n34
  );


  buf
  g81
  (
    n59,
    n34
  );


  not
  g82
  (
    n103,
    n39
  );


  buf
  g83
  (
    n53,
    n43
  );


  buf
  g84
  (
    n113,
    n43
  );


  not
  g85
  (
    n57,
    n41
  );


  buf
  g86
  (
    n100,
    n37
  );


  buf
  g87
  (
    n76,
    n45
  );


  buf
  g88
  (
    n79,
    n37
  );


  not
  g89
  (
    n116,
    n39
  );


  not
  g90
  (
    n65,
    n41
  );


  not
  g91
  (
    n61,
    n38
  );


  not
  g92
  (
    n119,
    n50
  );


  not
  g93
  (
    n120,
    n50
  );


  buf
  g94
  (
    n127,
    n120
  );


  not
  g95
  (
    n121,
    n119
  );


  not
  g96
  (
    n126,
    n120
  );


  not
  g97
  (
    n128,
    n120
  );


  buf
  g98
  (
    n124,
    n120
  );


  not
  g99
  (
    n125,
    n119
  );


  not
  g100
  (
    n123,
    n119
  );


  not
  g101
  (
    n122,
    n119
  );


  xnor
  g102
  (
    n133,
    n123,
    n19
  );


  or
  g103
  (
    n150,
    n14,
    n16,
    n22,
    n15
  );


  or
  g104
  (
    n129,
    n2,
    n4,
    n19,
    n124
  );


  nor
  g105
  (
    n153,
    n20,
    n21,
    n16,
    n5
  );


  xnor
  g106
  (
    n143,
    n16,
    n122,
    n7,
    n12
  );


  nand
  g107
  (
    n154,
    n6,
    n19,
    n24,
    n10
  );


  nand
  g108
  (
    n149,
    n127,
    n18,
    n23,
    n6
  );


  and
  g109
  (
    n132,
    n126,
    n9,
    n25,
    n121
  );


  or
  g110
  (
    n140,
    n14,
    n16,
    n20,
    n5
  );


  xor
  g111
  (
    n141,
    n17,
    n11,
    n24,
    n2
  );


  nor
  g112
  (
    n142,
    n17,
    n123,
    n13,
    n12
  );


  and
  g113
  (
    n157,
    n4,
    n7,
    n123
  );


  xor
  g114
  (
    n131,
    n124,
    n15,
    n21,
    n6
  );


  nor
  g115
  (
    n152,
    n14,
    n121,
    n3,
    n21
  );


  nand
  g116
  (
    n134,
    n121,
    n22,
    n9,
    n25
  );


  nor
  g117
  (
    n130,
    n128,
    n127,
    n22
  );


  nor
  g118
  (
    n159,
    n8,
    n3,
    n126,
    n25
  );


  and
  g119
  (
    n158,
    n128,
    n128,
    n124,
    n8
  );


  nor
  g120
  (
    n147,
    n125,
    n125,
    n13,
    n20
  );


  and
  g121
  (
    n148,
    n9,
    n2,
    n18,
    n10
  );


  and
  g122
  (
    n137,
    n24,
    n125,
    n124,
    n4
  );


  nor
  g123
  (
    n136,
    n10,
    n18,
    n6,
    n13
  );


  nor
  g124
  (
    n151,
    n125,
    n15,
    n23,
    n126
  );


  or
  g125
  (
    n156,
    n14,
    n15,
    n5,
    n127
  );


  nand
  g126
  (
    n139,
    n24,
    n10,
    n11,
    n12
  );


  nor
  g127
  (
    n160,
    n9,
    n11,
    n18,
    n23
  );


  xnor
  g128
  (
    n135,
    n8,
    n128,
    n19,
    n21
  );


  nor
  g129
  (
    n155,
    n123,
    n122,
    n22,
    n8
  );


  or
  g130
  (
    n146,
    n3,
    n122,
    n23,
    n13
  );


  or
  g131
  (
    n145,
    n11,
    n122,
    n7,
    n3
  );


  and
  g132
  (
    n144,
    n20,
    n121,
    n12,
    n126
  );


  nand
  g133
  (
    n138,
    n4,
    n17,
    n5
  );


  not
  g134
  (
    n183,
    n138
  );


  buf
  g135
  (
    n172,
    n144
  );


  buf
  g136
  (
    n162,
    n131
  );


  buf
  g137
  (
    n193,
    n137
  );


  not
  g138
  (
    n188,
    n133
  );


  buf
  g139
  (
    n168,
    n138
  );


  not
  g140
  (
    n164,
    n134
  );


  buf
  g141
  (
    n173,
    n144
  );


  not
  g142
  (
    n166,
    n135
  );


  buf
  g143
  (
    n175,
    n139
  );


  not
  g144
  (
    n192,
    n133
  );


  buf
  g145
  (
    n169,
    n140
  );


  buf
  g146
  (
    n181,
    n134
  );


  not
  g147
  (
    n191,
    n139
  );


  not
  g148
  (
    n194,
    n139
  );


  not
  g149
  (
    n189,
    n135
  );


  not
  g150
  (
    n184,
    n137
  );


  buf
  g151
  (
    n199,
    n143
  );


  not
  g152
  (
    n197,
    n132
  );


  not
  g153
  (
    n177,
    n138
  );


  not
  g154
  (
    n161,
    n130
  );


  not
  g155
  (
    n176,
    n143
  );


  buf
  g156
  (
    n178,
    n141
  );


  not
  g157
  (
    n174,
    n140
  );


  not
  g158
  (
    n195,
    n137
  );


  buf
  g159
  (
    n198,
    n143
  );


  not
  g160
  (
    n179,
    n131
  );


  buf
  g161
  (
    n167,
    n129
  );


  buf
  g162
  (
    n170,
    n141
  );


  not
  g163
  (
    n171,
    n140
  );


  not
  g164
  (
    n187,
    n129
  );


  buf
  g165
  (
    n180,
    n141
  );


  not
  g166
  (
    n163,
    n136
  );


  not
  g167
  (
    n165,
    n142
  );


  buf
  g168
  (
    n196,
    n142
  );


  buf
  g169
  (
    n182,
    n142
  );


  not
  g170
  (
    n186,
    n136
  );


  not
  g171
  (
    n185,
    n132
  );


  buf
  g172
  (
    n190,
    n130
  );


  buf
  g173
  (
    n213,
    n166
  );


  buf
  g174
  (
    n205,
    n177
  );


  not
  g175
  (
    n214,
    n162
  );


  not
  g176
  (
    n200,
    n180
  );


  not
  g177
  (
    n203,
    n176
  );


  not
  g178
  (
    n217,
    n167
  );


  not
  g179
  (
    n210,
    n172
  );


  buf
  g180
  (
    n204,
    n174
  );


  buf
  g181
  (
    n215,
    n178
  );


  not
  g182
  (
    n202,
    n171
  );


  buf
  g183
  (
    n207,
    n165
  );


  buf
  g184
  (
    n206,
    n161
  );


  not
  g185
  (
    n212,
    n163
  );


  not
  g186
  (
    n216,
    n173
  );


  not
  g187
  (
    n209,
    n164
  );


  buf
  g188
  (
    n201,
    n175
  );


  not
  g189
  (
    n218,
    n170
  );


  buf
  g190
  (
    n211,
    n168
  );


  buf
  g191
  (
    n208,
    n169
  );


  not
  g192
  (
    n219,
    n179
  );


  nand
  g193
  (
    n227,
    n62,
    n105,
    n71,
    n58
  );


  xnor
  g194
  (
    n244,
    n70,
    n71,
    n55,
    n100
  );


  nor
  g195
  (
    n256,
    n91,
    n77,
    n69,
    n102
  );


  nand
  g196
  (
    n285,
    n101,
    n104,
    n102
  );


  nor
  g197
  (
    n225,
    n52,
    n212,
    n82,
    n77
  );


  nor
  g198
  (
    n286,
    n218,
    n87,
    n216,
    n52
  );


  or
  g199
  (
    n279,
    n55,
    n91,
    n97
  );


  and
  g200
  (
    n271,
    n84,
    n213,
    n100,
    n54
  );


  xnor
  g201
  (
    n240,
    n99,
    n209,
    n206,
    n71
  );


  xor
  g202
  (
    n230,
    n70,
    n93,
    n83,
    n200
  );


  nor
  g203
  (
    n234,
    n63,
    n77,
    n200,
    n211
  );


  nand
  g204
  (
    n263,
    n206,
    n58,
    n205,
    n55
  );


  nor
  g205
  (
    n291,
    n53,
    n86,
    n76,
    n66
  );


  nand
  g206
  (
    n270,
    n79,
    n72,
    n203,
    n73
  );


  xnor
  g207
  (
    n242,
    n94,
    n207,
    n92,
    n83
  );


  xor
  g208
  (
    n224,
    n55,
    n204,
    n217,
    n69
  );


  or
  g209
  (
    n232,
    n78,
    n77,
    n81,
    n202
  );


  or
  g210
  (
    n282,
    n86,
    n75,
    n98,
    n208
  );


  nor
  g211
  (
    n251,
    n214,
    n82,
    n93,
    n209
  );


  nor
  g212
  (
    n220,
    n67,
    n68,
    n62,
    n51
  );


  and
  g213
  (
    n264,
    n216,
    n201,
    n79,
    n209
  );


  nand
  g214
  (
    n284,
    n104,
    n200,
    n215,
    n217
  );


  xnor
  g215
  (
    n257,
    n82,
    n213,
    n210,
    n88
  );


  or
  g216
  (
    n236,
    n103,
    n98,
    n96,
    n93
  );


  and
  g217
  (
    n238,
    n75,
    n101,
    n67,
    n91
  );


  xor
  g218
  (
    n235,
    n202,
    n210,
    n74,
    n87
  );


  nor
  g219
  (
    n267,
    n83,
    n78,
    n97,
    n213
  );


  or
  g220
  (
    n258,
    n69,
    n80,
    n201
  );


  xor
  g221
  (
    n249,
    n64,
    n63,
    n203,
    n96
  );


  or
  g222
  (
    n274,
    n204,
    n88,
    n58,
    n53
  );


  xnor
  g223
  (
    n239,
    n70,
    n89,
    n74,
    n214
  );


  xnor
  g224
  (
    n287,
    n68,
    n78,
    n76,
    n63
  );


  xnor
  g225
  (
    n229,
    n54,
    n80,
    n86,
    n98
  );


  xor
  g226
  (
    n283,
    n90,
    n60,
    n61,
    n89
  );


  xnor
  g227
  (
    n243,
    n94,
    n68,
    n203,
    n62
  );


  xnor
  g228
  (
    n290,
    n67,
    n79,
    n66,
    n50
  );


  nor
  g229
  (
    n288,
    n104,
    n99,
    n66,
    n65
  );


  xor
  g230
  (
    n278,
    n202,
    n96,
    n94,
    n92
  );


  xor
  g231
  (
    n277,
    n61,
    n99,
    n215,
    n85
  );


  and
  g232
  (
    n241,
    n211,
    n69,
    n52,
    n206
  );


  nand
  g233
  (
    n265,
    n84,
    n88,
    n207,
    n59
  );


  xnor
  g234
  (
    n226,
    n56,
    n210,
    n87,
    n205
  );


  xnor
  g235
  (
    n228,
    n53,
    n51,
    n90,
    n101
  );


  nand
  g236
  (
    n254,
    n65,
    n68,
    n89,
    n64
  );


  xnor
  g237
  (
    n262,
    n61,
    n103,
    n207,
    n209
  );


  and
  g238
  (
    n247,
    n76,
    n66,
    n205,
    n57
  );


  or
  g239
  (
    n248,
    n73,
    n95,
    n212,
    n91
  );


  xor
  g240
  (
    n269,
    n51,
    n78,
    n211,
    n81
  );


  xor
  g241
  (
    n281,
    n74,
    n64,
    n103,
    n216
  );


  xor
  g242
  (
    n280,
    n67,
    n201,
    n92,
    n64
  );


  nand
  g243
  (
    n289,
    n202,
    n81,
    n74,
    n102
  );


  xor
  g244
  (
    n273,
    n57,
    n97,
    n211,
    n76
  );


  nor
  g245
  (
    n246,
    n52,
    n53,
    n70,
    n96
  );


  nor
  g246
  (
    n255,
    n61,
    n50,
    n84,
    n72
  );


  or
  g247
  (
    n266,
    n72,
    n82,
    n204,
    n213
  );


  or
  g248
  (
    n252,
    n101,
    n98,
    n65,
    n73
  );


  or
  g249
  (
    n237,
    n56,
    n206,
    n60,
    n217
  );


  xor
  g250
  (
    n259,
    n57,
    n56,
    n100,
    n212
  );


  xnor
  g251
  (
    n233,
    n85,
    n99,
    n62,
    n92
  );


  xor
  g252
  (
    n272,
    n63,
    n57,
    n207,
    n60
  );


  nand
  g253
  (
    n260,
    n100,
    n90,
    n84,
    n75
  );


  xor
  g254
  (
    n268,
    n95,
    n58,
    n208,
    n83
  );


  nand
  g255
  (
    n231,
    n73,
    n200,
    n212,
    n87
  );


  and
  g256
  (
    n276,
    n72,
    n59,
    n95,
    n80
  );


  xor
  g257
  (
    n275,
    n94,
    n203,
    n56,
    n88
  );


  xor
  g258
  (
    n292,
    n216,
    n208,
    n95,
    n60
  );


  or
  g259
  (
    n253,
    n75,
    n90,
    n86,
    n217
  );


  nor
  g260
  (
    n223,
    n54,
    n93,
    n59,
    n214
  );


  nand
  g261
  (
    n261,
    n79,
    n85,
    n51,
    n208
  );


  xor
  g262
  (
    n250,
    n215,
    n210,
    n81,
    n205
  );


  nand
  g263
  (
    n222,
    n89,
    n54,
    n103,
    n85
  );


  nor
  g264
  (
    n221,
    n71,
    n59,
    n204,
    n215
  );


  xnor
  g265
  (
    n245,
    n65,
    n201,
    n104,
    n214
  );


  xor
  g266
  (
    n330,
    n251,
    n226,
    n230,
    n236
  );


  nand
  g267
  (
    n307,
    n257,
    n259,
    n220,
    n264
  );


  nand
  g268
  (
    n318,
    n231,
    n263,
    n250,
    n239
  );


  xnor
  g269
  (
    n333,
    n246,
    n244,
    n226,
    n222
  );


  or
  g270
  (
    n301,
    n234,
    n244,
    n252,
    n245
  );


  nand
  g271
  (
    KeyWire_0_30,
    n269,
    n105,
    n224,
    n222
  );


  nor
  g272
  (
    n310,
    n223,
    n248,
    n259,
    n241
  );


  xnor
  g273
  (
    n335,
    n268,
    n245,
    n238,
    n264
  );


  nand
  g274
  (
    n327,
    n225,
    n233,
    n226,
    n238
  );


  nand
  g275
  (
    n293,
    n259,
    n256,
    n248,
    n224
  );


  or
  g276
  (
    n300,
    n246,
    n268,
    n238,
    n260
  );


  xor
  g277
  (
    n297,
    n242,
    n265,
    n222,
    n251
  );


  xnor
  g278
  (
    n305,
    n243,
    n236,
    n231,
    n230
  );


  nand
  g279
  (
    n324,
    n240,
    n220,
    n225,
    n247
  );


  nor
  g280
  (
    n337,
    n255,
    n232,
    n267,
    n230
  );


  nor
  g281
  (
    n334,
    n251,
    n247,
    n268,
    n242
  );


  and
  g282
  (
    n323,
    n248,
    n266,
    n240,
    n227
  );


  nand
  g283
  (
    n299,
    n239,
    n241,
    n252,
    n221
  );


  xor
  g284
  (
    n304,
    n253,
    n223,
    n249,
    n235
  );


  and
  g285
  (
    n338,
    n223,
    n261,
    n254,
    n266
  );


  xnor
  g286
  (
    n314,
    n243,
    n237,
    n228,
    n220
  );


  or
  g287
  (
    n325,
    n256,
    n233,
    n232,
    n227
  );


  xor
  g288
  (
    n328,
    n224,
    n229,
    n256,
    n263
  );


  nor
  g289
  (
    n326,
    n249,
    n225,
    n228,
    n241
  );


  nand
  g290
  (
    n336,
    n224,
    n257,
    n235,
    n265
  );


  nor
  g291
  (
    n306,
    n254,
    n267,
    n232
  );


  nand
  g292
  (
    n298,
    n246,
    n260,
    n242,
    n254
  );


  or
  g293
  (
    n295,
    n234,
    n254,
    n255,
    n253
  );


  xor
  g294
  (
    n340,
    n229,
    n256,
    n245,
    n240
  );


  or
  g295
  (
    n315,
    n264,
    n243,
    n250,
    n237
  );


  or
  g296
  (
    n339,
    n262,
    n234,
    n221,
    n259
  );


  or
  g297
  (
    n320,
    n261,
    n236,
    n239,
    n244
  );


  xnor
  g298
  (
    n341,
    n255,
    n262,
    n269,
    n223
  );


  and
  g299
  (
    n322,
    n220,
    n238,
    n263,
    n239
  );


  nand
  g300
  (
    n311,
    n262,
    n265,
    n250,
    n235
  );


  or
  g301
  (
    n329,
    n225,
    n249,
    n231,
    n262
  );


  xnor
  g302
  (
    n342,
    n253,
    n248,
    n257,
    n236
  );


  nand
  g303
  (
    n321,
    n226,
    n227,
    n229,
    n255
  );


  nor
  g304
  (
    n313,
    n233,
    n221,
    n261,
    n266
  );


  nand
  g305
  (
    n302,
    n234,
    n258,
    n260
  );


  and
  g306
  (
    n331,
    n249,
    n229,
    n222,
    n252
  );


  nor
  g307
  (
    n319,
    n258,
    n241,
    n232,
    n231
  );


  nand
  g308
  (
    n309,
    n235,
    n258,
    n265
  );


  or
  g309
  (
    n303,
    n267,
    n266,
    n221,
    n263
  );


  xor
  g310
  (
    n296,
    n230,
    n227,
    n233,
    n244
  );


  xor
  g311
  (
    n294,
    n237,
    n245,
    n246,
    n243
  );


  xor
  g312
  (
    n312,
    n264,
    n247,
    n242,
    n105
  );


  nand
  g313
  (
    n316,
    n228,
    n251,
    n261,
    n250
  );


  and
  g314
  (
    n317,
    n237,
    n257,
    n252,
    n228
  );


  xnor
  g315
  (
    n308,
    n268,
    n240,
    n253,
    n247
  );


  xor
  g316
  (
    n362,
    n306,
    n307,
    n145
  );


  and
  g317
  (
    n356,
    n148,
    n153,
    n304,
    n108
  );


  and
  g318
  (
    n349,
    n307,
    n106,
    n302,
    n107
  );


  nand
  g319
  (
    n360,
    n146,
    n146,
    n300,
    n105
  );


  or
  g320
  (
    n348,
    n152,
    n305,
    n301,
    n151
  );


  xnor
  g321
  (
    n363,
    n271,
    n294,
    n272,
    n106
  );


  nor
  g322
  (
    n343,
    n271,
    n303,
    n153,
    n270
  );


  or
  g323
  (
    n353,
    n272,
    n300,
    n271,
    n270
  );


  or
  g324
  (
    n345,
    n106,
    n303,
    n302,
    n151
  );


  nor
  g325
  (
    n354,
    n148,
    n149,
    n107,
    n106
  );


  nor
  g326
  (
    n357,
    n108,
    n270,
    n301,
    n150
  );


  nor
  g327
  (
    n361,
    n154,
    n155,
    n150,
    n298
  );


  and
  g328
  (
    n347,
    n155,
    n299,
    n308,
    n272
  );


  nor
  g329
  (
    n351,
    n297,
    n147,
    n151,
    n269
  );


  xnor
  g330
  (
    n346,
    n147,
    n146,
    n108,
    n152
  );


  xnor
  g331
  (
    n355,
    n296,
    n155,
    n152,
    n145
  );


  nand
  g332
  (
    n344,
    n149,
    n153,
    n270,
    n154
  );


  xor
  g333
  (
    n359,
    n306,
    n107,
    n218,
    n108
  );


  xnor
  g334
  (
    n364,
    n299,
    n305,
    n154,
    n269
  );


  and
  g335
  (
    n352,
    n271,
    n149,
    n144,
    n150
  );


  xor
  g336
  (
    n358,
    n145,
    n272,
    n147,
    n293
  );


  or
  g337
  (
    n350,
    n148,
    n107,
    n295,
    n304
  );


  not
  g338
  (
    n374,
    n360
  );


  not
  g339
  (
    n370,
    n361
  );


  buf
  g340
  (
    n375,
    n351
  );


  not
  g341
  (
    n371,
    n345
  );


  not
  g342
  (
    n373,
    n349
  );


  buf
  g343
  (
    n376,
    n348
  );


  not
  g344
  (
    n372,
    n357
  );


  buf
  g345
  (
    n366,
    n364
  );


  not
  g346
  (
    n368,
    n354
  );


  not
  g347
  (
    n382,
    n353
  );


  buf
  g348
  (
    n369,
    n363
  );


  buf
  g349
  (
    n381,
    n355
  );


  buf
  g350
  (
    n379,
    n346
  );


  buf
  g351
  (
    n378,
    n358
  );


  not
  g352
  (
    n367,
    n356
  );


  buf
  g353
  (
    n384,
    n347
  );


  buf
  g354
  (
    n377,
    n362
  );


  buf
  g355
  (
    n383,
    n350
  );


  not
  g356
  (
    n380,
    n359
  );


  not
  g357
  (
    n365,
    n352
  );


  buf
  g358
  (
    n388,
    n365
  );


  buf
  g359
  (
    n387,
    n365
  );


  not
  g360
  (
    n386,
    n366
  );


  buf
  g361
  (
    n385,
    n366
  );


  buf
  g362
  (
    n395,
    n219
  );


  not
  g363
  (
    n392,
    n385
  );


  buf
  g364
  (
    n394,
    n385
  );


  buf
  g365
  (
    n396,
    n387
  );


  not
  g366
  (
    n401,
    n387
  );


  not
  g367
  (
    n391,
    n387
  );


  buf
  g368
  (
    n399,
    n388
  );


  not
  g369
  (
    n389,
    n385
  );


  not
  g370
  (
    n400,
    n218
  );


  buf
  g371
  (
    n390,
    n387
  );


  buf
  g372
  (
    n398,
    n386
  );


  not
  g373
  (
    n393,
    n386
  );


  buf
  g374
  (
    n403,
    n386
  );


  not
  g375
  (
    n397,
    n388
  );


  and
  g376
  (
    n402,
    n385,
    n386,
    n218,
    n388
  );


  not
  g377
  (
    n407,
    n389
  );


  buf
  g378
  (
    n404,
    n389
  );


  buf
  g379
  (
    n405,
    n389
  );


  not
  g380
  (
    n406,
    n389
  );


  buf
  g381
  (
    n411,
    n406
  );


  buf
  g382
  (
    n415,
    n407
  );


  not
  g383
  (
    n418,
    n405
  );


  buf
  g384
  (
    n419,
    n404
  );


  buf
  g385
  (
    n410,
    n406
  );


  not
  g386
  (
    n409,
    n406
  );


  buf
  g387
  (
    n412,
    n405
  );


  buf
  g388
  (
    n421,
    n404
  );


  buf
  g389
  (
    n420,
    n405
  );


  not
  g390
  (
    n408,
    n404
  );


  not
  g391
  (
    n422,
    n406
  );


  buf
  g392
  (
    n416,
    n405
  );


  buf
  g393
  (
    n413,
    n407
  );


  buf
  g394
  (
    n417,
    n407
  );


  buf
  g395
  (
    n414,
    n407
  );


  not
  g396
  (
    n423,
    n417
  );


  not
  g397
  (
    n434,
    n109
  );


  buf
  g398
  (
    n424,
    n111
  );


  buf
  g399
  (
    n429,
    n414
  );


  not
  g400
  (
    n430,
    n415
  );


  not
  g401
  (
    n425,
    n111
  );


  buf
  g402
  (
    n431,
    n413
  );


  not
  g403
  (
    n428,
    n110
  );


  nor
  g404
  (
    n427,
    n411,
    n109,
    n110
  );


  nand
  g405
  (
    n433,
    n408,
    n409,
    n111
  );


  xnor
  g406
  (
    n426,
    n110,
    n416,
    n410
  );


  nand
  g407
  (
    n432,
    n412,
    n110,
    n109,
    n417
  );


  not
  g408
  (
    n444,
    n429
  );


  not
  g409
  (
    n440,
    n424
  );


  buf
  g410
  (
    n443,
    n423
  );


  buf
  g411
  (
    n439,
    n426
  );


  not
  g412
  (
    n435,
    n427
  );


  buf
  g413
  (
    n447,
    n424
  );


  not
  g414
  (
    n436,
    n423
  );


  buf
  g415
  (
    n438,
    n425
  );


  buf
  g416
  (
    n437,
    n425
  );


  not
  g417
  (
    n445,
    n428
  );


  not
  g418
  (
    n442,
    n428
  );


  not
  g419
  (
    n446,
    n427
  );


  not
  g420
  (
    n441,
    n426
  );


  or
  g421
  (
    n450,
    n435,
    n438
  );


  xnor
  g422
  (
    n453,
    n437,
    n435,
    n440
  );


  and
  g423
  (
    n451,
    n439,
    n438,
    n436,
    n437
  );


  nor
  g424
  (
    n449,
    n436,
    n438,
    n440,
    n439
  );


  xor
  g425
  (
    n452,
    n439,
    n438,
    n437,
    n436
  );


  or
  g426
  (
    n454,
    n436,
    n440,
    n439
  );


  or
  g427
  (
    n448,
    n435,
    n112,
    n437
  );


  buf
  g428
  (
    n467,
    n400
  );


  not
  g429
  (
    n478,
    n454
  );


  buf
  g430
  (
    n458,
    n451
  );


  buf
  g431
  (
    n463,
    n395
  );


  not
  g432
  (
    n476,
    n399
  );


  buf
  g433
  (
    n471,
    n397
  );


  buf
  g434
  (
    n475,
    n391
  );


  buf
  g435
  (
    n457,
    n401
  );


  buf
  g436
  (
    n470,
    n398
  );


  and
  g437
  (
    n477,
    n390,
    n391,
    n399
  );


  nor
  g438
  (
    n474,
    n450,
    n399,
    n394,
    n390
  );


  and
  g439
  (
    n466,
    n398,
    n451,
    n394,
    n397
  );


  xor
  g440
  (
    n455,
    n26,
    n392,
    n454
  );


  xnor
  g441
  (
    n460,
    n392,
    n451,
    n391,
    n394
  );


  nand
  g442
  (
    n469,
    n453,
    n396,
    n449,
    n393
  );


  xor
  g443
  (
    n461,
    n26,
    n450,
    n400,
    n396
  );


  xnor
  g444
  (
    n464,
    n395,
    n392,
    n450,
    n452
  );


  or
  g445
  (
    KeyWire_0_2,
    n395,
    n398,
    n401
  );


  or
  g446
  (
    n480,
    n449,
    n393,
    n396
  );


  and
  g447
  (
    KeyWire_0_4,
    n397,
    n402,
    n25,
    n454
  );


  nand
  g448
  (
    n456,
    n401,
    n396,
    n392,
    n448
  );


  or
  g449
  (
    n465,
    n26,
    n449,
    n393,
    n450
  );


  nand
  g450
  (
    n473,
    n452,
    n395,
    n399,
    n390
  );


  nor
  g451
  (
    KeyWire_0_3,
    n453,
    n391,
    n452,
    n397
  );


  and
  g452
  (
    n472,
    n453,
    n448,
    n451,
    n449
  );


  and
  g453
  (
    n481,
    n452,
    n394,
    n400,
    n390
  );


  nand
  g454
  (
    n459,
    n398,
    n453,
    n400,
    n448
  );


  not
  g455
  (
    n497,
    n460
  );


  not
  g456
  (
    n484,
    n456
  );


  buf
  g457
  (
    n496,
    n457
  );


  buf
  g458
  (
    n498,
    n455
  );


  not
  g459
  (
    n489,
    n458
  );


  buf
  g460
  (
    n492,
    n159
  );


  not
  g461
  (
    n495,
    n157
  );


  buf
  g462
  (
    n494,
    n458
  );


  buf
  g463
  (
    n493,
    n456
  );


  not
  g464
  (
    n491,
    n160
  );


  xnor
  g465
  (
    n485,
    n459,
    n158,
    n31,
    n458
  );


  nor
  g466
  (
    n482,
    n157,
    n457,
    n160
  );


  nand
  g467
  (
    n488,
    n157,
    n459,
    n160,
    n159
  );


  nor
  g468
  (
    n487,
    n158,
    n460,
    n31,
    n156
  );


  xor
  g469
  (
    n483,
    n158,
    n159,
    n456,
    n455
  );


  nand
  g470
  (
    n499,
    n459,
    n156,
    n457,
    n458
  );


  nand
  g471
  (
    n486,
    n456,
    n112,
    n459,
    n26
  );


  nand
  g472
  (
    n490,
    n460,
    n156,
    n455
  );


  or
  g473
  (
    n505,
    n487,
    n49,
    n186,
    n491
  );


  xor
  g474
  (
    n515,
    n488,
    n49,
    n420,
    n182
  );


  nand
  g475
  (
    n509,
    n482,
    n493,
    n184,
    n491
  );


  nor
  g476
  (
    n500,
    n493,
    n487,
    n195,
    n193
  );


  and
  g477
  (
    n516,
    n194,
    n493,
    n492,
    n486
  );


  xnor
  g478
  (
    n504,
    n487,
    n196,
    n492,
    n418
  );


  or
  g479
  (
    n508,
    n492,
    n483,
    n421,
    n489
  );


  or
  g480
  (
    n517,
    n191,
    n484,
    n492
  );


  xnor
  g481
  (
    n514,
    n419,
    n199,
    n490,
    n482
  );


  and
  g482
  (
    n501,
    n490,
    n484,
    n420,
    n485
  );


  nand
  g483
  (
    n506,
    n486,
    n489,
    n418
  );


  xor
  g484
  (
    n502,
    n491,
    n483,
    n484
  );


  xnor
  g485
  (
    n510,
    n198,
    n489,
    n488,
    n421
  );


  xor
  g486
  (
    n507,
    n483,
    n485,
    n490,
    n482
  );


  nor
  g487
  (
    n511,
    n486,
    n183,
    n422
  );


  nand
  g488
  (
    n512,
    n419,
    n490,
    n486,
    n487
  );


  xor
  g489
  (
    n513,
    n185,
    n49,
    n187,
    n482
  );


  nand
  g490
  (
    n503,
    n493,
    n188,
    n491,
    n189
  );


  nand
  g491
  (
    n518,
    n181,
    n488,
    n485,
    n190
  );


  and
  g492
  (
    n519,
    n488,
    n197,
    n192,
    n485
  );


  not
  g493
  (
    n520,
    n501
  );


  buf
  g494
  (
    n522,
    n500
  );


  buf
  g495
  (
    n523,
    n500
  );


  buf
  g496
  (
    n524,
    n502
  );


  not
  g497
  (
    n521,
    n501
  );


  nand
  g498
  (
    n529,
    n273,
    n521,
    n275,
    n276
  );


  xor
  g499
  (
    n540,
    n114,
    n114,
    n273,
    n278
  );


  nand
  g500
  (
    n528,
    n279,
    n113,
    n116,
    n115
  );


  xnor
  g501
  (
    n525,
    n278,
    n117,
    n522
  );


  and
  g502
  (
    n526,
    n276,
    n279,
    n523,
    n278
  );


  xor
  g503
  (
    n533,
    n524,
    n279,
    n277,
    n280
  );


  or
  g504
  (
    n527,
    n523,
    n275,
    n118,
    n274
  );


  xor
  g505
  (
    n535,
    n276,
    n114,
    n116,
    n273
  );


  or
  g506
  (
    n538,
    n277,
    n112,
    n115,
    n278
  );


  or
  g507
  (
    n539,
    n277,
    n113,
    n523,
    n520
  );


  and
  g508
  (
    n536,
    n117,
    n273,
    n523,
    n520
  );


  xnor
  g509
  (
    n534,
    n275,
    n277,
    n116,
    n274
  );


  and
  g510
  (
    n537,
    n274,
    n118,
    n280,
    n115
  );


  xnor
  g511
  (
    n541,
    n521,
    n522,
    n274,
    n524
  );


  or
  g512
  (
    n542,
    n275,
    n116,
    n522,
    n117
  );


  nand
  g513
  (
    n531,
    n279,
    n118,
    n113,
    n521
  );


  xnor
  g514
  (
    n530,
    n113,
    n520,
    n522
  );


  or
  g515
  (
    n532,
    n521,
    n114,
    n115,
    n276
  );


  not
  g516
  (
    n574,
    n541
  );


  not
  g517
  (
    n577,
    n320
  );


  not
  g518
  (
    KeyWire_0_10,
    n319
  );


  buf
  g519
  (
    n567,
    n335
  );


  not
  g520
  (
    n569,
    n339
  );


  not
  g521
  (
    n571,
    n538
  );


  not
  g522
  (
    n557,
    n526
  );


  not
  g523
  (
    n547,
    n321
  );


  buf
  g524
  (
    n545,
    n528
  );


  buf
  g525
  (
    n563,
    n542
  );


  buf
  g526
  (
    n553,
    n337
  );


  buf
  g527
  (
    n562,
    n330
  );


  not
  g528
  (
    n565,
    n534
  );


  nor
  g529
  (
    n548,
    n539,
    n532,
    n318
  );


  or
  g530
  (
    n549,
    n336,
    n527,
    n316,
    n533
  );


  xnor
  g531
  (
    n568,
    n327,
    n525,
    n535,
    n542
  );


  xor
  g532
  (
    n572,
    n526,
    n535,
    n323,
    n540
  );


  or
  g533
  (
    n551,
    n528,
    n328,
    n333,
    n325
  );


  and
  g534
  (
    n564,
    n311,
    n317,
    n324,
    n332
  );


  and
  g535
  (
    n575,
    n525,
    n539,
    n531,
    n322
  );


  and
  g536
  (
    n556,
    n334,
    n331,
    n324,
    n310
  );


  nor
  g537
  (
    n558,
    n309,
    n311,
    n334,
    n313
  );


  and
  g538
  (
    n576,
    n339,
    n529,
    n541,
    n320
  );


  nand
  g539
  (
    n554,
    n317,
    n325,
    n527,
    n536
  );


  xnor
  g540
  (
    n543,
    n321,
    n315,
    n537,
    n314
  );


  xnor
  g541
  (
    n561,
    n331,
    n327,
    n330,
    n341
  );


  nand
  g542
  (
    n573,
    n333,
    n341,
    n338,
    n540
  );


  xnor
  g543
  (
    n555,
    n531,
    n310,
    n316,
    n342
  );


  xnor
  g544
  (
    n560,
    n337,
    n322,
    n309,
    n340
  );


  xnor
  g545
  (
    n544,
    n319,
    n335,
    n312,
    n313
  );


  or
  g546
  (
    n578,
    n533,
    n318,
    n537,
    n529
  );


  xor
  g547
  (
    n566,
    n329,
    n340,
    n534,
    n326
  );


  and
  g548
  (
    n559,
    n336,
    n314,
    n312,
    n329
  );


  or
  g549
  (
    n570,
    n338,
    n328,
    n536,
    n538
  );


  nor
  g550
  (
    n550,
    n530,
    n315,
    n532,
    n323
  );


  xor
  g551
  (
    n546,
    n308,
    n530,
    n326,
    n332
  );


  buf
  g552
  (
    n579,
    n543
  );


  buf
  g553
  (
    n580,
    n543
  );


  buf
  g554
  (
    n585,
    n495
  );


  buf
  g555
  (
    n581,
    n367
  );


  buf
  g556
  (
    n584,
    n494
  );


  buf
  g557
  (
    n588,
    n494
  );


  and
  g558
  (
    n586,
    n494,
    n580
  );


  or
  g559
  (
    n587,
    n580,
    n579
  );


  or
  g560
  (
    n582,
    n494,
    n579
  );


  or
  g561
  (
    n583,
    n367,
    n580,
    n495
  );


  buf
  g562
  (
    n589,
    n588
  );


  not
  g563
  (
    n590,
    n586
  );


  not
  g564
  (
    n591,
    n587
  );


  xor
  g565
  (
    n595,
    n590,
    n284,
    n286,
    n282
  );


  or
  g566
  (
    KeyWire_0_31,
    n280,
    n219,
    n282,
    n590
  );


  nor
  g567
  (
    n593,
    n282,
    n281,
    n285,
    n284
  );


  xnor
  g568
  (
    n601,
    n286,
    n284,
    n589,
    n283
  );


  nor
  g569
  (
    n600,
    n280,
    n589,
    n283,
    n281
  );


  or
  g570
  (
    n592,
    n590,
    n285
  );


  nand
  g571
  (
    n599,
    n591,
    n284,
    n281,
    n285
  );


  nor
  g572
  (
    n598,
    n283,
    n589,
    n219
  );


  nor
  g573
  (
    n597,
    n219,
    n283,
    n286
  );


  nand
  g574
  (
    n596,
    n287,
    n591,
    n282,
    n281
  );


  or
  g575
  (
    KeyWire_0_12,
    n289,
    n288
  );


  xor
  g576
  (
    n609,
    n593,
    n544
  );


  xnor
  g577
  (
    n611,
    n593,
    n287
  );


  xor
  g578
  (
    n608,
    n592,
    n287
  );


  and
  g579
  (
    n605,
    n289,
    n288
  );


  xor
  g580
  (
    n606,
    n592,
    n290,
    n288,
    n594
  );


  nor
  g581
  (
    n604,
    n290,
    n289,
    n592
  );


  and
  g582
  (
    n602,
    n290,
    n291,
    n288,
    n593
  );


  xnor
  g583
  (
    n607,
    n287,
    n291,
    n594,
    n544
  );


  nand
  g584
  (
    n610,
    n544,
    n544,
    n594,
    n543
  );


  or
  g585
  (
    n612,
    n543,
    n290,
    n289,
    n593
  );


  or
  g586
  (
    n615,
    n550,
    n548
  );


  nor
  g587
  (
    n614,
    n550,
    n603
  );


  xnor
  g588
  (
    n617,
    n546,
    n604
  );


  xor
  g589
  (
    n616,
    n605,
    n602,
    n551,
    n549
  );


  or
  g590
  (
    n621,
    n603,
    n547,
    n549,
    n552
  );


  nor
  g591
  (
    n619,
    n549,
    n548,
    n602
  );


  nand
  g592
  (
    n620,
    n551,
    n545,
    n603
  );


  or
  g593
  (
    n622,
    n545,
    n604,
    n602,
    n550
  );


  and
  g594
  (
    n613,
    n547,
    n602,
    n551,
    n550
  );


  nand
  g595
  (
    n618,
    n548,
    n546,
    n549
  );


  xnor
  g596
  (
    n623,
    n604,
    n603,
    n547,
    n545
  );


  xor
  g597
  (
    n624,
    n547,
    n546,
    n604,
    n551
  );


  xor
  g598
  (
    n636,
    n614,
    n373,
    n374,
    n381
  );


  or
  g599
  (
    n646,
    n554,
    n432,
    n614,
    n622
  );


  and
  g600
  (
    n653,
    n381,
    n552,
    n371,
    n621
  );


  nor
  g601
  (
    n651,
    n554,
    n432,
    n370,
    n623
  );


  nand
  g602
  (
    n631,
    n429,
    n433,
    n618,
    n623
  );


  xor
  g603
  (
    n628,
    n613,
    n431,
    n372,
    n623
  );


  xnor
  g604
  (
    n643,
    n429,
    n372,
    n624,
    n616
  );


  xor
  g605
  (
    n642,
    n617,
    n616,
    n430,
    n369
  );


  xnor
  g606
  (
    n625,
    n615,
    n382,
    n379,
    n613
  );


  and
  g607
  (
    n627,
    n368,
    n380,
    n379,
    n552
  );


  or
  g608
  (
    n648,
    n614,
    n618,
    n613,
    n620
  );


  nor
  g609
  (
    n640,
    n434,
    n615,
    n379,
    n621
  );


  xnor
  g610
  (
    n649,
    n374,
    n618,
    n619,
    n552
  );


  and
  g611
  (
    n629,
    n373,
    n619,
    n620,
    n432
  );


  nor
  g612
  (
    n630,
    n376,
    n382,
    n378,
    n380
  );


  nor
  g613
  (
    n635,
    n431,
    n623,
    n553,
    n430
  );


  xor
  g614
  (
    KeyWire_0_22,
    n613,
    n375,
    n624
  );


  and
  g615
  (
    n626,
    n555,
    n622,
    n383,
    n378
  );


  and
  g616
  (
    n652,
    n377,
    n618,
    n378,
    n615
  );


  nor
  g617
  (
    n637,
    n381,
    n615,
    n605,
    n554
  );


  nand
  g618
  (
    n647,
    n553,
    n382,
    n621,
    n380
  );


  xnor
  g619
  (
    n650,
    n619,
    n616,
    n553,
    n370
  );


  and
  g620
  (
    n632,
    n617,
    n554,
    n624,
    n377
  );


  xor
  g621
  (
    n638,
    n375,
    n433,
    n368,
    n431
  );


  xnor
  g622
  (
    n634,
    n614,
    n434,
    n430,
    n377
  );


  and
  g623
  (
    n645,
    n616,
    n376,
    n434,
    n382
  );


  xnor
  g624
  (
    n639,
    n620,
    n622,
    n371,
    n621
  );


  and
  g625
  (
    n633,
    n622,
    n369,
    n553,
    n433
  );


  xnor
  g626
  (
    n641,
    n619,
    n620,
    n617
  );


  nand
  g627
  (
    n660,
    n443,
    n445,
    n626,
    n627
  );


  nand
  g628
  (
    n661,
    n447,
    n442,
    n445
  );


  nand
  g629
  (
    n654,
    n447,
    n441,
    n626
  );


  nand
  g630
  (
    n659,
    n625,
    n444,
    n446
  );


  xor
  g631
  (
    n655,
    n447,
    n444,
    n442,
    n441
  );


  nand
  g632
  (
    n662,
    n441,
    n446,
    n443,
    n625
  );


  and
  g633
  (
    n658,
    n446,
    n443,
    n444,
    n626
  );


  nand
  g634
  (
    n657,
    n442,
    n626,
    n445,
    n625
  );


  or
  g635
  (
    n656,
    n443,
    n625,
    n446,
    n445
  );


  xor
  g636
  (
    n668,
    n655,
    n606,
    n607
  );


  and
  g637
  (
    n667,
    n591,
    n661,
    n555
  );


  nand
  g638
  (
    n666,
    n658,
    n403,
    n591
  );


  xnor
  g639
  (
    n670,
    n388,
    n657,
    n595,
    n660
  );


  or
  g640
  (
    n665,
    n606,
    n403,
    n402
  );


  nand
  g641
  (
    n672,
    n656,
    n605,
    n662,
    n556
  );


  xnor
  g642
  (
    n664,
    n556,
    n607,
    n595,
    n402
  );


  xnor
  g643
  (
    n673,
    n606,
    n662,
    n555,
    n596
  );


  and
  g644
  (
    n663,
    n654,
    n605,
    n596,
    n607
  );


  and
  g645
  (
    n671,
    n403,
    n555,
    n659,
    n606
  );


  xor
  g646
  (
    n669,
    n661,
    n594,
    n595
  );


  buf
  g647
  (
    n681,
    n609
  );


  not
  g648
  (
    n677,
    n663
  );


  or
  g649
  (
    n676,
    n665,
    n664
  );


  nor
  g650
  (
    n678,
    n609,
    n667,
    n608,
    n610
  );


  nand
  g651
  (
    n680,
    n610,
    n607,
    n608,
    n596
  );


  or
  g652
  (
    n679,
    n610,
    n665,
    n666,
    n596
  );


  nor
  g653
  (
    n675,
    n608,
    n597,
    n609
  );


  nand
  g654
  (
    n674,
    n608,
    n609,
    n664,
    n666
  );


  not
  g655
  (
    n684,
    n674
  );


  buf
  g656
  (
    n683,
    n674
  );


  not
  g657
  (
    n689,
    n675
  );


  buf
  g658
  (
    n686,
    n674
  );


  not
  g659
  (
    n682,
    n675
  );


  buf
  g660
  (
    n687,
    n610
  );


  buf
  g661
  (
    n688,
    n675
  );


  xor
  g662
  (
    n685,
    n675,
    n674
  );


  not
  g663
  (
    n695,
    n682
  );


  buf
  g664
  (
    n692,
    n683
  );


  not
  g665
  (
    n691,
    n682
  );


  buf
  g666
  (
    n690,
    n683
  );


  not
  g667
  (
    n693,
    n682
  );


  not
  g668
  (
    n696,
    n683
  );


  not
  g669
  (
    n694,
    n682
  );


  xnor
  g670
  (
    n715,
    n647,
    n629,
    n636,
    n696
  );


  xor
  g671
  (
    n700,
    n646,
    n645,
    n629,
    n691
  );


  xnor
  g672
  (
    n710,
    n694,
    n630,
    n631,
    n641
  );


  xor
  g673
  (
    KeyWire_0_29,
    n628,
    n647,
    n696,
    n644
  );


  and
  g674
  (
    n711,
    n638,
    n630,
    n632,
    n635
  );


  and
  g675
  (
    n719,
    n634,
    n646,
    n644,
    n638
  );


  and
  g676
  (
    n712,
    n643,
    n632,
    n638
  );


  xor
  g677
  (
    n704,
    n695,
    n642,
    n647
  );


  nand
  g678
  (
    n697,
    n635,
    n636,
    n695
  );


  xnor
  g679
  (
    n717,
    n695,
    n640,
    n690
  );


  xnor
  g680
  (
    n718,
    n636,
    n694,
    n691,
    n648
  );


  nand
  g681
  (
    n699,
    n637,
    n646,
    n690,
    n694
  );


  nor
  g682
  (
    n707,
    n640,
    n630,
    n639,
    n634
  );


  xor
  g683
  (
    n702,
    n631,
    n693,
    n646,
    n642
  );


  nand
  g684
  (
    n714,
    n692,
    n627,
    n637,
    n644
  );


  nand
  g685
  (
    n705,
    n645,
    n693,
    n641,
    n635
  );


  xnor
  g686
  (
    n723,
    n643,
    n631,
    n639
  );


  nor
  g687
  (
    n722,
    n633,
    n692,
    n628,
    n637
  );


  and
  g688
  (
    n709,
    n690,
    n645,
    n693,
    n637
  );


  xor
  g689
  (
    KeyWire_0_14,
    n694,
    n644,
    n691
  );


  nor
  g690
  (
    n721,
    n633,
    n640,
    n690,
    n692
  );


  nand
  g691
  (
    n713,
    n693,
    n629,
    n635,
    n641
  );


  and
  g692
  (
    n701,
    n629,
    n628,
    n627,
    n639
  );


  nor
  g693
  (
    n724,
    n643,
    n642,
    n628,
    n634
  );


  nand
  g694
  (
    n703,
    n692,
    n634,
    n696,
    n627
  );


  nor
  g695
  (
    n706,
    n696,
    n643,
    n645,
    n630
  );


  nand
  g696
  (
    n720,
    n641,
    n642,
    n695,
    n632
  );


  nand
  g697
  (
    n698,
    n638,
    n639,
    n633
  );


  not
  g698
  (
    n749,
    n718
  );


  not
  g699
  (
    n779,
    n716
  );


  not
  g700
  (
    n769,
    n711
  );


  buf
  g701
  (
    n807,
    n706
  );


  not
  g702
  (
    n735,
    n697
  );


  buf
  g703
  (
    n815,
    n713
  );


  not
  g704
  (
    n745,
    n705
  );


  buf
  g705
  (
    n795,
    n704
  );


  buf
  g706
  (
    n777,
    n712
  );


  not
  g707
  (
    n763,
    n709
  );


  buf
  g708
  (
    n743,
    n698
  );


  buf
  g709
  (
    n809,
    n705
  );


  not
  g710
  (
    n762,
    n697
  );


  not
  g711
  (
    n792,
    n718
  );


  buf
  g712
  (
    n797,
    n710
  );


  buf
  g713
  (
    n747,
    n707
  );


  not
  g714
  (
    n803,
    n711
  );


  buf
  g715
  (
    n789,
    n704
  );


  not
  g716
  (
    n725,
    n706
  );


  buf
  g717
  (
    n742,
    n715
  );


  buf
  g718
  (
    n727,
    n705
  );


  not
  g719
  (
    n755,
    n709
  );


  not
  g720
  (
    n758,
    n719
  );


  not
  g721
  (
    n778,
    n712
  );


  not
  g722
  (
    n812,
    n710
  );


  buf
  g723
  (
    n774,
    n718
  );


  not
  g724
  (
    n808,
    n697
  );


  not
  g725
  (
    n772,
    n717
  );


  not
  g726
  (
    n730,
    n716
  );


  buf
  g727
  (
    n757,
    n712
  );


  not
  g728
  (
    n731,
    n697
  );


  buf
  g729
  (
    n787,
    n719
  );


  not
  g730
  (
    n768,
    n707
  );


  buf
  g731
  (
    n726,
    n700
  );


  not
  g732
  (
    n733,
    n699
  );


  not
  g733
  (
    n810,
    n702
  );


  not
  g734
  (
    n765,
    n710
  );


  not
  g735
  (
    n802,
    n715
  );


  not
  g736
  (
    n756,
    n703
  );


  not
  g737
  (
    n784,
    n715
  );


  not
  g738
  (
    n744,
    n703
  );


  not
  g739
  (
    n816,
    n714
  );


  buf
  g740
  (
    n782,
    n719
  );


  not
  g741
  (
    n748,
    n698
  );


  not
  g742
  (
    n739,
    n716
  );


  not
  g743
  (
    n728,
    n713
  );


  not
  g744
  (
    n740,
    n702
  );


  buf
  g745
  (
    n767,
    n715
  );


  buf
  g746
  (
    n732,
    n708
  );


  buf
  g747
  (
    n783,
    n714
  );


  not
  g748
  (
    n805,
    n711
  );


  not
  g749
  (
    n785,
    n712
  );


  not
  g750
  (
    n776,
    n708
  );


  not
  g751
  (
    n736,
    n718
  );


  not
  g752
  (
    n766,
    n702
  );


  buf
  g753
  (
    n814,
    n709
  );


  not
  g754
  (
    n801,
    n706
  );


  buf
  g755
  (
    n770,
    n711
  );


  buf
  g756
  (
    n729,
    n717
  );


  buf
  g757
  (
    n791,
    n716
  );


  buf
  g758
  (
    n759,
    n705
  );


  not
  g759
  (
    n780,
    n701
  );


  buf
  g760
  (
    n800,
    n714
  );


  buf
  g761
  (
    n737,
    n708
  );


  buf
  g762
  (
    n813,
    n704
  );


  buf
  g763
  (
    n746,
    n719
  );


  not
  g764
  (
    n760,
    n704
  );


  not
  g765
  (
    n806,
    n717
  );


  buf
  g766
  (
    n799,
    n698
  );


  not
  g767
  (
    KeyWire_0_28,
    n700
  );


  not
  g768
  (
    n741,
    n713
  );


  not
  g769
  (
    n793,
    n717
  );


  not
  g770
  (
    n788,
    n703
  );


  not
  g771
  (
    n750,
    n698
  );


  buf
  g772
  (
    n753,
    n703
  );


  buf
  g773
  (
    n752,
    n710
  );


  not
  g774
  (
    n798,
    n707
  );


  buf
  g775
  (
    n761,
    n699
  );


  buf
  g776
  (
    n804,
    n708
  );


  buf
  g777
  (
    n764,
    n699
  );


  not
  g778
  (
    KeyWire_0_1,
    n706
  );


  not
  g779
  (
    n773,
    n701
  );


  buf
  g780
  (
    n751,
    n700
  );


  not
  g781
  (
    n738,
    n699
  );


  buf
  g782
  (
    n775,
    n701
  );


  buf
  g783
  (
    n754,
    n713
  );


  buf
  g784
  (
    n786,
    n701
  );


  buf
  g785
  (
    n796,
    n700
  );


  buf
  g786
  (
    n771,
    n714
  );


  not
  g787
  (
    n734,
    n709
  );


  buf
  g788
  (
    n794,
    n707
  );


  not
  g789
  (
    n781,
    n702
  );


  nor
  g790
  (
    n826,
    n561,
    n565,
    n563,
    n558
  );


  nand
  g791
  (
    n829,
    n728,
    n726,
    n564,
    n566
  );


  xor
  g792
  (
    n823,
    n557,
    n560,
    n565,
    n725
  );


  or
  g793
  (
    n820,
    n556,
    n565,
    n559,
    n726
  );


  nor
  g794
  (
    n825,
    n560,
    n560,
    n562,
    n563
  );


  xor
  g795
  (
    KeyWire_0_11,
    n563,
    n556,
    n725,
    n562
  );


  nand
  g796
  (
    n827,
    n560,
    n558,
    n557
  );


  nor
  g797
  (
    n824,
    n561,
    n558,
    n563,
    n564
  );


  nand
  g798
  (
    n828,
    n559,
    n727,
    n565,
    n561
  );


  xor
  g799
  (
    n817,
    n725,
    n727,
    n562
  );


  xor
  g800
  (
    n818,
    n726,
    n558,
    n564,
    n559
  );


  xor
  g801
  (
    n821,
    n725,
    n564,
    n557,
    n727
  );


  nor
  g802
  (
    n819,
    n726,
    n559,
    n727,
    n561
  );


  buf
  g803
  (
    n831,
    n817
  );


  nand
  g804
  (
    n830,
    n818,
    n676
  );


  buf
  g805
  (
    n833,
    n831
  );


  not
  g806
  (
    n835,
    n830
  );


  buf
  g807
  (
    n836,
    n831
  );


  buf
  g808
  (
    n832,
    n831
  );


  buf
  g809
  (
    n837,
    n830
  );


  not
  g810
  (
    n838,
    n831
  );


  not
  g811
  (
    n834,
    n830
  );


  buf
  g812
  (
    n839,
    n830
  );


  not
  g813
  (
    n850,
    n835
  );


  not
  g814
  (
    n848,
    n836
  );


  buf
  g815
  (
    n845,
    n834
  );


  buf
  g816
  (
    n843,
    n837
  );


  buf
  g817
  (
    n842,
    n833
  );


  not
  g818
  (
    n847,
    n832
  );


  not
  g819
  (
    n846,
    n835
  );


  buf
  g820
  (
    n849,
    n834
  );


  not
  g821
  (
    n841,
    n833
  );


  buf
  g822
  (
    n844,
    n832
  );


  not
  g823
  (
    n840,
    n836
  );


  not
  g824
  (
    n856,
    n840
  );


  not
  g825
  (
    n851,
    n841
  );


  not
  g826
  (
    n855,
    n840
  );


  not
  g827
  (
    n852,
    n841
  );


  not
  g828
  (
    n857,
    n840
  );


  buf
  g829
  (
    n853,
    n841
  );


  not
  g830
  (
    n854,
    n840
  );


  buf
  g831
  (
    n864,
    n855
  );


  buf
  g832
  (
    n880,
    n854
  );


  buf
  g833
  (
    n877,
    n855
  );


  buf
  g834
  (
    n876,
    n852
  );


  buf
  g835
  (
    n875,
    n851
  );


  not
  g836
  (
    n862,
    n853
  );


  buf
  g837
  (
    n874,
    n853
  );


  buf
  g838
  (
    n867,
    n854
  );


  buf
  g839
  (
    n859,
    n855
  );


  not
  g840
  (
    n868,
    n852
  );


  not
  g841
  (
    n858,
    n852
  );


  not
  g842
  (
    n866,
    n854
  );


  not
  g843
  (
    n872,
    n852
  );


  buf
  g844
  (
    n879,
    n854
  );


  not
  g845
  (
    n865,
    n853
  );


  buf
  g846
  (
    n873,
    n853
  );


  not
  g847
  (
    n860,
    n851
  );


  buf
  g848
  (
    n869,
    n856
  );


  buf
  g849
  (
    n863,
    n851
  );


  buf
  g850
  (
    n871,
    n851
  );


  buf
  g851
  (
    n878,
    n855
  );


  not
  g852
  (
    n870,
    n856
  );


  not
  g853
  (
    KeyWire_0_6,
    n856
  );


  xor
  g854
  (
    n885,
    n567,
    n571,
    n568
  );


  xnor
  g855
  (
    n887,
    n567,
    n566,
    n858
  );


  nor
  g856
  (
    KeyWire_0_19,
    n859,
    n570,
    n568
  );


  or
  g857
  (
    n886,
    n342,
    n859,
    n569
  );


  and
  g858
  (
    n884,
    n567,
    n570,
    n858
  );


  and
  g859
  (
    n881,
    n571,
    n858,
    n569
  );


  xor
  g860
  (
    n883,
    n570,
    n569,
    n568,
    n566
  );


  xnor
  g861
  (
    n888,
    n858,
    n859,
    n567,
    n571
  );


  or
  g862
  (
    n889,
    n885,
    n648,
    n651,
    n649
  );


  nand
  g863
  (
    n896,
    n649,
    n887,
    n652,
    n611
  );


  or
  g864
  (
    n893,
    n888,
    n652,
    n881
  );


  and
  g865
  (
    n894,
    n653,
    n650,
    n648,
    n883
  );


  xnor
  g866
  (
    n892,
    n886,
    n653,
    n882,
    n649
  );


  xor
  g867
  (
    n895,
    n652,
    n653,
    n884,
    n650
  );


  xor
  g868
  (
    n891,
    n650,
    n651,
    n653,
    n649
  );


  and
  g869
  (
    n890,
    n650,
    n648,
    n651
  );


  nand
  g870
  (
    n900,
    n677,
    n678
  );


  xnor
  g871
  (
    n898,
    n677,
    n678,
    n676
  );


  nand
  g872
  (
    n899,
    n676,
    n889,
    n678
  );


  xor
  g873
  (
    n897,
    n889,
    n677
  );


  nand
  g874
  (
    n904,
    n669,
    n598,
    n678
  );


  nor
  g875
  (
    n907,
    n668,
    n898,
    n601,
    n600
  );


  nand
  g876
  (
    n906,
    n897,
    n897,
    n680,
    n898
  );


  nor
  g877
  (
    n909,
    n599,
    n600,
    n679,
    n898
  );


  xor
  g878
  (
    n901,
    n669,
    n897,
    n601,
    n679
  );


  xor
  g879
  (
    n908,
    n680,
    n680,
    n899,
    n597
  );


  xor
  g880
  (
    n911,
    n899,
    n599,
    n668,
    n601
  );


  or
  g881
  (
    n905,
    n898,
    n897,
    n600
  );


  nor
  g882
  (
    n903,
    n598,
    n667,
    n899,
    n680
  );


  xor
  g883
  (
    n910,
    n601,
    n599,
    n597
  );


  nor
  g884
  (
    n902,
    n670,
    n679,
    n598
  );


  nand
  g885
  (
    n914,
    n611,
    n906
  );


  not
  g886
  (
    n912,
    n681
  );


  nor
  g887
  (
    n915,
    n681,
    n907
  );


  nand
  g888
  (
    n916,
    n681,
    n903
  );


  or
  g889
  (
    n913,
    n905,
    n904
  );


  or
  g890
  (
    n917,
    n912,
    n685,
    n686
  );


  and
  g891
  (
    n920,
    n684,
    n685
  );


  and
  g892
  (
    n918,
    n686,
    n913,
    n684,
    n683
  );


  xnor
  g893
  (
    n919,
    n611,
    n914,
    n684,
    n913
  );


  buf
  g894
  (
    n921,
    n919
  );


  xor
  g895
  (
    n922,
    n118,
    n918
  );


  xnor
  g896
  (
    n923,
    n917,
    n920
  );


  buf
  g897
  (
    n924,
    n921
  );


  nand
  g898
  (
    n928,
    n673,
    n900
  );


  xnor
  g899
  (
    n927,
    n671,
    n672,
    n924
  );


  and
  g900
  (
    n925,
    n900,
    n899,
    n672,
    n924
  );


  xor
  g901
  (
    n926,
    n670,
    n900,
    n671,
    n924
  );


  buf
  g902
  (
    n929,
    n925
  );


  nor
  g903
  (
    n930,
    n687,
    n688
  );


  or
  g904
  (
    n933,
    n929,
    n686,
    n687,
    n688
  );


  xnor
  g905
  (
    n932,
    n929,
    n929,
    n687,
    n686
  );


  xor
  g906
  (
    n931,
    n929,
    n688,
    n689
  );


  not
  g907
  (
    n935,
    n931
  );


  buf
  g908
  (
    n936,
    n931
  );


  not
  g909
  (
    n937,
    n930
  );


  buf
  g910
  (
    n938,
    n930
  );


  not
  g911
  (
    n934,
    n930
  );


  buf
  g912
  (
    n939,
    n930
  );


  nor
  g913
  (
    n958,
    n847,
    n496,
    n843
  );


  nor
  g914
  (
    n953,
    n934,
    n849,
    n843,
    n496
  );


  and
  g915
  (
    n960,
    n849,
    n923,
    n921,
    n292
  );


  nor
  g916
  (
    n963,
    n922,
    n292,
    n939,
    n845
  );


  and
  g917
  (
    n951,
    n923,
    n846,
    n922,
    n937
  );


  xor
  g918
  (
    n940,
    n939,
    n496,
    n937,
    n843
  );


  nor
  g919
  (
    n943,
    n848,
    n495,
    n934,
    n937
  );


  and
  g920
  (
    n944,
    n844,
    n935,
    n850,
    n291
  );


  xor
  g921
  (
    n959,
    n841,
    n922,
    n498
  );


  nor
  g922
  (
    n947,
    n848,
    n499,
    n845,
    n291
  );


  xnor
  g923
  (
    n946,
    n842,
    n934,
    n935,
    n937
  );


  and
  g924
  (
    n942,
    n938,
    n499,
    n847,
    n850
  );


  nand
  g925
  (
    n954,
    n497,
    n922,
    n292
  );


  xnor
  g926
  (
    n961,
    n850,
    n846,
    n936,
    n923
  );


  and
  g927
  (
    n956,
    n842,
    n935,
    n936,
    n921
  );


  nor
  g928
  (
    n952,
    n499,
    n939,
    n498,
    n935
  );


  and
  g929
  (
    n945,
    n498,
    n939,
    n497,
    n921
  );


  xnor
  g930
  (
    n955,
    n845,
    n934,
    n936,
    n495
  );


  nand
  g931
  (
    n950,
    n923,
    n938,
    n845,
    n849
  );


  xnor
  g932
  (
    n957,
    n847,
    n938,
    n848,
    n850
  );


  nor
  g933
  (
    n948,
    n936,
    n844,
    n846,
    n842
  );


  xnor
  g934
  (
    n962,
    n499,
    n848,
    n497
  );


  and
  g935
  (
    n949,
    n938,
    n844,
    n842,
    n847
  );


  nor
  g936
  (
    n941,
    n846,
    n844,
    n849,
    n843
  );


  buf
  g937
  (
    n1009,
    n958
  );


  buf
  g938
  (
    n1047,
    n505
  );


  buf
  g939
  (
    n1024,
    n723
  );


  not
  g940
  (
    n980,
    n724
  );


  not
  g941
  (
    n1012,
    n955
  );


  not
  g942
  (
    n1006,
    n952
  );


  not
  g943
  (
    n1008,
    n516
  );


  not
  g944
  (
    n1044,
    n513
  );


  buf
  g945
  (
    n1049,
    n942
  );


  not
  g946
  (
    n1027,
    n944
  );


  not
  g947
  (
    n1040,
    n959
  );


  buf
  g948
  (
    n998,
    n941
  );


  buf
  g949
  (
    n990,
    n950
  );


  not
  g950
  (
    n1055,
    n506
  );


  not
  g951
  (
    n1004,
    n953
  );


  not
  g952
  (
    n981,
    n949
  );


  buf
  g953
  (
    n988,
    n945
  );


  not
  g954
  (
    n978,
    n503
  );


  buf
  g955
  (
    n1052,
    n857
  );


  not
  g956
  (
    n984,
    n512
  );


  not
  g957
  (
    n968,
    n951
  );


  not
  g958
  (
    n1018,
    n956
  );


  buf
  g959
  (
    n966,
    n508
  );


  not
  g960
  (
    n1005,
    n910
  );


  not
  g961
  (
    n974,
    n940
  );


  not
  g962
  (
    n967,
    n723
  );


  buf
  g963
  (
    n1002,
    n949
  );


  not
  g964
  (
    n965,
    n942
  );


  buf
  g965
  (
    n1041,
    n946
  );


  not
  g966
  (
    n997,
    n611
  );


  not
  g967
  (
    n1042,
    n957
  );


  not
  g968
  (
    n1051,
    n953
  );


  not
  g969
  (
    n1026,
    n961
  );


  buf
  g970
  (
    n1032,
    n504
  );


  not
  g971
  (
    n1050,
    n941
  );


  not
  g972
  (
    n986,
    n960
  );


  not
  g973
  (
    n1036,
    n509
  );


  not
  g974
  (
    n1003,
    n953
  );


  buf
  g975
  (
    n992,
    n515
  );


  buf
  g976
  (
    n1016,
    n957
  );


  buf
  g977
  (
    n983,
    n943
  );


  buf
  g978
  (
    n987,
    n689
  );


  buf
  g979
  (
    n1010,
    n952
  );


  buf
  g980
  (
    n969,
    n948
  );


  not
  g981
  (
    n1014,
    n952
  );


  buf
  g982
  (
    n1059,
    n508
  );


  buf
  g983
  (
    n970,
    n514
  );


  not
  g984
  (
    n1025,
    n949
  );


  buf
  g985
  (
    n993,
    n510
  );


  not
  g986
  (
    n1030,
    n857
  );


  not
  g987
  (
    n1011,
    n958
  );


  not
  g988
  (
    n1021,
    n506
  );


  buf
  g989
  (
    n1045,
    n954
  );


  buf
  g990
  (
    n1022,
    n948
  );


  buf
  g991
  (
    n985,
    n952
  );


  not
  g992
  (
    n1019,
    n947
  );


  buf
  g993
  (
    n1037,
    n959
  );


  buf
  g994
  (
    n991,
    n857
  );


  not
  g995
  (
    n989,
    n954
  );


  buf
  g996
  (
    n1029,
    n908
  );


  not
  g997
  (
    n964,
    n941
  );


  not
  g998
  (
    n1023,
    n511
  );


  buf
  g999
  (
    n1034,
    n612
  );


  buf
  g1000
  (
    n1013,
    n956
  );


  not
  g1001
  (
    n1028,
    n943
  );


  buf
  g1002
  (
    n1058,
    n960
  );


  buf
  g1003
  (
    n1057,
    n962
  );


  not
  g1004
  (
    n1031,
    n507
  );


  buf
  g1005
  (
    n1033,
    n941
  );


  buf
  g1006
  (
    n1035,
    n945
  );


  not
  g1007
  (
    n1039,
    n503
  );


  buf
  g1008
  (
    n982,
    n515
  );


  or
  g1009
  (
    n1007,
    n940,
    n509,
    n721,
    n722
  );


  xor
  g1010
  (
    n999,
    n954,
    n958,
    n857,
    n957
  );


  and
  g1011
  (
    n1046,
    n961,
    n950,
    n945,
    n944
  );


  xnor
  g1012
  (
    n1020,
    n961,
    n512,
    n723,
    n940
  );


  xnor
  g1013
  (
    n971,
    n504,
    n962,
    n510
  );


  nor
  g1014
  (
    n977,
    n946,
    n948,
    n954,
    n911
  );


  xor
  g1015
  (
    n1053,
    n962,
    n956,
    n951,
    n728
  );


  or
  g1016
  (
    n1043,
    n957,
    n721,
    n612,
    n909
  );


  xor
  g1017
  (
    n995,
    n960,
    n447,
    n940,
    n950
  );


  xor
  g1018
  (
    n1017,
    n856,
    n946,
    n505,
    n944
  );


  or
  g1019
  (
    n1001,
    n518,
    n947,
    n963,
    n961
  );


  or
  g1020
  (
    n979,
    n518,
    n723,
    n948,
    n721
  );


  nor
  g1021
  (
    n975,
    n943,
    n963,
    n612,
    n959
  );


  nand
  g1022
  (
    n1048,
    n955,
    n724,
    n514,
    n507
  );


  nor
  g1023
  (
    n1015,
    n955,
    n950,
    n722,
    n511
  );


  nand
  g1024
  (
    n996,
    n943,
    n942,
    n519,
    n949
  );


  xnor
  g1025
  (
    n1054,
    n942,
    n502,
    n720,
    n689
  );


  and
  g1026
  (
    n1000,
    n963,
    n953,
    n513,
    n720
  );


  xnor
  g1027
  (
    n1056,
    n722,
    n517,
    n963,
    n955
  );


  nand
  g1028
  (
    n976,
    n944,
    n720,
    n951,
    n724
  );


  nand
  g1029
  (
    n972,
    n724,
    n947,
    n945,
    n958
  );


  xnor
  g1030
  (
    n973,
    n612,
    n722,
    n959,
    n960
  );


  and
  g1031
  (
    n994,
    n516,
    n720,
    n956,
    n947
  );


  or
  g1032
  (
    n1038,
    n951,
    n517,
    n721,
    n946
  );


  nand
  g1033
  (
    n1220,
    n796,
    n925
  );


  xor
  g1034
  (
    n1222,
    n751,
    n1036
  );


  xor
  g1035
  (
    n1287,
    n730,
    n808
  );


  and
  g1036
  (
    KeyWire_0_15,
    n765,
    n764
  );


  xor
  g1037
  (
    n1296,
    n1023,
    n1041
  );


  xor
  g1038
  (
    n1146,
    n741,
    n799
  );


  and
  g1039
  (
    n1214,
    n760,
    n1051
  );


  and
  g1040
  (
    n1138,
    n814,
    n471
  );


  xnor
  g1041
  (
    n1212,
    n753,
    n477
  );


  and
  g1042
  (
    KeyWire_0_7,
    n783,
    n751
  );


  xnor
  g1043
  (
    n1128,
    n780,
    n786
  );


  xnor
  g1044
  (
    n1251,
    n1034,
    n791
  );


  xnor
  g1045
  (
    n1260,
    n927,
    n803
  );


  nand
  g1046
  (
    n1211,
    n1033,
    n914
  );


  nor
  g1047
  (
    n1142,
    n758,
    n808
  );


  nand
  g1048
  (
    n1088,
    n860,
    n747
  );


  xnor
  g1049
  (
    n1154,
    n971,
    n1046
  );


  xnor
  g1050
  (
    n1118,
    n974,
    n1011
  );


  xnor
  g1051
  (
    n1283,
    n807,
    n1003
  );


  nand
  g1052
  (
    n1217,
    n752,
    n806
  );


  xor
  g1053
  (
    n1240,
    n1039,
    n1009
  );


  nor
  g1054
  (
    n1186,
    n965,
    n742
  );


  or
  g1055
  (
    n1136,
    n1027,
    n870,
    n1031
  );


  and
  g1056
  (
    n1095,
    n478,
    n1031,
    n1051,
    n1026
  );


  xnor
  g1057
  (
    n1074,
    n740,
    n760,
    n979,
    n964
  );


  and
  g1058
  (
    n1278,
    n477,
    n1053,
    n975,
    n978
  );


  nand
  g1059
  (
    n1170,
    n739,
    n981,
    n746,
    n788
  );


  and
  g1060
  (
    n1120,
    n778,
    n972,
    n973,
    n728
  );


  xnor
  g1061
  (
    n1158,
    n791,
    n774,
    n1030,
    n736
  );


  nand
  g1062
  (
    n1275,
    n1044,
    n1017,
    n980,
    n729
  );


  nand
  g1063
  (
    n1221,
    n868,
    n1022,
    n1025,
    n791
  );


  nor
  g1064
  (
    n1255,
    n731,
    n744,
    n803,
    n877
  );


  and
  g1065
  (
    n1270,
    n1008,
    n748,
    n757,
    n774
  );


  nand
  g1066
  (
    n1235,
    n870,
    n819,
    n777,
    n478
  );


  nor
  g1067
  (
    n1234,
    n1044,
    n998,
    n990,
    n1022
  );


  and
  g1068
  (
    n1151,
    n777,
    n793,
    n464,
    n742
  );


  xor
  g1069
  (
    n1267,
    n469,
    n993,
    n977,
    n779
  );


  or
  g1070
  (
    n1078,
    n794,
    n809,
    n763,
    n766
  );


  nand
  g1071
  (
    n1086,
    n826,
    n1055,
    n475,
    n738
  );


  nand
  g1072
  (
    n1064,
    n1043,
    n1053,
    n1002,
    n968
  );


  nand
  g1073
  (
    n1139,
    n767,
    n1022,
    n1040,
    n810
  );


  or
  g1074
  (
    n1273,
    n871,
    n969,
    n735,
    n1052
  );


  nand
  g1075
  (
    n1153,
    n797,
    n974,
    n1056,
    n1036
  );


  xor
  g1076
  (
    n1197,
    n782,
    n811,
    n996,
    n1006
  );


  xnor
  g1077
  (
    n1266,
    n731,
    n741,
    n864,
    n1049
  );


  xnor
  g1078
  (
    n1203,
    n481,
    n768,
    n808,
    n875
  );


  or
  g1079
  (
    n1104,
    n808,
    n1001,
    n813,
    n1026
  );


  xnor
  g1080
  (
    n1070,
    n736,
    n1027,
    n872,
    n867
  );


  nor
  g1081
  (
    n1143,
    n1019,
    n873,
    n747,
    n1057
  );


  or
  g1082
  (
    n1168,
    n1019,
    n980,
    n749,
    n990
  );


  and
  g1083
  (
    n1236,
    n794,
    n769,
    n766,
    n472
  );


  nand
  g1084
  (
    n1259,
    n1054,
    n463,
    n986,
    n789
  );


  and
  g1085
  (
    n1124,
    n775,
    n797,
    n816,
    n784
  );


  nor
  g1086
  (
    n1130,
    n788,
    n770,
    n797,
    n465
  );


  and
  g1087
  (
    n1119,
    n1034,
    n758,
    n785,
    n873
  );


  nand
  g1088
  (
    n1167,
    n749,
    n733,
    n1031,
    n761
  );


  xnor
  g1089
  (
    n1081,
    n928,
    n984,
    n783,
    n729
  );


  nor
  g1090
  (
    n1094,
    n1012,
    n733,
    n927,
    n822
  );


  xor
  g1091
  (
    n1258,
    n999,
    n1019,
    n765,
    n784
  );


  or
  g1092
  (
    n1091,
    n776,
    n1055,
    n478,
    n524
  );


  or
  g1093
  (
    n1152,
    n777,
    n770,
    n807,
    n767
  );


  nand
  g1094
  (
    n1286,
    n986,
    n869,
    n768,
    n990
  );


  nor
  g1095
  (
    n1297,
    n737,
    n750,
    n812
  );


  or
  g1096
  (
    n1210,
    n1018,
    n967,
    n741,
    n467
  );


  or
  g1097
  (
    n1106,
    n798,
    n813,
    n983,
    n824
  );


  or
  g1098
  (
    n1096,
    n971,
    n739,
    n976,
    n863
  );


  xor
  g1099
  (
    n1272,
    n860,
    n1015,
    n967,
    n1041
  );


  xnor
  g1100
  (
    n1125,
    n1008,
    n473,
    n926,
    n970
  );


  nor
  g1101
  (
    n1245,
    n972,
    n1048,
    n1032,
    n768
  );


  xor
  g1102
  (
    n1108,
    n1012,
    n1011,
    n875,
    n984
  );


  xnor
  g1103
  (
    n1162,
    n777,
    n782,
    n785,
    n765
  );


  or
  g1104
  (
    n1145,
    n987,
    n731,
    n973,
    n773
  );


  xor
  g1105
  (
    n1198,
    n974,
    n751,
    n1007,
    n1059
  );


  nand
  g1106
  (
    n1116,
    n916,
    n476,
    n1040,
    n968
  );


  and
  g1107
  (
    n1061,
    n1037,
    n734,
    n798,
    n1016
  );


  nand
  g1108
  (
    n1131,
    n759,
    n748,
    n1040,
    n1026
  );


  xnor
  g1109
  (
    n1292,
    n964,
    n864,
    n863,
    n801
  );


  nor
  g1110
  (
    n1298,
    n983,
    n763,
    n775,
    n865
  );


  xnor
  g1111
  (
    n1175,
    n759,
    n872,
    n1010,
    n978
  );


  xor
  g1112
  (
    n1279,
    n748,
    n968,
    n807,
    n471
  );


  xnor
  g1113
  (
    n1159,
    n827,
    n1000,
    n873,
    n987
  );


  and
  g1114
  (
    n1102,
    n828,
    n466,
    n756,
    n462
  );


  nor
  g1115
  (
    n1242,
    n994,
    n1034,
    n730,
    n737
  );


  and
  g1116
  (
    n1177,
    n875,
    n1042,
    n472,
    n475
  );


  and
  g1117
  (
    n1093,
    n764,
    n993,
    n467,
    n1030
  );


  nor
  g1118
  (
    n1063,
    n972,
    n789,
    n1057,
    n1009
  );


  nand
  g1119
  (
    n1201,
    n762,
    n1050,
    n755,
    n735
  );


  and
  g1120
  (
    n1176,
    n793,
    n975,
    n973,
    n997
  );


  xor
  g1121
  (
    n1190,
    n926,
    n995,
    n782
  );


  and
  g1122
  (
    n1157,
    n964,
    n755,
    n1000,
    n786
  );


  and
  g1123
  (
    n1299,
    n786,
    n810,
    n1014,
    n468
  );


  and
  g1124
  (
    n1179,
    n877,
    n729,
    n799,
    n1014
  );


  nand
  g1125
  (
    n1281,
    n992,
    n754,
    n792,
    n1034
  );


  and
  g1126
  (
    n1288,
    n1037,
    n827,
    n991,
    n795
  );


  nor
  g1127
  (
    n1300,
    n770,
    n781,
    n991,
    n1007
  );


  nor
  g1128
  (
    n1276,
    n1004,
    n965,
    n976,
    n986
  );


  nand
  g1129
  (
    n1226,
    n994,
    n1018,
    n925,
    n1024
  );


  and
  g1130
  (
    n1105,
    n813,
    n468,
    n970,
    n820
  );


  or
  g1131
  (
    n1092,
    n799,
    n475,
    n469,
    n871
  );


  nand
  g1132
  (
    n1204,
    n814,
    n1052,
    n1045,
    n794
  );


  and
  g1133
  (
    n1219,
    n968,
    n460,
    n1037,
    n1050
  );


  nand
  g1134
  (
    n1182,
    n1016,
    n916,
    n803,
    n481
  );


  nor
  g1135
  (
    n1223,
    n739,
    n969,
    n1039,
    n473
  );


  xor
  g1136
  (
    n1254,
    n1025,
    n739,
    n1033,
    n1054
  );


  and
  g1137
  (
    n1230,
    n759,
    n1016,
    n1020,
    n740
  );


  and
  g1138
  (
    n1293,
    n985,
    n468,
    n761,
    n473
  );


  nand
  g1139
  (
    n1077,
    n800,
    n1001,
    n1035,
    n997
  );


  xnor
  g1140
  (
    n1225,
    n1006,
    n985,
    n1015,
    n868
  );


  xor
  g1141
  (
    n1079,
    n1039,
    n1011,
    n1029,
    n480
  );


  nand
  g1142
  (
    n1140,
    n806,
    n795,
    n740,
    n748
  );


  xor
  g1143
  (
    n1196,
    n787,
    n976,
    n757,
    n465
  );


  and
  g1144
  (
    n1295,
    n476,
    n733,
    n471,
    n1025
  );


  xor
  g1145
  (
    n1246,
    n772,
    n471,
    n866,
    n760
  );


  xor
  g1146
  (
    n1087,
    n975,
    n880,
    n754,
    n928
  );


  nand
  g1147
  (
    n1249,
    n472,
    n801,
    n790,
    n1046
  );


  nor
  g1148
  (
    n1269,
    n1047,
    n805,
    n997,
    n769
  );


  xnor
  g1149
  (
    n1183,
    n980,
    n470,
    n996,
    n813
  );


  or
  g1150
  (
    n1189,
    n1026,
    n1005,
    n1045,
    n781
  );


  or
  g1151
  (
    n1231,
    n1018,
    n809,
    n816
  );


  xor
  g1152
  (
    n1213,
    n1010,
    n870,
    n823,
    n466
  );


  or
  g1153
  (
    n1285,
    n771,
    n743,
    n879,
    n964
  );


  nand
  g1154
  (
    n1248,
    n781,
    n481,
    n1004,
    n1044
  );


  xor
  g1155
  (
    n1277,
    n735,
    n809,
    n1002,
    n1006
  );


  or
  g1156
  (
    n1180,
    n1031,
    n469,
    n794,
    n989
  );


  nand
  g1157
  (
    n1261,
    n992,
    n815,
    n792,
    n872
  );


  and
  g1158
  (
    n1257,
    n743,
    n998,
    n971,
    n761
  );


  xnor
  g1159
  (
    n1244,
    n740,
    n749,
    n461,
    n1025
  );


  nand
  g1160
  (
    n1173,
    n1020,
    n765,
    n868,
    n805
  );


  xnor
  g1161
  (
    n1228,
    n774,
    n769,
    n736,
    n987
  );


  nand
  g1162
  (
    n1290,
    n979,
    n877,
    n473,
    n474
  );


  or
  g1163
  (
    n1265,
    n779,
    n747,
    n782,
    n788
  );


  and
  g1164
  (
    n1218,
    n762,
    n1033,
    n1044,
    n1013
  );


  nand
  g1165
  (
    n1137,
    n993,
    n1003,
    n780,
    n746
  );


  xor
  g1166
  (
    n1181,
    n1003,
    n1038,
    n1058,
    n477
  );


  or
  g1167
  (
    n1150,
    n772,
    n478,
    n1013,
    n1054
  );


  nand
  g1168
  (
    n1155,
    n750,
    n970,
    n804,
    n982
  );


  xor
  g1169
  (
    n1171,
    n977,
    n800,
    n804,
    n469
  );


  xor
  g1170
  (
    n1156,
    n735,
    n992,
    n783,
    n1014
  );


  xor
  g1171
  (
    n1282,
    n1056,
    n874,
    n1004,
    n1014
  );


  xnor
  g1172
  (
    n1103,
    n775,
    n744,
    n987,
    n1029
  );


  or
  g1173
  (
    n1147,
    n1007,
    n863,
    n880,
    n994
  );


  or
  g1174
  (
    n1085,
    n798,
    n1007,
    n1011,
    n785
  );


  and
  g1175
  (
    n1185,
    n866,
    n811,
    n815,
    n464
  );


  nand
  g1176
  (
    n1135,
    n737,
    n1035,
    n861,
    n474
  );


  nor
  g1177
  (
    n1187,
    n988,
    n1032,
    n1022,
    n756
  );


  nand
  g1178
  (
    n1099,
    n738,
    n762,
    n756,
    n1013
  );


  nand
  g1179
  (
    n1083,
    n1057,
    n1012,
    n874,
    n998
  );


  xor
  g1180
  (
    n1060,
    n1043,
    n860,
    n790,
    n828
  );


  nor
  g1181
  (
    n1301,
    n1012,
    n995,
    n795,
    n772
  );


  nor
  g1182
  (
    n1284,
    n746,
    n767,
    n989,
    n790
  );


  nor
  g1183
  (
    n1229,
    n1030,
    n742,
    n745,
    n871
  );


  or
  g1184
  (
    n1280,
    n1046,
    n1005,
    n1027,
    n778
  );


  and
  g1185
  (
    n1098,
    n1032,
    n1043,
    n466,
    n479
  );


  xnor
  g1186
  (
    n1090,
    n476,
    n738,
    n925,
    n461
  );


  or
  g1187
  (
    n1264,
    n878,
    n755,
    n811,
    n1023
  );


  or
  g1188
  (
    n1164,
    n879,
    n752,
    n1023,
    n1010
  );


  or
  g1189
  (
    n1208,
    n1016,
    n728,
    n1005,
    n1028
  );


  or
  g1190
  (
    n1134,
    n814,
    n1005,
    n1046,
    n798
  );


  or
  g1191
  (
    n1294,
    n966,
    n984,
    n866,
    n1000
  );


  nand
  g1192
  (
    n1227,
    n758,
    n928,
    n988,
    n1059
  );


  xnor
  g1193
  (
    n1233,
    n1059,
    n743,
    n784,
    n983
  );


  xnor
  g1194
  (
    n1305,
    n1036,
    n991,
    n801,
    n981
  );


  or
  g1195
  (
    n1205,
    n1053,
    n775,
    n732,
    n472
  );


  and
  g1196
  (
    n1289,
    n811,
    n480,
    n872,
    n965
  );


  and
  g1197
  (
    n1065,
    n876,
    n821,
    n1004,
    n1024
  );


  xnor
  g1198
  (
    n1241,
    n752,
    n470,
    n755,
    n731
  );


  xnor
  g1199
  (
    n1112,
    n793,
    n874,
    n768,
    n879
  );


  nand
  g1200
  (
    n1192,
    n869,
    n879,
    n464,
    n754
  );


  xor
  g1201
  (
    n1115,
    n995,
    n1038,
    n734,
    n1018
  );


  or
  g1202
  (
    n1263,
    n759,
    n971,
    n771,
    n760
  );


  nor
  g1203
  (
    n1268,
    n1052,
    n975,
    n730,
    n1003
  );


  nor
  g1204
  (
    n1113,
    n867,
    n978,
    n464,
    n1047
  );


  xnor
  g1205
  (
    n1243,
    n792,
    n1032,
    n806,
    n1015
  );


  nand
  g1206
  (
    n1148,
    n1051,
    n474,
    n1002,
    n738
  );


  and
  g1207
  (
    n1123,
    n999,
    n876,
    n985,
    n787
  );


  nand
  g1208
  (
    n1133,
    n804,
    n461,
    n789,
    n729
  );


  nand
  g1209
  (
    n1066,
    n997,
    n877,
    n763,
    n1008
  );


  or
  g1210
  (
    n1252,
    n1036,
    n861,
    n1040,
    n462
  );


  nand
  g1211
  (
    n1206,
    n470,
    n1024,
    n815,
    n465
  );


  and
  g1212
  (
    n1160,
    n747,
    n757,
    n800,
    n1048
  );


  or
  g1213
  (
    n1216,
    n1035,
    n733,
    n988,
    n796
  );


  or
  g1214
  (
    n1144,
    n927,
    n862,
    n810,
    n1002
  );


  and
  g1215
  (
    n1306,
    n462,
    n734,
    n977,
    n976
  );


  nor
  g1216
  (
    n1161,
    n1042,
    n1027,
    n1041,
    n1028
  );


  nand
  g1217
  (
    n1178,
    n873,
    n773,
    n793,
    n812
  );


  xor
  g1218
  (
    n1224,
    n800,
    n480,
    n479,
    n1057
  );


  xor
  g1219
  (
    n1109,
    n1058,
    n778,
    n992,
    n756
  );


  or
  g1220
  (
    n1237,
    n970,
    n876,
    n999,
    n802
  );


  nor
  g1221
  (
    n1100,
    n799,
    n788,
    n779,
    n926
  );


  xor
  g1222
  (
    n1184,
    n994,
    n465,
    n1021,
    n461
  );


  xnor
  g1223
  (
    n1122,
    n1049,
    n776,
    n814,
    n730
  );


  xnor
  g1224
  (
    n1166,
    n1053,
    n1055,
    n1045,
    n753
  );


  nand
  g1225
  (
    n1068,
    n466,
    n736,
    n1050,
    n825
  );


  and
  g1226
  (
    n1250,
    n990,
    n973,
    n870,
    n880
  );


  xnor
  g1227
  (
    n1274,
    n1035,
    n1030,
    n743,
    n915
  );


  and
  g1228
  (
    n1084,
    n771,
    n766,
    n974,
    n753
  );


  and
  g1229
  (
    n1117,
    n774,
    n988,
    n989,
    n773
  );


  nor
  g1230
  (
    n1126,
    n865,
    n1013,
    n757,
    n986
  );


  nor
  g1231
  (
    n1207,
    n982,
    n878,
    n479,
    n791
  );


  xor
  g1232
  (
    n1072,
    n1045,
    n1029,
    n861,
    n862
  );


  nor
  g1233
  (
    n1163,
    n862,
    n762,
    n734,
    n816
  );


  xor
  g1234
  (
    n1238,
    n1017,
    n778,
    n737,
    n732
  );


  nor
  g1235
  (
    n1062,
    n801,
    n480,
    n752,
    n754
  );


  nor
  g1236
  (
    n1215,
    n751,
    n1039,
    n467,
    n780
  );


  xnor
  g1237
  (
    n1239,
    n481,
    n983,
    n766,
    n744
  );


  nand
  g1238
  (
    n1076,
    n1047,
    n773,
    n772,
    n1019
  );


  xnor
  g1239
  (
    n1127,
    n875,
    n744,
    n1052,
    n866
  );


  or
  g1240
  (
    n1169,
    n1009,
    n880,
    n865,
    n764
  );


  or
  g1241
  (
    n1071,
    n761,
    n1041,
    n783,
    n470
  );


  or
  g1242
  (
    n1101,
    n796,
    n864,
    n874,
    n795
  );


  xor
  g1243
  (
    n1082,
    n1049,
    n996,
    n1021,
    n780
  );


  xor
  g1244
  (
    n1209,
    n979,
    n806,
    n1009,
    n797
  );


  nand
  g1245
  (
    n1304,
    n867,
    n1017,
    n796,
    n732
  );


  or
  g1246
  (
    n1193,
    n861,
    n746,
    n479,
    n785
  );


  nand
  g1247
  (
    n1302,
    n862,
    n981,
    n776,
    n477
  );


  xor
  g1248
  (
    n1110,
    n1056,
    n977,
    n803,
    n928
  );


  and
  g1249
  (
    n1303,
    n804,
    n468,
    n750,
    n745
  );


  and
  g1250
  (
    n1195,
    n763,
    n991,
    n1047,
    n462
  );


  nand
  g1251
  (
    n1256,
    n810,
    n1029,
    n969,
    n1037
  );


  nor
  g1252
  (
    n1129,
    n989,
    n463,
    n1008,
    n802
  );


  or
  g1253
  (
    n1172,
    n787,
    n1006,
    n770,
    n1042
  );


  nor
  g1254
  (
    KeyWire_0_18,
    n1010,
    n863,
    n815,
    n1021
  );


  xor
  g1255
  (
    n1271,
    n467,
    n476,
    n475,
    n1058
  );


  xor
  g1256
  (
    n1097,
    n1017,
    n865,
    n1051,
    n792
  );


  xor
  g1257
  (
    n1200,
    n878,
    n802,
    n1059,
    n965
  );


  nand
  g1258
  (
    n1080,
    n784,
    n1042,
    n1043,
    n980
  );


  and
  g1259
  (
    n1089,
    n871,
    n878,
    n742,
    n776
  );


  or
  g1260
  (
    n1141,
    n985,
    n979,
    n967,
    n789
  );


  xnor
  g1261
  (
    n1253,
    n966,
    n1038,
    n1050,
    n745
  );


  xnor
  g1262
  (
    n1188,
    n1048,
    n1028,
    n1054,
    n1058
  );


  nand
  g1263
  (
    n1132,
    n1028,
    n1038,
    n1001,
    n1020
  );


  or
  g1264
  (
    n1262,
    n1033,
    n876,
    n982,
    n967
  );


  xnor
  g1265
  (
    KeyWire_0_5,
    n981,
    n978,
    n463,
    n750
  );


  nand
  g1266
  (
    n1232,
    n805,
    n1001,
    n998,
    n966
  );


  xnor
  g1267
  (
    n1073,
    n972,
    n749,
    n829,
    n779
  );


  or
  g1268
  (
    n1114,
    n829,
    n1056,
    n787,
    n732
  );


  nor
  g1269
  (
    n1107,
    n745,
    n982,
    n1024,
    n758
  );


  xor
  g1270
  (
    n1202,
    n869,
    n864,
    n868,
    n1021
  );


  xor
  g1271
  (
    n1247,
    n790,
    n969,
    n1020,
    n1023
  );


  and
  g1272
  (
    n1191,
    n915,
    n1049,
    n802,
    n764
  );


  or
  g1273
  (
    n1067,
    n993,
    n1055,
    n767,
    n996
  );


  nor
  g1274
  (
    n1199,
    n805,
    n741,
    n1015,
    n807
  );


  xnor
  g1275
  (
    n1165,
    n753,
    n1048,
    n1000,
    n771
  );


  xnor
  g1276
  (
    n1075,
    n769,
    n786,
    n809,
    n867
  );


  nand
  g1277
  (
    n1121,
    n860,
    n781,
    n999,
    n927
  );


  xnor
  g1278
  (
    n1111,
    n812,
    n966,
    n524,
    n984
  );


  xor
  g1279
  (
    n1174,
    n869,
    n474,
    n926,
    n463
  );


  buf
  g1280
  (
    n1308,
    n1240
  );


  buf
  g1281
  (
    n1389,
    n1138
  );


  buf
  g1282
  (
    KeyWire_0_27,
    n1128
  );


  not
  g1283
  (
    n1558,
    n1257
  );


  not
  g1284
  (
    n1321,
    n1288
  );


  not
  g1285
  (
    n1435,
    n1111
  );


  not
  g1286
  (
    n1366,
    n1074
  );


  buf
  g1287
  (
    n1469,
    n1161
  );


  not
  g1288
  (
    n1332,
    n1276
  );


  not
  g1289
  (
    n1313,
    n1266
  );


  not
  g1290
  (
    n1404,
    n1151
  );


  buf
  g1291
  (
    n1531,
    n1075
  );


  not
  g1292
  (
    n1382,
    n1300
  );


  buf
  g1293
  (
    n1523,
    n1144
  );


  not
  g1294
  (
    n1380,
    n1109
  );


  not
  g1295
  (
    n1360,
    n1180
  );


  buf
  g1296
  (
    n1470,
    n1146
  );


  not
  g1297
  (
    n1559,
    n1134
  );


  buf
  g1298
  (
    n1471,
    n1235
  );


  not
  g1299
  (
    n1311,
    n1231
  );


  buf
  g1300
  (
    n1438,
    n1263
  );


  buf
  g1301
  (
    n1526,
    n1205
  );


  not
  g1302
  (
    n1467,
    n1237
  );


  not
  g1303
  (
    n1393,
    n1215
  );


  not
  g1304
  (
    n1455,
    n1199
  );


  not
  g1305
  (
    n1554,
    n1167
  );


  buf
  g1306
  (
    n1362,
    n1260
  );


  buf
  g1307
  (
    n1461,
    n1264
  );


  buf
  g1308
  (
    n1540,
    n1133
  );


  buf
  g1309
  (
    n1319,
    n1140
  );


  not
  g1310
  (
    n1529,
    n1084
  );


  buf
  g1311
  (
    n1549,
    n1254
  );


  nand
  g1312
  (
    n1532,
    n1079,
    n1148,
    n1197,
    n1068
  );


  xor
  g1313
  (
    n1449,
    n1137,
    n1156,
    n1284,
    n1268
  );


  or
  g1314
  (
    n1342,
    n1298,
    n1283,
    n1121,
    n1295
  );


  or
  g1315
  (
    n1309,
    n1109,
    n1137,
    n1071,
    n1274
  );


  nor
  g1316
  (
    n1545,
    n1099,
    n1157,
    n1084,
    n1135
  );


  nand
  g1317
  (
    KeyWire_0_8,
    n1211,
    n1223,
    n1065,
    n1124
  );


  xor
  g1318
  (
    n1326,
    n1196,
    n1070,
    n1078,
    n1245
  );


  and
  g1319
  (
    n1562,
    n1262,
    n1283,
    n1167,
    n1163
  );


  xnor
  g1320
  (
    n1436,
    n1150,
    n1183,
    n1195,
    n1086
  );


  nor
  g1321
  (
    n1394,
    n1217,
    n1226,
    n1131,
    n1138
  );


  and
  g1322
  (
    n1421,
    n1244,
    n1153,
    n1173,
    n1094
  );


  xor
  g1323
  (
    n1424,
    n1152,
    n1272,
    n1090,
    n1236
  );


  xnor
  g1324
  (
    n1507,
    n1079,
    n1089,
    n1287,
    n1066
  );


  nand
  g1325
  (
    n1476,
    n1299,
    n1196,
    n1263,
    n1118
  );


  and
  g1326
  (
    n1355,
    n1249,
    n1253,
    n1297,
    n1237
  );


  or
  g1327
  (
    n1350,
    n1127,
    n1234,
    n1258
  );


  xor
  g1328
  (
    n1553,
    n1220,
    n1151,
    n1228,
    n1067
  );


  nand
  g1329
  (
    n1493,
    n1227,
    n1302,
    n1175,
    n1177
  );


  nor
  g1330
  (
    n1506,
    n1213,
    n1241,
    n1261,
    n1165
  );


  and
  g1331
  (
    n1511,
    n1277,
    n1114,
    n1129,
    n1074
  );


  nor
  g1332
  (
    n1518,
    n1110,
    n1238,
    n1136,
    n1098
  );


  xor
  g1333
  (
    n1427,
    n1246,
    n1215,
    n1120,
    n1230
  );


  nor
  g1334
  (
    KeyWire_0_25,
    n1096,
    n1091,
    n1080,
    n1109
  );


  nor
  g1335
  (
    n1398,
    n1227,
    n1200,
    n1279,
    n1271
  );


  xor
  g1336
  (
    n1503,
    n1076,
    n1156,
    n1181,
    n1180
  );


  xnor
  g1337
  (
    n1333,
    n1274,
    n383,
    n1112,
    n1252
  );


  nand
  g1338
  (
    n1539,
    n1300,
    n1107,
    n1213,
    n1285
  );


  nand
  g1339
  (
    n1397,
    n1280,
    n1243,
    n1162,
    n1089
  );


  and
  g1340
  (
    n1315,
    n1277,
    n1256,
    n1159,
    n1244
  );


  or
  g1341
  (
    n1433,
    n1125,
    n1192,
    n1225,
    n1258
  );


  xnor
  g1342
  (
    n1445,
    n1218,
    n1123,
    n1087,
    n1165
  );


  nand
  g1343
  (
    n1542,
    n1287,
    n1123,
    n1147,
    n1260
  );


  nor
  g1344
  (
    n1384,
    n1182,
    n1256,
    n1270,
    n1244
  );


  and
  g1345
  (
    n1330,
    n1091,
    n1108,
    n1168,
    n1107
  );


  xor
  g1346
  (
    n1430,
    n1082,
    n383,
    n1132,
    n1240
  );


  or
  g1347
  (
    n1481,
    n1161,
    n1242,
    n1072,
    n1208
  );


  xnor
  g1348
  (
    n1387,
    n1151,
    n1204,
    n1306,
    n1291
  );


  nor
  g1349
  (
    n1499,
    n1305,
    n1113,
    n1231,
    n1239
  );


  xnor
  g1350
  (
    n1361,
    n1243,
    n1213,
    n1166,
    n1188
  );


  or
  g1351
  (
    n1405,
    n1114,
    n1144,
    n1197,
    n1302
  );


  nor
  g1352
  (
    n1563,
    n1114,
    n1113,
    n1206,
    n1153
  );


  xor
  g1353
  (
    n1533,
    n1201,
    n1179,
    n1183,
    n1253
  );


  or
  g1354
  (
    n1391,
    n1141,
    n1174,
    n1116,
    n1086
  );


  and
  g1355
  (
    n1579,
    n1116,
    n1158,
    n1123,
    n1198
  );


  nor
  g1356
  (
    n1419,
    n1157,
    n1262,
    n1217,
    n1242
  );


  nor
  g1357
  (
    n1410,
    n1191,
    n1157,
    n1108,
    n1229
  );


  and
  g1358
  (
    n1347,
    n1199,
    n1203,
    n1118,
    n1116
  );


  nor
  g1359
  (
    n1411,
    n1201,
    n1250,
    n1135,
    n1192
  );


  xnor
  g1360
  (
    n1402,
    n1085,
    n1092,
    n1270,
    n1292
  );


  xnor
  g1361
  (
    n1462,
    n1069,
    n1094,
    n1253,
    n1087
  );


  nor
  g1362
  (
    n1385,
    n1074,
    n1219,
    n1239,
    n1184
  );


  xnor
  g1363
  (
    n1541,
    n1161,
    n1200,
    n1181,
    n1223
  );


  or
  g1364
  (
    n1498,
    n1235,
    n1088,
    n1198,
    n1077
  );


  xor
  g1365
  (
    n1336,
    n1067,
    n1084,
    n1247,
    n1121
  );


  xor
  g1366
  (
    n1475,
    n1288,
    n1146,
    n1190,
    n1278
  );


  xnor
  g1367
  (
    n1464,
    n1219,
    n1280,
    n1248,
    n1063
  );


  or
  g1368
  (
    n1508,
    n1267,
    n1131,
    n1107,
    n1268
  );


  xnor
  g1369
  (
    n1544,
    n1063,
    n1249,
    n1164,
    n1066
  );


  nand
  g1370
  (
    n1426,
    n1238,
    n1168,
    n1273,
    n1288
  );


  and
  g1371
  (
    n1474,
    n1155,
    n1208,
    n1201,
    n1083
  );


  and
  g1372
  (
    n1431,
    n1145,
    n1126,
    n1159,
    n1282
  );


  or
  g1373
  (
    n1552,
    n1219,
    n1064,
    n1274,
    n1246
  );


  nor
  g1374
  (
    n1524,
    n1242,
    n1297,
    n1102,
    n1196
  );


  nand
  g1375
  (
    n1337,
    n1090,
    n1080,
    n1194,
    n1101
  );


  and
  g1376
  (
    n1452,
    n1252,
    n1240,
    n1145,
    n384
  );


  or
  g1377
  (
    n1519,
    n1261,
    n1106,
    n1073,
    n1174
  );


  xor
  g1378
  (
    n1514,
    n1099,
    n1272,
    n1297,
    n1237
  );


  nand
  g1379
  (
    n1496,
    n1190,
    n1185,
    n1125,
    n1106
  );


  xnor
  g1380
  (
    n1458,
    n1200,
    n1241,
    n1230,
    n1216
  );


  xor
  g1381
  (
    n1509,
    n1285,
    n1120,
    n1261,
    n1138
  );


  nand
  g1382
  (
    n1550,
    n1170,
    n1194,
    n1188,
    n1183
  );


  nand
  g1383
  (
    n1392,
    n1098,
    n1269,
    n1125,
    n1102
  );


  nor
  g1384
  (
    n1517,
    n1154,
    n1192,
    n1067,
    n1107
  );


  nor
  g1385
  (
    n1569,
    n1201,
    n1133,
    n1117,
    n1247
  );


  xor
  g1386
  (
    n1513,
    n1143,
    n1179,
    n1257,
    n1076
  );


  xor
  g1387
  (
    n1463,
    n1185,
    n1066,
    n1159,
    n1182
  );


  xor
  g1388
  (
    n1368,
    n1186,
    n1206,
    n1130,
    n1235
  );


  nand
  g1389
  (
    n1369,
    n1170,
    n1230,
    n920,
    n1147
  );


  or
  g1390
  (
    n1459,
    n1303,
    n1078,
    n1113,
    n1148
  );


  xnor
  g1391
  (
    n1345,
    n1132,
    n1293,
    n1245,
    n1147
  );


  nand
  g1392
  (
    n1510,
    n1222,
    n1149,
    n1099,
    n384
  );


  and
  g1393
  (
    n1422,
    n1194,
    n1287,
    n1187,
    n1096
  );


  nor
  g1394
  (
    n1497,
    n1243,
    n1286,
    n1177,
    n1209
  );


  and
  g1395
  (
    n1441,
    n1068,
    n1291,
    n1062,
    n1224
  );


  xnor
  g1396
  (
    n1423,
    n1251,
    n1142,
    n1265,
    n1192
  );


  nor
  g1397
  (
    n1327,
    n1122,
    n1304,
    n1284,
    n1241
  );


  xor
  g1398
  (
    n1555,
    n1160,
    n1093,
    n1130,
    n1184
  );


  xnor
  g1399
  (
    n1372,
    n1286,
    n1179,
    n1080,
    n1139
  );


  xor
  g1400
  (
    n1371,
    n1149,
    n1221,
    n1156,
    n1129
  );


  or
  g1401
  (
    n1395,
    n1068,
    n1223,
    n1144,
    n1097
  );


  nand
  g1402
  (
    n1334,
    n1116,
    n1221,
    n1260,
    n1272
  );


  xor
  g1403
  (
    n1451,
    n1236,
    n1169,
    n1136,
    n1127
  );


  xor
  g1404
  (
    n1495,
    n1207,
    n1121,
    n1145,
    n1218
  );


  and
  g1405
  (
    n1364,
    n1178,
    n1112,
    n1180,
    n1195
  );


  and
  g1406
  (
    n1515,
    n1292,
    n1160,
    n1187,
    n1166
  );


  xor
  g1407
  (
    n1340,
    n1189,
    n1181,
    n1092,
    n1229
  );


  xnor
  g1408
  (
    n1348,
    n1293,
    n1072,
    n1210,
    n1105
  );


  and
  g1409
  (
    n1521,
    n1073,
    n1176,
    n1072,
    n1247
  );


  xnor
  g1410
  (
    n1388,
    n1265,
    n1249,
    n1291,
    n1119
  );


  nor
  g1411
  (
    n1446,
    n1226,
    n1276,
    n1068,
    n1193
  );


  nand
  g1412
  (
    n1359,
    n1209,
    n1141,
    n1185,
    n1132
  );


  and
  g1413
  (
    n1516,
    n1134,
    n1232,
    n1158,
    n1203
  );


  and
  g1414
  (
    n1460,
    n1101,
    n1170,
    n1139,
    n1305
  );


  nand
  g1415
  (
    n1386,
    n1274,
    n1161,
    n1259,
    n1097
  );


  and
  g1416
  (
    n1416,
    n1094,
    n1062,
    n1105,
    n1087
  );


  or
  g1417
  (
    n1370,
    n1297,
    n1062,
    n1126,
    n1230
  );


  xor
  g1418
  (
    n1434,
    n1065,
    n1182,
    n1174,
    n1271
  );


  nand
  g1419
  (
    n1341,
    n1132,
    n1158,
    n1195,
    n1060
  );


  xnor
  g1420
  (
    n1534,
    n1233,
    n1173,
    n1067,
    n1212
  );


  xor
  g1421
  (
    n1489,
    n1242,
    n1293,
    n1185,
    n1222
  );


  xor
  g1422
  (
    n1314,
    n1100,
    n1252,
    n1130
  );


  and
  g1423
  (
    n1453,
    n1146,
    n1220,
    n1258,
    n1268
  );


  nor
  g1424
  (
    n1478,
    n1115,
    n1071,
    n1255,
    n1102
  );


  and
  g1425
  (
    n1329,
    n1289,
    n1106,
    n1164,
    n1118
  );


  and
  g1426
  (
    n1354,
    n1304,
    n1103,
    n1289,
    n1251
  );


  nor
  g1427
  (
    n1535,
    n1154,
    n1191,
    n1141,
    n384
  );


  xor
  g1428
  (
    n1406,
    n1133,
    n1244,
    n1255,
    n1305
  );


  and
  g1429
  (
    n1358,
    n1220,
    n1104,
    n1163,
    n1137
  );


  and
  g1430
  (
    n1324,
    n1216,
    n1187,
    n1102,
    n1124
  );


  nand
  g1431
  (
    n1543,
    n1082,
    n1250,
    n1226,
    n1290
  );


  nor
  g1432
  (
    n1573,
    n1191,
    n1301,
    n1106,
    n1264
  );


  and
  g1433
  (
    n1491,
    n1060,
    n1183,
    n1177,
    n1202
  );


  or
  g1434
  (
    n1556,
    n1069,
    n1256,
    n1228,
    n1113
  );


  or
  g1435
  (
    n1568,
    n1120,
    n1064,
    n1247,
    n1281
  );


  nor
  g1436
  (
    n1429,
    n1159,
    n1225,
    n1117,
    n1143
  );


  xor
  g1437
  (
    n1572,
    n1141,
    n1061,
    n1212,
    n1198
  );


  and
  g1438
  (
    n1413,
    n1283,
    n1253,
    n1304,
    n1294
  );


  or
  g1439
  (
    n1420,
    n1088,
    n1290,
    n1281,
    n1162
  );


  and
  g1440
  (
    n1363,
    n1282,
    n1063,
    n1232,
    n1119
  );


  xnor
  g1441
  (
    n1378,
    n1166,
    n1135,
    n1172,
    n1296
  );


  and
  g1442
  (
    n1440,
    n1270,
    n1172,
    n1276,
    n1126
  );


  xnor
  g1443
  (
    n1318,
    n1099,
    n1264,
    n1181,
    n1169
  );


  xnor
  g1444
  (
    n1567,
    n1173,
    n1154,
    n1196,
    n1142
  );


  nand
  g1445
  (
    n1418,
    n1240,
    n1269,
    n1117,
    n1090
  );


  xor
  g1446
  (
    n1400,
    n1136,
    n1140,
    n1286,
    n1302
  );


  nor
  g1447
  (
    n1343,
    n1296,
    n1218,
    n1206,
    n1108
  );


  xnor
  g1448
  (
    n1357,
    n1150,
    n1257,
    n1228,
    n1109
  );


  nand
  g1449
  (
    n1409,
    n1124,
    n1207,
    n1233,
    n1178
  );


  nand
  g1450
  (
    n1396,
    n1177,
    n1203,
    n1301,
    n1122
  );


  nor
  g1451
  (
    n1483,
    n1287,
    n1214,
    n1199,
    n1137
  );


  xnor
  g1452
  (
    n1548,
    n1093,
    n1223,
    n1126,
    n1077
  );


  nor
  g1453
  (
    n1525,
    n1088,
    n1168,
    n1241,
    n1163
  );


  and
  g1454
  (
    n1328,
    n1092,
    n1093,
    n1303,
    n1284
  );


  or
  g1455
  (
    n1379,
    n1164,
    n1202,
    n1197,
    n1128
  );


  xnor
  g1456
  (
    n1320,
    n1302,
    n1063,
    n1271,
    n1128
  );


  xnor
  g1457
  (
    n1401,
    n1269,
    n1277,
    n1245,
    n1284
  );


  and
  g1458
  (
    n1335,
    n1204,
    n1152,
    n1138,
    n1232
  );


  or
  g1459
  (
    n1492,
    n1211,
    n1277,
    n1071,
    n1095
  );


  xor
  g1460
  (
    n1323,
    n1150,
    n1189,
    n1110,
    n1205
  );


  xnor
  g1461
  (
    n1505,
    n1145,
    n1162,
    n1200,
    n1255
  );


  or
  g1462
  (
    n1415,
    n1104,
    n1217,
    n1119,
    n1259
  );


  nor
  g1463
  (
    n1557,
    n1081,
    n1156,
    n1189,
    n1142
  );


  and
  g1464
  (
    n1450,
    n1209,
    n1073,
    n1133,
    n1293
  );


  nor
  g1465
  (
    n1528,
    n1283,
    n1085,
    n1298,
    n1266
  );


  xnor
  g1466
  (
    n1376,
    n1248,
    n1152,
    n1202,
    n1255
  );


  xor
  g1467
  (
    n1447,
    n1254,
    n1186,
    n1194,
    n1215
  );


  and
  g1468
  (
    n1536,
    n1245,
    n1300,
    n1062,
    n1152
  );


  xnor
  g1469
  (
    n1479,
    n1295,
    n1088,
    n1198,
    n1261
  );


  and
  g1470
  (
    n1578,
    n1215,
    n1306,
    n1081,
    n1281
  );


  nand
  g1471
  (
    n1351,
    n1135,
    n1288,
    n1292,
    n1127
  );


  nor
  g1472
  (
    n1381,
    n1103,
    n1290,
    n1060,
    n1154
  );


  xor
  g1473
  (
    n1399,
    n1075,
    n1273,
    n1224,
    n1290
  );


  xor
  g1474
  (
    KeyWire_0_21,
    n1258,
    n1285,
    n1262,
    n1212
  );


  xnor
  g1475
  (
    n1353,
    n1221,
    n1268,
    n1096,
    n1231
  );


  xor
  g1476
  (
    n1331,
    n1301,
    n1105,
    n1134,
    n1171
  );


  xnor
  g1477
  (
    n1490,
    n1146,
    n1238,
    n1218,
    n1119
  );


  and
  g1478
  (
    n1575,
    n1220,
    n1172,
    n1083,
    n1264
  );


  nand
  g1479
  (
    n1317,
    n1139,
    n1094,
    n1144,
    n1272
  );


  nor
  g1480
  (
    n1546,
    n1279,
    n1115,
    n1140,
    n1081
  );


  nand
  g1481
  (
    n1407,
    n1259,
    n1233,
    n1164,
    n1235
  );


  xor
  g1482
  (
    n1504,
    n1280,
    n1060,
    n1263,
    n1298
  );


  nand
  g1483
  (
    n1383,
    n1279,
    n1248,
    n1305,
    n1299
  );


  nand
  g1484
  (
    n1472,
    n1147,
    n1279,
    n1123,
    n1121
  );


  xor
  g1485
  (
    n1365,
    n1153,
    n1208,
    n1143,
    n1176
  );


  nand
  g1486
  (
    n1468,
    n1173,
    n1167,
    n1128,
    n1289
  );


  nand
  g1487
  (
    n1346,
    n1069,
    n1289,
    n1210,
    n1082
  );


  nand
  g1488
  (
    n1560,
    n1216,
    n1098,
    n1101,
    n1072
  );


  nor
  g1489
  (
    n1375,
    n1226,
    n1188,
    n1239,
    n1285
  );


  nand
  g1490
  (
    n1456,
    n1100,
    n1219,
    n1083,
    n1065
  );


  xnor
  g1491
  (
    n1487,
    n1112,
    n1296,
    n1122,
    n1103
  );


  xor
  g1492
  (
    n1316,
    n1275,
    n1148,
    n1108,
    n1224
  );


  xnor
  g1493
  (
    n1571,
    n1282,
    n1267,
    n1263,
    n1103
  );


  nand
  g1494
  (
    n1344,
    n1187,
    n1160,
    n1275,
    n1251
  );


  or
  g1495
  (
    n1356,
    n1061,
    n1155,
    n1086,
    n1204
  );


  or
  g1496
  (
    n1530,
    n1171,
    n1077,
    n1061,
    n1097
  );


  and
  g1497
  (
    n1482,
    n1234,
    n1131,
    n1080,
    n1158
  );


  nor
  g1498
  (
    n1564,
    n1249,
    n1186,
    n1180,
    n1184
  );


  or
  g1499
  (
    n1520,
    n1211,
    n1165,
    n1246
  );


  and
  g1500
  (
    n1439,
    n1097,
    n1134,
    n1171,
    n1176
  );


  xnor
  g1501
  (
    n1325,
    n1120,
    n1076,
    n1095,
    n1083
  );


  nand
  g1502
  (
    n1484,
    n1079,
    n1214,
    n1127,
    n1236
  );


  xor
  g1503
  (
    n1465,
    n1246,
    n1155,
    n1100,
    n1257
  );


  or
  g1504
  (
    n1454,
    n1221,
    n1157,
    n1193,
    n1111
  );


  xor
  g1505
  (
    n1570,
    n1175,
    n1273,
    n1098,
    n1066
  );


  xnor
  g1506
  (
    n1537,
    n1225,
    n1298,
    n1281,
    n1278
  );


  nor
  g1507
  (
    n1577,
    n1078,
    n1292,
    n1254,
    n1216
  );


  xor
  g1508
  (
    n1473,
    n1095,
    n1266,
    n1124,
    n384
  );


  xor
  g1509
  (
    n1551,
    n1114,
    n1295,
    n1213,
    n1250
  );


  xnor
  g1510
  (
    n1339,
    n1095,
    n1110,
    n1299,
    n1303
  );


  and
  g1511
  (
    n1432,
    n1271,
    n1210,
    n1122,
    n1278
  );


  xor
  g1512
  (
    n1485,
    n1208,
    n1197,
    n1260,
    n1212
  );


  xnor
  g1513
  (
    n1502,
    n1199,
    n1090,
    n1174,
    n1282
  );


  nand
  g1514
  (
    n1312,
    n1193,
    n1096,
    n1205,
    n1118
  );


  xor
  g1515
  (
    n1428,
    n1176,
    n1294,
    n1093,
    n1267
  );


  nor
  g1516
  (
    n1374,
    n1087,
    n1301,
    n1206,
    n1250
  );


  and
  g1517
  (
    n1367,
    n1195,
    n1085,
    n1104,
    n1092
  );


  xnor
  g1518
  (
    n1377,
    n1191,
    n383,
    n1243,
    n1294
  );


  nand
  g1519
  (
    n1310,
    n1150,
    n1104,
    n1233,
    n1236
  );


  nand
  g1520
  (
    n1574,
    n1205,
    n1294,
    n1125,
    n1175
  );


  or
  g1521
  (
    n1488,
    n1139,
    n1075,
    n1178
  );


  xor
  g1522
  (
    n1486,
    n1079,
    n1115,
    n1225,
    n1193
  );


  nand
  g1523
  (
    n1566,
    n1214,
    n1209,
    n1112,
    n1136
  );


  nor
  g1524
  (
    n1494,
    n1175,
    n1148,
    n1064,
    n1149
  );


  nor
  g1525
  (
    n1480,
    n1172,
    n1278,
    n1207,
    n1265
  );


  xnor
  g1526
  (
    n1442,
    n1222,
    n1086,
    n1071,
    n1295
  );


  nor
  g1527
  (
    n1417,
    n1232,
    n1091,
    n1184,
    n1169
  );


  or
  g1528
  (
    n1373,
    n1069,
    n1229,
    n1276,
    n1160
  );


  nand
  g1529
  (
    n1477,
    n1214,
    n1267,
    n1115,
    n1117
  );


  nand
  g1530
  (
    n1338,
    n1190,
    n1286,
    n1182,
    n1169
  );


  nand
  g1531
  (
    n1403,
    n1190,
    n1142,
    n1306,
    n1155
  );


  nor
  g1532
  (
    n1527,
    n1070,
    n1073,
    n1303,
    n1131
  );


  and
  g1533
  (
    n1512,
    n1234,
    n1227,
    n1084,
    n1153
  );


  xor
  g1534
  (
    n1565,
    n1188,
    n1186,
    n1251,
    n1291
  );


  nand
  g1535
  (
    n1414,
    n1081,
    n1070,
    n1170,
    n1280
  );


  and
  g1536
  (
    n1448,
    n1254,
    n1082,
    n1256,
    n1167
  );


  nor
  g1537
  (
    n1576,
    n1168,
    n1076,
    n1130,
    n1275
  );


  and
  g1538
  (
    n1444,
    n1179,
    n1269,
    n1151,
    n1065
  );


  nand
  g1539
  (
    n1443,
    n1238,
    n1202,
    n1304,
    n1273
  );


  nand
  g1540
  (
    n1437,
    n1129,
    n1227,
    n1189,
    n1077
  );


  or
  g1541
  (
    n1408,
    n1228,
    n1149,
    n1231,
    n1265
  );


  and
  g1542
  (
    n1522,
    n1270,
    n1143,
    n1110,
    n1306
  );


  xor
  g1543
  (
    n1352,
    n1275,
    n1140,
    n1248,
    n1171
  );


  xor
  g1544
  (
    n1390,
    n1259,
    n1074,
    n1129,
    n1204
  );


  xor
  g1545
  (
    n1466,
    n1111,
    n1111,
    n1211,
    n1217
  );


  and
  g1546
  (
    n1425,
    n1061,
    n1070,
    n1166,
    n1224
  );


  xnor
  g1547
  (
    n1547,
    n1178,
    n1239,
    n1296,
    n1105
  );


  or
  g1548
  (
    KeyWire_0_0,
    n1299,
    n1163,
    n1064,
    n1089
  );


  xnor
  g1549
  (
    n1349,
    n1162,
    n1089,
    n1300,
    n1085
  );


  xnor
  g1550
  (
    n1561,
    n1091,
    n1262,
    n1229,
    n1237
  );


  xor
  g1551
  (
    KeyWire_0_16,
    n1222,
    n1203,
    n1100,
    n1210
  );


  xor
  g1552
  (
    n1500,
    n1101,
    n1266,
    n1207,
    n1078
  );


  and
  g1553
  (
    n1744,
    n1374,
    n1329,
    n1424,
    n1332
  );


  xor
  g1554
  (
    n1800,
    n1534,
    n1578,
    n1438,
    n1511
  );


  xnor
  g1555
  (
    n1630,
    n1481,
    n1350,
    n1508,
    n1392
  );


  xnor
  g1556
  (
    n1634,
    n1500,
    n890,
    n574,
    n1501
  );


  and
  g1557
  (
    n1819,
    n1430,
    n1347,
    n1441,
    n1449
  );


  nor
  g1558
  (
    n1802,
    n573,
    n1359,
    n1532,
    n1500
  );


  or
  g1559
  (
    n1769,
    n1566,
    n1491,
    n1324,
    n1490
  );


  nand
  g1560
  (
    n1623,
    n1460,
    n1351,
    n1572,
    n1493
  );


  nand
  g1561
  (
    n1659,
    n1518,
    n837,
    n1407,
    n932
  );


  xor
  g1562
  (
    n1696,
    n1473,
    n1570,
    n1482,
    n1438
  );


  xnor
  g1563
  (
    n1700,
    n1313,
    n1440,
    n1348,
    n1373
  );


  and
  g1564
  (
    n1821,
    n1533,
    n1308,
    n1340,
    n1422
  );


  nand
  g1565
  (
    n1805,
    n1318,
    n1493,
    n1484,
    n1540
  );


  xor
  g1566
  (
    n1589,
    n1377,
    n1570,
    n1453,
    n1360
  );


  and
  g1567
  (
    n1711,
    n1426,
    n1525,
    n1326,
    n1370
  );


  or
  g1568
  (
    n1799,
    n1567,
    n1307,
    n1527,
    n1543
  );


  or
  g1569
  (
    n1772,
    n1519,
    n1413,
    n1456,
    n1327
  );


  nor
  g1570
  (
    n1703,
    n1525,
    n1472,
    n1452,
    n1446
  );


  nor
  g1571
  (
    n1639,
    n1358,
    n1466,
    n1387
  );


  xnor
  g1572
  (
    n1822,
    n1498,
    n1353,
    n1496,
    n1394
  );


  or
  g1573
  (
    n1682,
    n1322,
    n1501,
    n1314,
    n890
  );


  nor
  g1574
  (
    n1732,
    n576,
    n890,
    n1390,
    n1448
  );


  xnor
  g1575
  (
    n1752,
    n1469,
    n1368,
    n896,
    n1369
  );


  xor
  g1576
  (
    n1653,
    n1423,
    n1523,
    n1417,
    n1421
  );


  nor
  g1577
  (
    n1719,
    n1330,
    n1450,
    n1492,
    n1478
  );


  xor
  g1578
  (
    n1833,
    n1401,
    n1409,
    n1382,
    n933
  );


  xor
  g1579
  (
    n1867,
    n1569,
    n1416,
    n1323,
    n1499
  );


  nand
  g1580
  (
    n1811,
    n1336,
    n1376,
    n1484,
    n1451
  );


  nand
  g1581
  (
    n1767,
    n932,
    n1523,
    n1397,
    n1334
  );


  xnor
  g1582
  (
    n1644,
    n1507,
    n1371,
    n1419,
    n891
  );


  xnor
  g1583
  (
    n1793,
    n1402,
    n1366,
    n1417,
    n1437
  );


  and
  g1584
  (
    n1681,
    n1561,
    n1313,
    n1444,
    n1550
  );


  xor
  g1585
  (
    n1585,
    n1392,
    n1479,
    n1476,
    n891
  );


  and
  g1586
  (
    n1725,
    n1308,
    n1543,
    n1314,
    n892
  );


  and
  g1587
  (
    n1824,
    n1437,
    n1515,
    n1520,
    n572
  );


  xnor
  g1588
  (
    n1771,
    n1309,
    n1436,
    n1535,
    n1392
  );


  xnor
  g1589
  (
    n1607,
    n1388,
    n1429,
    n1484,
    n1332
  );


  or
  g1590
  (
    n1704,
    n1561,
    n1367,
    n1320,
    n1509
  );


  xnor
  g1591
  (
    n1794,
    n1447,
    n1512,
    n1548,
    n1483
  );


  nor
  g1592
  (
    n1587,
    n1557,
    n1521,
    n1549,
    n1314
  );


  xor
  g1593
  (
    n1816,
    n1324,
    n1517,
    n1572,
    n1328
  );


  nand
  g1594
  (
    n1830,
    n1506,
    n1446,
    n1386,
    n1518
  );


  xnor
  g1595
  (
    n1803,
    n1550,
    n1488,
    n1532,
    n1377
  );


  nand
  g1596
  (
    n1736,
    n1490,
    n1375,
    n1355,
    n1465
  );


  nor
  g1597
  (
    n1746,
    n1481,
    n1559,
    n1431,
    n1429
  );


  and
  g1598
  (
    n1668,
    n894,
    n1308,
    n1465,
    n1505
  );


  nor
  g1599
  (
    n1810,
    n1434,
    n1530,
    n1546,
    n1459
  );


  nor
  g1600
  (
    n1633,
    n1551,
    n1509,
    n1526,
    n1530
  );


  and
  g1601
  (
    n1707,
    n1552,
    n1533,
    n1372,
    n895
  );


  nand
  g1602
  (
    n1602,
    n1500,
    n1382,
    n1528,
    n1345
  );


  xnor
  g1603
  (
    n1597,
    n1390,
    n1424,
    n1391,
    n892
  );


  nand
  g1604
  (
    n1678,
    n1382,
    n1495,
    n1497,
    n1578
  );


  nor
  g1605
  (
    n1795,
    n1361,
    n1502,
    n1523,
    n1407
  );


  xnor
  g1606
  (
    n1599,
    n1312,
    n1462,
    n578,
    n1424
  );


  nor
  g1607
  (
    n1658,
    n1346,
    n1411,
    n1486,
    n1525
  );


  and
  g1608
  (
    n1777,
    n1439,
    n1410,
    n1375
  );


  or
  g1609
  (
    n1642,
    n1362,
    n1552,
    n1535,
    n1517
  );


  and
  g1610
  (
    n1825,
    n1399,
    n1326,
    n1475,
    n1565
  );


  and
  g1611
  (
    n1685,
    n1348,
    n1376,
    n1488,
    n1455
  );


  xnor
  g1612
  (
    n1701,
    n578,
    n1477,
    n1514,
    n1329
  );


  nand
  g1613
  (
    n1837,
    n577,
    n1389,
    n1350,
    n1548
  );


  xor
  g1614
  (
    n1817,
    n1337,
    n1510,
    n1328,
    n1420
  );


  nand
  g1615
  (
    n1868,
    n1359,
    n1445,
    n1497,
    n1381
  );


  nand
  g1616
  (
    n1806,
    n1572,
    n1348,
    n1421,
    n1442
  );


  xor
  g1617
  (
    n1665,
    n1382,
    n1344,
    n1506,
    n1557
  );


  xnor
  g1618
  (
    n1790,
    n1363,
    n1390,
    n573,
    n1564
  );


  and
  g1619
  (
    n1751,
    n1485,
    n1563,
    n1410,
    n1560
  );


  xor
  g1620
  (
    n1595,
    n1443,
    n1473,
    n574,
    n1451
  );


  nand
  g1621
  (
    n1672,
    n573,
    n1426,
    n1508,
    n1311
  );


  nor
  g1622
  (
    n1846,
    n1535,
    n1335,
    n1442,
    n1504
  );


  and
  g1623
  (
    n1600,
    n1553,
    n1474,
    n1453,
    n1457
  );


  nor
  g1624
  (
    n1737,
    n1464,
    n1403,
    n1457,
    n1566
  );


  xnor
  g1625
  (
    n1814,
    n574,
    n1432,
    n1428,
    n1423
  );


  nor
  g1626
  (
    n1712,
    n1409,
    n1487,
    n1385,
    n1448
  );


  and
  g1627
  (
    n1588,
    n1393,
    n1364,
    n1379,
    n1477
  );


  nor
  g1628
  (
    n1733,
    n1458,
    n1357,
    n1424,
    n1516
  );


  nand
  g1629
  (
    n1766,
    n1547,
    n575,
    n1387,
    n1579
  );


  xnor
  g1630
  (
    n1679,
    n1322,
    n1459,
    n1476,
    n1345
  );


  and
  g1631
  (
    n1852,
    n1500,
    n1510,
    n1356,
    n1524
  );


  nand
  g1632
  (
    n1862,
    n1313,
    n893,
    n1349,
    n1377
  );


  nand
  g1633
  (
    n1775,
    n519,
    n1349,
    n1384,
    n1413
  );


  or
  g1634
  (
    n1859,
    n1445,
    n1340,
    n1425,
    n1528
  );


  or
  g1635
  (
    n1738,
    n1349,
    n1388,
    n1330,
    n1383
  );


  or
  g1636
  (
    n1845,
    n1418,
    n1434,
    n839,
    n1560
  );


  xor
  g1637
  (
    n1723,
    n1421,
    n1404,
    n1567,
    n1405
  );


  nor
  g1638
  (
    n1742,
    n892,
    n1570,
    n578,
    n1365
  );


  nor
  g1639
  (
    n1706,
    n1401,
    n1482,
    n1569,
    n1522
  );


  and
  g1640
  (
    n1680,
    n1540,
    n1557,
    n1403,
    n1561
  );


  or
  g1641
  (
    n1693,
    n1441,
    n1480,
    n1432,
    n1310
  );


  or
  g1642
  (
    n1662,
    n1438,
    n1336,
    n1341,
    n1467
  );


  xnor
  g1643
  (
    n1618,
    n1537,
    n1354,
    n1331,
    n1516
  );


  nor
  g1644
  (
    n1843,
    n1521,
    n1520,
    n1423,
    n1353
  );


  and
  g1645
  (
    n1850,
    n1319,
    n1556,
    n1413,
    n1509
  );


  nor
  g1646
  (
    n1645,
    n1354,
    n1342,
    n1571,
    n1544
  );


  or
  g1647
  (
    n1776,
    n1538,
    n1393,
    n1435,
    n1489
  );


  and
  g1648
  (
    n1643,
    n1546,
    n1351,
    n1541,
    n1448
  );


  xnor
  g1649
  (
    n1603,
    n1568,
    n575,
    n1497,
    n1474
  );


  xor
  g1650
  (
    n1605,
    n1431,
    n1434,
    n1464,
    n1456
  );


  nand
  g1651
  (
    n1606,
    n1325,
    n1449,
    n1317,
    n894
  );


  and
  g1652
  (
    n1760,
    n1519,
    n894,
    n1435,
    n1406
  );


  and
  g1653
  (
    n1783,
    n1539,
    n1475,
    n1334,
    n1573
  );


  nor
  g1654
  (
    n1650,
    n1579,
    n894,
    n1384,
    n1344
  );


  xor
  g1655
  (
    n1628,
    n1455,
    n1474,
    n896,
    n895
  );


  and
  g1656
  (
    n1646,
    n1312,
    n1487,
    n1550,
    n1386
  );


  xor
  g1657
  (
    n1781,
    n1398,
    n1323,
    n1475,
    n1449
  );


  xor
  g1658
  (
    n1652,
    n1391,
    n1537,
    n1512,
    n1576
  );


  or
  g1659
  (
    n1692,
    n1415,
    n1507,
    n1394,
    n1471
  );


  nand
  g1660
  (
    n1592,
    n1453,
    n1562,
    n1428,
    n1343
  );


  xnor
  g1661
  (
    n1861,
    n1577,
    n1464,
    n1339,
    n1377
  );


  nor
  g1662
  (
    n1609,
    n1406,
    n1451,
    n1357,
    n1474
  );


  nor
  g1663
  (
    n1834,
    n1331,
    n1502,
    n1454,
    n1340
  );


  xnor
  g1664
  (
    n1674,
    n1515,
    n1398,
    n1431,
    n1459
  );


  nor
  g1665
  (
    n1840,
    n1565,
    n1394,
    n1521,
    n1308
  );


  and
  g1666
  (
    n1581,
    n1357,
    n1491,
    n1378,
    n1526
  );


  xnor
  g1667
  (
    n1669,
    n1488,
    n1538,
    n933,
    n1460
  );


  xor
  g1668
  (
    n1582,
    n1540,
    n1476,
    n1325,
    n1549
  );


  nor
  g1669
  (
    n1677,
    n838,
    n1510,
    n1536,
    n1559
  );


  and
  g1670
  (
    n1813,
    n575,
    n1447,
    n1410,
    n1517
  );


  xor
  g1671
  (
    n1841,
    n1473,
    n1522,
    n1562,
    n1416
  );


  nand
  g1672
  (
    n1695,
    n1438,
    n1573,
    n1459,
    n893
  );


  xnor
  g1673
  (
    n1715,
    n1499,
    n1490,
    n1495,
    n1469
  );


  nor
  g1674
  (
    n1773,
    n1501,
    n1443,
    n1333,
    n1433
  );


  nor
  g1675
  (
    n1735,
    n1518,
    n1538,
    n1475,
    n1436
  );


  and
  g1676
  (
    n1670,
    n1523,
    n1454,
    n1504,
    n1565
  );


  nor
  g1677
  (
    n1747,
    n1540,
    n1462,
    n1564,
    n1575
  );


  xnor
  g1678
  (
    n1820,
    n1326,
    n1408,
    n1351,
    n1532
  );


  xnor
  g1679
  (
    n1676,
    n1338,
    n1526,
    n1473,
    n1336
  );


  xor
  g1680
  (
    n1641,
    n1396,
    n1414,
    n1397,
    n1420
  );


  xor
  g1681
  (
    n1801,
    n1502,
    n1321,
    n1339,
    n1355
  );


  and
  g1682
  (
    n1762,
    n1490,
    n1564,
    n1310,
    n1361
  );


  xor
  g1683
  (
    n1717,
    n1427,
    n1419,
    n1343,
    n1526
  );


  nand
  g1684
  (
    n1694,
    n1573,
    n1384,
    n1560,
    n1546
  );


  nand
  g1685
  (
    n1750,
    n1543,
    n1361,
    n1320,
    n1426
  );


  and
  g1686
  (
    n1656,
    n1577,
    n1368,
    n1451,
    n1567
  );


  and
  g1687
  (
    n1661,
    n838,
    n1342,
    n1461,
    n1419
  );


  xnor
  g1688
  (
    n1763,
    n1409,
    n1393,
    n1310,
    n578
  );


  and
  g1689
  (
    n1815,
    n1449,
    n1436,
    n1485,
    n1497
  );


  nor
  g1690
  (
    n1624,
    n1531,
    n1483,
    n1560,
    n573
  );


  and
  g1691
  (
    n1727,
    n1338,
    n1486,
    n1427,
    n1533
  );


  and
  g1692
  (
    n1586,
    n1503,
    n1575,
    n1541,
    n1524
  );


  nor
  g1693
  (
    n1853,
    n1452,
    n1386,
    n1539,
    n1553
  );


  or
  g1694
  (
    KeyWire_0_17,
    n1319,
    n1458,
    n1554,
    n1568
  );


  nor
  g1695
  (
    n1686,
    n1481,
    n1381,
    n1426,
    n1374
  );


  nor
  g1696
  (
    n1621,
    n1326,
    n1576,
    n1470,
    n1555
  );


  xor
  g1697
  (
    n1590,
    n1487,
    n895,
    n1368,
    n1317
  );


  xnor
  g1698
  (
    n1691,
    n1408,
    n1528,
    n1323,
    n1516
  );


  and
  g1699
  (
    n1828,
    n1579,
    n1401,
    n1416,
    n1362
  );


  or
  g1700
  (
    n1739,
    n1492,
    n1360,
    n1430,
    n1354
  );


  and
  g1701
  (
    n1774,
    n1576,
    n1480,
    n1339,
    n1341
  );


  nor
  g1702
  (
    n1856,
    n1470,
    n1322,
    n895,
    n1339
  );


  nand
  g1703
  (
    n1638,
    n1443,
    n1551,
    n1318,
    n1324
  );


  and
  g1704
  (
    n1864,
    n1328,
    n1385,
    n1374,
    n1536
  );


  xor
  g1705
  (
    n1870,
    n1343,
    n1415,
    n1376,
    n1528
  );


  or
  g1706
  (
    n1710,
    n1446,
    n1442,
    n838,
    n1435
  );


  and
  g1707
  (
    n1610,
    n1401,
    n1409,
    n1360,
    n1547
  );


  xnor
  g1708
  (
    n1619,
    n1338,
    n1389,
    n1317,
    n1513
  );


  nor
  g1709
  (
    n1847,
    n1489,
    n1520,
    n1579,
    n1388
  );


  xor
  g1710
  (
    n1797,
    n1411,
    n1463,
    n1545,
    n1309
  );


  or
  g1711
  (
    n1616,
    n1414,
    n1545,
    n1566,
    n1494
  );


  xor
  g1712
  (
    n1629,
    n1332,
    n1316,
    n574,
    n1445
  );


  xnor
  g1713
  (
    n1855,
    n1545,
    n1400,
    n1392,
    n1467
  );


  and
  g1714
  (
    n1756,
    n1364,
    n1519,
    n1422,
    n1335
  );


  xnor
  g1715
  (
    n1611,
    n1408,
    n1538,
    n1492,
    n1372
  );


  or
  g1716
  (
    n1731,
    n1544,
    n1469,
    n1563,
    n1455
  );


  xor
  g1717
  (
    n1649,
    n1399,
    n1320,
    n1334,
    n1380
  );


  and
  g1718
  (
    n1689,
    n1429,
    n1450,
    n1327,
    n1547
  );


  nand
  g1719
  (
    n1831,
    n1327,
    n1376,
    n572,
    n1406
  );


  or
  g1720
  (
    n1614,
    n1329,
    n1551,
    n1525,
    n1548
  );


  xor
  g1721
  (
    n1789,
    n1330,
    n1468,
    n576,
    n1553
  );


  nor
  g1722
  (
    n1697,
    n1390,
    n1350,
    n1577,
    n1503
  );


  nand
  g1723
  (
    n1858,
    n1346,
    n1552,
    n1406,
    n1405
  );


  xor
  g1724
  (
    n1613,
    n1330,
    n1356,
    n1333,
    n1443
  );


  nor
  g1725
  (
    n1748,
    n1373,
    n1555,
    n1558,
    n893
  );


  and
  g1726
  (
    n1709,
    n839,
    n1539,
    n1468,
    n1574
  );


  or
  g1727
  (
    n1796,
    n1437,
    n1345,
    n1395
  );


  xor
  g1728
  (
    n1730,
    n1558,
    n1378,
    n1435,
    n1367
  );


  xor
  g1729
  (
    n1758,
    n1562,
    n1463,
    n1324,
    n1461
  );


  or
  g1730
  (
    n1836,
    n1428,
    n1384,
    n1466,
    n1472
  );


  or
  g1731
  (
    n1713,
    n1353,
    n1400,
    n1335,
    n1450
  );


  or
  g1732
  (
    n1596,
    n1344,
    n1379,
    n1369,
    n1458
  );


  or
  g1733
  (
    n1604,
    n1387,
    n1554,
    n1405,
    n1454
  );


  nand
  g1734
  (
    n1708,
    n933,
    n1421,
    n1529,
    n1480
  );


  and
  g1735
  (
    n1625,
    n1527,
    n1489,
    n1486,
    n1547
  );


  or
  g1736
  (
    n1734,
    n1400,
    n1311,
    n1542,
    n1491
  );


  xnor
  g1737
  (
    n1749,
    n1441,
    n1457,
    n1420,
    n1439
  );


  xor
  g1738
  (
    n1770,
    n1411,
    n839,
    n1544,
    n1571
  );


  xor
  g1739
  (
    n1745,
    n576,
    n1472,
    n1517,
    n1450
  );


  or
  g1740
  (
    n1838,
    n1510,
    n1398,
    n1512,
    n1530
  );


  xnor
  g1741
  (
    n1740,
    n1337,
    n1444,
    n1504,
    n1531
  );


  nor
  g1742
  (
    n1826,
    n1371,
    n1363,
    n1375,
    n1309
  );


  or
  g1743
  (
    n1714,
    n1320,
    n1513,
    n1389,
    n1454
  );


  or
  g1744
  (
    n1648,
    n1479,
    n1425,
    n1575,
    n1358
  );


  or
  g1745
  (
    n1728,
    n577,
    n1312,
    n1403,
    n1316
  );


  nand
  g1746
  (
    n1754,
    n891,
    n1478,
    n1400,
    n1493
  );


  xor
  g1747
  (
    n1807,
    n1559,
    n1502,
    n1576,
    n1433
  );


  xor
  g1748
  (
    n1791,
    n1412,
    n1553,
    n1428,
    n1319
  );


  or
  g1749
  (
    n1808,
    n1558,
    n1356,
    n1367,
    n1552
  );


  or
  g1750
  (
    n1753,
    n1314,
    n1417,
    n1381,
    n1372
  );


  xor
  g1751
  (
    n1809,
    n1504,
    n1507,
    n1493,
    n1352
  );


  xnor
  g1752
  (
    n1617,
    n1341,
    n1506,
    n1399,
    n1350
  );


  xor
  g1753
  (
    n1743,
    n1395,
    n1312,
    n1447,
    n1534
  );


  nor
  g1754
  (
    n1835,
    n1519,
    n1429,
    n1530,
    n1568
  );


  nor
  g1755
  (
    n1779,
    n1403,
    n1422,
    n1506,
    n1571
  );


  xnor
  g1756
  (
    n1851,
    n1495,
    n1368,
    n1524,
    n1557
  );


  or
  g1757
  (
    n1675,
    n1427,
    n1397,
    n1505,
    n1344
  );


  nand
  g1758
  (
    n1726,
    n1542,
    n1532,
    n893,
    n1380
  );


  xor
  g1759
  (
    n1765,
    n1355,
    n1381,
    n1533,
    n1492
  );


  nor
  g1760
  (
    n1718,
    n1468,
    n1336,
    n1529,
    n1337
  );


  nor
  g1761
  (
    n1785,
    n1374,
    n1514,
    n1539,
    n1564
  );


  or
  g1762
  (
    n1757,
    n1542,
    n1432,
    n1531,
    n1325
  );


  xor
  g1763
  (
    n1612,
    n1555,
    n1516,
    n1534,
    n1480
  );


  and
  g1764
  (
    n1673,
    n1363,
    n1352,
    n1496,
    n572
  );


  xnor
  g1765
  (
    n1854,
    n1462,
    n1489,
    n1499,
    n1383
  );


  nand
  g1766
  (
    n1721,
    n1444,
    n1542,
    n1529,
    n1463
  );


  xnor
  g1767
  (
    n1812,
    n1361,
    n1405,
    n931,
    n1558
  );


  xnor
  g1768
  (
    n1651,
    n1496,
    n1373,
    n1575,
    n1494
  );


  or
  g1769
  (
    n1702,
    n1466,
    n1541,
    n1444,
    n1452
  );


  and
  g1770
  (
    n1844,
    n1383,
    n1570,
    n1453,
    n1520
  );


  or
  g1771
  (
    n1655,
    n1495,
    n1394,
    n932,
    n1378
  );


  xnor
  g1772
  (
    n1755,
    n1359,
    n1329,
    n1486,
    n1499
  );


  xor
  g1773
  (
    n1804,
    n1472,
    n1470,
    n1554,
    n1307
  );


  xnor
  g1774
  (
    n1663,
    n1566,
    n1476,
    n1546,
    n1549
  );


  xor
  g1775
  (
    n1705,
    n1307,
    n1574,
    n1440,
    n1358
  );


  and
  g1776
  (
    n1601,
    n1527,
    n1545,
    n1574,
    n1536
  );


  nor
  g1777
  (
    n1580,
    n1370,
    n1402,
    n1408,
    n1505
  );


  nor
  g1778
  (
    n1782,
    n1507,
    n1485,
    n1543,
    n1503
  );


  xor
  g1779
  (
    n1632,
    n1464,
    n1332,
    n1379,
    n1440
  );


  and
  g1780
  (
    n1583,
    n1346,
    n1529,
    n1511,
    n1439
  );


  and
  g1781
  (
    n1584,
    n1353,
    n1416,
    n1311,
    n1514
  );


  xor
  g1782
  (
    n1591,
    n1430,
    n1430,
    n1369,
    n1373
  );


  nor
  g1783
  (
    n1666,
    n1423,
    n1404,
    n1569
  );


  and
  g1784
  (
    n1784,
    n1563,
    n1310,
    n1315,
    n1527
  );


  xnor
  g1785
  (
    n1780,
    n1544,
    n1452,
    n1331,
    n1567
  );


  xnor
  g1786
  (
    n1827,
    n1341,
    n576,
    n1360,
    n1327
  );


  xnor
  g1787
  (
    n1626,
    n1554,
    n1561,
    n1370,
    n1508
  );


  xnor
  g1788
  (
    n1622,
    n1491,
    n1317,
    n1415,
    n1541
  );


  nand
  g1789
  (
    n1688,
    n1534,
    n1461,
    n1448,
    n1348
  );


  xor
  g1790
  (
    n1832,
    n1346,
    n1402,
    n575,
    n1549
  );


  xnor
  g1791
  (
    n1698,
    n1501,
    n1521,
    n1396,
    n1383
  );


  and
  g1792
  (
    n1741,
    n1458,
    n839,
    n1375,
    n1537
  );


  and
  g1793
  (
    n1722,
    n1334,
    n1323,
    n1465,
    n1363
  );


  or
  g1794
  (
    n1857,
    n1425,
    n1347,
    n1389
  );


  nand
  g1795
  (
    n1720,
    n1471,
    n1563,
    n1371,
    n1511
  );


  xnor
  g1796
  (
    n1863,
    n1321,
    n1387,
    n1442,
    n896
  );


  and
  g1797
  (
    n1871,
    n1439,
    n1412,
    n1407,
    n1414
  );


  and
  g1798
  (
    n1866,
    n1418,
    n1365,
    n1307,
    n890
  );


  xor
  g1799
  (
    n1839,
    n577,
    n1569,
    n1488,
    n1515
  );


  nor
  g1800
  (
    n1690,
    n1311,
    n1397,
    n1509,
    n1455
  );


  xnor
  g1801
  (
    n1860,
    n1366,
    n1469,
    n1396,
    n1367
  );


  nand
  g1802
  (
    n1654,
    n1467,
    n1573,
    n1518,
    n1372
  );


  xor
  g1803
  (
    n1684,
    n1309,
    n1366,
    n1340,
    n1440
  );


  nand
  g1804
  (
    n1823,
    n1359,
    n1402,
    n1337,
    n1522
  );


  nand
  g1805
  (
    n1627,
    n1477,
    n1577,
    n1318,
    n1333
  );


  xor
  g1806
  (
    n1593,
    n1432,
    n1418,
    n1370,
    n1524
  );


  or
  g1807
  (
    n1761,
    n1388,
    n1462,
    n1318,
    n1481
  );


  xnor
  g1808
  (
    n1598,
    n1380,
    n1364,
    n1537,
    n892
  );


  or
  g1809
  (
    n1667,
    n1420,
    n1498,
    n1511,
    n1419
  );


  xor
  g1810
  (
    n1786,
    n891,
    n1555,
    n1354,
    n1395
  );


  xor
  g1811
  (
    n1647,
    n1535,
    n1496,
    n1483,
    n1393
  );


  nor
  g1812
  (
    n1657,
    n1418,
    n838,
    n1559,
    n1460
  );


  nand
  g1813
  (
    n1842,
    n1556,
    n1365,
    n1471,
    n1380
  );


  nand
  g1814
  (
    n1631,
    n1494,
    n1378,
    n1562,
    n1358
  );


  and
  g1815
  (
    n1635,
    n1485,
    n1445,
    n1417,
    n1347
  );


  nand
  g1816
  (
    n1849,
    n1433,
    n1484,
    n1362,
    n1512
  );


  and
  g1817
  (
    n1594,
    n1479,
    n1513,
    n1333,
    n1508
  );


  or
  g1818
  (
    n1792,
    n1471,
    n1398,
    n1487,
    n1422
  );


  and
  g1819
  (
    n1829,
    n1433,
    n1379,
    n1391,
    n1513
  );


  or
  g1820
  (
    n1818,
    n1482,
    n1335,
    n1404,
    n1365
  );


  xnor
  g1821
  (
    n1764,
    n1470,
    n1446,
    n1321,
    n932
  );


  xnor
  g1822
  (
    n1787,
    n1436,
    n1434,
    n1571,
    n1399
  );


  and
  g1823
  (
    n1778,
    n1550,
    n1331,
    n1396,
    n1441
  );


  nor
  g1824
  (
    n1664,
    n1460,
    n1412,
    n1578,
    n1551
  );


  nand
  g1825
  (
    n1615,
    n1461,
    n1456,
    n1352,
    n1463
  );


  xor
  g1826
  (
    n1788,
    n1386,
    n1356,
    n1565,
    n1556
  );


  xor
  g1827
  (
    n1636,
    n1316,
    n1322,
    n1342,
    n1531
  );


  nor
  g1828
  (
    n1683,
    n1572,
    n1574,
    n1568,
    n1415
  );


  nand
  g1829
  (
    n1865,
    n1457,
    n1315,
    n1556,
    n1316
  );


  xor
  g1830
  (
    n1699,
    n1342,
    n1395,
    n1479,
    n1548
  );


  and
  g1831
  (
    n1798,
    n1362,
    n1385,
    n1427,
    n1413
  );


  and
  g1832
  (
    n1869,
    n1351,
    n1514,
    n933,
    n1498
  );


  xnor
  g1833
  (
    n1848,
    n1468,
    n1447,
    n1425,
    n1371
  );


  nor
  g1834
  (
    n1660,
    n1522,
    n1503,
    n1391,
    n1482
  );


  or
  g1835
  (
    n1608,
    n1478,
    n1357,
    n1536,
    n1366
  );


  or
  g1836
  (
    n1716,
    n1338,
    n1505,
    n1407,
    n1321
  );


  and
  g1837
  (
    n1724,
    n1414,
    n1498,
    n1319,
    n1369
  );


  nor
  g1838
  (
    KeyWire_0_20,
    n572,
    n1349,
    n1467,
    n1355
  );


  xnor
  g1839
  (
    n1759,
    n1315,
    n1465,
    n577,
    n1412
  );


  or
  g1840
  (
    n1768,
    n1483,
    n1431,
    n1352,
    n1313
  );


  xor
  g1841
  (
    n1729,
    n1494,
    n1411,
    n1456,
    n1578
  );


  nor
  g1842
  (
    n1671,
    n1315,
    n1325,
    n1437,
    n1515
  );


  xor
  g1843
  (
    n1620,
    n1328,
    n1478,
    n896,
    n1364
  );


  xor
  g1844
  (
    n1687,
    n1385,
    n1343,
    n1477,
    n931
  );


  and
  g1845
  (
    n1895,
    n1629,
    n1620,
    n1858,
    n1733
  );


  nand
  g1846
  (
    n1947,
    n1632,
    n1818,
    n1702,
    n1787
  );


  xor
  g1847
  (
    n1880,
    n1671,
    n1738,
    n1868,
    n1743
  );


  and
  g1848
  (
    n1873,
    n1694,
    n1707,
    n1768,
    n1624
  );


  nor
  g1849
  (
    n1876,
    n1730,
    n1845,
    n1658,
    n1762
  );


  and
  g1850
  (
    n1942,
    n1710,
    n1754,
    n1667,
    n1584
  );


  nand
  g1851
  (
    n1936,
    n1831,
    n1806,
    n1808,
    n1597
  );


  and
  g1852
  (
    n1881,
    n1869,
    n1598,
    n1824,
    n1809
  );


  xor
  g1853
  (
    n1905,
    n1682,
    n1812,
    n1633,
    n1613
  );


  nor
  g1854
  (
    n1919,
    n1719,
    n1863,
    n1697,
    n1708
  );


  nand
  g1855
  (
    n1914,
    n1656,
    n1616,
    n1588,
    n1766
  );


  xor
  g1856
  (
    n1911,
    n1760,
    n1870,
    n1692,
    n1590
  );


  xor
  g1857
  (
    n1877,
    n1820,
    n1861,
    n1581,
    n1706
  );


  xnor
  g1858
  (
    n1918,
    n1592,
    n1867,
    n1735,
    n1614
  );


  xor
  g1859
  (
    n1922,
    n1783,
    n1644,
    n1746,
    n1799
  );


  xor
  g1860
  (
    n1927,
    n1777,
    n1716,
    n1744,
    n1674
  );


  or
  g1861
  (
    KeyWire_0_23,
    n1622,
    n1654,
    n1804,
    n1837
  );


  nor
  g1862
  (
    n1884,
    n1625,
    n1759,
    n1749,
    n1859
  );


  nor
  g1863
  (
    n1883,
    n1753,
    n1862,
    n1819,
    n1689
  );


  nand
  g1864
  (
    n1920,
    n1854,
    n1770,
    n1758,
    n1627
  );


  xnor
  g1865
  (
    n1916,
    n1636,
    n1803,
    n1607,
    n1615
  );


  or
  g1866
  (
    n1900,
    n1639,
    n1717,
    n1647,
    n1871
  );


  nor
  g1867
  (
    n1938,
    n1830,
    n1619,
    n1868,
    n1790
  );


  nand
  g1868
  (
    n1909,
    n1847,
    n1684,
    n1652,
    n1609
  );


  xnor
  g1869
  (
    n1890,
    n1591,
    n1792,
    n1797,
    n1839
  );


  or
  g1870
  (
    n1878,
    n1670,
    n1623,
    n1666,
    n1685
  );


  and
  g1871
  (
    n1917,
    n1763,
    n1686,
    n1649,
    n1778
  );


  or
  g1872
  (
    n1872,
    n1605,
    n1688,
    n1648,
    n1596
  );


  and
  g1873
  (
    n1925,
    n1834,
    n1829,
    n1822,
    n1860
  );


  xor
  g1874
  (
    n1886,
    n1608,
    n1638,
    n1755,
    n1793
  );


  nor
  g1875
  (
    n1875,
    n1864,
    n1813,
    n1828,
    n1791
  );


  xor
  g1876
  (
    n1906,
    n1736,
    n1677,
    n1725,
    n1861
  );


  nand
  g1877
  (
    n1929,
    n1678,
    n1805,
    n1765,
    n1798
  );


  xnor
  g1878
  (
    n1874,
    n1600,
    n1643,
    n1665,
    n1756
  );


  nand
  g1879
  (
    n1907,
    n1595,
    n1826,
    n1865,
    n1618
  );


  or
  g1880
  (
    n1926,
    n1626,
    n1860,
    n1673,
    n1601
  );


  or
  g1881
  (
    n1894,
    n1723,
    n1764,
    n1724,
    n1767
  );


  nand
  g1882
  (
    n1932,
    n1659,
    n1720,
    n1850,
    n1796
  );


  nand
  g1883
  (
    n1891,
    n1788,
    n1705,
    n1664,
    n1711
  );


  xor
  g1884
  (
    n1892,
    n1775,
    n1780,
    n1662,
    n1641
  );


  xor
  g1885
  (
    n1928,
    n1864,
    n1807,
    n1801,
    n1602
  );


  xnor
  g1886
  (
    n1879,
    n1811,
    n1867,
    n1739,
    n1838
  );


  nand
  g1887
  (
    n1887,
    n1630,
    n1776,
    n1851,
    n1751
  );


  and
  g1888
  (
    n1933,
    n1748,
    n1729,
    n1679,
    n1696
  );


  nor
  g1889
  (
    n1885,
    n1668,
    n1631,
    n1709,
    n1782
  );


  nor
  g1890
  (
    n1937,
    n1795,
    n1715,
    n1774,
    n1681
  );


  xnor
  g1891
  (
    n1902,
    n1842,
    n1853,
    n1810,
    n1669
  );


  or
  g1892
  (
    n1896,
    n1866,
    n1721,
    n1732,
    n1741
  );


  xnor
  g1893
  (
    n1903,
    n1683,
    n1855,
    n1701,
    n1773
  );


  xor
  g1894
  (
    n1930,
    n1712,
    n1752,
    n1769,
    n1734
  );


  xnor
  g1895
  (
    KeyWire_0_13,
    n1663,
    n1660,
    n1698,
    n1650
  );


  xor
  g1896
  (
    n1935,
    n1599,
    n1593,
    n1635,
    n1761
  );


  xor
  g1897
  (
    n1940,
    n1779,
    n1676,
    n1821,
    n1651
  );


  xnor
  g1898
  (
    n1939,
    n1825,
    n1852,
    n1589,
    n1833
  );


  xnor
  g1899
  (
    n1899,
    n1628,
    n1640,
    n1646,
    n1718
  );


  or
  g1900
  (
    n1888,
    n1750,
    n1789,
    n1675,
    n1869
  );


  xor
  g1901
  (
    n1944,
    n1841,
    n1587,
    n1781,
    n1785
  );


  or
  g1902
  (
    n1908,
    n1657,
    n1815,
    n1672,
    n1606
  );


  or
  g1903
  (
    n1941,
    n1661,
    n1604,
    n1690,
    n1863
  );


  xor
  g1904
  (
    n1934,
    n1726,
    n1827,
    n1836,
    n1642
  );


  xnor
  g1905
  (
    n1921,
    n1794,
    n1586,
    n1848,
    n1653
  );


  nor
  g1906
  (
    n1945,
    n1687,
    n1727,
    n1634,
    n1594
  );


  xor
  g1907
  (
    n1924,
    n1832,
    n1757,
    n1870,
    n1772
  );


  nand
  g1908
  (
    n1904,
    n1731,
    n1742,
    n1728,
    n1802
  );


  or
  g1909
  (
    n1912,
    n1617,
    n1645,
    n1611,
    n1699
  );


  or
  g1910
  (
    n1923,
    n1680,
    n1582,
    n1612,
    n1814
  );


  and
  g1911
  (
    n1897,
    n1722,
    n1817,
    n1691,
    n1700
  );


  xnor
  g1912
  (
    n1915,
    n1823,
    n1857,
    n1737,
    n1816
  );


  xnor
  g1913
  (
    n1913,
    n1747,
    n1637,
    n1714,
    n1703
  );


  xnor
  g1914
  (
    KeyWire_0_24,
    n1784,
    n1849,
    n1846,
    n1603
  );


  xor
  g1915
  (
    n1898,
    n1844,
    n1800,
    n1871,
    n1856
  );


  and
  g1916
  (
    n1931,
    n1695,
    n1740,
    n1693,
    n1840
  );


  or
  g1917
  (
    n1946,
    n1583,
    n1585,
    n1862,
    n1843
  );


  xor
  g1918
  (
    n1901,
    n1835,
    n1859,
    n1610,
    n1745
  );


  xnor
  g1919
  (
    n1943,
    n1865,
    n1771,
    n1621,
    n1655
  );


  and
  g1920
  (
    n1889,
    n1866,
    n1786,
    n1713,
    n1704
  );


  nor
  g1921
  (
    n1949,
    n1931,
    n1897,
    n1909,
    n1947
  );


  xor
  g1922
  (
    n1948,
    n1912,
    n1900,
    n1941,
    n1927
  );


  nor
  g1923
  (
    n1956,
    n1902,
    n1892,
    n1944,
    n1914
  );


  xnor
  g1924
  (
    n1960,
    n1946,
    n1911,
    n1913,
    n1918
  );


  nor
  g1925
  (
    n1951,
    n1926,
    n1928,
    n1878,
    n1891
  );


  and
  g1926
  (
    n1961,
    n1923,
    n1920,
    n1894,
    n1935
  );


  xor
  g1927
  (
    n1950,
    n1945,
    n1908,
    n1929,
    n1938
  );


  nor
  g1928
  (
    n1954,
    n1936,
    n1917,
    n1939,
    n1876
  );


  and
  g1929
  (
    n1957,
    n1906,
    n1919,
    n1925,
    n1903
  );


  nand
  g1930
  (
    n1962,
    n1890,
    n1880,
    n1901,
    n1887
  );


  xnor
  g1931
  (
    n1952,
    n1937,
    n1895,
    n1883,
    n1899
  );


  and
  g1932
  (
    n1964,
    n1921,
    n1874,
    n1877,
    n1943
  );


  and
  g1933
  (
    n1965,
    n1886,
    n1930,
    n1910,
    n1942
  );


  and
  g1934
  (
    n1955,
    n1873,
    n1889,
    n1924,
    n1932
  );


  or
  g1935
  (
    n1958,
    n1885,
    n1888,
    n1884,
    n1905
  );


  or
  g1936
  (
    n1963,
    n1916,
    n1904,
    n1933,
    n1881
  );


  or
  g1937
  (
    n1959,
    n1898,
    n1875,
    n1896,
    n1922
  );


  nand
  g1938
  (
    n1953,
    n1907,
    n1872,
    n1934,
    n1915
  );


  or
  g1939
  (
    n1966,
    n1940,
    n1893,
    n1882,
    n1879
  );


  xnor
  KeyGate_0_0
  (
    n1307,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n811,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n479,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n462,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n468,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1149,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n861,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1194,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1538,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n36,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n552,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n822,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n603,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1882,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n716,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1291,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1457,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1637,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n1069,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n882,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n1640,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1322,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n644,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1910,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1893,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1412,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n54,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1501,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n790,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n708,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n332,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n594,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


