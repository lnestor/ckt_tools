

module Stat_183_517
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n122,
  n171,
  n124,
  n178,
  n160,
  n125,
  n165,
  n177,
  n130,
  n208,
  n204,
  n192,
  n199,
  n203,
  n205,
  n198,
  n200,
  n197,
  n201,
  n195,
  n196,
  n209,
  n194,
  n207,
  n206,
  n202,
  n193
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n122;output n171;output n124;output n178;output n160;output n125;output n165;output n177;output n130;output n208;output n204;output n192;output n199;output n203;output n205;output n198;output n200;output n197;output n201;output n195;output n196;output n209;output n194;output n207;output n206;output n202;output n193;
  wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n123;wire n126;wire n127;wire n128;wire n129;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n161;wire n162;wire n163;wire n164;wire n166;wire n167;wire n168;wire n169;wire n170;wire n172;wire n173;wire n174;wire n175;wire n176;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyWire_0_38;wire KeyNOTWire_0_38;wire KeyWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyWire_0_42;wire KeyNOTWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyNOTWire_0_44;wire KeyWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyWire_0_48;wire KeyNOTWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyNOTWire_0_51;wire KeyWire_0_52;wire KeyNOTWire_0_52;wire KeyWire_0_53;wire KeyNOTWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyNOTWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyNOTWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyNOTWire_0_62;wire KeyWire_0_63;

  not
  g0
  (
    KeyWire_0_23,
    n8
  );


  not
  g1
  (
    KeyWire_0_53,
    n23
  );


  not
  g2
  (
    n64,
    n10
  );


  buf
  g3
  (
    n72,
    n1
  );


  buf
  g4
  (
    KeyWire_0_48,
    n17
  );


  not
  g5
  (
    n73,
    n9
  );


  not
  g6
  (
    n80,
    n14
  );


  not
  g7
  (
    n91,
    n8
  );


  buf
  g8
  (
    n77,
    n4
  );


  buf
  g9
  (
    n79,
    n19
  );


  buf
  g10
  (
    KeyWire_0_43,
    n10
  );


  not
  g11
  (
    KeyWire_0_19,
    n11
  );


  buf
  g12
  (
    n47,
    n19
  );


  not
  g13
  (
    KeyWire_0_29,
    n7
  );


  not
  g14
  (
    KeyWire_0_4,
    n5
  );


  buf
  g15
  (
    n90,
    n20
  );


  not
  g16
  (
    KeyWire_0_42,
    n4
  );


  not
  g17
  (
    n97,
    n23
  );


  not
  g18
  (
    n55,
    n7
  );


  not
  g19
  (
    n86,
    n12
  );


  not
  g20
  (
    n30,
    n3
  );


  buf
  g21
  (
    n84,
    n1
  );


  not
  g22
  (
    n70,
    n9
  );


  not
  g23
  (
    KeyWire_0_41,
    n20
  );


  buf
  g24
  (
    KeyWire_0_5,
    n13
  );


  not
  g25
  (
    n69,
    n14
  );


  not
  g26
  (
    KeyWire_0_56,
    n22
  );


  buf
  g27
  (
    n32,
    n24
  );


  not
  g28
  (
    n58,
    n6
  );


  buf
  g29
  (
    KeyWire_0_15,
    n20
  );


  not
  g30
  (
    n42,
    n2
  );


  buf
  g31
  (
    n76,
    n11
  );


  buf
  g32
  (
    n49,
    n3
  );


  buf
  g33
  (
    KeyWire_0_2,
    n16
  );


  not
  g34
  (
    KeyWire_0_45,
    n17
  );


  not
  g35
  (
    KeyWire_0_34,
    n22
  );


  not
  g36
  (
    KeyWire_0_27,
    n11
  );


  buf
  g37
  (
    n59,
    n6
  );


  buf
  g38
  (
    n33,
    n2
  );


  buf
  g39
  (
    n63,
    n5
  );


  not
  g40
  (
    n62,
    n8
  );


  not
  g41
  (
    n36,
    n14
  );


  buf
  g42
  (
    n96,
    n15
  );


  buf
  g43
  (
    KeyWire_0_44,
    n21
  );


  not
  g44
  (
    n39,
    n1
  );


  not
  g45
  (
    KeyWire_0_54,
    n6
  );


  not
  g46
  (
    n68,
    n5
  );


  not
  g47
  (
    KeyWire_0_52,
    n13
  );


  not
  g48
  (
    n44,
    n13
  );


  buf
  g49
  (
    KeyWire_0_60,
    n18
  );


  buf
  g50
  (
    n88,
    n10
  );


  buf
  g51
  (
    KeyWire_0_58,
    n7
  );


  buf
  g52
  (
    KeyWire_0_25,
    n3
  );


  buf
  g53
  (
    KeyWire_0_7,
    n4
  );


  buf
  g54
  (
    n60,
    n9
  );


  not
  g55
  (
    KeyWire_0_17,
    n18
  );


  not
  g56
  (
    n35,
    n15
  );


  buf
  g57
  (
    n48,
    n17
  );


  buf
  g58
  (
    n52,
    n16
  );


  not
  g59
  (
    n67,
    n23
  );


  buf
  g60
  (
    KeyWire_0_1,
    n16
  );


  buf
  g61
  (
    n95,
    n18
  );


  buf
  g62
  (
    n89,
    n15
  );


  buf
  g63
  (
    n82,
    n12
  );


  not
  g64
  (
    n98,
    n21
  );


  buf
  g65
  (
    n81,
    n12
  );


  buf
  g66
  (
    n31,
    n24
  );


  buf
  g67
  (
    n46,
    n2
  );


  not
  g68
  (
    KeyWire_0_57,
    n22
  );


  not
  g69
  (
    n94,
    n21
  );


  not
  g70
  (
    n93,
    n24
  );


  buf
  g71
  (
    n85,
    n19
  );


  not
  g72
  (
    n109,
    n30
  );


  not
  g73
  (
    n110,
    n29
  );


  not
  g74
  (
    KeyWire_0_11,
    n33
  );


  buf
  g75
  (
    n106,
    n34
  );


  buf
  g76
  (
    n115,
    n31
  );


  not
  g77
  (
    n118,
    n26
  );


  not
  g78
  (
    n108,
    n28
  );


  buf
  g79
  (
    n119,
    n27
  );


  not
  g80
  (
    KeyWire_0_37,
    n25
  );


  not
  g81
  (
    n107,
    n30
  );


  not
  g82
  (
    KeyWire_0_12,
    n26
  );


  buf
  g83
  (
    n105,
    n26
  );


  buf
  g84
  (
    KeyWire_0_9,
    n29
  );


  buf
  g85
  (
    n120,
    n25
  );


  buf
  g86
  (
    n100,
    n31
  );


  not
  g87
  (
    KeyWire_0_51,
    n32
  );


  buf
  g88
  (
    n101,
    n27
  );


  buf
  g89
  (
    n117,
    n31
  );


  buf
  g90
  (
    n103,
    n33
  );


  buf
  g91
  (
    KeyWire_0_63,
    n32
  );


  xnor
  g92
  (
    KeyWire_0_3,
    n30,
    n27,
    n32,
    n28
  );


  nor
  g93
  (
    n113,
    n33,
    n28,
    n25,
    n29
  );


  and
  g94
  (
    n128,
    n49,
    n116,
    n95
  );


  or
  g95
  (
    KeyWire_0_13,
    n42,
    n94,
    n113,
    n107
  );


  or
  g96
  (
    n160,
    n51,
    n69,
    n100,
    n60
  );


  or
  g97
  (
    n138,
    n83,
    n60,
    n79,
    n42
  );


  xnor
  g98
  (
    KeyWire_0_40,
    n61,
    n66,
    n79,
    n56
  );


  nor
  g99
  (
    KeyWire_0_14,
    n79,
    n94,
    n103,
    n73
  );


  and
  g100
  (
    KeyWire_0_26,
    n82,
    n86,
    n109,
    n93
  );


  nor
  g101
  (
    n137,
    n50,
    n72,
    n41,
    n45
  );


  xor
  g102
  (
    n124,
    n51,
    n55,
    n57,
    n117
  );


  nand
  g103
  (
    KeyWire_0_38,
    n104,
    n108,
    n77,
    n41
  );


  nand
  g104
  (
    KeyWire_0_16,
    n72,
    n54,
    n53,
    n47
  );


  nor
  g105
  (
    n184,
    n43,
    n48,
    n40,
    n117
  );


  and
  g106
  (
    n182,
    n62,
    n80,
    n53,
    n82
  );


  xnor
  g107
  (
    KeyWire_0_46,
    n113,
    n85,
    n64,
    n115
  );


  xor
  g108
  (
    n125,
    n36,
    n72,
    n78,
    n89
  );


  or
  g109
  (
    KeyWire_0_18,
    n81,
    n82,
    n69,
    n84
  );


  xor
  g110
  (
    n172,
    n46,
    n114,
    n115,
    n108
  );


  or
  g111
  (
    n122,
    n77,
    n68,
    n80,
    n78
  );


  and
  g112
  (
    n139,
    n50,
    n43,
    n99,
    n68
  );


  and
  g113
  (
    n157,
    n93,
    n110,
    n100,
    n92
  );


  nand
  g114
  (
    n135,
    n87,
    n88,
    n71,
    n99
  );


  or
  g115
  (
    n156,
    n86,
    n111,
    n87,
    n73
  );


  and
  g116
  (
    n178,
    n96,
    n76,
    n36,
    n52
  );


  nor
  g117
  (
    KeyWire_0_49,
    n100,
    n38,
    n92,
    n34
  );


  xor
  g118
  (
    n153,
    n112,
    n93,
    n47,
    n89
  );


  or
  g119
  (
    KeyWire_0_30,
    n103,
    n58,
    n88,
    n85
  );


  xnor
  g120
  (
    KeyWire_0_61,
    n112,
    n96,
    n75,
    n99
  );


  or
  g121
  (
    n162,
    n83,
    n49,
    n67,
    n35
  );


  xnor
  g122
  (
    n155,
    n101,
    n84,
    n60,
    n61
  );


  or
  g123
  (
    KeyWire_0_36,
    n103,
    n53,
    n106,
    n49
  );


  nand
  g124
  (
    n130,
    n59,
    n54,
    n62,
    n104
  );


  nand
  g125
  (
    KeyWire_0_33,
    n106,
    n107,
    n105,
    n114
  );


  nor
  g126
  (
    n133,
    n78,
    n120,
    n70,
    n59
  );


  xnor
  g127
  (
    n127,
    n68,
    n57,
    n46,
    n64
  );


  xnor
  g128
  (
    KeyWire_0_22,
    n35,
    n67,
    n76,
    n91
  );


  nor
  g129
  (
    KeyWire_0_28,
    n111,
    n39,
    n63,
    n44
  );


  xor
  g130
  (
    n123,
    n112,
    n88,
    n44,
    n38
  );


  and
  g131
  (
    n152,
    n81,
    n71,
    n111,
    n65
  );


  nor
  g132
  (
    n163,
    n74,
    n66,
    n118,
    n51
  );


  xor
  g133
  (
    KeyWire_0_62,
    n90,
    n90,
    n39,
    n84
  );


  nor
  g134
  (
    n143,
    n59,
    n104,
    n118,
    n63
  );


  nor
  g135
  (
    KeyWire_0_35,
    n108,
    n62,
    n113,
    n52
  );


  xnor
  g136
  (
    n183,
    n97,
    n87,
    n55,
    n98
  );


  nor
  g137
  (
    KeyWire_0_31,
    n58,
    n63,
    n119,
    n55
  );


  nand
  g138
  (
    n129,
    n44,
    n95,
    n98,
    n97
  );


  xor
  g139
  (
    n141,
    n102,
    n75,
    n71,
    n45
  );


  nand
  g140
  (
    KeyWire_0_39,
    n74,
    n80,
    n118,
    n101
  );


  xor
  g141
  (
    n168,
    n102,
    n95,
    n61,
    n40
  );


  or
  g142
  (
    KeyWire_0_20,
    n36,
    n57,
    n109,
    n120
  );


  xnor
  g143
  (
    KeyWire_0_21,
    n90,
    n86,
    n47,
    n117
  );


  nor
  g144
  (
    KeyWire_0_6,
    n83,
    n56,
    n75,
    n98
  );


  xnor
  g145
  (
    n131,
    n119,
    n74,
    n39,
    n69
  );


  xor
  g146
  (
    KeyWire_0_47,
    n64,
    n35,
    n38,
    n34
  );


  xor
  g147
  (
    n148,
    n107,
    n102,
    n37,
    n65
  );


  and
  g148
  (
    n176,
    n54,
    n94,
    n45,
    n89
  );


  xor
  g149
  (
    n173,
    n48,
    n110,
    n81
  );


  or
  g150
  (
    n170,
    n76,
    n97,
    n92,
    n109
  );


  or
  g151
  (
    n146,
    n91,
    n105,
    n66,
    n40
  );


  and
  g152
  (
    n174,
    n46,
    n37,
    n65,
    n77
  );


  nand
  g153
  (
    n159,
    n67,
    n50,
    n115,
    n91
  );


  and
  g154
  (
    n132,
    n114,
    n73,
    n116,
    n96
  );


  or
  g155
  (
    KeyWire_0_50,
    n58,
    n42,
    n119,
    n56
  );


  or
  g156
  (
    n161,
    n101,
    n37,
    n70,
    n106
  );


  nand
  g157
  (
    n150,
    n85,
    n105,
    n48,
    n52
  );


  nand
  g158
  (
    n167,
    n41,
    n116,
    n70,
    n43
  );


  buf
  g159
  (
    n191,
    n131
  );


  buf
  g160
  (
    n186,
    n132
  );


  buf
  g161
  (
    n190,
    n120
  );


  not
  g162
  (
    n189,
    n134
  );


  buf
  g163
  (
    n188,
    n133
  );


  or
  g164
  (
    KeyWire_0_24,
    n135,
    n130
  );


  nor
  g165
  (
    KeyWire_0_8,
    n139,
    n164,
    n150,
    n191
  );


  nand
  g166
  (
    n208,
    n190,
    n143,
    n159,
    n191
  );


  xor
  g167
  (
    KeyWire_0_0,
    n187,
    n187,
    n144,
    n178
  );


  xor
  g168
  (
    n200,
    n176,
    n188,
    n163,
    n160
  );


  or
  g169
  (
    n194,
    n165,
    n138,
    n167,
    n181
  );


  xnor
  g170
  (
    KeyWire_0_55,
    n166,
    n189,
    n171,
    n186
  );


  nor
  g171
  (
    n207,
    n172,
    n157,
    n151,
    n174
  );


  or
  g172
  (
    KeyWire_0_10,
    n190,
    n191,
    n185,
    n155
  );


  nor
  g173
  (
    n205,
    n187,
    n145,
    n190,
    n149
  );


  or
  g174
  (
    n201,
    n189,
    n185,
    n175,
    n156
  );


  xor
  g175
  (
    KeyWire_0_59,
    n148,
    n184,
    n146
  );


  or
  g176
  (
    n203,
    n140,
    n185,
    n162,
    n137
  );


  nand
  g177
  (
    n197,
    n184,
    n189,
    n186,
    n153
  );


  nor
  g178
  (
    KeyWire_0_32,
    n173,
    n169,
    n186,
    n161
  );


  xor
  g179
  (
    n196,
    n188,
    n136,
    n147,
    n177
  );


  xor
  g180
  (
    n204,
    n179,
    n142,
    n141,
    n154
  );


  or
  g181
  (
    n199,
    n158,
    n182,
    n170,
    n152
  );


  nor
  g182
  (
    n193,
    n168,
    n188,
    n183,
    n180
  );


  xnor
  KeyGate_0_0
  (
    n195,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n75,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n83,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n116,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n37,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n66,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n136,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n43,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n206,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n102,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n209,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n111,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n99,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n142,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n147,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n53,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n126,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n51,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n134,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n57,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n121,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n185,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n165,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n54,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n187,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n45,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n151,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n38,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n164,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n50,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n175,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n180,
    keyIn_0_31,
    KeyWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n192,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n144,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n40,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n140,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n145,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n114,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n179,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n181,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n149,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n78,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n41,
    KeyNOTWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n56,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n87,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    n92,
    keyIn_0_45,
    KeyWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n158,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n177,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n28,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n171,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n154,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n104,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n27,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n61,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n29,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n198,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n71,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n65,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n34,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n202,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n74,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n166,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n169,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n112,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule


