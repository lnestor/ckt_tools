

module Stat_114_49
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n130,
  n118,
  n131,
  n123,
  n115,
  n117,
  n114,
  n120,
  n128,
  n121,
  n119,
  n126,
  n129,
  n124,
  n116,
  n125,
  n127,
  n122,
  n113,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n130;
  output n118;
  output n131;
  output n123;
  output n115;
  output n117;
  output n114;
  output n120;
  output n128;
  output n121;
  output n119;
  output n126;
  output n129;
  output n124;
  output n116;
  output n125;
  output n127;
  output n122;
  output n113;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n32,
    n17
  );


  buf
  g1
  (
    n26,
    n7
  );


  buf
  g2
  (
    n20,
    n11
  );


  not
  g3
  (
    n24,
    n6
  );


  not
  g4
  (
    n18,
    n9
  );


  buf
  g5
  (
    n25,
    n17
  );


  buf
  g6
  (
    n23,
    n12
  );


  buf
  g7
  (
    n28,
    n15
  );


  buf
  g8
  (
    n30,
    n14
  );


  not
  g9
  (
    n35,
    n13
  );


  buf
  g10
  (
    n27,
    n10
  );


  not
  g11
  (
    n22,
    n16
  );


  buf
  g12
  (
    n34,
    n5
  );


  not
  g13
  (
    n33,
    n3
  );


  buf
  g14
  (
    n21,
    n1
  );


  buf
  g15
  (
    KeyWire_0_5,
    n4
  );


  buf
  g16
  (
    n31,
    n2
  );


  buf
  g17
  (
    n29,
    n8
  );


  not
  g18
  (
    n41,
    n31
  );


  buf
  g19
  (
    n63,
    n34
  );


  not
  g20
  (
    n43,
    n24
  );


  not
  g21
  (
    n65,
    n20
  );


  buf
  g22
  (
    n52,
    n27
  );


  not
  g23
  (
    n39,
    n35
  );


  not
  g24
  (
    KeyWire_0_4,
    n19
  );


  buf
  g25
  (
    n49,
    n26
  );


  not
  g26
  (
    n42,
    n24
  );


  buf
  g27
  (
    n45,
    n35
  );


  not
  g28
  (
    n36,
    n27
  );


  not
  g29
  (
    KeyWire_0_1,
    n29
  );


  not
  g30
  (
    n72,
    n30
  );


  buf
  g31
  (
    n50,
    n35
  );


  not
  g32
  (
    n60,
    n31
  );


  not
  g33
  (
    n70,
    n33
  );


  buf
  g34
  (
    n55,
    n22
  );


  not
  g35
  (
    n44,
    n18
  );


  not
  g36
  (
    n66,
    n29
  );


  not
  g37
  (
    n61,
    n23
  );


  not
  g38
  (
    n37,
    n22
  );


  buf
  g39
  (
    n68,
    n18
  );


  not
  g40
  (
    n40,
    n34
  );


  not
  g41
  (
    n47,
    n28
  );


  not
  g42
  (
    KeyWire_0_7,
    n34
  );


  buf
  g43
  (
    n69,
    n25
  );


  not
  g44
  (
    n38,
    n30
  );


  buf
  g45
  (
    n58,
    n20
  );


  buf
  g46
  (
    n51,
    n19
  );


  buf
  g47
  (
    n57,
    n33
  );


  buf
  g48
  (
    n73,
    n28
  );


  buf
  g49
  (
    n62,
    n23
  );


  buf
  g50
  (
    n54,
    n32
  );


  not
  g51
  (
    n46,
    n21
  );


  not
  g52
  (
    n67,
    n26
  );


  not
  g53
  (
    KeyWire_0_12,
    n21
  );


  buf
  g54
  (
    n53,
    n32
  );


  not
  g55
  (
    KeyWire_0_9,
    n25
  );


  not
  g56
  (
    n76,
    n49
  );


  not
  g57
  (
    n104,
    n68
  );


  buf
  g58
  (
    KeyWire_0_14,
    n39
  );


  buf
  g59
  (
    n107,
    n38
  );


  buf
  g60
  (
    KeyWire_0_11,
    n55
  );


  buf
  g61
  (
    n106,
    n43
  );


  not
  g62
  (
    KeyWire_0_13,
    n37
  );


  buf
  g63
  (
    n92,
    n42
  );


  buf
  g64
  (
    n90,
    n51
  );


  not
  g65
  (
    n75,
    n65
  );


  buf
  g66
  (
    n83,
    n66
  );


  not
  g67
  (
    n112,
    n60
  );


  not
  g68
  (
    n103,
    n64
  );


  buf
  g69
  (
    n91,
    n53
  );


  buf
  g70
  (
    n78,
    n69
  );


  not
  g71
  (
    n93,
    n40
  );


  buf
  g72
  (
    n97,
    n72
  );


  not
  g73
  (
    n96,
    n36
  );


  buf
  g74
  (
    n85,
    n46
  );


  buf
  g75
  (
    n98,
    n48
  );


  not
  g76
  (
    n79,
    n71
  );


  buf
  g77
  (
    n88,
    n57
  );


  buf
  g78
  (
    n105,
    n73
  );


  buf
  g79
  (
    n89,
    n58
  );


  not
  g80
  (
    n99,
    n61
  );


  buf
  g81
  (
    n101,
    n41
  );


  buf
  g82
  (
    n102,
    n54
  );


  not
  g83
  (
    n86,
    n59
  );


  not
  g84
  (
    n77,
    n52
  );


  not
  g85
  (
    n84,
    n67
  );


  not
  g86
  (
    KeyWire_0_0,
    n73
  );


  not
  g87
  (
    n80,
    n63
  );


  buf
  g88
  (
    KeyWire_0_8,
    n62
  );


  buf
  g89
  (
    n109,
    n56
  );


  buf
  g90
  (
    n82,
    n50
  );


  not
  g91
  (
    n111,
    n70
  );


  not
  g92
  (
    KeyWire_0_6,
    n44
  );


  buf
  g93
  (
    n81,
    n45
  );


  not
  g94
  (
    n95,
    n47
  );


  not
  g95
  (
    n115,
    n88
  );


  buf
  g96
  (
    n123,
    n108
  );


  not
  g97
  (
    n129,
    n107
  );


  buf
  g98
  (
    n124,
    n106
  );


  buf
  g99
  (
    n119,
    n75
  );


  buf
  g100
  (
    KeyWire_0_3,
    n100
  );


  buf
  g101
  (
    n126,
    n98
  );


  buf
  g102
  (
    n131,
    n78
  );


  not
  g103
  (
    n125,
    n82
  );


  not
  g104
  (
    KeyWire_0_2,
    n93
  );


  not
  g105
  (
    n127,
    n110
  );


  not
  g106
  (
    n121,
    n94
  );


  xnor
  g107
  (
    n116,
    n105,
    n101,
    n92
  );


  xor
  g108
  (
    n130,
    n102,
    n109,
    n87,
    n96
  );


  and
  g109
  (
    KeyWire_0_10,
    n91,
    n97,
    n77,
    n99
  );


  xor
  g110
  (
    n114,
    n80,
    n90,
    n76,
    n79
  );


  nor
  g111
  (
    n117,
    n74,
    n111,
    n95,
    n83
  );


  nand
  g112
  (
    n113,
    n81,
    n104,
    n112,
    n86
  );


  or
  g113
  (
    KeyWire_0_15,
    n84,
    n103,
    n89,
    n85
  );


  xor
  KeyGate_0_0
  (
    n110,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n48,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n120,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n128,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n64,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n19,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n108,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n56,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n87,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n59,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n118,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n74,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n71,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n94,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n100,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n122,
    KeyNOTWire_0_15
  );


endmodule

