

module Stat_3000_303
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2547,
  n2535,
  n2540,
  n2543,
  n2556,
  n2555,
  n2550,
  n2530,
  n2554,
  n2537,
  n2546,
  n2557,
  n2558,
  n2622,
  n2620,
  n2615,
  n2616,
  n2612,
  n2606,
  n2623,
  n2613,
  n2608,
  n2614,
  n2610,
  n2607,
  n2618,
  n2617,
  n2611,
  n2619,
  n3031,
  n3032,
  n3030,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n2547;
  output n2535;
  output n2540;
  output n2543;
  output n2556;
  output n2555;
  output n2550;
  output n2530;
  output n2554;
  output n2537;
  output n2546;
  output n2557;
  output n2558;
  output n2622;
  output n2620;
  output n2615;
  output n2616;
  output n2612;
  output n2606;
  output n2623;
  output n2613;
  output n2608;
  output n2614;
  output n2610;
  output n2607;
  output n2618;
  output n2617;
  output n2611;
  output n2619;
  output n3031;
  output n3032;
  output n3030;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2536;
  wire n2538;
  wire n2539;
  wire n2541;
  wire n2542;
  wire n2544;
  wire n2545;
  wire n2548;
  wire n2549;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2609;
  wire n2621;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n77,
    n12
  );


  buf
  g1
  (
    n120,
    n13
  );


  not
  g2
  (
    n111,
    n23
  );


  not
  g3
  (
    n86,
    n8
  );


  not
  g4
  (
    n75,
    n1
  );


  buf
  g5
  (
    n142,
    n6
  );


  buf
  g6
  (
    n99,
    n30
  );


  not
  g7
  (
    n54,
    n11
  );


  buf
  g8
  (
    n73,
    n11
  );


  not
  g9
  (
    n44,
    n25
  );


  not
  g10
  (
    n93,
    n24
  );


  buf
  g11
  (
    n70,
    n32
  );


  not
  g12
  (
    n82,
    n5
  );


  not
  g13
  (
    n55,
    n29
  );


  not
  g14
  (
    n38,
    n26
  );


  buf
  g15
  (
    n96,
    n2
  );


  not
  g16
  (
    n127,
    n9
  );


  not
  g17
  (
    n159,
    n4
  );


  buf
  g18
  (
    n144,
    n24
  );


  buf
  g19
  (
    n110,
    n19
  );


  not
  g20
  (
    n63,
    n24
  );


  buf
  g21
  (
    n42,
    n12
  );


  not
  g22
  (
    n89,
    n27
  );


  buf
  g23
  (
    n81,
    n16
  );


  buf
  g24
  (
    n104,
    n4
  );


  buf
  g25
  (
    n138,
    n19
  );


  not
  g26
  (
    n91,
    n5
  );


  not
  g27
  (
    n118,
    n16
  );


  buf
  g28
  (
    n98,
    n31
  );


  buf
  g29
  (
    n69,
    n12
  );


  buf
  g30
  (
    n122,
    n9
  );


  buf
  g31
  (
    n78,
    n18
  );


  buf
  g32
  (
    n43,
    n21
  );


  not
  g33
  (
    n153,
    n16
  );


  buf
  g34
  (
    n156,
    n26
  );


  not
  g35
  (
    n79,
    n2
  );


  buf
  g36
  (
    n74,
    n11
  );


  not
  g37
  (
    n76,
    n3
  );


  not
  g38
  (
    n102,
    n20
  );


  not
  g39
  (
    n45,
    n10
  );


  buf
  g40
  (
    n129,
    n8
  );


  not
  g41
  (
    KeyWire_0_8,
    n25
  );


  buf
  g42
  (
    n139,
    n6
  );


  buf
  g43
  (
    n158,
    n18
  );


  not
  g44
  (
    n67,
    n20
  );


  buf
  g45
  (
    n115,
    n12
  );


  not
  g46
  (
    n126,
    n11
  );


  not
  g47
  (
    n136,
    n4
  );


  not
  g48
  (
    n90,
    n29
  );


  buf
  g49
  (
    n57,
    n28
  );


  buf
  g50
  (
    n160,
    n29
  );


  not
  g51
  (
    n58,
    n30
  );


  buf
  g52
  (
    n152,
    n28
  );


  buf
  g53
  (
    n53,
    n13
  );


  not
  g54
  (
    n113,
    n4
  );


  not
  g55
  (
    n92,
    n23
  );


  not
  g56
  (
    n56,
    n1
  );


  not
  g57
  (
    n64,
    n15
  );


  buf
  g58
  (
    n124,
    n31
  );


  not
  g59
  (
    n140,
    n14
  );


  not
  g60
  (
    n148,
    n3
  );


  not
  g61
  (
    n59,
    n24
  );


  not
  g62
  (
    n151,
    n16
  );


  buf
  g63
  (
    n134,
    n17
  );


  buf
  g64
  (
    n123,
    n15
  );


  buf
  g65
  (
    n112,
    n14
  );


  not
  g66
  (
    n101,
    n22
  );


  not
  g67
  (
    n141,
    n9
  );


  buf
  g68
  (
    n155,
    n20
  );


  not
  g69
  (
    n71,
    n13
  );


  buf
  g70
  (
    n133,
    n28
  );


  not
  g71
  (
    n36,
    n9
  );


  not
  g72
  (
    n109,
    n22
  );


  not
  g73
  (
    n50,
    n28
  );


  buf
  g74
  (
    n150,
    n1
  );


  not
  g75
  (
    n146,
    n7
  );


  buf
  g76
  (
    n40,
    n19
  );


  not
  g77
  (
    n85,
    n23
  );


  not
  g78
  (
    n83,
    n26
  );


  not
  g79
  (
    n106,
    n6
  );


  not
  g80
  (
    n108,
    n21
  );


  not
  g81
  (
    n47,
    n10
  );


  buf
  g82
  (
    n65,
    n31
  );


  buf
  g83
  (
    n107,
    n2
  );


  not
  g84
  (
    n95,
    n8
  );


  buf
  g85
  (
    n157,
    n30
  );


  buf
  g86
  (
    n60,
    n32
  );


  not
  g87
  (
    n121,
    n30
  );


  buf
  g88
  (
    n39,
    n26
  );


  buf
  g89
  (
    n145,
    n21
  );


  buf
  g90
  (
    n52,
    n25
  );


  buf
  g91
  (
    n137,
    n27
  );


  not
  g92
  (
    n103,
    n10
  );


  buf
  g93
  (
    n66,
    n13
  );


  not
  g94
  (
    n143,
    n2
  );


  not
  g95
  (
    n149,
    n15
  );


  buf
  g96
  (
    n135,
    n22
  );


  not
  g97
  (
    n61,
    n8
  );


  not
  g98
  (
    n68,
    n15
  );


  buf
  g99
  (
    n62,
    n5
  );


  buf
  g100
  (
    n125,
    n7
  );


  buf
  g101
  (
    n72,
    n32
  );


  buf
  g102
  (
    n105,
    n14
  );


  buf
  g103
  (
    n34,
    n14
  );


  buf
  g104
  (
    n46,
    n7
  );


  buf
  g105
  (
    n87,
    n27
  );


  not
  g106
  (
    n37,
    n19
  );


  not
  g107
  (
    n51,
    n32
  );


  buf
  g108
  (
    n88,
    n17
  );


  buf
  g109
  (
    n116,
    n22
  );


  buf
  g110
  (
    n128,
    n17
  );


  not
  g111
  (
    n94,
    n1
  );


  not
  g112
  (
    n100,
    n7
  );


  buf
  g113
  (
    n33,
    n20
  );


  buf
  g114
  (
    n119,
    n18
  );


  buf
  g115
  (
    n84,
    n31
  );


  buf
  g116
  (
    n49,
    n17
  );


  not
  g117
  (
    n131,
    n29
  );


  buf
  g118
  (
    n147,
    n10
  );


  not
  g119
  (
    n114,
    n18
  );


  not
  g120
  (
    n80,
    n21
  );


  not
  g121
  (
    n154,
    n23
  );


  buf
  g122
  (
    n97,
    n27
  );


  not
  g123
  (
    n130,
    n25
  );


  buf
  g124
  (
    n48,
    n3
  );


  buf
  g125
  (
    n132,
    n5
  );


  buf
  g126
  (
    n117,
    n6
  );


  not
  g127
  (
    n41,
    n3
  );


  not
  g128
  (
    n502,
    n100
  );


  not
  g129
  (
    n519,
    n67
  );


  buf
  g130
  (
    n439,
    n66
  );


  buf
  g131
  (
    n646,
    n77
  );


  not
  g132
  (
    n433,
    n55
  );


  buf
  g133
  (
    n565,
    n144
  );


  buf
  g134
  (
    n462,
    n129
  );


  buf
  g135
  (
    n185,
    n121
  );


  not
  g136
  (
    KeyWire_0_10,
    n91
  );


  not
  g137
  (
    n541,
    n68
  );


  buf
  g138
  (
    n238,
    n112
  );


  buf
  g139
  (
    n322,
    n111
  );


  buf
  g140
  (
    n272,
    n149
  );


  buf
  g141
  (
    n212,
    n126
  );


  buf
  g142
  (
    n279,
    n156
  );


  buf
  g143
  (
    n328,
    n142
  );


  not
  g144
  (
    n177,
    n90
  );


  not
  g145
  (
    n280,
    n89
  );


  not
  g146
  (
    n299,
    n35
  );


  not
  g147
  (
    n626,
    n106
  );


  buf
  g148
  (
    n388,
    n104
  );


  not
  g149
  (
    n363,
    n116
  );


  buf
  g150
  (
    n297,
    n155
  );


  buf
  g151
  (
    n550,
    n151
  );


  buf
  g152
  (
    n513,
    n118
  );


  buf
  g153
  (
    n447,
    n47
  );


  buf
  g154
  (
    n430,
    n44
  );


  buf
  g155
  (
    n524,
    n94
  );


  not
  g156
  (
    n494,
    n113
  );


  buf
  g157
  (
    n567,
    n143
  );


  buf
  g158
  (
    n507,
    n75
  );


  buf
  g159
  (
    n469,
    n100
  );


  not
  g160
  (
    n426,
    n42
  );


  not
  g161
  (
    n618,
    n116
  );


  not
  g162
  (
    n243,
    n141
  );


  not
  g163
  (
    n351,
    n152
  );


  buf
  g164
  (
    n568,
    n158
  );


  not
  g165
  (
    n254,
    n134
  );


  not
  g166
  (
    n471,
    n69
  );


  not
  g167
  (
    n650,
    n85
  );


  buf
  g168
  (
    n558,
    n65
  );


  not
  g169
  (
    n384,
    n46
  );


  buf
  g170
  (
    n183,
    n156
  );


  not
  g171
  (
    n162,
    n57
  );


  buf
  g172
  (
    n395,
    n119
  );


  not
  g173
  (
    n429,
    n131
  );


  not
  g174
  (
    n544,
    n88
  );


  not
  g175
  (
    n509,
    n101
  );


  not
  g176
  (
    n308,
    n39
  );


  buf
  g177
  (
    n397,
    n72
  );


  not
  g178
  (
    n521,
    n112
  );


  not
  g179
  (
    n240,
    n151
  );


  buf
  g180
  (
    n444,
    n48
  );


  not
  g181
  (
    n383,
    n70
  );


  not
  g182
  (
    n540,
    n119
  );


  buf
  g183
  (
    KeyWire_0_0,
    n109
  );


  buf
  g184
  (
    KeyWire_0_7,
    n139
  );


  not
  g185
  (
    n459,
    n50
  );


  not
  g186
  (
    n312,
    n133
  );


  buf
  g187
  (
    n520,
    n36
  );


  not
  g188
  (
    n233,
    n60
  );


  buf
  g189
  (
    n579,
    n65
  );


  buf
  g190
  (
    n268,
    n95
  );


  buf
  g191
  (
    n294,
    n138
  );


  buf
  g192
  (
    n659,
    n90
  );


  buf
  g193
  (
    n473,
    n81
  );


  not
  g194
  (
    n636,
    n130
  );


  buf
  g195
  (
    n499,
    n134
  );


  not
  g196
  (
    n249,
    n108
  );


  buf
  g197
  (
    n324,
    n158
  );


  buf
  g198
  (
    n493,
    n140
  );


  buf
  g199
  (
    n236,
    n117
  );


  not
  g200
  (
    n203,
    n60
  );


  buf
  g201
  (
    n518,
    n96
  );


  buf
  g202
  (
    n464,
    n56
  );


  not
  g203
  (
    n375,
    n159
  );


  not
  g204
  (
    n194,
    n101
  );


  buf
  g205
  (
    n653,
    n51
  );


  not
  g206
  (
    n581,
    n51
  );


  buf
  g207
  (
    n370,
    n123
  );


  buf
  g208
  (
    n246,
    n49
  );


  not
  g209
  (
    n443,
    n152
  );


  buf
  g210
  (
    n537,
    n72
  );


  buf
  g211
  (
    n169,
    n147
  );


  buf
  g212
  (
    n605,
    n96
  );


  not
  g213
  (
    n197,
    n126
  );


  buf
  g214
  (
    n633,
    n34
  );


  buf
  g215
  (
    n530,
    n148
  );


  buf
  g216
  (
    n274,
    n133
  );


  buf
  g217
  (
    n529,
    n78
  );


  buf
  g218
  (
    n296,
    n115
  );


  buf
  g219
  (
    n615,
    n124
  );


  buf
  g220
  (
    n237,
    n141
  );


  not
  g221
  (
    n623,
    n139
  );


  buf
  g222
  (
    n330,
    n104
  );


  buf
  g223
  (
    n526,
    n82
  );


  not
  g224
  (
    n594,
    n40
  );


  not
  g225
  (
    n412,
    n83
  );


  not
  g226
  (
    n476,
    n57
  );


  buf
  g227
  (
    n580,
    n133
  );


  not
  g228
  (
    n463,
    n59
  );


  not
  g229
  (
    n259,
    n57
  );


  not
  g230
  (
    n391,
    n104
  );


  not
  g231
  (
    n173,
    n142
  );


  buf
  g232
  (
    n217,
    n64
  );


  not
  g233
  (
    n457,
    n58
  );


  buf
  g234
  (
    n298,
    n106
  );


  buf
  g235
  (
    n442,
    n42
  );


  not
  g236
  (
    n250,
    n153
  );


  buf
  g237
  (
    n420,
    n74
  );


  not
  g238
  (
    n461,
    n119
  );


  not
  g239
  (
    n198,
    n87
  );


  not
  g240
  (
    n584,
    n94
  );


  buf
  g241
  (
    n367,
    n102
  );


  buf
  g242
  (
    n491,
    n61
  );


  buf
  g243
  (
    n434,
    n45
  );


  buf
  g244
  (
    n453,
    n54
  );


  not
  g245
  (
    n368,
    n38
  );


  not
  g246
  (
    n230,
    n46
  );


  buf
  g247
  (
    n588,
    n71
  );


  not
  g248
  (
    n352,
    n87
  );


  buf
  g249
  (
    n546,
    n154
  );


  buf
  g250
  (
    n649,
    n51
  );


  buf
  g251
  (
    n621,
    n157
  );


  buf
  g252
  (
    n566,
    n108
  );


  not
  g253
  (
    n508,
    n71
  );


  not
  g254
  (
    n415,
    n42
  );


  buf
  g255
  (
    n394,
    n43
  );


  not
  g256
  (
    n641,
    n66
  );


  not
  g257
  (
    n392,
    n120
  );


  buf
  g258
  (
    n510,
    n125
  );


  not
  g259
  (
    n320,
    n61
  );


  not
  g260
  (
    n496,
    n62
  );


  not
  g261
  (
    n340,
    n151
  );


  not
  g262
  (
    n480,
    n86
  );


  not
  g263
  (
    n332,
    n64
  );


  buf
  g264
  (
    n602,
    n111
  );


  not
  g265
  (
    n390,
    n102
  );


  not
  g266
  (
    n314,
    n114
  );


  buf
  g267
  (
    n451,
    n110
  );


  buf
  g268
  (
    n532,
    n123
  );


  not
  g269
  (
    n571,
    n54
  );


  not
  g270
  (
    n338,
    n91
  );


  not
  g271
  (
    n593,
    n134
  );


  buf
  g272
  (
    n396,
    n153
  );


  buf
  g273
  (
    n305,
    n42
  );


  buf
  g274
  (
    n306,
    n56
  );


  buf
  g275
  (
    n423,
    n111
  );


  buf
  g276
  (
    n564,
    n101
  );


  buf
  g277
  (
    n293,
    n148
  );


  not
  g278
  (
    n591,
    n79
  );


  buf
  g279
  (
    n263,
    n108
  );


  buf
  g280
  (
    n582,
    n127
  );


  buf
  g281
  (
    n643,
    n96
  );


  not
  g282
  (
    n321,
    n140
  );


  not
  g283
  (
    n450,
    n52
  );


  not
  g284
  (
    n168,
    n136
  );


  buf
  g285
  (
    n525,
    n116
  );


  not
  g286
  (
    n589,
    n149
  );


  buf
  g287
  (
    n552,
    n158
  );


  buf
  g288
  (
    n247,
    n78
  );


  buf
  g289
  (
    n355,
    n154
  );


  not
  g290
  (
    n231,
    n53
  );


  buf
  g291
  (
    n292,
    n153
  );


  buf
  g292
  (
    n422,
    n46
  );


  not
  g293
  (
    n516,
    n105
  );


  buf
  g294
  (
    n199,
    n126
  );


  not
  g295
  (
    n536,
    n36
  );


  buf
  g296
  (
    n278,
    n34
  );


  not
  g297
  (
    n614,
    n53
  );


  buf
  g298
  (
    n317,
    n144
  );


  not
  g299
  (
    n481,
    n152
  );


  not
  g300
  (
    n576,
    n48
  );


  not
  g301
  (
    n213,
    n98
  );


  not
  g302
  (
    n210,
    n81
  );


  buf
  g303
  (
    n583,
    n92
  );


  buf
  g304
  (
    n627,
    n60
  );


  not
  g305
  (
    n346,
    n123
  );


  buf
  g306
  (
    n440,
    n125
  );


  not
  g307
  (
    n492,
    n149
  );


  not
  g308
  (
    n304,
    n151
  );


  not
  g309
  (
    n281,
    n99
  );


  buf
  g310
  (
    n282,
    n157
  );


  buf
  g311
  (
    n219,
    n74
  );


  buf
  g312
  (
    n616,
    n144
  );


  not
  g313
  (
    KeyWire_0_3,
    n63
  );


  buf
  g314
  (
    n474,
    n80
  );


  not
  g315
  (
    n319,
    n102
  );


  buf
  g316
  (
    n189,
    n109
  );


  not
  g317
  (
    n495,
    n63
  );


  buf
  g318
  (
    KeyWire_0_26,
    n94
  );


  not
  g319
  (
    n629,
    n70
  );


  not
  g320
  (
    n642,
    n69
  );


  not
  g321
  (
    n232,
    n140
  );


  buf
  g322
  (
    n331,
    n143
  );


  buf
  g323
  (
    n190,
    n65
  );


  not
  g324
  (
    n348,
    n84
  );


  not
  g325
  (
    n287,
    n103
  );


  buf
  g326
  (
    n467,
    n115
  );


  buf
  g327
  (
    n271,
    n117
  );


  buf
  g328
  (
    n204,
    n138
  );


  buf
  g329
  (
    n229,
    n154
  );


  not
  g330
  (
    n235,
    n41
  );


  buf
  g331
  (
    n586,
    n92
  );


  buf
  g332
  (
    n645,
    n127
  );


  not
  g333
  (
    n349,
    n122
  );


  buf
  g334
  (
    n180,
    n45
  );


  buf
  g335
  (
    KeyWire_0_19,
    n110
  );


  not
  g336
  (
    n610,
    n75
  );


  not
  g337
  (
    n477,
    n85
  );


  buf
  g338
  (
    n631,
    n53
  );


  not
  g339
  (
    n211,
    n142
  );


  not
  g340
  (
    n399,
    n70
  );


  not
  g341
  (
    n561,
    n106
  );


  buf
  g342
  (
    n178,
    n156
  );


  not
  g343
  (
    n652,
    n86
  );


  not
  g344
  (
    n551,
    n94
  );


  buf
  g345
  (
    n245,
    n76
  );


  not
  g346
  (
    n512,
    n35
  );


  buf
  g347
  (
    n562,
    n117
  );


  buf
  g348
  (
    n613,
    n43
  );


  buf
  g349
  (
    n625,
    n47
  );


  buf
  g350
  (
    n360,
    n100
  );


  buf
  g351
  (
    n470,
    n92
  );


  buf
  g352
  (
    n624,
    n38
  );


  buf
  g353
  (
    n489,
    n118
  );


  not
  g354
  (
    n606,
    n127
  );


  buf
  g355
  (
    n654,
    n101
  );


  not
  g356
  (
    n667,
    n120
  );


  not
  g357
  (
    n417,
    n150
  );


  buf
  g358
  (
    n644,
    n74
  );


  buf
  g359
  (
    n468,
    n39
  );


  not
  g360
  (
    n585,
    n53
  );


  not
  g361
  (
    n325,
    n79
  );


  not
  g362
  (
    n448,
    n55
  );


  not
  g363
  (
    n380,
    n112
  );


  buf
  g364
  (
    n161,
    n46
  );


  not
  g365
  (
    n339,
    n90
  );


  not
  g366
  (
    n234,
    n121
  );


  buf
  g367
  (
    n424,
    n43
  );


  not
  g368
  (
    n270,
    n49
  );


  not
  g369
  (
    n454,
    n126
  );


  not
  g370
  (
    n445,
    n69
  );


  buf
  g371
  (
    n377,
    n38
  );


  not
  g372
  (
    n534,
    n97
  );


  not
  g373
  (
    n220,
    n70
  );


  not
  g374
  (
    n260,
    n144
  );


  buf
  g375
  (
    n214,
    n128
  );


  buf
  g376
  (
    n456,
    n81
  );


  buf
  g377
  (
    n358,
    n139
  );


  not
  g378
  (
    n506,
    n120
  );


  not
  g379
  (
    n170,
    n68
  );


  not
  g380
  (
    n309,
    n107
  );


  buf
  g381
  (
    n342,
    n44
  );


  buf
  g382
  (
    n172,
    n79
  );


  buf
  g383
  (
    n611,
    n130
  );


  buf
  g384
  (
    n206,
    n65
  );


  buf
  g385
  (
    KeyWire_0_25,
    n97
  );


  not
  g386
  (
    n441,
    n147
  );


  buf
  g387
  (
    n539,
    n130
  );


  not
  g388
  (
    n577,
    n107
  );


  not
  g389
  (
    n553,
    n34
  );


  not
  g390
  (
    n431,
    n89
  );


  not
  g391
  (
    n374,
    n87
  );


  not
  g392
  (
    n258,
    n122
  );


  buf
  g393
  (
    n478,
    n157
  );


  not
  g394
  (
    n575,
    n54
  );


  not
  g395
  (
    n665,
    n109
  );


  not
  g396
  (
    n224,
    n155
  );


  not
  g397
  (
    n592,
    n116
  );


  buf
  g398
  (
    n216,
    n145
  );


  not
  g399
  (
    n658,
    n103
  );


  buf
  g400
  (
    n285,
    n83
  );


  buf
  g401
  (
    n404,
    n155
  );


  buf
  g402
  (
    n400,
    n41
  );


  not
  g403
  (
    n378,
    n140
  );


  buf
  g404
  (
    n570,
    n120
  );


  not
  g405
  (
    n475,
    n150
  );


  not
  g406
  (
    n598,
    n75
  );


  not
  g407
  (
    n261,
    n54
  );


  buf
  g408
  (
    n628,
    n91
  );


  not
  g409
  (
    n501,
    n59
  );


  buf
  g410
  (
    n514,
    n61
  );


  buf
  g411
  (
    n344,
    n59
  );


  not
  g412
  (
    n596,
    n131
  );


  not
  g413
  (
    n256,
    n113
  );


  not
  g414
  (
    n657,
    n125
  );


  not
  g415
  (
    n239,
    n100
  );


  buf
  g416
  (
    n277,
    n124
  );


  not
  g417
  (
    n488,
    n63
  );


  buf
  g418
  (
    n490,
    n78
  );


  buf
  g419
  (
    n302,
    n104
  );


  buf
  g420
  (
    n187,
    n137
  );


  buf
  g421
  (
    n336,
    n105
  );


  buf
  g422
  (
    n164,
    n107
  );


  buf
  g423
  (
    n373,
    n87
  );


  not
  g424
  (
    n381,
    n78
  );


  buf
  g425
  (
    n630,
    n135
  );


  not
  g426
  (
    n295,
    n61
  );


  not
  g427
  (
    n563,
    n33
  );


  not
  g428
  (
    n307,
    n103
  );


  buf
  g429
  (
    n333,
    n114
  );


  buf
  g430
  (
    n313,
    n71
  );


  not
  g431
  (
    n604,
    n98
  );


  buf
  g432
  (
    n289,
    n112
  );


  not
  g433
  (
    n315,
    n89
  );


  not
  g434
  (
    n484,
    n135
  );


  not
  g435
  (
    n218,
    n58
  );


  buf
  g436
  (
    n635,
    n118
  );


  buf
  g437
  (
    n634,
    n156
  );


  not
  g438
  (
    n387,
    n84
  );


  not
  g439
  (
    n301,
    n37
  );


  not
  g440
  (
    n413,
    n108
  );


  buf
  g441
  (
    n372,
    n138
  );


  buf
  g442
  (
    n222,
    n58
  );


  not
  g443
  (
    n337,
    n145
  );


  not
  g444
  (
    n175,
    n148
  );


  not
  g445
  (
    n662,
    n129
  );


  not
  g446
  (
    n371,
    n37
  );


  not
  g447
  (
    n416,
    n59
  );


  not
  g448
  (
    n291,
    n76
  );


  not
  g449
  (
    n522,
    n97
  );


  buf
  g450
  (
    n538,
    n45
  );


  not
  g451
  (
    n223,
    n77
  );


  not
  g452
  (
    n438,
    n122
  );


  not
  g453
  (
    n418,
    n38
  );


  buf
  g454
  (
    n555,
    n136
  );


  not
  g455
  (
    n226,
    n113
  );


  buf
  g456
  (
    n221,
    n85
  );


  not
  g457
  (
    n265,
    n118
  );


  buf
  g458
  (
    n326,
    n80
  );


  not
  g459
  (
    n407,
    n82
  );


  not
  g460
  (
    n466,
    n95
  );


  buf
  g461
  (
    n632,
    n33
  );


  not
  g462
  (
    n446,
    n74
  );


  not
  g463
  (
    n425,
    n69
  );


  buf
  g464
  (
    n225,
    n111
  );


  not
  g465
  (
    n410,
    n75
  );


  buf
  g466
  (
    n533,
    n35
  );


  buf
  g467
  (
    n465,
    n159
  );


  not
  g468
  (
    n253,
    n64
  );


  buf
  g469
  (
    n345,
    n86
  );


  not
  g470
  (
    n455,
    n40
  );


  buf
  g471
  (
    n300,
    n49
  );


  buf
  g472
  (
    n207,
    n73
  );


  not
  g473
  (
    n334,
    n68
  );


  not
  g474
  (
    n640,
    n76
  );


  buf
  g475
  (
    n365,
    n34
  );


  not
  g476
  (
    n612,
    n77
  );


  buf
  g477
  (
    n242,
    n106
  );


  not
  g478
  (
    n188,
    n132
  );


  not
  g479
  (
    n609,
    n131
  );


  buf
  g480
  (
    n528,
    n95
  );


  not
  g481
  (
    n421,
    n88
  );


  not
  g482
  (
    n487,
    n84
  );


  buf
  g483
  (
    n354,
    n135
  );


  buf
  g484
  (
    n398,
    n83
  );


  buf
  g485
  (
    n485,
    n155
  );


  not
  g486
  (
    n347,
    n83
  );


  not
  g487
  (
    n497,
    n150
  );


  buf
  g488
  (
    n176,
    n146
  );


  not
  g489
  (
    n248,
    n136
  );


  not
  g490
  (
    n181,
    n47
  );


  buf
  g491
  (
    n639,
    n49
  );


  buf
  g492
  (
    n341,
    n133
  );


  not
  g493
  (
    n531,
    n81
  );


  not
  g494
  (
    n366,
    n36
  );


  not
  g495
  (
    n167,
    n145
  );


  buf
  g496
  (
    n428,
    n153
  );


  buf
  g497
  (
    n449,
    n89
  );


  not
  g498
  (
    n405,
    n114
  );


  not
  g499
  (
    n600,
    n136
  );


  not
  g500
  (
    n436,
    n88
  );


  not
  g501
  (
    n267,
    n80
  );


  buf
  g502
  (
    n437,
    n68
  );


  not
  g503
  (
    n385,
    n98
  );


  not
  g504
  (
    n482,
    n135
  );


  not
  g505
  (
    n503,
    n57
  );


  buf
  g506
  (
    n208,
    n105
  );


  not
  g507
  (
    n376,
    n113
  );


  buf
  g508
  (
    n663,
    n158
  );


  buf
  g509
  (
    n472,
    n37
  );


  buf
  g510
  (
    n200,
    n63
  );


  buf
  g511
  (
    n329,
    n137
  );


  buf
  g512
  (
    n393,
    n62
  );


  buf
  g513
  (
    n559,
    n58
  );


  not
  g514
  (
    n569,
    n102
  );


  not
  g515
  (
    n595,
    n47
  );


  not
  g516
  (
    n403,
    n125
  );


  buf
  g517
  (
    n479,
    n148
  );


  buf
  g518
  (
    n661,
    n110
  );


  not
  g519
  (
    n527,
    n124
  );


  buf
  g520
  (
    n353,
    n76
  );


  not
  g521
  (
    n406,
    n137
  );


  not
  g522
  (
    n323,
    n50
  );


  buf
  g523
  (
    n554,
    n154
  );


  buf
  g524
  (
    n574,
    n115
  );


  buf
  g525
  (
    n523,
    n109
  );


  buf
  g526
  (
    n542,
    n85
  );


  buf
  g527
  (
    n290,
    n122
  );


  buf
  g528
  (
    n273,
    n37
  );


  buf
  g529
  (
    n486,
    n67
  );


  buf
  g530
  (
    n311,
    n159
  );


  not
  g531
  (
    n251,
    n146
  );


  not
  g532
  (
    n362,
    n93
  );


  buf
  g533
  (
    n607,
    n142
  );


  not
  g534
  (
    n227,
    n79
  );


  not
  g535
  (
    n166,
    n132
  );


  buf
  g536
  (
    n379,
    n129
  );


  not
  g537
  (
    n411,
    n132
  );


  not
  g538
  (
    n432,
    n43
  );


  not
  g539
  (
    n364,
    n143
  );


  buf
  g540
  (
    n572,
    n152
  );


  not
  g541
  (
    n517,
    n50
  );


  not
  g542
  (
    n483,
    n107
  );


  buf
  g543
  (
    n435,
    n77
  );


  not
  g544
  (
    n182,
    n119
  );


  buf
  g545
  (
    n460,
    n127
  );


  buf
  g546
  (
    n587,
    n33
  );


  buf
  g547
  (
    n327,
    n51
  );


  not
  g548
  (
    n597,
    n121
  );


  not
  g549
  (
    n335,
    n130
  );


  not
  g550
  (
    n288,
    n150
  );


  buf
  g551
  (
    n419,
    n73
  );


  buf
  g552
  (
    n201,
    n39
  );


  not
  g553
  (
    n504,
    n96
  );


  not
  g554
  (
    n557,
    n132
  );


  buf
  g555
  (
    n195,
    n73
  );


  buf
  g556
  (
    n452,
    n103
  );


  not
  g557
  (
    n310,
    n56
  );


  not
  g558
  (
    n275,
    n67
  );


  buf
  g559
  (
    n427,
    n97
  );


  not
  g560
  (
    n414,
    n41
  );


  buf
  g561
  (
    n620,
    n90
  );


  not
  g562
  (
    n556,
    n128
  );


  not
  g563
  (
    n241,
    n145
  );


  not
  g564
  (
    n651,
    n117
  );


  buf
  g565
  (
    n191,
    n56
  );


  not
  g566
  (
    n343,
    n138
  );


  not
  g567
  (
    n401,
    n137
  );


  buf
  g568
  (
    n386,
    n52
  );


  buf
  g569
  (
    n244,
    n66
  );


  not
  g570
  (
    n202,
    n55
  );


  buf
  g571
  (
    n498,
    n40
  );


  not
  g572
  (
    n389,
    n52
  );


  buf
  g573
  (
    n603,
    n141
  );


  buf
  g574
  (
    n560,
    n72
  );


  buf
  g575
  (
    n637,
    n129
  );


  not
  g576
  (
    n276,
    n52
  );


  buf
  g577
  (
    n547,
    n45
  );


  not
  g578
  (
    n660,
    n72
  );


  buf
  g579
  (
    n257,
    n36
  );


  buf
  g580
  (
    n283,
    n82
  );


  not
  g581
  (
    n573,
    n124
  );


  buf
  g582
  (
    n638,
    n41
  );


  buf
  g583
  (
    n171,
    n123
  );


  not
  g584
  (
    n228,
    n67
  );


  not
  g585
  (
    n601,
    n134
  );


  buf
  g586
  (
    n664,
    n99
  );


  not
  g587
  (
    n548,
    n62
  );


  buf
  g588
  (
    n543,
    n48
  );


  buf
  g589
  (
    n209,
    n39
  );


  not
  g590
  (
    n359,
    n82
  );


  buf
  g591
  (
    n656,
    n114
  );


  buf
  g592
  (
    n402,
    n64
  );


  buf
  g593
  (
    n179,
    n80
  );


  not
  g594
  (
    n255,
    n131
  );


  not
  g595
  (
    n369,
    n93
  );


  buf
  g596
  (
    n578,
    n62
  );


  not
  g597
  (
    n262,
    n143
  );


  not
  g598
  (
    n545,
    n139
  );


  not
  g599
  (
    n382,
    n99
  );


  not
  g600
  (
    n617,
    n86
  );


  not
  g601
  (
    KeyWire_0_20,
    n121
  );


  not
  g602
  (
    n655,
    n40
  );


  not
  g603
  (
    n266,
    n95
  );


  not
  g604
  (
    n196,
    n35
  );


  not
  g605
  (
    n269,
    n93
  );


  buf
  g606
  (
    n186,
    n50
  );


  buf
  g607
  (
    n409,
    n60
  );


  buf
  g608
  (
    n647,
    n44
  );


  not
  g609
  (
    n316,
    n146
  );


  not
  g610
  (
    n619,
    n92
  );


  not
  g611
  (
    n535,
    n149
  );


  buf
  g612
  (
    n608,
    n147
  );


  not
  g613
  (
    n500,
    n99
  );


  not
  g614
  (
    n590,
    n71
  );


  buf
  g615
  (
    n163,
    n128
  );


  buf
  g616
  (
    n284,
    n105
  );


  not
  g617
  (
    n549,
    n73
  );


  not
  g618
  (
    n192,
    n33
  );


  not
  g619
  (
    n165,
    n66
  );


  not
  g620
  (
    n264,
    n88
  );


  not
  g621
  (
    n622,
    n146
  );


  not
  g622
  (
    n666,
    n115
  );


  not
  g623
  (
    n205,
    n110
  );


  not
  g624
  (
    n357,
    n84
  );


  not
  g625
  (
    n361,
    n91
  );


  not
  g626
  (
    n193,
    n128
  );


  buf
  g627
  (
    n408,
    n157
  );


  buf
  g628
  (
    n356,
    n141
  );


  buf
  g629
  (
    n318,
    n55
  );


  buf
  g630
  (
    n458,
    n147
  );


  buf
  g631
  (
    n515,
    n48
  );


  buf
  g632
  (
    n184,
    n93
  );


  not
  g633
  (
    n303,
    n98
  );


  buf
  g634
  (
    n505,
    n44
  );


  not
  g635
  (
    n861,
    n315
  );


  not
  g636
  (
    n1255,
    n477
  );


  not
  g637
  (
    n1039,
    n394
  );


  buf
  g638
  (
    n1080,
    n523
  );


  not
  g639
  (
    n1587,
    n494
  );


  not
  g640
  (
    n706,
    n526
  );


  buf
  g641
  (
    n1240,
    n473
  );


  not
  g642
  (
    n959,
    n476
  );


  not
  g643
  (
    n1775,
    n173
  );


  not
  g644
  (
    n1202,
    n376
  );


  not
  g645
  (
    n876,
    n517
  );


  buf
  g646
  (
    n1075,
    n314
  );


  not
  g647
  (
    n1428,
    n251
  );


  buf
  g648
  (
    n1346,
    n465
  );


  not
  g649
  (
    n995,
    n373
  );


  not
  g650
  (
    n1375,
    n497
  );


  buf
  g651
  (
    n1623,
    n230
  );


  buf
  g652
  (
    n1792,
    n465
  );


  buf
  g653
  (
    n1810,
    n174
  );


  not
  g654
  (
    n1624,
    n345
  );


  not
  g655
  (
    n1292,
    n590
  );


  buf
  g656
  (
    n1464,
    n383
  );


  not
  g657
  (
    n870,
    n546
  );


  not
  g658
  (
    n1189,
    n554
  );


  buf
  g659
  (
    n668,
    n268
  );


  buf
  g660
  (
    n799,
    n423
  );


  not
  g661
  (
    n1563,
    n623
  );


  buf
  g662
  (
    n1174,
    n404
  );


  buf
  g663
  (
    n989,
    n202
  );


  buf
  g664
  (
    n1246,
    n464
  );


  not
  g665
  (
    n1211,
    n628
  );


  buf
  g666
  (
    n961,
    n573
  );


  buf
  g667
  (
    n1008,
    n611
  );


  not
  g668
  (
    n1207,
    n184
  );


  not
  g669
  (
    n775,
    n295
  );


  buf
  g670
  (
    n1197,
    n568
  );


  not
  g671
  (
    n747,
    n347
  );


  buf
  g672
  (
    n1590,
    n205
  );


  buf
  g673
  (
    n1708,
    n174
  );


  not
  g674
  (
    n1093,
    n200
  );


  not
  g675
  (
    n1697,
    n638
  );


  not
  g676
  (
    n994,
    n276
  );


  not
  g677
  (
    n1423,
    n417
  );


  not
  g678
  (
    n919,
    n612
  );


  not
  g679
  (
    n925,
    n601
  );


  not
  g680
  (
    n765,
    n177
  );


  buf
  g681
  (
    n1715,
    n537
  );


  not
  g682
  (
    n699,
    n470
  );


  buf
  g683
  (
    n1151,
    n299
  );


  buf
  g684
  (
    n1191,
    n268
  );


  buf
  g685
  (
    n1723,
    n630
  );


  not
  g686
  (
    n1293,
    n373
  );


  not
  g687
  (
    n1339,
    n175
  );


  buf
  g688
  (
    n874,
    n488
  );


  buf
  g689
  (
    n1507,
    n296
  );


  buf
  g690
  (
    n1824,
    n175
  );


  buf
  g691
  (
    n852,
    n491
  );


  not
  g692
  (
    n1645,
    n350
  );


  buf
  g693
  (
    n1314,
    n592
  );


  not
  g694
  (
    n1062,
    n508
  );


  not
  g695
  (
    n1785,
    n469
  );


  buf
  g696
  (
    n943,
    n494
  );


  buf
  g697
  (
    n1466,
    n293
  );


  buf
  g698
  (
    n783,
    n428
  );


  buf
  g699
  (
    n682,
    n285
  );


  not
  g700
  (
    n975,
    n377
  );


  not
  g701
  (
    n1817,
    n563
  );


  not
  g702
  (
    n1446,
    n164
  );


  not
  g703
  (
    n938,
    n219
  );


  not
  g704
  (
    n1456,
    n462
  );


  buf
  g705
  (
    n1578,
    n176
  );


  buf
  g706
  (
    n1130,
    n352
  );


  buf
  g707
  (
    n1070,
    n422
  );


  not
  g708
  (
    n1606,
    n218
  );


  buf
  g709
  (
    n1262,
    n503
  );


  buf
  g710
  (
    n1634,
    n602
  );


  not
  g711
  (
    n1582,
    n182
  );


  buf
  g712
  (
    n1562,
    n335
  );


  buf
  g713
  (
    n1795,
    n228
  );


  buf
  g714
  (
    n937,
    n398
  );


  not
  g715
  (
    n676,
    n234
  );


  not
  g716
  (
    n1381,
    n195
  );


  not
  g717
  (
    n1443,
    n311
  );


  buf
  g718
  (
    n809,
    n565
  );


  buf
  g719
  (
    n1169,
    n563
  );


  not
  g720
  (
    n900,
    n465
  );


  buf
  g721
  (
    n1317,
    n389
  );


  buf
  g722
  (
    n1395,
    n233
  );


  buf
  g723
  (
    n1717,
    n416
  );


  buf
  g724
  (
    n974,
    n471
  );


  not
  g725
  (
    n1689,
    n559
  );


  buf
  g726
  (
    n978,
    n269
  );


  not
  g727
  (
    n1179,
    n392
  );


  buf
  g728
  (
    n709,
    n374
  );


  buf
  g729
  (
    n792,
    n174
  );


  buf
  g730
  (
    n781,
    n525
  );


  not
  g731
  (
    n1672,
    n413
  );


  not
  g732
  (
    n1004,
    n518
  );


  buf
  g733
  (
    n1682,
    n638
  );


  not
  g734
  (
    n1777,
    n498
  );


  not
  g735
  (
    n1569,
    n199
  );


  not
  g736
  (
    n960,
    n640
  );


  not
  g737
  (
    n1765,
    n229
  );


  buf
  g738
  (
    n1121,
    n506
  );


  not
  g739
  (
    n776,
    n591
  );


  buf
  g740
  (
    n1750,
    n326
  );


  buf
  g741
  (
    n1639,
    n427
  );


  buf
  g742
  (
    n1372,
    n490
  );


  buf
  g743
  (
    n1519,
    n647
  );


  buf
  g744
  (
    n1050,
    n354
  );


  not
  g745
  (
    n794,
    n319
  );


  buf
  g746
  (
    n1148,
    n515
  );


  buf
  g747
  (
    n1033,
    n550
  );


  not
  g748
  (
    n1140,
    n324
  );


  not
  g749
  (
    n1437,
    n198
  );


  not
  g750
  (
    n1745,
    n369
  );


  buf
  g751
  (
    n993,
    n271
  );


  buf
  g752
  (
    n1132,
    n618
  );


  buf
  g753
  (
    n823,
    n433
  );


  buf
  g754
  (
    n1595,
    n213
  );


  buf
  g755
  (
    n894,
    n563
  );


  buf
  g756
  (
    n845,
    n484
  );


  not
  g757
  (
    n1095,
    n340
  );


  not
  g758
  (
    n1641,
    n223
  );


  not
  g759
  (
    n1532,
    n508
  );


  buf
  g760
  (
    n1340,
    n268
  );


  not
  g761
  (
    n1297,
    n186
  );


  buf
  g762
  (
    n1405,
    n606
  );


  buf
  g763
  (
    n1009,
    n462
  );


  not
  g764
  (
    n1352,
    n442
  );


  not
  g765
  (
    n904,
    n233
  );


  not
  g766
  (
    n1489,
    n514
  );


  buf
  g767
  (
    n1244,
    n635
  );


  buf
  g768
  (
    n681,
    n504
  );


  not
  g769
  (
    n1125,
    n506
  );


  buf
  g770
  (
    n1823,
    n316
  );


  not
  g771
  (
    n1284,
    n353
  );


  buf
  g772
  (
    n1632,
    n214
  );


  buf
  g773
  (
    n914,
    n557
  );


  buf
  g774
  (
    n1205,
    n354
  );


  not
  g775
  (
    n1758,
    n485
  );


  buf
  g776
  (
    n1473,
    n294
  );


  buf
  g777
  (
    n1001,
    n384
  );


  not
  g778
  (
    n1753,
    n404
  );


  buf
  g779
  (
    n908,
    n348
  );


  buf
  g780
  (
    n1005,
    n629
  );


  not
  g781
  (
    n853,
    n388
  );


  buf
  g782
  (
    n1161,
    n589
  );


  not
  g783
  (
    n1213,
    n306
  );


  not
  g784
  (
    n933,
    n629
  );


  buf
  g785
  (
    n1392,
    n575
  );


  buf
  g786
  (
    n1360,
    n425
  );


  not
  g787
  (
    n1143,
    n214
  );


  not
  g788
  (
    n918,
    n262
  );


  buf
  g789
  (
    n996,
    n170
  );


  buf
  g790
  (
    n1173,
    n249
  );


  buf
  g791
  (
    n935,
    n191
  );


  buf
  g792
  (
    n1442,
    n542
  );


  buf
  g793
  (
    n915,
    n319
  );


  not
  g794
  (
    n1522,
    n376
  );


  not
  g795
  (
    n1520,
    n214
  );


  not
  g796
  (
    n757,
    n470
  );


  buf
  g797
  (
    n1509,
    n267
  );


  buf
  g798
  (
    n1110,
    n424
  );


  buf
  g799
  (
    n1105,
    n431
  );


  buf
  g800
  (
    n748,
    n519
  );


  buf
  g801
  (
    n1270,
    n535
  );


  not
  g802
  (
    n1335,
    n346
  );


  not
  g803
  (
    n905,
    n280
  );


  not
  g804
  (
    n1705,
    n430
  );


  buf
  g805
  (
    n1759,
    n222
  );


  buf
  g806
  (
    n768,
    n244
  );


  not
  g807
  (
    n910,
    n406
  );


  not
  g808
  (
    n916,
    n554
  );


  not
  g809
  (
    n684,
    n592
  );


  buf
  g810
  (
    n820,
    n558
  );


  buf
  g811
  (
    n1784,
    n475
  );


  not
  g812
  (
    n711,
    n553
  );


  not
  g813
  (
    n818,
    n287
  );


  not
  g814
  (
    n761,
    n371
  );


  not
  g815
  (
    n1396,
    n644
  );


  not
  g816
  (
    n1113,
    n512
  );


  buf
  g817
  (
    n931,
    n351
  );


  not
  g818
  (
    n1277,
    n582
  );


  not
  g819
  (
    n1323,
    n485
  );


  buf
  g820
  (
    n1282,
    n428
  );


  buf
  g821
  (
    n1341,
    n646
  );


  buf
  g822
  (
    n1751,
    n499
  );


  not
  g823
  (
    n1348,
    n484
  );


  buf
  g824
  (
    n1794,
    n644
  );


  not
  g825
  (
    n1625,
    n538
  );


  buf
  g826
  (
    n1067,
    n321
  );


  buf
  g827
  (
    n1788,
    n461
  );


  not
  g828
  (
    n1159,
    n356
  );


  buf
  g829
  (
    n1772,
    n534
  );


  buf
  g830
  (
    n976,
    n240
  );


  buf
  g831
  (
    n1028,
    n250
  );


  buf
  g832
  (
    n1731,
    n331
  );


  buf
  g833
  (
    n1478,
    n163
  );


  not
  g834
  (
    n858,
    n621
  );


  buf
  g835
  (
    n1412,
    n363
  );


  not
  g836
  (
    n1101,
    n648
  );


  buf
  g837
  (
    n1180,
    n168
  );


  buf
  g838
  (
    n1783,
    n379
  );


  buf
  g839
  (
    n1414,
    n400
  );


  not
  g840
  (
    n1579,
    n401
  );


  not
  g841
  (
    n692,
    n265
  );


  not
  g842
  (
    n1576,
    n205
  );


  buf
  g843
  (
    n1188,
    n480
  );


  buf
  g844
  (
    n1376,
    n308
  );


  not
  g845
  (
    n1328,
    n623
  );


  buf
  g846
  (
    n1424,
    n354
  );


  not
  g847
  (
    n1727,
    n339
  );


  not
  g848
  (
    n1721,
    n265
  );


  buf
  g849
  (
    n1081,
    n198
  );


  buf
  g850
  (
    n1704,
    n227
  );


  not
  g851
  (
    n895,
    n532
  );


  not
  g852
  (
    n1126,
    n523
  );


  buf
  g853
  (
    n839,
    n298
  );


  buf
  g854
  (
    n1716,
    n453
  );


  not
  g855
  (
    n1542,
    n506
  );


  not
  g856
  (
    n966,
    n348
  );


  not
  g857
  (
    n932,
    n593
  );


  buf
  g858
  (
    n1020,
    n566
  );


  not
  g859
  (
    n1178,
    n275
  );


  buf
  g860
  (
    n1411,
    n247
  );


  not
  g861
  (
    n1153,
    n524
  );


  buf
  g862
  (
    n741,
    n278
  );


  buf
  g863
  (
    n1048,
    n403
  );


  buf
  g864
  (
    n929,
    n429
  );


  buf
  g865
  (
    n1329,
    n641
  );


  buf
  g866
  (
    n927,
    n562
  );


  buf
  g867
  (
    n1118,
    n575
  );


  buf
  g868
  (
    n1170,
    n198
  );


  buf
  g869
  (
    n1511,
    n259
  );


  not
  g870
  (
    n1680,
    n382
  );


  not
  g871
  (
    n784,
    n628
  );


  buf
  g872
  (
    n1799,
    n493
  );


  buf
  g873
  (
    n1540,
    n417
  );


  not
  g874
  (
    n1397,
    n337
  );


  not
  g875
  (
    n702,
    n330
  );


  not
  g876
  (
    n728,
    n599
  );


  buf
  g877
  (
    n1552,
    n553
  );


  not
  g878
  (
    n1796,
    n368
  );


  buf
  g879
  (
    n678,
    n614
  );


  not
  g880
  (
    n1218,
    n510
  );


  buf
  g881
  (
    n1308,
    n436
  );


  buf
  g882
  (
    n1150,
    n372
  );


  not
  g883
  (
    n669,
    n288
  );


  buf
  g884
  (
    n689,
    n385
  );


  not
  g885
  (
    n875,
    n446
  );


  buf
  g886
  (
    n963,
    n181
  );


  buf
  g887
  (
    n1377,
    n266
  );


  buf
  g888
  (
    n672,
    n543
  );


  not
  g889
  (
    n1065,
    n409
  );


  not
  g890
  (
    n1220,
    n485
  );


  buf
  g891
  (
    n1768,
    n290
  );


  buf
  g892
  (
    n1002,
    n451
  );


  buf
  g893
  (
    n1195,
    n472
  );


  buf
  g894
  (
    n1800,
    n546
  );


  not
  g895
  (
    n1049,
    n347
  );


  not
  g896
  (
    n1198,
    n204
  );


  not
  g897
  (
    n1684,
    n212
  );


  buf
  g898
  (
    n1612,
    n495
  );


  buf
  g899
  (
    n1107,
    n393
  );


  buf
  g900
  (
    n713,
    n346
  );


  not
  g901
  (
    n1807,
    n252
  );


  not
  g902
  (
    n1802,
    n568
  );


  not
  g903
  (
    n1670,
    n266
  );


  buf
  g904
  (
    n1383,
    n163
  );


  buf
  g905
  (
    n1815,
    n174
  );


  buf
  g906
  (
    n981,
    n440
  );


  buf
  g907
  (
    n1116,
    n604
  );


  buf
  g908
  (
    n1458,
    n303
  );


  not
  g909
  (
    n1103,
    n343
  );


  buf
  g910
  (
    n737,
    n211
  );


  not
  g911
  (
    n1015,
    n488
  );


  not
  g912
  (
    n1508,
    n629
  );


  buf
  g913
  (
    n685,
    n597
  );


  not
  g914
  (
    n671,
    n396
  );


  not
  g915
  (
    n1157,
    n251
  );


  not
  g916
  (
    n1671,
    n464
  );


  not
  g917
  (
    n1237,
    n637
  );


  not
  g918
  (
    KeyWire_0_30,
    n483
  );


  not
  g919
  (
    n1321,
    n301
  );


  buf
  g920
  (
    n1057,
    n236
  );


  buf
  g921
  (
    n1779,
    n456
  );


  not
  g922
  (
    n913,
    n302
  );


  not
  g923
  (
    n1633,
    n423
  );


  not
  g924
  (
    n1215,
    n591
  );


  buf
  g925
  (
    n1322,
    n501
  );


  buf
  g926
  (
    n1530,
    n357
  );


  not
  g927
  (
    n1433,
    n418
  );


  buf
  g928
  (
    n1295,
    n329
  );


  not
  g929
  (
    n1762,
    n478
  );


  buf
  g930
  (
    n1604,
    n597
  );


  buf
  g931
  (
    n1011,
    n321
  );


  buf
  g932
  (
    n1755,
    n480
  );


  buf
  g933
  (
    n1764,
    n272
  );


  not
  g934
  (
    n1460,
    n315
  );


  not
  g935
  (
    n1034,
    n474
  );


  not
  g936
  (
    n1256,
    n263
  );


  buf
  g937
  (
    n1462,
    n500
  );


  not
  g938
  (
    n1131,
    n189
  );


  buf
  g939
  (
    n850,
    n186
  );


  buf
  g940
  (
    n1556,
    n225
  );


  buf
  g941
  (
    KeyWire_0_16,
    n408
  );


  buf
  g942
  (
    n1588,
    n377
  );


  buf
  g943
  (
    n1371,
    n275
  );


  not
  g944
  (
    n1500,
    n408
  );


  buf
  g945
  (
    n1338,
    n573
  );


  not
  g946
  (
    n1659,
    n437
  );


  buf
  g947
  (
    n1431,
    n201
  );


  buf
  g948
  (
    n1575,
    n605
  );


  buf
  g949
  (
    n1259,
    n290
  );


  not
  g950
  (
    n1248,
    n218
  );


  not
  g951
  (
    n1361,
    n405
  );


  buf
  g952
  (
    n766,
    n179
  );


  not
  g953
  (
    n700,
    n163
  );


  not
  g954
  (
    n881,
    n334
  );


  not
  g955
  (
    n769,
    n627
  );


  buf
  g956
  (
    n836,
    n310
  );


  not
  g957
  (
    n1778,
    n270
  );


  not
  g958
  (
    n1754,
    n364
  );


  buf
  g959
  (
    n841,
    n242
  );


  buf
  g960
  (
    n1117,
    n637
  );


  not
  g961
  (
    n1822,
    n373
  );


  not
  g962
  (
    n1390,
    n613
  );


  not
  g963
  (
    n888,
    n503
  );


  not
  g964
  (
    n834,
    n382
  );


  not
  g965
  (
    n716,
    n519
  );


  buf
  g966
  (
    n1186,
    n393
  );


  buf
  g967
  (
    n1076,
    n486
  );


  buf
  g968
  (
    n1052,
    n579
  );


  not
  g969
  (
    n1123,
    n633
  );


  buf
  g970
  (
    n1108,
    n172
  );


  buf
  g971
  (
    n832,
    n280
  );


  not
  g972
  (
    n865,
    n326
  );


  not
  g973
  (
    n1221,
    n219
  );


  not
  g974
  (
    n871,
    n322
  );


  not
  g975
  (
    n1642,
    n169
  );


  buf
  g976
  (
    n1681,
    n378
  );


  not
  g977
  (
    n1082,
    n524
  );


  buf
  g978
  (
    n1538,
    n243
  );


  not
  g979
  (
    n1531,
    n421
  );


  not
  g980
  (
    n827,
    n341
  );


  buf
  g981
  (
    n1319,
    n487
  );


  not
  g982
  (
    n1688,
    n239
  );


  not
  g983
  (
    n1266,
    n337
  );


  buf
  g984
  (
    n1289,
    n377
  );


  buf
  g985
  (
    n730,
    n188
  );


  buf
  g986
  (
    n864,
    n305
  );


  not
  g987
  (
    n1739,
    n196
  );


  not
  g988
  (
    n1469,
    n307
  );


  buf
  g989
  (
    n1212,
    n288
  );


  buf
  g990
  (
    n764,
    n617
  );


  buf
  g991
  (
    n877,
    n360
  );


  not
  g992
  (
    n1662,
    n483
  );


  buf
  g993
  (
    n1550,
    n381
  );


  not
  g994
  (
    n800,
    n300
  );


  buf
  g995
  (
    n773,
    n390
  );


  not
  g996
  (
    n1133,
    n391
  );


  buf
  g997
  (
    n1204,
    n557
  );


  buf
  g998
  (
    n1769,
    n559
  );


  not
  g999
  (
    n1746,
    n218
  );


  not
  g1000
  (
    n1679,
    n298
  );


  buf
  g1001
  (
    n1445,
    n616
  );


  buf
  g1002
  (
    n987,
    n244
  );


  not
  g1003
  (
    n1744,
    n301
  );


  buf
  g1004
  (
    n1182,
    n204
  );


  not
  g1005
  (
    n1363,
    n482
  );


  buf
  g1006
  (
    n1463,
    n236
  );


  buf
  g1007
  (
    n1331,
    n414
  );


  not
  g1008
  (
    n1031,
    n319
  );


  buf
  g1009
  (
    n1012,
    n166
  );


  buf
  g1010
  (
    n1577,
    n245
  );


  not
  g1011
  (
    n719,
    n338
  );


  not
  g1012
  (
    n1206,
    n368
  );


  not
  g1013
  (
    n1393,
    n285
  );


  not
  g1014
  (
    n808,
    n287
  );


  not
  g1015
  (
    n920,
    n412
  );


  buf
  g1016
  (
    n1429,
    n589
  );


  buf
  g1017
  (
    n1102,
    n463
  );


  buf
  g1018
  (
    n1096,
    n552
  );


  buf
  g1019
  (
    n1610,
    n509
  );


  buf
  g1020
  (
    KeyWire_0_21,
    n258
  );


  buf
  g1021
  (
    n829,
    n556
  );


  not
  g1022
  (
    n1527,
    n439
  );


  not
  g1023
  (
    n1030,
    n422
  );


  not
  g1024
  (
    n1042,
    n181
  );


  not
  g1025
  (
    n1249,
    n583
  );


  not
  g1026
  (
    n917,
    n248
  );


  not
  g1027
  (
    n1674,
    n427
  );


  buf
  g1028
  (
    n1242,
    n436
  );


  buf
  g1029
  (
    n683,
    n615
  );


  not
  g1030
  (
    n892,
    n517
  );


  buf
  g1031
  (
    n695,
    n403
  );


  not
  g1032
  (
    n1185,
    n363
  );


  buf
  g1033
  (
    n1597,
    n617
  );


  buf
  g1034
  (
    n1155,
    n323
  );


  buf
  g1035
  (
    n1719,
    n203
  );


  not
  g1036
  (
    n1086,
    n620
  );


  buf
  g1037
  (
    n824,
    n595
  );


  not
  g1038
  (
    n1692,
    n579
  );


  not
  g1039
  (
    n1487,
    n291
  );


  buf
  g1040
  (
    n1814,
    n200
  );


  buf
  g1041
  (
    n1074,
    n603
  );


  not
  g1042
  (
    n797,
    n214
  );


  buf
  g1043
  (
    n1264,
    n616
  );


  buf
  g1044
  (
    n1358,
    n561
  );


  buf
  g1045
  (
    n1555,
    n325
  );


  buf
  g1046
  (
    n1658,
    n271
  );


  not
  g1047
  (
    n1752,
    n373
  );


  not
  g1048
  (
    n1693,
    n631
  );


  not
  g1049
  (
    n1265,
    n610
  );


  not
  g1050
  (
    n1801,
    n607
  );


  not
  g1051
  (
    n1279,
    n398
  );


  not
  g1052
  (
    n1236,
    n448
  );


  buf
  g1053
  (
    n750,
    n571
  );


  buf
  g1054
  (
    n805,
    n318
  );


  buf
  g1055
  (
    n743,
    n620
  );


  not
  g1056
  (
    n1541,
    n328
  );


  buf
  g1057
  (
    n1687,
    n593
  );


  not
  g1058
  (
    n1083,
    n375
  );


  not
  g1059
  (
    n704,
    n197
  );


  not
  g1060
  (
    n1468,
    n249
  );


  not
  g1061
  (
    n1496,
    n514
  );


  buf
  g1062
  (
    n1621,
    n277
  );


  buf
  g1063
  (
    n674,
    n578
  );


  not
  g1064
  (
    n705,
    n638
  );


  not
  g1065
  (
    n759,
    n384
  );


  not
  g1066
  (
    n868,
    n317
  );


  not
  g1067
  (
    n1379,
    n585
  );


  buf
  g1068
  (
    n1722,
    n383
  );


  not
  g1069
  (
    n1092,
    n216
  );


  buf
  g1070
  (
    n811,
    n444
  );


  not
  g1071
  (
    n1183,
    n641
  );


  not
  g1072
  (
    n847,
    n343
  );


  not
  g1073
  (
    n1490,
    n578
  );


  buf
  g1074
  (
    n1480,
    n620
  );


  not
  g1075
  (
    n1017,
    n555
  );


  not
  g1076
  (
    n1686,
    n293
  );


  buf
  g1077
  (
    n1055,
    n568
  );


  buf
  g1078
  (
    n1320,
    n507
  );


  not
  g1079
  (
    n1683,
    n418
  );


  not
  g1080
  (
    n867,
    n161
  );


  buf
  g1081
  (
    n1200,
    n420
  );


  not
  g1082
  (
    n1544,
    n290
  );


  buf
  g1083
  (
    n733,
    n172
  );


  not
  g1084
  (
    n1325,
    n199
  );


  not
  g1085
  (
    n1023,
    n179
  );


  buf
  g1086
  (
    n1664,
    n534
  );


  not
  g1087
  (
    n1286,
    n473
  );


  buf
  g1088
  (
    n1225,
    n425
  );


  not
  g1089
  (
    n901,
    n449
  );


  not
  g1090
  (
    n1056,
    n545
  );


  buf
  g1091
  (
    n970,
    n535
  );


  not
  g1092
  (
    n760,
    n469
  );


  buf
  g1093
  (
    n762,
    n204
  );


  not
  g1094
  (
    n1134,
    n618
  );


  not
  g1095
  (
    n1710,
    n215
  );


  not
  g1096
  (
    n1163,
    n469
  );


  not
  g1097
  (
    n1482,
    n484
  );


  not
  g1098
  (
    n1233,
    n461
  );


  not
  g1099
  (
    n1391,
    n213
  );


  buf
  g1100
  (
    n1732,
    n277
  );


  buf
  g1101
  (
    n1401,
    n651
  );


  not
  g1102
  (
    n983,
    n326
  );


  buf
  g1103
  (
    n1058,
    n294
  );


  buf
  g1104
  (
    n1425,
    n515
  );


  not
  g1105
  (
    n1069,
    n341
  );


  not
  g1106
  (
    n942,
    n604
  );


  not
  g1107
  (
    n736,
    n379
  );


  buf
  g1108
  (
    n1440,
    n627
  );


  not
  g1109
  (
    n1027,
    n197
  );


  not
  g1110
  (
    n1029,
    n500
  );


  buf
  g1111
  (
    n947,
    n182
  );


  buf
  g1112
  (
    n1811,
    n614
  );


  buf
  g1113
  (
    n1452,
    n605
  );


  buf
  g1114
  (
    n945,
    n397
  );


  buf
  g1115
  (
    n1347,
    n550
  );


  buf
  g1116
  (
    n988,
    n439
  );


  not
  g1117
  (
    n1094,
    n452
  );


  buf
  g1118
  (
    n1332,
    n178
  );


  buf
  g1119
  (
    n1294,
    n399
  );


  not
  g1120
  (
    n701,
    n561
  );


  not
  g1121
  (
    n1374,
    n380
  );


  buf
  g1122
  (
    n1145,
    n220
  );


  not
  g1123
  (
    n1770,
    n240
  );


  not
  g1124
  (
    n1354,
    n255
  );


  not
  g1125
  (
    n1757,
    n545
  );


  not
  g1126
  (
    n675,
    n520
  );


  not
  g1127
  (
    n751,
    n256
  );


  buf
  g1128
  (
    n721,
    n481
  );


  not
  g1129
  (
    n789,
    n445
  );


  buf
  g1130
  (
    n1702,
    n632
  );


  buf
  g1131
  (
    n869,
    n526
  );


  not
  g1132
  (
    n1327,
    n518
  );


  buf
  g1133
  (
    n1491,
    n377
  );


  not
  g1134
  (
    n1650,
    n414
  );


  buf
  g1135
  (
    n1038,
    n324
  );


  buf
  g1136
  (
    n1495,
    n251
  );


  buf
  g1137
  (
    n1304,
    n204
  );


  buf
  g1138
  (
    n1761,
    n491
  );


  not
  g1139
  (
    n854,
    n570
  );


  not
  g1140
  (
    n1434,
    n257
  );


  buf
  g1141
  (
    n880,
    n235
  );


  buf
  g1142
  (
    n1137,
    n386
  );


  buf
  g1143
  (
    n1647,
    n609
  );


  buf
  g1144
  (
    n1616,
    n454
  );


  buf
  g1145
  (
    n1690,
    n571
  );


  not
  g1146
  (
    n878,
    n253
  );


  buf
  g1147
  (
    n1296,
    n379
  );


  buf
  g1148
  (
    n1615,
    n624
  );


  not
  g1149
  (
    KeyWire_0_29,
    n217
  );


  buf
  g1150
  (
    n1476,
    n587
  );


  buf
  g1151
  (
    n1515,
    n362
  );


  buf
  g1152
  (
    n1063,
    n353
  );


  buf
  g1153
  (
    n1644,
    n260
  );


  buf
  g1154
  (
    n1479,
    n332
  );


  not
  g1155
  (
    n1591,
    n290
  );


  not
  g1156
  (
    n1553,
    n292
  );


  buf
  g1157
  (
    n1535,
    n472
  );


  buf
  g1158
  (
    n1694,
    n456
  );


  buf
  g1159
  (
    n822,
    n261
  );


  not
  g1160
  (
    n744,
    n567
  );


  buf
  g1161
  (
    n896,
    n491
  );


  not
  g1162
  (
    n670,
    n338
  );


  not
  g1163
  (
    n1127,
    n614
  );


  buf
  g1164
  (
    n1380,
    n335
  );


  not
  g1165
  (
    n1114,
    n634
  );


  buf
  g1166
  (
    n1366,
    n415
  );


  not
  g1167
  (
    n887,
    n222
  );


  not
  g1168
  (
    n1164,
    n570
  );


  not
  g1169
  (
    n1510,
    n341
  );


  not
  g1170
  (
    n862,
    n613
  );


  buf
  g1171
  (
    n1536,
    n368
  );


  not
  g1172
  (
    n1021,
    n336
  );


  buf
  g1173
  (
    n1600,
    n230
  );


  buf
  g1174
  (
    n1275,
    n642
  );


  buf
  g1175
  (
    n795,
    n545
  );


  not
  g1176
  (
    n810,
    n569
  );


  buf
  g1177
  (
    n1386,
    n338
  );


  not
  g1178
  (
    n957,
    n430
  );


  not
  g1179
  (
    n1657,
    n162
  );


  not
  g1180
  (
    n1646,
    n256
  );


  buf
  g1181
  (
    n746,
    n344
  );


  buf
  g1182
  (
    n1635,
    n630
  );


  buf
  g1183
  (
    n1006,
    n248
  );


  not
  g1184
  (
    n735,
    n578
  );


  not
  g1185
  (
    n1747,
    n626
  );


  not
  g1186
  (
    n1333,
    n184
  );


  not
  g1187
  (
    n785,
    n654
  );


  buf
  g1188
  (
    n1402,
    n375
  );


  not
  g1189
  (
    n1669,
    n309
  );


  buf
  g1190
  (
    n1791,
    n632
  );


  buf
  g1191
  (
    n1741,
    n511
  );


  not
  g1192
  (
    n1272,
    n582
  );


  not
  g1193
  (
    n1100,
    n482
  );


  buf
  g1194
  (
    n720,
    n431
  );


  not
  g1195
  (
    n1247,
    n641
  );


  not
  g1196
  (
    n1656,
    n387
  );


  buf
  g1197
  (
    n1141,
    n234
  );


  buf
  g1198
  (
    n844,
    n414
  );


  buf
  g1199
  (
    n802,
    n206
  );


  not
  g1200
  (
    n1059,
    n316
  );


  not
  g1201
  (
    n703,
    n441
  );


  buf
  g1202
  (
    n696,
    n329
  );


  buf
  g1203
  (
    n1809,
    n357
  );


  not
  g1204
  (
    n752,
    n619
  );


  buf
  g1205
  (
    n969,
    n502
  );


  not
  g1206
  (
    n677,
    n478
  );


  buf
  g1207
  (
    n1450,
    n362
  );


  buf
  g1208
  (
    n1149,
    n653
  );


  not
  g1209
  (
    n1276,
    n454
  );


  buf
  g1210
  (
    KeyWire_0_1,
    n592
  );


  buf
  g1211
  (
    n1120,
    n624
  );


  buf
  g1212
  (
    n1607,
    n596
  );


  buf
  g1213
  (
    n690,
    n453
  );


  not
  g1214
  (
    n1586,
    n494
  );


  not
  g1215
  (
    n1477,
    n240
  );


  buf
  g1216
  (
    n1699,
    n586
  );


  buf
  g1217
  (
    n754,
    n510
  );


  buf
  g1218
  (
    n1585,
    n388
  );


  not
  g1219
  (
    n1628,
    n426
  );


  buf
  g1220
  (
    n1337,
    n355
  );


  buf
  g1221
  (
    n803,
    n209
  );


  buf
  g1222
  (
    n1162,
    n598
  );


  buf
  g1223
  (
    n1298,
    n315
  );


  not
  g1224
  (
    n1449,
    n374
  );


  buf
  g1225
  (
    n886,
    n584
  );


  buf
  g1226
  (
    n1136,
    n623
  );


  buf
  g1227
  (
    n1609,
    n553
  );


  buf
  g1228
  (
    n673,
    n352
  );


  buf
  g1229
  (
    n1649,
    n312
  );


  not
  g1230
  (
    n1573,
    n171
  );


  buf
  g1231
  (
    n1617,
    n655
  );


  buf
  g1232
  (
    n967,
    n221
  );


  not
  g1233
  (
    n1524,
    n270
  );


  not
  g1234
  (
    n882,
    n212
  );


  not
  g1235
  (
    n1330,
    n429
  );


  not
  g1236
  (
    n782,
    n383
  );


  buf
  g1237
  (
    n1003,
    n215
  );


  not
  g1238
  (
    n1806,
    n399
  );


  buf
  g1239
  (
    n710,
    n320
  );


  buf
  g1240
  (
    n1700,
    n305
  );


  not
  g1241
  (
    n1711,
    n555
  );


  not
  g1242
  (
    n1740,
    n239
  );


  not
  g1243
  (
    n1720,
    n474
  );


  buf
  g1244
  (
    n1280,
    n634
  );


  not
  g1245
  (
    n731,
    n625
  );


  not
  g1246
  (
    n1516,
    n217
  );


  not
  g1247
  (
    n985,
    n314
  );


  buf
  g1248
  (
    n826,
    n551
  );


  not
  g1249
  (
    n1305,
    n289
  );


  buf
  g1250
  (
    n926,
    n196
  );


  buf
  g1251
  (
    n1436,
    n206
  );


  buf
  g1252
  (
    n1040,
    n654
  );


  buf
  g1253
  (
    n954,
    n408
  );


  not
  g1254
  (
    n771,
    n438
  );


  not
  g1255
  (
    n1701,
    n577
  );


  not
  g1256
  (
    n1685,
    n320
  );


  buf
  g1257
  (
    n1201,
    n490
  );


  buf
  g1258
  (
    n1344,
    n471
  );


  not
  g1259
  (
    n1819,
    n342
  );


  not
  g1260
  (
    n1362,
    n407
  );


  buf
  g1261
  (
    n1051,
    n601
  );


  not
  g1262
  (
    n842,
    n351
  );


  not
  g1263
  (
    n838,
    n463
  );


  buf
  g1264
  (
    n1345,
    n442
  );


  buf
  g1265
  (
    n1253,
    n376
  );


  not
  g1266
  (
    n1064,
    n619
  );


  buf
  g1267
  (
    n1349,
    n523
  );


  not
  g1268
  (
    n1565,
    n543
  );


  not
  g1269
  (
    n1526,
    n255
  );


  buf
  g1270
  (
    n1813,
    n541
  );


  not
  g1271
  (
    n1167,
    n246
  );


  buf
  g1272
  (
    n977,
    n193
  );


  not
  g1273
  (
    n1353,
    n621
  );


  not
  g1274
  (
    n1651,
    n477
  );


  not
  g1275
  (
    n1413,
    n317
  );


  not
  g1276
  (
    n1512,
    n183
  );


  not
  g1277
  (
    n1250,
    n237
  );


  buf
  g1278
  (
    n1097,
    n448
  );


  not
  g1279
  (
    n1318,
    n492
  );


  buf
  g1280
  (
    n1568,
    n630
  );


  not
  g1281
  (
    n788,
    n604
  );


  buf
  g1282
  (
    n1426,
    n261
  );


  not
  g1283
  (
    n1176,
    n465
  );


  not
  g1284
  (
    n1138,
    n355
  );


  buf
  g1285
  (
    n1528,
    n556
  );


  not
  g1286
  (
    n1427,
    n173
  );


  buf
  g1287
  (
    n855,
    n325
  );


  not
  g1288
  (
    n1663,
    n530
  );


  buf
  g1289
  (
    n1767,
    n300
  );


  not
  g1290
  (
    n1691,
    n183
  );


  not
  g1291
  (
    n738,
    n322
  );


  buf
  g1292
  (
    n1394,
    n254
  );


  buf
  g1293
  (
    n1399,
    n341
  );


  not
  g1294
  (
    n1252,
    n566
  );


  buf
  g1295
  (
    n1439,
    n224
  );


  buf
  g1296
  (
    n790,
    n266
  );


  buf
  g1297
  (
    n911,
    n567
  );


  not
  g1298
  (
    n1144,
    n413
  );


  not
  g1299
  (
    n891,
    n549
  );


  not
  g1300
  (
    n1175,
    n295
  );


  not
  g1301
  (
    n1283,
    n184
  );


  not
  g1302
  (
    n1668,
    n378
  );


  not
  g1303
  (
    n948,
    n339
  );


  not
  g1304
  (
    n1326,
    n612
  );


  buf
  g1305
  (
    n1493,
    n334
  );


  not
  g1306
  (
    n1045,
    n522
  );


  buf
  g1307
  (
    n902,
    n522
  );


  buf
  g1308
  (
    n1514,
    n180
  );


  buf
  g1309
  (
    n909,
    n211
  );


  buf
  g1310
  (
    n923,
    n412
  );


  buf
  g1311
  (
    n1551,
    n400
  );


  buf
  g1312
  (
    n1486,
    n261
  );


  buf
  g1313
  (
    n815,
    n317
  );


  not
  g1314
  (
    n1407,
    n305
  );


  not
  g1315
  (
    n1087,
    n511
  );


  buf
  g1316
  (
    n1226,
    n428
  );


  buf
  g1317
  (
    n1315,
    n259
  );


  not
  g1318
  (
    n1611,
    n588
  );


  buf
  g1319
  (
    n778,
    n206
  );


  not
  g1320
  (
    n1453,
    n417
  );


  buf
  g1321
  (
    n1598,
    n203
  );


  not
  g1322
  (
    n1521,
    n478
  );


  not
  g1323
  (
    n939,
    n496
  );


  not
  g1324
  (
    n786,
    n384
  );


  buf
  g1325
  (
    n1698,
    n650
  );


  buf
  g1326
  (
    n1019,
    n455
  );


  buf
  g1327
  (
    n1334,
    n530
  );


  buf
  g1328
  (
    n715,
    n296
  );


  not
  g1329
  (
    n1384,
    n203
  );


  buf
  g1330
  (
    n1229,
    n185
  );


  not
  g1331
  (
    n1457,
    n333
  );


  buf
  g1332
  (
    KeyWire_0_14,
    n245
  );


  not
  g1333
  (
    n1037,
    n569
  );


  not
  g1334
  (
    n1287,
    n395
  );


  not
  g1335
  (
    n1288,
    n273
  );


  buf
  g1336
  (
    n1085,
    n489
  );


  not
  g1337
  (
    n1454,
    n513
  );


  not
  g1338
  (
    n1438,
    n441
  );


  not
  g1339
  (
    n1599,
    n529
  );


  buf
  g1340
  (
    n1032,
    n602
  );


  buf
  g1341
  (
    n1224,
    n536
  );


  not
  g1342
  (
    n1422,
    n522
  );


  not
  g1343
  (
    n1415,
    n247
  );


  buf
  g1344
  (
    n1158,
    n640
  );


  not
  g1345
  (
    n1734,
    n242
  );


  not
  g1346
  (
    n1278,
    n421
  );


  not
  g1347
  (
    n1467,
    n323
  );


  not
  g1348
  (
    n1409,
    n292
  );


  buf
  g1349
  (
    n707,
    n572
  );


  buf
  g1350
  (
    n1084,
    n361
  );


  not
  g1351
  (
    n1593,
    n208
  );


  not
  g1352
  (
    n1342,
    n639
  );


  not
  g1353
  (
    n722,
    n543
  );


  not
  g1354
  (
    n1547,
    n495
  );


  buf
  g1355
  (
    n1821,
    n244
  );


  buf
  g1356
  (
    n1025,
    n161
  );


  buf
  g1357
  (
    n944,
    n209
  );


  buf
  g1358
  (
    n884,
    n511
  );


  buf
  g1359
  (
    n724,
    n242
  );


  not
  g1360
  (
    n1124,
    n628
  );


  not
  g1361
  (
    n817,
    n408
  );


  not
  g1362
  (
    n1627,
    n434
  );


  buf
  g1363
  (
    n1790,
    n646
  );


  not
  g1364
  (
    n1089,
    n331
  );


  not
  g1365
  (
    n843,
    n235
  );


  buf
  g1366
  (
    n903,
    n487
  );


  not
  g1367
  (
    n906,
    n172
  );


  not
  g1368
  (
    n1351,
    n539
  );


  buf
  g1369
  (
    n955,
    n456
  );


  not
  g1370
  (
    n1228,
    n526
  );


  not
  g1371
  (
    n727,
    n384
  );


  buf
  g1372
  (
    n1567,
    n400
  );


  buf
  g1373
  (
    n807,
    n440
  );


  not
  g1374
  (
    n1142,
    n633
  );


  not
  g1375
  (
    n1618,
    n212
  );


  not
  g1376
  (
    n1355,
    n475
  );


  not
  g1377
  (
    n739,
    n359
  );


  not
  g1378
  (
    n1350,
    n649
  );


  not
  g1379
  (
    n922,
    n379
  );


  not
  g1380
  (
    n1104,
    n603
  );


  not
  g1381
  (
    n1403,
    n472
  );


  buf
  g1382
  (
    n1274,
    n556
  );


  not
  g1383
  (
    n1196,
    n259
  );


  not
  g1384
  (
    n837,
    n547
  );


  not
  g1385
  (
    n1077,
    n514
  );


  buf
  g1386
  (
    n883,
    n323
  );


  not
  g1387
  (
    n1494,
    n310
  );


  not
  g1388
  (
    n1336,
    n573
  );


  buf
  g1389
  (
    n1300,
    n636
  );


  not
  g1390
  (
    n962,
    n342
  );


  not
  g1391
  (
    n840,
    n445
  );


  buf
  g1392
  (
    n1122,
    n570
  );


  buf
  g1393
  (
    n1184,
    n468
  );


  not
  g1394
  (
    n1417,
    n539
  );


  buf
  g1395
  (
    n687,
    n396
  );


  not
  g1396
  (
    n1492,
    n281
  );


  buf
  g1397
  (
    n856,
    n577
  );


  buf
  g1398
  (
    n1517,
    n232
  );


  not
  g1399
  (
    n1234,
    n566
  );


  not
  g1400
  (
    n1267,
    n450
  );


  buf
  g1401
  (
    n1261,
    n170
  );


  buf
  g1402
  (
    n812,
    n333
  );


  buf
  g1403
  (
    n1637,
    n390
  );


  buf
  g1404
  (
    n1303,
    n236
  );


  not
  g1405
  (
    n1073,
    n564
  );


  not
  g1406
  (
    n899,
    n490
  );


  not
  g1407
  (
    n1543,
    n499
  );


  not
  g1408
  (
    n1068,
    n577
  );


  buf
  g1409
  (
    KeyWire_0_27,
    n476
  );


  buf
  g1410
  (
    n1614,
    n643
  );


  buf
  g1411
  (
    n848,
    n600
  );


  not
  g1412
  (
    n1678,
    n328
  );


  buf
  g1413
  (
    n1506,
    n576
  );


  not
  g1414
  (
    n1564,
    n263
  );


  not
  g1415
  (
    n688,
    n587
  );


  not
  g1416
  (
    n1018,
    n329
  );


  buf
  g1417
  (
    n1448,
    n647
  );


  buf
  g1418
  (
    n1594,
    n380
  );


  buf
  g1419
  (
    n1416,
    n358
  );


  buf
  g1420
  (
    n1066,
    n329
  );


  buf
  g1421
  (
    n1060,
    n444
  );


  buf
  g1422
  (
    n1388,
    n418
  );


  buf
  g1423
  (
    n1099,
    n195
  );


  buf
  g1424
  (
    n1475,
    n651
  );


  not
  g1425
  (
    n1760,
    n498
  );


  buf
  g1426
  (
    n1441,
    n304
  );


  buf
  g1427
  (
    n1660,
    n543
  );


  not
  g1428
  (
    n1465,
    n547
  );


  not
  g1429
  (
    n1654,
    n213
  );


  not
  g1430
  (
    n1738,
    n386
  );


  buf
  g1431
  (
    n816,
    n538
  );


  not
  g1432
  (
    n992,
    n431
  );


  not
  g1433
  (
    n1398,
    n345
  );


  buf
  g1434
  (
    n729,
    n358
  );


  not
  g1435
  (
    n1418,
    n563
  );


  not
  g1436
  (
    n698,
    n438
  );


  not
  g1437
  (
    n1290,
    n403
  );


  not
  g1438
  (
    n1385,
    n395
  );


  buf
  g1439
  (
    n1420,
    n529
  );


  buf
  g1440
  (
    n1281,
    n380
  );


  buf
  g1441
  (
    n1648,
    n376
  );


  not
  g1442
  (
    n1497,
    n483
  );


  buf
  g1443
  (
    n1773,
    n271
  );


  buf
  g1444
  (
    n1171,
    n265
  );


  buf
  g1445
  (
    n924,
    n360
  );


  buf
  g1446
  (
    n726,
    n162
  );


  buf
  g1447
  (
    n1111,
    n381
  );


  buf
  g1448
  (
    n1000,
    n505
  );


  not
  g1449
  (
    n828,
    n312
  );


  not
  g1450
  (
    n1210,
    n300
  );


  buf
  g1451
  (
    n1470,
    n468
  );


  not
  g1452
  (
    n857,
    n471
  );


  buf
  g1453
  (
    n1603,
    n281
  );


  not
  g1454
  (
    n1112,
    n194
  );


  buf
  g1455
  (
    n1245,
    n221
  );


  not
  g1456
  (
    n1581,
    n426
  );


  not
  g1457
  (
    n796,
    n502
  );


  not
  g1458
  (
    n859,
    n188
  );


  not
  g1459
  (
    n1419,
    n590
  );


  not
  g1460
  (
    n941,
    n173
  );


  not
  g1461
  (
    n889,
    n468
  );


  not
  g1462
  (
    n1620,
    n608
  );


  buf
  g1463
  (
    n1602,
    n537
  );


  buf
  g1464
  (
    n1559,
    n542
  );


  not
  g1465
  (
    n1776,
    n458
  );


  not
  g1466
  (
    n958,
    n426
  );


  not
  g1467
  (
    n912,
    n259
  );


  not
  g1468
  (
    n1724,
    n582
  );


  not
  g1469
  (
    n1596,
    n366
  );


  buf
  g1470
  (
    n1343,
    n453
  );


  not
  g1471
  (
    n1216,
    n635
  );


  not
  g1472
  (
    n1046,
    n345
  );


  buf
  g1473
  (
    n1177,
    n471
  );


  not
  g1474
  (
    n1024,
    n645
  );


  not
  g1475
  (
    n866,
    n428
  );


  not
  g1476
  (
    n717,
    n601
  );


  buf
  g1477
  (
    n1572,
    n225
  );


  buf
  g1478
  (
    n679,
    n561
  );


  not
  g1479
  (
    n1115,
    n318
  );


  not
  g1480
  (
    n1373,
    n243
  );


  buf
  g1481
  (
    n1156,
    n413
  );


  not
  g1482
  (
    n780,
    n610
  );


  buf
  g1483
  (
    n745,
    n549
  );


  not
  g1484
  (
    n1119,
    n411
  );


  not
  g1485
  (
    n1707,
    n570
  );


  buf
  g1486
  (
    n952,
    n639
  );


  buf
  g1487
  (
    n1222,
    n481
  );


  buf
  g1488
  (
    n1356,
    n402
  );


  not
  g1489
  (
    n1561,
    n636
  );


  not
  g1490
  (
    n1797,
    n267
  );


  buf
  g1491
  (
    n846,
    n520
  );


  buf
  g1492
  (
    n708,
    n541
  );


  not
  g1493
  (
    n1311,
    n645
  );


  buf
  g1494
  (
    n1619,
    n164
  );


  buf
  g1495
  (
    n1309,
    n437
  );


  buf
  g1496
  (
    n1273,
    n198
  );


  not
  g1497
  (
    n714,
    n215
  );


  buf
  g1498
  (
    n734,
    n306
  );


  buf
  g1499
  (
    n725,
    n538
  );


  buf
  g1500
  (
    n1539,
    n502
  );


  buf
  g1501
  (
    n1444,
    n305
  );


  not
  g1502
  (
    n956,
    n528
  );


  buf
  g1503
  (
    n1299,
    n626
  );


  not
  g1504
  (
    n1435,
    n552
  );


  not
  g1505
  (
    n1152,
    n464
  );


  not
  g1506
  (
    n965,
    n309
  );


  not
  g1507
  (
    n686,
    n366
  );


  not
  g1508
  (
    n1816,
    n297
  );


  buf
  g1509
  (
    n1774,
    n558
  );


  not
  g1510
  (
    n1172,
    n598
  );


  buf
  g1511
  (
    n758,
    n183
  );


  not
  g1512
  (
    n1088,
    n649
  );


  buf
  g1513
  (
    n1243,
    n632
  );


  buf
  g1514
  (
    n1365,
    n411
  );


  not
  g1515
  (
    n1047,
    n588
  );


  buf
  g1516
  (
    n1165,
    n205
  );


  not
  g1517
  (
    n1459,
    n524
  );


  nor
  g1518
  (
    n1502,
    n425,
    n595,
    n479,
    n327
  );


  nor
  g1519
  (
    n1504,
    n427,
    n224,
    n583,
    n429
  );


  or
  g1520
  (
    n1378,
    n325,
    n447,
    n411,
    n650
  );


  or
  g1521
  (
    n1803,
    n310,
    n586,
    n165,
    n459
  );


  or
  g1522
  (
    n1820,
    n626,
    n256,
    n302,
    n624
  );


  nand
  g1523
  (
    n1655,
    n348,
    n607,
    n262,
    n626
  );


  xnor
  g1524
  (
    n1227,
    n442,
    n179,
    n371,
    n372
  );


  nor
  g1525
  (
    n1523,
    n313,
    n361,
    n311,
    n242
  );


  xnor
  g1526
  (
    n1798,
    n601,
    n403,
    n278,
    n547
  );


  or
  g1527
  (
    n1622,
    n631,
    n292,
    n633,
    n642
  );


  xnor
  g1528
  (
    n1192,
    n342,
    n279,
    n161,
    n577
  );


  or
  g1529
  (
    n1673,
    n420,
    n535,
    n588,
    n607
  );


  and
  g1530
  (
    n1484,
    n390,
    n650,
    n556,
    n193
  );


  nor
  g1531
  (
    n1601,
    n274,
    n336,
    n191,
    n518
  );


  or
  g1532
  (
    n973,
    n187,
    n254,
    n286,
    n353
  );


  xnor
  g1533
  (
    n851,
    n455,
    n285,
    n317,
    n549
  );


  and
  g1534
  (
    n1793,
    n284,
    n479,
    n313,
    n263
  );


  nand
  g1535
  (
    n1230,
    n569,
    n653,
    n414,
    n189
  );


  and
  g1536
  (
    n986,
    n438,
    n283,
    n574,
    n571
  );


  xor
  g1537
  (
    n1718,
    n625,
    n402,
    n567,
    n594
  );


  xnor
  g1538
  (
    n1041,
    n499,
    n201,
    n530,
    n251
  );


  xnor
  g1539
  (
    n1251,
    n419,
    n628,
    n479,
    n266
  );


  xor
  g1540
  (
    n1560,
    n423,
    n324,
    n534,
    n513
  );


  nand
  g1541
  (
    n1804,
    n221,
    n487,
    n449,
    n375
  );


  or
  g1542
  (
    n1194,
    n511,
    n378,
    n167,
    n476
  );


  nor
  g1543
  (
    n1054,
    n169,
    n618,
    n596,
    n299
  );


  xnor
  g1544
  (
    n697,
    n433,
    n176,
    n544,
    n572
  );


  or
  g1545
  (
    n1780,
    n439,
    n194,
    n189,
    n272
  );


  xor
  g1546
  (
    n1696,
    n652,
    n642,
    n551,
    n276
  );


  and
  g1547
  (
    n756,
    n602,
    n225,
    n230,
    n301
  );


  or
  g1548
  (
    n1667,
    n596,
    n644,
    n569,
    n579
  );


  nand
  g1549
  (
    n1166,
    n585,
    n308,
    n433,
    n434
  );


  nand
  g1550
  (
    n1726,
    n435,
    n187,
    n407,
    n397
  );


  and
  g1551
  (
    n1675,
    n457,
    n525,
    n531,
    n217
  );


  xor
  g1552
  (
    n1013,
    n381,
    n382,
    n166,
    n306
  );


  nor
  g1553
  (
    n1302,
    n385,
    n593,
    n209,
    n559
  );


  or
  g1554
  (
    n732,
    n594,
    n178,
    n606,
    n238
  );


  or
  g1555
  (
    n885,
    n606,
    n450,
    n283,
    n269
  );


  and
  g1556
  (
    n1079,
    n247,
    n578,
    n396,
    n427
  );


  xor
  g1557
  (
    n1291,
    n231,
    n619,
    n284,
    n207
  );


  xnor
  g1558
  (
    n1461,
    n492,
    n207,
    n355,
    n525
  );


  nor
  g1559
  (
    n793,
    n366,
    n327,
    n537,
    n277
  );


  nand
  g1560
  (
    n1713,
    n455,
    n542,
    n581,
    n401
  );


  and
  g1561
  (
    n1091,
    n630,
    n631,
    n293,
    n389
  );


  nor
  g1562
  (
    n1285,
    n622,
    n340,
    n548,
    n478
  );


  and
  g1563
  (
    n1430,
    n231,
    n344,
    n226,
    n298
  );


  nand
  g1564
  (
    n830,
    n327,
    n624,
    n232,
    n291
  );


  and
  g1565
  (
    n1254,
    n378,
    n322,
    n589,
    n190
  );


  xnor
  g1566
  (
    n1574,
    n638,
    n603,
    n369,
    n264
  );


  xor
  g1567
  (
    n1357,
    n356,
    n529,
    n413,
    n623
  );


  nand
  g1568
  (
    n1203,
    n366,
    n466,
    n510,
    n299
  );


  and
  g1569
  (
    n819,
    n422,
    n345,
    n207,
    n536
  );


  nor
  g1570
  (
    n1733,
    n652,
    n600,
    n580,
    n596
  );


  nand
  g1571
  (
    n1808,
    n367,
    n229,
    n503,
    n321
  );


  or
  g1572
  (
    n1306,
    n576,
    n269,
    n216,
    n201
  );


  and
  g1573
  (
    n1232,
    n552,
    n246,
    n310,
    n575
  );


  nor
  g1574
  (
    n940,
    n337,
    n392,
    n164,
    n292
  );


  xnor
  g1575
  (
    n1557,
    n536,
    n446,
    n210,
    n364
  );


  nand
  g1576
  (
    n1035,
    n486,
    n330,
    n535,
    n190
  );


  nor
  g1577
  (
    n1763,
    n279,
    n265,
    n544,
    n222
  );


  or
  g1578
  (
    n1219,
    n392,
    n289,
    n469,
    n581
  );


  nor
  g1579
  (
    n1078,
    n322,
    n587,
    n179,
    n604
  );


  nand
  g1580
  (
    n1257,
    n168,
    n512,
    n201,
    n275
  );


  nor
  g1581
  (
    n772,
    n255,
    n412,
    n531,
    n434
  );


  nor
  g1582
  (
    n991,
    n472,
    n391,
    n448,
    n394
  );


  xnor
  g1583
  (
    n1007,
    n481,
    n332,
    n276,
    n621
  );


  xnor
  g1584
  (
    n1187,
    n241,
    n200,
    n330,
    n497
  );


  nor
  g1585
  (
    n1789,
    n475,
    n258,
    n452,
    n171
  );


  nor
  g1586
  (
    n1231,
    n599,
    n582,
    n166,
    n436
  );


  xnor
  g1587
  (
    n1653,
    n579,
    n540,
    n600,
    n435
  );


  xnor
  g1588
  (
    n1359,
    n416,
    n598,
    n496,
    n554
  );


  nand
  g1589
  (
    n1129,
    n437,
    n621,
    n223,
    n612
  );


  xnor
  g1590
  (
    n897,
    n406,
    n336,
    n231,
    n386
  );


  and
  g1591
  (
    n777,
    n296,
    n616,
    n459,
    n289
  );


  and
  g1592
  (
    n801,
    n217,
    n486,
    n456,
    n531
  );


  nor
  g1593
  (
    n833,
    n272,
    n491,
    n410,
    n190
  );


  xnor
  g1594
  (
    n1665,
    n466,
    n526,
    n451,
    n459
  );


  nor
  g1595
  (
    n814,
    n436,
    n477,
    n264,
    n608
  );


  xor
  g1596
  (
    n1580,
    n245,
    n519,
    n497,
    n381
  );


  xnor
  g1597
  (
    KeyWire_0_24,
    n525,
    n237,
    n316,
    n637
  );


  nor
  g1598
  (
    n898,
    n260,
    n533,
    n399,
    n499
  );


  or
  g1599
  (
    n1534,
    n243,
    n625,
    n239,
    n565
  );


  xnor
  g1600
  (
    n1406,
    n387,
    n443,
    n249,
    n257
  );


  xor
  g1601
  (
    n997,
    n512,
    n312,
    n218,
    n580
  );


  xor
  g1602
  (
    n1571,
    n182,
    n344,
    n370,
    n274
  );


  xor
  g1603
  (
    n1548,
    n615,
    n655,
    n303,
    n622
  );


  xor
  g1604
  (
    n1818,
    n308,
    n177,
    n287,
    n350
  );


  and
  g1605
  (
    n1382,
    n515,
    n617,
    n516,
    n281
  );


  or
  g1606
  (
    n680,
    n397,
    n335,
    n627,
    n258
  );


  or
  g1607
  (
    n990,
    n250,
    n457,
    n343,
    n181
  );


  nand
  g1608
  (
    n1471,
    n540,
    n644,
    n178,
    n432
  );


  xnor
  g1609
  (
    n1584,
    n383,
    n500,
    n326,
    n476
  );


  nand
  g1610
  (
    n1369,
    n561,
    n280,
    n580,
    n278
  );


  nor
  g1611
  (
    n1260,
    n576,
    n597,
    n206,
    n572
  );


  nand
  g1612
  (
    n742,
    n516,
    n548,
    n406,
    n559
  );


  nand
  g1613
  (
    n1503,
    n387,
    n356,
    n461,
    n286
  );


  nand
  g1614
  (
    n1643,
    n252,
    n464,
    n339,
    n500
  );


  xnor
  g1615
  (
    n972,
    n541,
    n421,
    n307,
    n550
  );


  xor
  g1616
  (
    n1630,
    n328,
    n283,
    n443,
    n299
  );


  nor
  g1617
  (
    n1748,
    n270,
    n192,
    n365,
    n226
  );


  or
  g1618
  (
    n936,
    n501,
    n404,
    n562,
    n275
  );


  or
  g1619
  (
    n1408,
    n537,
    n333,
    n348,
    n532
  );


  nor
  g1620
  (
    n1570,
    n521,
    n180,
    n241,
    n334
  );


  xor
  g1621
  (
    n1737,
    n169,
    n342,
    n363,
    n296
  );


  xnor
  g1622
  (
    n1677,
    n304,
    n531,
    n510,
    n279
  );


  nand
  g1623
  (
    n1652,
    n489,
    n466,
    n223,
    n177
  );


  nand
  g1624
  (
    n1258,
    n279,
    n397,
    n226,
    n202
  );


  nor
  g1625
  (
    n1629,
    n234,
    n216,
    n304,
    n232
  );


  and
  g1626
  (
    n1214,
    n283,
    n501,
    n170,
    n619
  );


  xnor
  g1627
  (
    n1014,
    n613,
    n555,
    n311,
    n512
  );


  nand
  g1628
  (
    n1268,
    n254,
    n431,
    n415,
    n493
  );


  xor
  g1629
  (
    n804,
    n371,
    n620,
    n564,
    n524
  );


  nor
  g1630
  (
    n873,
    n288,
    n430,
    n211,
    n406
  );


  xor
  g1631
  (
    n1071,
    n462,
    n297,
    n518,
    n484
  );


  nor
  g1632
  (
    n1451,
    n584,
    n460,
    n547,
    n235
  );


  xnor
  g1633
  (
    n1782,
    n565,
    n467,
    n231,
    n560
  );


  xnor
  g1634
  (
    n1676,
    n398,
    n639,
    n380,
    n482
  );


  nor
  g1635
  (
    n1199,
    n653,
    n210,
    n513,
    n649
  );


  and
  g1636
  (
    n1589,
    n517,
    n508,
    n339,
    n392
  );


  xor
  g1637
  (
    n1709,
    n412,
    n294,
    n607,
    n504
  );


  xnor
  g1638
  (
    n863,
    n594,
    n548,
    n612,
    n241
  );


  or
  g1639
  (
    n1310,
    n492,
    n162,
    n208,
    n199
  );


  xnor
  g1640
  (
    n1098,
    n191,
    n303,
    n652,
    n309
  );


  and
  g1641
  (
    n1209,
    n350,
    n432,
    n605,
    n232
  );


  nand
  g1642
  (
    n835,
    n568,
    n505,
    n470,
    n590
  );


  nand
  g1643
  (
    n1756,
    n252,
    n447,
    n184,
    n215
  );


  xor
  g1644
  (
    n1546,
    n458,
    n261,
    n479,
    n622
  );


  nand
  g1645
  (
    n1147,
    n364,
    n627,
    n586,
    n433
  );


  xnor
  g1646
  (
    n779,
    n186,
    n407,
    n370,
    n185
  );


  xnor
  g1647
  (
    n1583,
    n355,
    n353,
    n338,
    n399
  );


  and
  g1648
  (
    n979,
    n521,
    n297,
    n239,
    n600
  );


  and
  g1649
  (
    n723,
    n643,
    n452,
    n180,
    n567
  );


  nor
  g1650
  (
    n1053,
    n424,
    n238,
    n222,
    n590
  );


  xor
  g1651
  (
    n890,
    n211,
    n219,
    n367,
    n417
  );


  nor
  g1652
  (
    n1533,
    n409,
    n445,
    n410,
    n282
  );


  xnor
  g1653
  (
    n1128,
    n293,
    n372,
    n460,
    n228
  );


  xnor
  g1654
  (
    n1217,
    n589,
    n445,
    n530,
    n313
  );


  nor
  g1655
  (
    n1537,
    n302,
    n527,
    n485,
    n365
  );


  or
  g1656
  (
    n1190,
    n391,
    n532,
    n552,
    n574
  );


  and
  g1657
  (
    n763,
    n191,
    n546,
    n225,
    n295
  );


  nor
  g1658
  (
    n1474,
    n246,
    n435,
    n520,
    n237
  );


  xnor
  g1659
  (
    n1271,
    n315,
    n424,
    n333,
    n409
  );


  and
  g1660
  (
    n1072,
    n502,
    n611,
    n219,
    n527
  );


  xor
  g1661
  (
    n1666,
    n203,
    n208,
    n457,
    n574
  );


  nand
  g1662
  (
    n1036,
    n420,
    n267,
    n425,
    n364
  );


  or
  g1663
  (
    n1061,
    n276,
    n354,
    n508,
    n474
  );


  or
  g1664
  (
    n1022,
    n611,
    n286,
    n487,
    n188
  );


  and
  g1665
  (
    n1370,
    n516,
    n352,
    n608,
    n520
  );


  nor
  g1666
  (
    n1109,
    n651,
    n196,
    n187,
    n220
  );


  and
  g1667
  (
    n1367,
    n193,
    n609,
    n583,
    n498
  );


  nor
  g1668
  (
    n813,
    n440,
    n635,
    n368,
    n646
  );


  nor
  g1669
  (
    n1044,
    n557,
    n303,
    n349,
    n540
  );


  or
  g1670
  (
    n1447,
    n302,
    n634,
    n356,
    n459
  );


  nand
  g1671
  (
    n1208,
    n539,
    n504,
    n374,
    n610
  );


  nand
  g1672
  (
    n1728,
    n253,
    n429,
    n480,
    n426
  );


  nor
  g1673
  (
    n872,
    n618,
    n581,
    n280,
    n282
  );


  or
  g1674
  (
    n787,
    n180,
    n481,
    n492,
    n393
  );


  nand
  g1675
  (
    n1160,
    n321,
    n572,
    n169,
    n385
  );


  nor
  g1676
  (
    n1239,
    n389,
    n462,
    n273,
    n529
  );


  and
  g1677
  (
    n770,
    n185,
    n467,
    n643,
    n374
  );


  and
  g1678
  (
    n1307,
    n274,
    n162,
    n419,
    n616
  );


  and
  g1679
  (
    n980,
    n447,
    n489,
    n171,
    n308
  );


  and
  g1680
  (
    n755,
    n212,
    n269,
    n295,
    n357
  );


  or
  g1681
  (
    n1135,
    n386,
    n586,
    n473,
    n654
  );


  nor
  g1682
  (
    n921,
    n194,
    n599,
    n645,
    n304
  );


  xor
  g1683
  (
    n1269,
    n495,
    n632,
    n647,
    n514
  );


  and
  g1684
  (
    n774,
    n444,
    n234,
    n306,
    n584
  );


  nand
  g1685
  (
    n1432,
    n244,
    n291,
    n410,
    n175
  );


  or
  g1686
  (
    n1529,
    n558,
    n415,
    n609,
    n221
  );


  or
  g1687
  (
    n1787,
    n634,
    n611,
    n546,
    n165
  );


  nand
  g1688
  (
    n767,
    n189,
    n595,
    n347,
    n549
  );


  nor
  g1689
  (
    n949,
    n617,
    n209,
    n346,
    n446
  );


  nor
  g1690
  (
    n1735,
    n393,
    n558,
    n307,
    n210
  );


  xor
  g1691
  (
    n1387,
    n328,
    n434,
    n301,
    n430
  );


  nand
  g1692
  (
    n831,
    n202,
    n496,
    n352,
    n401
  );


  nand
  g1693
  (
    KeyWire_0_12,
    n182,
    n362,
    n263,
    n648
  );


  xor
  g1694
  (
    n1483,
    n396,
    n493,
    n506,
    n460
  );


  xnor
  g1695
  (
    n1313,
    n318,
    n359,
    n648,
    n226
  );


  xnor
  g1696
  (
    n1786,
    n281,
    n260,
    n337,
    n324
  );


  or
  g1697
  (
    n1742,
    n551,
    n457,
    n167,
    n314
  );


  and
  g1698
  (
    n712,
    n172,
    n585,
    n202,
    n521
  );


  nor
  g1699
  (
    n1703,
    n551,
    n187,
    n161,
    n631
  );


  or
  g1700
  (
    n821,
    n452,
    n205,
    n360,
    n422
  );


  and
  g1701
  (
    n1605,
    n193,
    n165,
    n451,
    n474
  );


  and
  g1702
  (
    n1193,
    n264,
    n536,
    n274,
    n553
  );


  nor
  g1703
  (
    n1518,
    n564,
    n423,
    n186,
    n323
  );


  or
  g1704
  (
    n1263,
    n402,
    n648,
    n208,
    n282
  );


  xnor
  g1705
  (
    n860,
    n513,
    n521,
    n298,
    n486
  );


  xor
  g1706
  (
    n1592,
    n420,
    n597,
    n249,
    n168
  );


  nand
  g1707
  (
    n1168,
    n260,
    n560,
    n228,
    n173
  );


  or
  g1708
  (
    n1016,
    n262,
    n507,
    n440,
    n200
  );


  xor
  g1709
  (
    n1636,
    n411,
    n517,
    n359,
    n650
  );


  xor
  g1710
  (
    n1640,
    n358,
    n320,
    n188,
    n641
  );


  and
  g1711
  (
    n791,
    n439,
    n196,
    n313,
    n336
  );


  nor
  g1712
  (
    n1410,
    n254,
    n639,
    n197,
    n560
  );


  or
  g1713
  (
    KeyWire_0_31,
    n591,
    n312,
    n235,
    n533
  );


  nor
  g1714
  (
    n879,
    n307,
    n635,
    n654,
    n245
  );


  nor
  g1715
  (
    n1181,
    n272,
    n164,
    n503,
    n571
  );


  and
  g1716
  (
    n1223,
    n183,
    n250,
    n194,
    n334
  );


  xnor
  g1717
  (
    n1400,
    n228,
    n360,
    n359,
    n605
  );


  nor
  g1718
  (
    n1026,
    n351,
    n167,
    n575,
    n584
  );


  xor
  g1719
  (
    n1771,
    n453,
    n177,
    n587,
    n437
  );


  or
  g1720
  (
    n1730,
    n647,
    n580,
    n603,
    n287
  );


  or
  g1721
  (
    n1805,
    n220,
    n370,
    n592,
    n248
  );


  nand
  g1722
  (
    n1736,
    n468,
    n583,
    n454,
    n444
  );


  nor
  g1723
  (
    n1301,
    n229,
    n176,
    n195,
    n314
  );


  nand
  g1724
  (
    n1661,
    n451,
    n488,
    n519,
    n541
  );


  nand
  g1725
  (
    n934,
    n458,
    n240,
    n297,
    n432
  );


  nand
  g1726
  (
    n1139,
    n599,
    n609,
    n340,
    n331
  );


  nor
  g1727
  (
    n930,
    n375,
    n418,
    n277,
    n560
  );


  and
  g1728
  (
    n1725,
    n573,
    n640,
    n501,
    n346
  );


  nor
  g1729
  (
    n1472,
    n496,
    n343,
    n419,
    n347
  );


  or
  g1730
  (
    n753,
    n230,
    n629,
    n614,
    n255
  );


  and
  g1731
  (
    n1501,
    n369,
    n432,
    n528,
    n227
  );


  xnor
  g1732
  (
    n1043,
    n532,
    n166,
    n527,
    n643
  );


  xor
  g1733
  (
    n1238,
    n319,
    n210,
    n365,
    n349
  );


  nand
  g1734
  (
    n1498,
    n424,
    n248,
    n574,
    n533
  );


  nor
  g1735
  (
    n1631,
    n564,
    n207,
    n483,
    n652
  );


  and
  g1736
  (
    n749,
    n349,
    n606,
    n490,
    n361
  );


  and
  g1737
  (
    n1505,
    n527,
    n223,
    n494,
    n224
  );


  xor
  g1738
  (
    n1324,
    n470,
    n441,
    n405,
    n350
  );


  xor
  g1739
  (
    n1421,
    n351,
    n497,
    n243,
    n516
  );


  xnor
  g1740
  (
    n1364,
    n258,
    n544,
    n185,
    n646
  );


  nor
  g1741
  (
    n1812,
    n264,
    n421,
    n488,
    n252
  );


  xor
  g1742
  (
    n1545,
    n382,
    n238,
    n405,
    n288
  );


  and
  g1743
  (
    n1714,
    n542,
    n388,
    n176,
    n163
  );


  nand
  g1744
  (
    n1608,
    n402,
    n199,
    n195,
    n224
  );


  xnor
  g1745
  (
    n1241,
    n475,
    n636,
    n220,
    n473
  );


  or
  g1746
  (
    n950,
    n608,
    n455,
    n522,
    n398
  );


  and
  g1747
  (
    n825,
    n409,
    n581,
    n372,
    n566
  );


  or
  g1748
  (
    n1695,
    n236,
    n395,
    n548,
    n545
  );


  nor
  g1749
  (
    n998,
    n534,
    n256,
    n523,
    n270
  );


  and
  g1750
  (
    n1488,
    n365,
    n410,
    n555,
    n253
  );


  xnor
  g1751
  (
    n1554,
    n229,
    n216,
    n404,
    n370
  );


  xnor
  g1752
  (
    n893,
    n362,
    n463,
    n369,
    n528
  );


  nor
  g1753
  (
    n1549,
    n441,
    n309,
    n238,
    n170
  );


  nor
  g1754
  (
    n984,
    n284,
    n285,
    n286,
    n507
  );


  and
  g1755
  (
    n964,
    n539,
    n168,
    n332,
    n320
  );


  xor
  g1756
  (
    n1154,
    n311,
    n388,
    n419,
    n443
  );


  or
  g1757
  (
    n946,
    n610,
    n450,
    n390,
    n192
  );


  or
  g1758
  (
    n1389,
    n538,
    n271,
    n594,
    n282
  );


  xnor
  g1759
  (
    n1712,
    n268,
    n330,
    n625,
    n615
  );


  xor
  g1760
  (
    n1749,
    n461,
    n171,
    n528,
    n227
  );


  xnor
  g1761
  (
    n1513,
    n482,
    n550,
    n262,
    n613
  );


  or
  g1762
  (
    n1638,
    n585,
    n653,
    n458,
    n467
  );


  xor
  g1763
  (
    n1146,
    n557,
    n257,
    n493,
    n247
  );


  nor
  g1764
  (
    n1312,
    n637,
    n640,
    n544,
    n395
  );


  and
  g1765
  (
    n968,
    n391,
    n416,
    n615,
    n332
  );


  or
  g1766
  (
    n971,
    n401,
    n257,
    n407,
    n450
  );


  or
  g1767
  (
    n1481,
    n505,
    n213,
    n463,
    n335
  );


  nor
  g1768
  (
    n1316,
    n331,
    n622,
    n294,
    n443
  );


  nor
  g1769
  (
    n907,
    n515,
    n233,
    n642,
    n387
  );


  and
  g1770
  (
    n1455,
    n227,
    n446,
    n449,
    n363
  );


  nand
  g1771
  (
    n1566,
    n540,
    n190,
    n554,
    n327
  );


  xor
  g1772
  (
    n849,
    n645,
    n454,
    n435,
    n509
  );


  nand
  g1773
  (
    n691,
    n636,
    n178,
    n371,
    n602
  );


  xor
  g1774
  (
    n806,
    n448,
    n344,
    n438,
    n361
  );


  xnor
  g1775
  (
    n740,
    n598,
    n651,
    n349,
    n340
  );


  xnor
  g1776
  (
    n1781,
    n588,
    n385,
    n278,
    n633
  );


  nor
  g1777
  (
    n1743,
    n477,
    n415,
    n367,
    n197
  );


  nand
  g1778
  (
    n1706,
    n467,
    n192,
    n509,
    n284
  );


  or
  g1779
  (
    n1404,
    n300,
    n498,
    n358,
    n253
  );


  and
  g1780
  (
    n1613,
    n316,
    n318,
    n405,
    n505
  );


  xnor
  g1781
  (
    n798,
    n165,
    n449,
    n325,
    n233
  );


  nand
  g1782
  (
    n1235,
    n291,
    n442,
    n591,
    n466
  );


  and
  g1783
  (
    n718,
    n181,
    n273,
    n655,
    n565
  );


  nor
  g1784
  (
    n1499,
    n367,
    n357,
    n495,
    n389
  );


  xnor
  g1785
  (
    n1090,
    n237,
    n562,
    n576,
    n593
  );


  nor
  g1786
  (
    n982,
    n562,
    n394,
    n246,
    n480
  );


  nand
  g1787
  (
    n928,
    n595,
    n267,
    n192,
    n507
  );


  or
  g1788
  (
    n1766,
    n289,
    n504,
    n273,
    n460
  );


  nand
  g1789
  (
    n693,
    n167,
    n416,
    n241,
    n394
  );


  nand
  g1790
  (
    n1485,
    n447,
    n509,
    n175,
    n649
  );


  and
  g1791
  (
    n1106,
    n250,
    n400,
    n533,
    n489
  );


  xnor
  g1792
  (
    n2167,
    n1010,
    n1224,
    n1423,
    n993
  );


  nand
  g1793
  (
    n1991,
    n1599,
    n1346,
    n920,
    n1652
  );


  xnor
  g1794
  (
    n2401,
    n1110,
    n1127,
    n879,
    n1004
  );


  xnor
  g1795
  (
    n1985,
    n1720,
    n1063,
    n1315,
    n1298
  );


  xnor
  g1796
  (
    n1939,
    n1352,
    n1182,
    n995,
    n1162
  );


  xor
  g1797
  (
    n2404,
    n728,
    n1670,
    n1190,
    n1653
  );


  xor
  g1798
  (
    n2067,
    n1149,
    n1482,
    n1558,
    n1277
  );


  xnor
  g1799
  (
    n2349,
    n1776,
    n1747,
    n1017,
    n1667
  );


  nor
  g1800
  (
    n1893,
    n882,
    n1591,
    n814,
    n1074
  );


  or
  g1801
  (
    n2279,
    n1139,
    n1402,
    n724,
    n913
  );


  nor
  g1802
  (
    n2094,
    n763,
    n970,
    n1763,
    n1270
  );


  nor
  g1803
  (
    n2319,
    n787,
    n1788,
    n1636,
    n863
  );


  nand
  g1804
  (
    n2307,
    n715,
    n1401,
    n1399,
    n1674
  );


  or
  g1805
  (
    n1858,
    n1162,
    n1570,
    n1700,
    n1720
  );


  nor
  g1806
  (
    n1965,
    n1572,
    n1123,
    n684,
    n1409
  );


  nor
  g1807
  (
    n2180,
    n1728,
    n1780,
    n1706,
    n1756
  );


  nor
  g1808
  (
    n1860,
    n1361,
    n1463,
    n790,
    n688
  );


  nand
  g1809
  (
    n2104,
    n1311,
    n1204,
    n1281,
    n994
  );


  nand
  g1810
  (
    n1867,
    n693,
    n1461,
    n1018,
    n1085
  );


  and
  g1811
  (
    n2131,
    n1737,
    n1383,
    n1476,
    n1802
  );


  nor
  g1812
  (
    n1992,
    n1673,
    n1296,
    n1660,
    n1569
  );


  nor
  g1813
  (
    n2092,
    n1316,
    n1435,
    n1765,
    n1497
  );


  nand
  g1814
  (
    n1877,
    n767,
    n694,
    n1092,
    n1714
  );


  nand
  g1815
  (
    n1978,
    n1661,
    n936,
    n1280
  );


  nor
  g1816
  (
    n2297,
    n948,
    n951,
    n1309,
    n1029
  );


  and
  g1817
  (
    n2204,
    n1750,
    n1399,
    n1414,
    n1606
  );


  nor
  g1818
  (
    n2158,
    n1659,
    n915,
    n1299,
    n1372
  );


  xor
  g1819
  (
    n2429,
    n1710,
    n1128,
    n1288,
    n1033
  );


  nor
  g1820
  (
    n2033,
    n1605,
    n1568,
    n1705,
    n737
  );


  and
  g1821
  (
    n2366,
    n881,
    n976,
    n973,
    n1163
  );


  and
  g1822
  (
    n2047,
    n1263,
    n964,
    n1108,
    n1580
  );


  xnor
  g1823
  (
    n2154,
    n869,
    n1725,
    n1473,
    n1660
  );


  xor
  g1824
  (
    n2281,
    n853,
    n1099,
    n1647,
    n835
  );


  or
  g1825
  (
    n2274,
    n1028,
    n1184,
    n752,
    n1239
  );


  nor
  g1826
  (
    n2075,
    n1329,
    n1654,
    n1196,
    n864
  );


  or
  g1827
  (
    n2382,
    n1746,
    n1210,
    n718,
    n1214
  );


  or
  g1828
  (
    n1879,
    n671,
    n1217,
    n1065,
    n1172
  );


  or
  g1829
  (
    n1863,
    n1732,
    n1761,
    n1413,
    n1426
  );


  nor
  g1830
  (
    n2150,
    n1549,
    n972,
    n1646,
    n1157
  );


  xor
  g1831
  (
    n2036,
    n1084,
    n1166,
    n1713,
    n1193
  );


  xnor
  g1832
  (
    n1862,
    n1558,
    n1066,
    n1602,
    n1719
  );


  and
  g1833
  (
    n2140,
    n1721,
    n681,
    n1258,
    n730
  );


  xnor
  g1834
  (
    n2034,
    n736,
    n1278,
    n1067,
    n1524
  );


  xnor
  g1835
  (
    n2009,
    n1607,
    n1807,
    n1671,
    n1088
  );


  xor
  g1836
  (
    n2258,
    n1311,
    n1770,
    n867,
    n1708
  );


  or
  g1837
  (
    n2270,
    n1547,
    n1058,
    n1715,
    n1210
  );


  nand
  g1838
  (
    n2433,
    n1195,
    n1491,
    n1169,
    n1725
  );


  or
  g1839
  (
    n2373,
    n967,
    n773,
    n917,
    n1706
  );


  or
  g1840
  (
    n2283,
    n1513,
    n1171,
    n1556,
    n1318
  );


  nor
  g1841
  (
    n2478,
    n878,
    n1603,
    n1698,
    n1783
  );


  nor
  g1842
  (
    n1894,
    n1049,
    n747,
    n792,
    n1060
  );


  and
  g1843
  (
    n1982,
    n1566,
    n1681,
    n747,
    n1195
  );


  xnor
  g1844
  (
    n2421,
    n1005,
    n1155,
    n922,
    n888
  );


  xor
  g1845
  (
    n2205,
    n801,
    n1755,
    n1328,
    n832
  );


  or
  g1846
  (
    n2458,
    n1608,
    n1215,
    n1055,
    n1443
  );


  or
  g1847
  (
    n2345,
    n844,
    n920,
    n1721,
    n676
  );


  nor
  g1848
  (
    n2407,
    n777,
    n1284,
    n760,
    n1213
  );


  xnor
  g1849
  (
    n1901,
    n799,
    n826,
    n1681,
    n1245
  );


  and
  g1850
  (
    n2346,
    n1382,
    n1537,
    n1373,
    n1015
  );


  nor
  g1851
  (
    n1848,
    n1440,
    n1338,
    n1793,
    n983
  );


  or
  g1852
  (
    n2317,
    n1714,
    n733,
    n1510,
    n809
  );


  nand
  g1853
  (
    n2077,
    n703,
    n935,
    n929,
    n1344
  );


  nor
  g1854
  (
    n2040,
    n1698,
    n1730,
    n1147,
    n1754
  );


  or
  g1855
  (
    n1948,
    n1643,
    n1803,
    n1563,
    n1470
  );


  and
  g1856
  (
    n2446,
    n1136,
    n1470,
    n1385,
    n746
  );


  nand
  g1857
  (
    n2237,
    n788,
    n1548,
    n1231,
    n1754
  );


  nand
  g1858
  (
    n2266,
    n1197,
    n996,
    n938,
    n727
  );


  nand
  g1859
  (
    n1968,
    n1567,
    n1760,
    n932,
    n1207
  );


  or
  g1860
  (
    n2300,
    n1289,
    n1496,
    n1574,
    n716
  );


  xor
  g1861
  (
    n2159,
    n924,
    n1675,
    n1116,
    n1799
  );


  nand
  g1862
  (
    n1938,
    n732,
    n1056,
    n1782,
    n1079
  );


  xnor
  g1863
  (
    n2151,
    n1691,
    n1689,
    n1271,
    n1560
  );


  nand
  g1864
  (
    n2189,
    n1376,
    n1680,
    n877,
    n910
  );


  nor
  g1865
  (
    n2017,
    n1080,
    n821,
    n1584,
    n818
  );


  xnor
  g1866
  (
    n2280,
    n717,
    n1431,
    n1481,
    n1489
  );


  nand
  g1867
  (
    n2112,
    n1654,
    n1287,
    n1408,
    n1104
  );


  xor
  g1868
  (
    n2100,
    n1133,
    n1046,
    n679,
    n719
  );


  xnor
  g1869
  (
    n2232,
    n1703,
    n1724,
    n1761,
    n1651
  );


  nand
  g1870
  (
    n2468,
    n1115,
    n1305,
    n1506,
    n1091
  );


  and
  g1871
  (
    n1933,
    n1229,
    n1120,
    n1717,
    n871
  );


  nor
  g1872
  (
    n2168,
    n1765,
    n1124,
    n1578,
    n1505
  );


  and
  g1873
  (
    n2249,
    n965,
    n1002,
    n1036,
    n1222
  );


  nand
  g1874
  (
    n2028,
    n1235,
    n745,
    n1518,
    n1714
  );


  and
  g1875
  (
    n2288,
    n1766,
    n885,
    n890,
    n1755
  );


  nand
  g1876
  (
    n1833,
    n1752,
    n1630,
    n902,
    n1352
  );


  nor
  g1877
  (
    n2002,
    n1290,
    n1782,
    n1469,
    n1665
  );


  xnor
  g1878
  (
    n2325,
    n1693,
    n1779,
    n1018,
    n1711
  );


  xor
  g1879
  (
    n2069,
    n1432,
    n1141,
    n1771,
    n1198
  );


  xor
  g1880
  (
    n1953,
    n1637,
    n1682,
    n808,
    n677
  );


  nor
  g1881
  (
    n2273,
    n859,
    n1650,
    n1274,
    n1032
  );


  nand
  g1882
  (
    n2343,
    n1684,
    n1508,
    n677,
    n1179
  );


  nor
  g1883
  (
    n1996,
    n1583,
    n1038,
    n991,
    n816
  );


  xnor
  g1884
  (
    n2103,
    n921,
    n756,
    n811,
    n1792
  );


  and
  g1885
  (
    n1840,
    n946,
    n1773,
    n918,
    n1056
  );


  xor
  g1886
  (
    n2060,
    n1652,
    n725,
    n1712,
    n1678
  );


  xor
  g1887
  (
    n2459,
    n943,
    n1079,
    n1696,
    n1702
  );


  and
  g1888
  (
    n2127,
    n1053,
    n911,
    n1451,
    n1722
  );


  nand
  g1889
  (
    n2099,
    n1713,
    n1643,
    n1742,
    n675
  );


  nor
  g1890
  (
    n2177,
    n1227,
    n1266,
    n1582,
    n1512
  );


  xor
  g1891
  (
    n2265,
    n1800,
    n1403,
    n1254,
    n1784
  );


  nor
  g1892
  (
    n1951,
    n1427,
    n1717,
    n1109,
    n766
  );


  xnor
  g1893
  (
    n2091,
    n1027,
    n941,
    n915,
    n1802
  );


  xnor
  g1894
  (
    n2096,
    n805,
    n1291,
    n1639,
    n963
  );


  xnor
  g1895
  (
    n2430,
    n1631,
    n1629,
    n722,
    n1548
  );


  xnor
  g1896
  (
    n2106,
    n1363,
    n1695,
    n916,
    n1450
  );


  nor
  g1897
  (
    n2064,
    n1302,
    n895,
    n872,
    n1248
  );


  xor
  g1898
  (
    n2448,
    n1753,
    n1792,
    n1452,
    n1806
  );


  xor
  g1899
  (
    n2275,
    n1788,
    n1607,
    n1716,
    n1606
  );


  nand
  g1900
  (
    n2409,
    n1719,
    n1100,
    n731,
    n1484
  );


  or
  g1901
  (
    n2367,
    n1553,
    n1060,
    n967,
    n1341
  );


  xnor
  g1902
  (
    n1825,
    n1253,
    n1402,
    n1708,
    n1778
  );


  nor
  g1903
  (
    n1842,
    n1667,
    n1447,
    n695,
    n1562
  );


  and
  g1904
  (
    n1969,
    n1700,
    n1522,
    n1622,
    n1458
  );


  and
  g1905
  (
    n1869,
    n1650,
    n1006,
    n1694,
    n1186
  );


  nor
  g1906
  (
    n1882,
    n1685,
    n1677,
    n1737,
    n676
  );


  nor
  g1907
  (
    n2334,
    n1794,
    n1091,
    n867,
    n822
  );


  nand
  g1908
  (
    n2065,
    n1680,
    n1760,
    n1235,
    n1726
  );


  or
  g1909
  (
    n1980,
    n1221,
    n1412,
    n1463,
    n1641
  );


  or
  g1910
  (
    n2013,
    n953,
    n1445,
    n1199,
    n770
  );


  nand
  g1911
  (
    n2330,
    n814,
    n862,
    n856,
    n1507
  );


  and
  g1912
  (
    n2139,
    n1702,
    n1136,
    n840,
    n1218
  );


  xnor
  g1913
  (
    n2415,
    n1501,
    n1161,
    n802,
    n1186
  );


  nand
  g1914
  (
    n2114,
    n1740,
    n1804,
    n1697,
    n1154
  );


  nor
  g1915
  (
    n1911,
    n876,
    n1809,
    n670,
    n1495
  );


  and
  g1916
  (
    n2257,
    n1165,
    n1752,
    n1723,
    n1007
  );


  nor
  g1917
  (
    n2161,
    n1692,
    n1272,
    n1734,
    n1093
  );


  and
  g1918
  (
    n2166,
    n1765,
    n1244,
    n1801,
    n1126
  );


  or
  g1919
  (
    n2244,
    n852,
    n1371,
    n1310,
    n1008
  );


  xnor
  g1920
  (
    n1891,
    n1042,
    n1571,
    n865,
    n1472
  );


  xor
  g1921
  (
    n2301,
    n1696,
    n1436,
    n1697,
    n1200
  );


  and
  g1922
  (
    KeyWire_0_15,
    n1188,
    n1328,
    n1357,
    n1275
  );


  and
  g1923
  (
    n2314,
    n1569,
    n1020,
    n876,
    n1090
  );


  nand
  g1924
  (
    n2015,
    n1262,
    n739,
    n1122,
    n902
  );


  nor
  g1925
  (
    n1915,
    n1743,
    n845,
    n704,
    n1171
  );


  and
  g1926
  (
    n2286,
    n1633,
    n1324,
    n1678,
    n1794
  );


  or
  g1927
  (
    n2160,
    n1773,
    n1158,
    n1807,
    n911
  );


  nor
  g1928
  (
    n2211,
    n861,
    n1705,
    n1798,
    n1710
  );


  or
  g1929
  (
    KeyWire_0_4,
    n1661,
    n1521,
    n740,
    n1390
  );


  xor
  g1930
  (
    n2181,
    n1515,
    n1174,
    n824,
    n1160
  );


  xnor
  g1931
  (
    n2145,
    n948,
    n1791,
    n1622,
    n1206
  );


  xor
  g1932
  (
    n2311,
    n1467,
    n997,
    n913,
    n1686
  );


  xor
  g1933
  (
    n2477,
    n673,
    n1783,
    n1030,
    n1394
  );


  and
  g1934
  (
    n2467,
    n1185,
    n1677,
    n1704,
    n819
  );


  xnor
  g1935
  (
    n2215,
    n972,
    n1754,
    n1798,
    n1121
  );


  xnor
  g1936
  (
    n2153,
    n1604,
    n853,
    n701,
    n1806
  );


  xor
  g1937
  (
    n2238,
    n1624,
    n1279,
    n1715,
    n1378
  );


  nand
  g1938
  (
    n2165,
    n1106,
    n1418,
    n1271,
    n1521
  );


  nand
  g1939
  (
    n2379,
    n1444,
    n1216,
    n1004,
    n1370
  );


  nand
  g1940
  (
    n2293,
    n748,
    n1597,
    n1595,
    n1524
  );


  xnor
  g1941
  (
    n1990,
    n1735,
    n1145,
    n1639,
    n1349
  );


  xor
  g1942
  (
    n2461,
    n1741,
    n1610,
    n1125,
    n1243
  );


  xor
  g1943
  (
    n2454,
    n1769,
    n851,
    n1540,
    n1624
  );


  nor
  g1944
  (
    n2149,
    n1247,
    n1718,
    n1301,
    n1130
  );


  xnor
  g1945
  (
    n1995,
    n1181,
    n1085,
    n1756,
    n898
  );


  or
  g1946
  (
    n2120,
    n684,
    n831,
    n1111,
    n1603
  );


  and
  g1947
  (
    n2394,
    n861,
    n1069,
    n1724,
    n1128
  );


  or
  g1948
  (
    n2287,
    n1379,
    n1726,
    n1219,
    n1728
  );


  and
  g1949
  (
    n2250,
    n931,
    n699,
    n873,
    n831
  );


  xor
  g1950
  (
    n1904,
    n1286,
    n1256,
    n1541,
    n1630
  );


  xnor
  g1951
  (
    n2289,
    n1176,
    n1668,
    n1780,
    n1181
  );


  or
  g1952
  (
    n2348,
    n1740,
    n870,
    n1806,
    n1687
  );


  xor
  g1953
  (
    n2347,
    n1102,
    n1337,
    n1189,
    n781
  );


  or
  g1954
  (
    n2246,
    n1700,
    n1441,
    n1440,
    n1739
  );


  xor
  g1955
  (
    n2217,
    n775,
    n1078,
    n1688,
    n882
  );


  or
  g1956
  (
    n1970,
    n855,
    n870,
    n1669,
    n1031
  );


  xnor
  g1957
  (
    n1878,
    n1137,
    n1106,
    n1321,
    n884
  );


  nand
  g1958
  (
    n1859,
    n1582,
    n929,
    n961,
    n1295
  );


  nor
  g1959
  (
    n2117,
    n1616,
    n1702,
    n1140,
    n1662
  );


  nand
  g1960
  (
    n1918,
    n1173,
    n987,
    n1071,
    n1763
  );


  nand
  g1961
  (
    n2318,
    n874,
    n1640,
    n885,
    n1672
  );


  xor
  g1962
  (
    n2046,
    n1237,
    n1531,
    n1491,
    n974
  );


  xnor
  g1963
  (
    n2377,
    n1594,
    n1342,
    n1082,
    n1208
  );


  and
  g1964
  (
    n2044,
    n1576,
    n1334,
    n796,
    n1714
  );


  nand
  g1965
  (
    n2162,
    n1642,
    n916,
    n1260,
    n1796
  );


  xor
  g1966
  (
    n2219,
    n1500,
    n1596,
    n1764,
    n1169
  );


  or
  g1967
  (
    n2210,
    n1044,
    n1314,
    n1590,
    n760
  );


  xnor
  g1968
  (
    n2371,
    n1322,
    n1117,
    n1702,
    n1420
  );


  xnor
  g1969
  (
    n2316,
    n1735,
    n1734,
    n1790,
    n1656
  );


  nand
  g1970
  (
    n2305,
    n1007,
    n1692,
    n782,
    n1148
  );


  or
  g1971
  (
    n2074,
    n1657,
    n1040,
    n720,
    n828
  );


  or
  g1972
  (
    n1832,
    n1648,
    n744,
    n959,
    n1778
  );


  nor
  g1973
  (
    n1937,
    n1775,
    n1441,
    n1081,
    n1645
  );


  nor
  g1974
  (
    n2133,
    n1388,
    n1509,
    n1294,
    n982
  );


  nor
  g1975
  (
    n2253,
    n904,
    n1333,
    n1503,
    n1377
  );


  nand
  g1976
  (
    n2245,
    n1116,
    n1444,
    n1013,
    n980
  );


  and
  g1977
  (
    n2375,
    n1211,
    n1746,
    n1585,
    n1058
  );


  or
  g1978
  (
    n2368,
    n1757,
    n1062,
    n1567,
    n1608
  );


  and
  g1979
  (
    n2358,
    n1059,
    n1014,
    n1617,
    n1149
  );


  or
  g1980
  (
    n2029,
    n1682,
    n829,
    n812,
    n1099
  );


  xnor
  g1981
  (
    n2406,
    n903,
    n1101,
    n1333,
    n1528
  );


  xnor
  g1982
  (
    KeyWire_0_17,
    n1806,
    n1762,
    n1589,
    n712
  );


  xor
  g1983
  (
    n2369,
    n845,
    n779,
    n1715,
    n1280
  );


  xnor
  g1984
  (
    n2474,
    n1750,
    n1097,
    n1492,
    n1679
  );


  xnor
  g1985
  (
    n1864,
    n1784,
    n852,
    n1593,
    n1805
  );


  or
  g1986
  (
    n2276,
    n1758,
    n1656,
    n1241,
    n1625
  );


  xnor
  g1987
  (
    n2422,
    n1142,
    n1110,
    n892,
    n1490
  );


  xor
  g1988
  (
    n2119,
    n811,
    n1768,
    n1687,
    n721
  );


  nand
  g1989
  (
    n2351,
    n1620,
    n778,
    n1781,
    n1386
  );


  or
  g1990
  (
    n1964,
    n1025,
    n1398,
    n764,
    n1150
  );


  nand
  g1991
  (
    n1857,
    n1103,
    n1076,
    n711,
    n1759
  );


  xor
  g1992
  (
    n2372,
    n729,
    n1564,
    n857,
    n1254
  );


  or
  g1993
  (
    n2105,
    n1335,
    n1515,
    n1680,
    n901
  );


  or
  g1994
  (
    n2445,
    n1037,
    n672,
    n160,
    n1632
  );


  nor
  g1995
  (
    n2386,
    n686,
    n1758,
    n798
  );


  nand
  g1996
  (
    n2291,
    n1729,
    n1487,
    n1763,
    n1648
  );


  nor
  g1997
  (
    n2437,
    n1022,
    n1459,
    n821,
    n699
  );


  xor
  g1998
  (
    n2227,
    n1797,
    n1127,
    n764,
    n856
  );


  nor
  g1999
  (
    n2271,
    n1729,
    n1660,
    n1698,
    n1172
  );


  or
  g2000
  (
    n2078,
    n956,
    n889,
    n1611,
    n1769
  );


  nand
  g2001
  (
    n1974,
    n687,
    n1326,
    n1760,
    n1488
  );


  and
  g2002
  (
    n1979,
    n1232,
    n1135,
    n1762,
    n1421
  );


  nor
  g2003
  (
    n1981,
    n1483,
    n159,
    n1379,
    n1080
  );


  and
  g2004
  (
    n1924,
    n1669,
    n1527,
    n1520,
    n669
  );


  nand
  g2005
  (
    n1889,
    n1320,
    n1107,
    n1690,
    n1323
  );


  and
  g2006
  (
    n1925,
    n1140,
    n1095,
    n1453,
    n1032
  );


  or
  g2007
  (
    n1926,
    n1711,
    n1244,
    n849,
    n886
  );


  xor
  g2008
  (
    n2285,
    n1670,
    n1800,
    n1400,
    n1205
  );


  xnor
  g2009
  (
    n2053,
    n1306,
    n1786,
    n761,
    n1623
  );


  or
  g2010
  (
    n2118,
    n1320,
    n1602,
    n1020,
    n1395
  );


  nor
  g2011
  (
    n1890,
    n1601,
    n1121,
    n838,
    n1448
  );


  nor
  g2012
  (
    n2396,
    n1759,
    n1466,
    n797,
    n919
  );


  or
  g2013
  (
    n1932,
    n1705,
    n1339,
    n1278,
    n802
  );


  xnor
  g2014
  (
    n1920,
    n970,
    n1745,
    n1693,
    n1755
  );


  nand
  g2015
  (
    n2255,
    n1447,
    n803,
    n1662,
    n1147
  );


  nand
  g2016
  (
    n2143,
    n894,
    n1476,
    n1474,
    n1560
  );


  and
  g2017
  (
    n2233,
    n1676,
    n700,
    n1775,
    n1406
  );


  xor
  g2018
  (
    n1975,
    n996,
    n1721,
    n1424,
    n790
  );


  or
  g2019
  (
    n1850,
    n1786,
    n1187,
    n1550,
    n1087
  );


  xor
  g2020
  (
    n2264,
    n813,
    n719,
    n1204,
    n1592
  );


  or
  g2021
  (
    n1836,
    n1246,
    n1264,
    n1098,
    n1439
  );


  nor
  g2022
  (
    n2121,
    n1626,
    n160,
    n693,
    n1801
  );


  xnor
  g2023
  (
    n1976,
    n1527,
    n1782,
    n976,
    n830
  );


  and
  g2024
  (
    n2023,
    n1583,
    n1711,
    n1734,
    n1146
  );


  nand
  g2025
  (
    n2327,
    n859,
    n1314,
    n1494,
    n941
  );


  nor
  g2026
  (
    n1913,
    n848,
    n1307,
    n1426,
    n1313
  );


  xor
  g2027
  (
    n2212,
    n1356,
    n1751,
    n1511
  );


  or
  g2028
  (
    n2142,
    n1749,
    n1808,
    n949,
    n748
  );


  or
  g2029
  (
    n2164,
    n864,
    n812,
    n1764,
    n1544
  );


  xnor
  g2030
  (
    n2335,
    n1760,
    n1375,
    n1716,
    n1668
  );


  or
  g2031
  (
    n1875,
    n1689,
    n1062,
    n994,
    n914
  );


  or
  g2032
  (
    n2365,
    n680,
    n795,
    n1739,
    n1766
  );


  nor
  g2033
  (
    n1854,
    n1772,
    n1799,
    n984,
    n1258
  );


  xor
  g2034
  (
    n2170,
    n1694,
    n1238,
    n1145,
    n1528
  );


  or
  g2035
  (
    n2236,
    n906,
    n1293,
    n1586,
    n1736
  );


  and
  g2036
  (
    n2397,
    n1507,
    n1250,
    n1362,
    n1478
  );


  nor
  g2037
  (
    n2176,
    n992,
    n1723,
    n1104,
    n1340
  );


  and
  g2038
  (
    n2455,
    n1807,
    n1805,
    n1665,
    n807
  );


  or
  g2039
  (
    n1898,
    n1677,
    n937,
    n951,
    n1132
  );


  nand
  g2040
  (
    KeyWire_0_5,
    n1347,
    n1468,
    n1485,
    n1297
  );


  xor
  g2041
  (
    n1952,
    n1794,
    n1298,
    n763,
    n1712
  );


  xor
  g2042
  (
    n2129,
    n1008,
    n906,
    n1693,
    n1178
  );


  xnor
  g2043
  (
    n1845,
    n800,
    n1353,
    n706,
    n1701
  );


  xnor
  g2044
  (
    n2269,
    n990,
    n1613,
    n773,
    n1655
  );


  xnor
  g2045
  (
    n1983,
    n1398,
    n1215,
    n1579,
    n1654
  );


  nand
  g2046
  (
    n2402,
    n945,
    n1764,
    n1485,
    n981
  );


  and
  g2047
  (
    n2169,
    n1598,
    n1368,
    n1113,
    n1807
  );


  or
  g2048
  (
    n2354,
    n1492,
    n1130,
    n1484,
    n1119
  );


  xnor
  g2049
  (
    n2294,
    n1074,
    n736,
    n1638,
    n1536
  );


  nand
  g2050
  (
    n2098,
    n1736,
    n1019,
    n1175,
    n872
  );


  or
  g2051
  (
    n2355,
    n1745,
    n1808,
    n1112,
    n1255
  );


  xor
  g2052
  (
    n1849,
    n1679,
    n1183,
    n1226,
    n1671
  );


  and
  g2053
  (
    n2247,
    n1581,
    n858,
    n1023,
    n1495
  );


  xnor
  g2054
  (
    n2398,
    n1308,
    n1511,
    n900,
    n1493
  );


  nand
  g2055
  (
    n2475,
    n762,
    n1034,
    n1778,
    n1772
  );


  nand
  g2056
  (
    n2376,
    n1799,
    n1737,
    n881,
    n1803
  );


  or
  g2057
  (
    n2030,
    n1563,
    n1425,
    n1417,
    n689
  );


  xnor
  g2058
  (
    n2333,
    n839,
    n1716,
    n825,
    n1688
  );


  and
  g2059
  (
    n1973,
    n1439,
    n1644,
    n1039,
    n723
  );


  nand
  g2060
  (
    n1945,
    n1407,
    n1785,
    n1457,
    n1437
  );


  and
  g2061
  (
    n2299,
    n1737,
    n1691,
    n1293,
    n1650
  );


  or
  g2062
  (
    n2399,
    n1774,
    n1135,
    n866,
    n1787
  );


  xor
  g2063
  (
    n1843,
    n1543,
    n1255,
    n1584,
    n1458
  );


  xor
  g2064
  (
    n2464,
    n923,
    n1695,
    n1749,
    n1770
  );


  or
  g2065
  (
    n2004,
    n1643,
    n1260,
    n682,
    n891
  );


  xnor
  g2066
  (
    n2082,
    n1801,
    n817,
    n1790,
    n850
  );


  and
  g2067
  (
    n1923,
    n1518,
    n780,
    n846,
    n1600
  );


  xnor
  g2068
  (
    n1886,
    n1800,
    n1330,
    n1430,
    n742
  );


  or
  g2069
  (
    n2195,
    n858,
    n1589,
    n1228,
    n1288
  );


  and
  g2070
  (
    n2007,
    n1705,
    n829,
    n999,
    n1261
  );


  nand
  g2071
  (
    n2037,
    n1064,
    n1216,
    n1796,
    n688
  );


  nor
  g2072
  (
    n2388,
    n1593,
    n965,
    n1227,
    n1403
  );


  nand
  g2073
  (
    n2138,
    n1378,
    n1792,
    n1075,
    n1389
  );


  or
  g2074
  (
    n1942,
    n1572,
    n716,
    n958
  );


  nor
  g2075
  (
    n2259,
    n989,
    n1720,
    n1732,
    n1797
  );


  xor
  g2076
  (
    n2073,
    n1561,
    n1752,
    n1367,
    n741
  );


  and
  g2077
  (
    n2192,
    n1415,
    n901,
    n1343,
    n935
  );


  xnor
  g2078
  (
    n2134,
    n1634,
    n1151,
    n1791,
    n1646
  );


  xor
  g2079
  (
    n2243,
    n679,
    n685,
    n1041,
    n1753
  );


  nor
  g2080
  (
    n1988,
    n1733,
    n1674,
    n758,
    n708
  );


  nor
  g2081
  (
    n1934,
    n791,
    n1638,
    n746,
    n1326
  );


  nand
  g2082
  (
    n1873,
    n1793,
    n1236,
    n1240,
    n1189
  );


  nor
  g2083
  (
    n2323,
    n1073,
    n749,
    n784,
    n722
  );


  or
  g2084
  (
    n2068,
    n1434,
    n721,
    n1448,
    n905
  );


  nand
  g2085
  (
    n1977,
    n960,
    n1587,
    n923,
    n841
  );


  or
  g2086
  (
    n2241,
    n1257,
    n1539,
    n1591,
    n1078
  );


  xor
  g2087
  (
    n2102,
    n1094,
    n1554,
    n1731,
    n1003
  );


  and
  g2088
  (
    n2443,
    n1779,
    n1449,
    n1516,
    n1220
  );


  xnor
  g2089
  (
    n1909,
    n1709,
    n1637,
    n1381,
    n1664
  );


  and
  g2090
  (
    n2393,
    n1552,
    n1761,
    n756,
    n1549
  );


  nand
  g2091
  (
    n2449,
    n828,
    n765,
    n1251,
    n1604
  );


  nor
  g2092
  (
    n2324,
    n999,
    n1767,
    n673,
    n1750
  );


  nand
  g2093
  (
    n2071,
    n1480,
    n1089,
    n681,
    n1095
  );


  xnor
  g2094
  (
    n1838,
    n1012,
    n1682,
    n1129,
    n1417
  );


  and
  g2095
  (
    n1941,
    n991,
    n1658,
    n1787,
    n984
  );


  nor
  g2096
  (
    n2048,
    n1040,
    n1044,
    n1708,
    n925
  );


  nor
  g2097
  (
    n1994,
    n698,
    n860,
    n1165,
    n1242
  );


  and
  g2098
  (
    n1881,
    n1057,
    n1354,
    n917,
    n1605
  );


  or
  g2099
  (
    n1826,
    n1357,
    n1619,
    n1276,
    n1573
  );


  nand
  g2100
  (
    n2444,
    n1674,
    n1026,
    n1005,
    n762
  );


  xnor
  g2101
  (
    n1958,
    n1552,
    n767,
    n1611,
    n1726
  );


  nand
  g2102
  (
    n2479,
    n1296,
    n1506,
    n734,
    n1386
  );


  nand
  g2103
  (
    n2408,
    n907,
    n1365,
    n1601,
    n1696
  );


  xor
  g2104
  (
    n2157,
    n1793,
    n1026,
    n1746,
    n1211
  );


  nand
  g2105
  (
    n2216,
    n1457,
    n891,
    n702,
    n1798
  );


  xnor
  g2106
  (
    n2405,
    n947,
    n1456,
    n1027,
    n1613
  );


  xor
  g2107
  (
    n2447,
    n1699,
    n1653,
    n1738,
    n1595
  );


  nor
  g2108
  (
    n1987,
    n1649,
    n1670,
    n1011,
    n1231
  );


  xnor
  g2109
  (
    n2172,
    n974,
    n1471,
    n1742,
    n695
  );


  nand
  g2110
  (
    n2469,
    n732,
    n1742,
    n1239,
    n1084
  );


  and
  g2111
  (
    n1967,
    n708,
    n1615,
    n1683,
    n1657
  );


  and
  g2112
  (
    n2124,
    n1483,
    n1517,
    n743,
    n932
  );


  xnor
  g2113
  (
    n2088,
    n900,
    n1218,
    n1238,
    n971
  );


  nor
  g2114
  (
    n2186,
    n1797,
    n1741,
    n1246,
    n1579
  );


  nor
  g2115
  (
    n2385,
    n1727,
    n1331,
    n1726,
    n1446
  );


  xor
  g2116
  (
    n2364,
    n770,
    n975,
    n1234,
    n1455
  );


  and
  g2117
  (
    n1855,
    n1002,
    n1187,
    n729,
    n1724
  );


  xnor
  g2118
  (
    n2050,
    n1765,
    n1592,
    n1113,
    n1684
  );


  and
  g2119
  (
    n2081,
    n1539,
    n938,
    n1598,
    n1054
  );


  or
  g2120
  (
    n2194,
    n1566,
    n1459,
    n1291,
    n1234
  );


  and
  g2121
  (
    n1884,
    n1771,
    n1384,
    n875,
    n1033
  );


  nor
  g2122
  (
    n2278,
    n1715,
    n1464,
    n842,
    n1735
  );


  nor
  g2123
  (
    n2038,
    n962,
    n1028,
    n1465,
    n921
  );


  or
  g2124
  (
    n2226,
    n730,
    n1725,
    n1285,
    n1658
  );


  and
  g2125
  (
    n2019,
    n1724,
    n1030,
    n1347,
    n1536
  );


  xor
  g2126
  (
    n1896,
    n1468,
    n1480,
    n1048,
    n709
  );


  and
  g2127
  (
    n2198,
    n926,
    n1356,
    n1400,
    n1615
  );


  and
  g2128
  (
    n2128,
    n1707,
    n1478,
    n1256,
    n1109
  );


  or
  g2129
  (
    KeyWire_0_28,
    n1361,
    n720,
    n1647,
    n1788
  );


  nand
  g2130
  (
    n2021,
    n1163,
    n1407,
    n1668,
    n1212
  );


  nand
  g2131
  (
    n2059,
    n1438,
    n1477,
    n969,
    n1795
  );


  xor
  g2132
  (
    n2235,
    n1370,
    n1785,
    n160,
    n1143
  );


  xnor
  g2133
  (
    n1986,
    n946,
    n1052,
    n1350,
    n1498
  );


  nand
  g2134
  (
    n2197,
    n1137,
    n1773,
    n1122,
    n774
  );


  xor
  g2135
  (
    n1935,
    n792,
    n880,
    n1687,
    n1358
  );


  xnor
  g2136
  (
    n1912,
    n1297,
    n1574,
    n1721,
    n1192
  );


  xor
  g2137
  (
    n2423,
    n1803,
    n1338,
    n1774,
    n1533
  );


  xor
  g2138
  (
    n1861,
    n980,
    n1695,
    n1442,
    n865
  );


  xor
  g2139
  (
    n1940,
    n1534,
    n899,
    n1224,
    n1077
  );


  xnor
  g2140
  (
    n2016,
    n927,
    n1717,
    n1662,
    n910
  );


  nand
  g2141
  (
    n2000,
    n1111,
    n1319,
    n1786,
    n804
  );


  nor
  g2142
  (
    n2132,
    n908,
    n1696,
    n928,
    n1642
  );


  or
  g2143
  (
    n2201,
    n934,
    n1191,
    n1767,
    n888
  );


  xor
  g2144
  (
    n1830,
    n1571,
    n1250,
    n956,
    n1594
  );


  nand
  g2145
  (
    n2027,
    n1655,
    n1374,
    n895,
    n731
  );


  and
  g2146
  (
    n2130,
    n1751,
    n1725,
    n816,
    n1777
  );


  nor
  g2147
  (
    n1851,
    n1299,
    n908,
    n1157,
    n1665
  );


  or
  g2148
  (
    n2039,
    n1279,
    n1188,
    n1488,
    n922
  );


  nand
  g2149
  (
    n1930,
    n1783,
    n1118,
    n1283,
    n933
  );


  or
  g2150
  (
    n1929,
    n1762,
    n1469,
    n1176,
    n1718
  );


  and
  g2151
  (
    n2190,
    n683,
    n979,
    n1701,
    n1789
  );


  nand
  g2152
  (
    n1883,
    n1270,
    n1644,
    n1153,
    n1228
  );


  nand
  g2153
  (
    n2026,
    n1406,
    n818,
    n1082,
    n1635
  );


  xnor
  g2154
  (
    n2182,
    n1798,
    n1736,
    n1427,
    n942
  );


  and
  g2155
  (
    n1962,
    n1262,
    n759,
    n1289,
    n1009
  );


  xnor
  g2156
  (
    n2178,
    n1042,
    n1324,
    n1553,
    n1559
  );


  or
  g2157
  (
    n2434,
    n1182,
    n1223,
    n1272,
    n1551
  );


  and
  g2158
  (
    n2087,
    n1317,
    n1596,
    n1368,
    n1362
  );


  nand
  g2159
  (
    n2248,
    n1131,
    n1413,
    n827,
    n1212
  );


  and
  g2160
  (
    n1835,
    n1519,
    n1692,
    n1269,
    n1164
  );


  xor
  g2161
  (
    n2184,
    n1632,
    n1656,
    n1083,
    n1401
  );


  or
  g2162
  (
    n1876,
    n817,
    n785,
    n1475,
    n789
  );


  nand
  g2163
  (
    n2020,
    n1733,
    n778,
    n1520,
    n1061
  );


  and
  g2164
  (
    n2043,
    n1519,
    n1034,
    n1221,
    n791
  );


  xnor
  g2165
  (
    n2308,
    n1126,
    n1739,
    n1684,
    n961
  );


  and
  g2166
  (
    n1910,
    n1343,
    n1257,
    n836,
    n1794
  );


  or
  g2167
  (
    n2072,
    n1695,
    n789,
    n1336,
    n1734
  );


  nand
  g2168
  (
    n2116,
    n1323,
    n1747,
    n728,
    n1344
  );


  or
  g2169
  (
    n2224,
    n1749,
    n1758,
    n1776,
    n883
  );


  and
  g2170
  (
    n1887,
    n1024,
    n1119,
    n875,
    n1669
  );


  nand
  g2171
  (
    n2010,
    n1088,
    n1676,
    n990,
    n1659
  );


  and
  g2172
  (
    n2356,
    n862,
    n1375,
    n674,
    n1683
  );


  and
  g2173
  (
    n2055,
    n1809,
    n1332,
    n1416,
    n1047
  );


  or
  g2174
  (
    n1984,
    n1727,
    n1284,
    n896,
    n1010
  );


  nor
  g2175
  (
    n1999,
    n1108,
    n1775,
    n1387,
    n1691
  );


  and
  g2176
  (
    n2076,
    n1740,
    n1532,
    n1003,
    n1707
  );


  or
  g2177
  (
    n2061,
    n1305,
    n925,
    n1404,
    n957
  );


  nand
  g2178
  (
    n2425,
    n847,
    n1681,
    n1662,
    n890
  );


  nand
  g2179
  (
    n2111,
    n1428,
    n989,
    n1546,
    n1555
  );


  or
  g2180
  (
    n2387,
    n1697,
    n1325,
    n777,
    n1118
  );


  xnor
  g2181
  (
    n2432,
    n954,
    n952,
    n1710,
    n1674
  );


  or
  g2182
  (
    n1829,
    n1396,
    n1384,
    n765,
    n713
  );


  or
  g2183
  (
    n2380,
    n1207,
    n1175,
    n1306,
    n1647
  );


  or
  g2184
  (
    n2251,
    n1446,
    n1265,
    n1796,
    n1486
  );


  nor
  g2185
  (
    n2320,
    n1259,
    n1428,
    n1454,
    n1161
  );


  xor
  g2186
  (
    n2095,
    n675,
    n815,
    n1573,
    n847
  );


  xor
  g2187
  (
    n2470,
    n739,
    n919,
    n1253,
    n1366
  );


  and
  g2188
  (
    n2453,
    n1649,
    n776,
    n1550,
    n962
  );


  nor
  g2189
  (
    n2101,
    n944,
    n1634,
    n1249,
    n1419
  );


  and
  g2190
  (
    n2451,
    n822,
    n1081,
    n1105,
    n973
  );


  xor
  g2191
  (
    n2115,
    n775,
    n907,
    n950,
    n771
  );


  and
  g2192
  (
    n2414,
    n1694,
    n1435,
    n786,
    n1740
  );


  xnor
  g2193
  (
    n2389,
    n1789,
    n1170,
    n1767,
    n1303
  );


  nand
  g2194
  (
    n2222,
    n1790,
    n1771,
    n1743,
    n1315
  );


  nand
  g2195
  (
    n2214,
    n1657,
    n1763,
    n1209,
    n1050
  );


  xor
  g2196
  (
    n2353,
    n692,
    n1661,
    n914,
    n949
  );


  and
  g2197
  (
    n2254,
    n857,
    n959,
    n1143,
    n1312
  );


  or
  g2198
  (
    n1868,
    n1070,
    n986,
    n1139,
    n1167
  );


  nand
  g2199
  (
    n2411,
    n683,
    n696,
    n1530,
    n1681
  );


  xnor
  g2200
  (
    n1971,
    n794,
    n1016,
    n768,
    n1599
  );


  xnor
  g2201
  (
    n2462,
    n705,
    n1535,
    n1466,
    n1281
  );


  or
  g2202
  (
    n2042,
    n1677,
    n725,
    n1048,
    n738
  );


  or
  g2203
  (
    n2199,
    n1718,
    n1129,
    n1073,
    n1077
  );


  or
  g2204
  (
    n2062,
    n833,
    n678,
    n1780,
    n1545
  );


  xor
  g2205
  (
    n2054,
    n1748,
    n755,
    n1068,
    n842
  );


  xnor
  g2206
  (
    n1959,
    n707,
    n1790,
    n1781,
    n1727
  );


  and
  g2207
  (
    n2086,
    n1383,
    n1731,
    n1267,
    n1679
  );


  and
  g2208
  (
    n2465,
    n1076,
    n808,
    n1644,
    n1259
  );


  xor
  g2209
  (
    n2079,
    n1093,
    n1423,
    n986,
    n1300
  );


  nand
  g2210
  (
    n2329,
    n1318,
    n1697,
    n1434,
    n1132
  );


  xnor
  g2211
  (
    n2144,
    n1245,
    n1666,
    n1064,
    n733
  );


  or
  g2212
  (
    n1944,
    n1772,
    n1142,
    n1196,
    n1252
  );


  and
  g2213
  (
    n2304,
    n1380,
    n1531,
    n1655,
    n1070
  );


  and
  g2214
  (
    n2126,
    n1192,
    n1199,
    n1363,
    n1351
  );


  xor
  g2215
  (
    n2374,
    n1355,
    n1804,
    n1000,
    n784
  );


  or
  g2216
  (
    n1847,
    n1031,
    n1114,
    n978,
    n1663
  );


  xnor
  g2217
  (
    KeyWire_0_11,
    n1226,
    n1086,
    n1501,
    n904
  );


  or
  g2218
  (
    n2361,
    n928,
    n1012,
    n1731,
    n1766
  );


  or
  g2219
  (
    n2262,
    n1001,
    n884,
    n1367,
    n1664
  );


  nand
  g2220
  (
    n2051,
    n1709,
    n1421,
    n1105,
    n1410
  );


  xnor
  g2221
  (
    n1936,
    n1585,
    n1138,
    n1243,
    n1523
  );


  nor
  g2222
  (
    n2084,
    n1739,
    n803,
    n1663,
    n1021
  );


  or
  g2223
  (
    n2225,
    n869,
    n1037,
    n1166,
    n1686
  );


  nor
  g2224
  (
    n2473,
    n1701,
    n889,
    n1094,
    n1738
  );


  xnor
  g2225
  (
    n2163,
    n1750,
    n1672,
    n1438,
    n883
  );


  nand
  g2226
  (
    n2298,
    n805,
    n1728,
    n1752,
    n1393
  );


  and
  g2227
  (
    n2331,
    n1678,
    n1360,
    n1371,
    n1282
  );


  nor
  g2228
  (
    n1998,
    n1452,
    n1201,
    n1433,
    n1011
  );


  xor
  g2229
  (
    n1905,
    n1201,
    n1445,
    n751,
    n1568
  );


  xor
  g2230
  (
    n2417,
    n1648,
    n1733,
    n1337,
    n711
  );


  nand
  g2231
  (
    n1888,
    n1770,
    n1230,
    n741,
    n1437
  );


  nor
  g2232
  (
    n2392,
    n715,
    n1633,
    n1787,
    n1312
  );


  and
  g2233
  (
    n2229,
    n1436,
    n937,
    n1290,
    n1397
  );


  xor
  g2234
  (
    n2457,
    n1364,
    n953,
    n1276,
    n1685
  );


  nand
  g2235
  (
    n2066,
    n1414,
    n160,
    n1387,
    n1036
  );


  xnor
  g2236
  (
    n1966,
    n1565,
    n1052,
    n868,
    n1197
  );


  and
  g2237
  (
    n1927,
    n1359,
    n840,
    n1538,
    n855
  );


  xnor
  g2238
  (
    n2427,
    n909,
    n686,
    n723,
    n1233
  );


  nand
  g2239
  (
    n2228,
    n783,
    n1757,
    n1623,
    n1653
  );


  nor
  g2240
  (
    n2303,
    n774,
    n1391,
    n806,
    n1802
  );


  xor
  g2241
  (
    n2041,
    n968,
    n950,
    n851,
    n1047
  );


  xor
  g2242
  (
    n2322,
    n1578,
    n780,
    n1667,
    n1789
  );


  or
  g2243
  (
    n2306,
    n1741,
    n1730,
    n1514,
    n1747
  );


  or
  g2244
  (
    n1831,
    n1626,
    n841,
    n1795,
    n1704
  );


  and
  g2245
  (
    n2209,
    n1510,
    n1788,
    n752,
    n1360
  );


  xor
  g2246
  (
    n1844,
    n1502,
    n1411,
    n1494,
    n690
  );


  and
  g2247
  (
    n2350,
    n1050,
    n1719,
    n1369,
    n1651
  );


  nor
  g2248
  (
    n2031,
    n1451,
    n1744,
    n1526,
    n1802
  );


  nor
  g2249
  (
    n2183,
    n1685,
    n1369,
    n1655,
    n1719
  );


  or
  g2250
  (
    n2292,
    n1743,
    n1557,
    n1273,
    n1489
  );


  xor
  g2251
  (
    n2272,
    n1385,
    n1575,
    n1462,
    n1659
  );


  and
  g2252
  (
    n2261,
    n1619,
    n1300,
    n893,
    n1680
  );


  nand
  g2253
  (
    n1957,
    n1693,
    n1393,
    n1014,
    n998
  );


  and
  g2254
  (
    n2390,
    n1222,
    n783,
    n697,
    n1731
  );


  xor
  g2255
  (
    n2123,
    n1461,
    n735,
    n924,
    n1660
  );


  nand
  g2256
  (
    n2342,
    n1699,
    n726,
    n1647,
    n1738
  );


  or
  g2257
  (
    n2263,
    n846,
    n1542,
    n1045,
    n1000
  );


  or
  g2258
  (
    n2313,
    n1287,
    n1049,
    n786,
    n1170
  );


  or
  g2259
  (
    n2234,
    n931,
    n1098,
    n1498,
    n1159
  );


  xor
  g2260
  (
    n2063,
    n844,
    n982,
    n1516,
    n1053
  );


  nand
  g2261
  (
    n1917,
    n1666,
    n1712,
    n1704,
    n1038
  );


  nor
  g2262
  (
    n1946,
    n712,
    n1230,
    n1504,
    n1194
  );


  nor
  g2263
  (
    n2420,
    n1394,
    n1141,
    n738,
    n1247
  );


  and
  g2264
  (
    n2022,
    n1152,
    n1703,
    n1673,
    n772
  );


  xor
  g2265
  (
    n2336,
    n979,
    n1631,
    n1723,
    n785
  );


  or
  g2266
  (
    n2125,
    n939,
    n1486,
    n1759,
    n969
  );


  nor
  g2267
  (
    n1902,
    n1331,
    n1473,
    n1178,
    n1167
  );


  xor
  g2268
  (
    n2284,
    n1041,
    n1781,
    n1474,
    n1508
  );


  nor
  g2269
  (
    n2155,
    n1522,
    n1627,
    n815,
    n897
  );


  and
  g2270
  (
    n2332,
    n1194,
    n1152,
    n781,
    n1409
  );


  xnor
  g2271
  (
    n1900,
    n709,
    n1679,
    n1614,
    n1791
  );


  xnor
  g2272
  (
    n2085,
    n1392,
    n1713,
    n1198,
    n1349
  );


  and
  g2273
  (
    n2413,
    n838,
    n1756,
    n926,
    n1784
  );


  and
  g2274
  (
    n2442,
    n957,
    n1223,
    n1525,
    n1411
  );


  nor
  g2275
  (
    n2426,
    n795,
    n1180,
    n1233,
    n892
  );


  and
  g2276
  (
    n2419,
    n801,
    n1408,
    n942,
    n1664
  );


  xor
  g2277
  (
    n2058,
    n1133,
    n1292,
    n1086,
    n886
  );


  or
  g2278
  (
    n1885,
    n1392,
    n1354,
    n834,
    n1778
  );


  xor
  g2279
  (
    n2049,
    n1177,
    n674,
    n940,
    n776
  );


  xor
  g2280
  (
    KeyWire_0_9,
    n1699,
    n1645,
    n1138,
    n754
  );


  xnor
  g2281
  (
    n2359,
    n1741,
    n1625,
    n1742,
    n1666
  );


  xnor
  g2282
  (
    n2418,
    n830,
    n879,
    n820,
    n1405
  );


  xor
  g2283
  (
    n2136,
    n1759,
    n1612,
    n1342,
    n1039
  );


  nor
  g2284
  (
    n2097,
    n1747,
    n1327,
    n1707,
    n1057
  );


  or
  g2285
  (
    n1955,
    n1072,
    n1418,
    n854,
    n1804
  );


  nand
  g2286
  (
    n1866,
    n745,
    n1538,
    n866,
    n1748
  );


  nand
  g2287
  (
    n2147,
    n687,
    n1770,
    n1663,
    n1751
  );


  xor
  g2288
  (
    n2179,
    n1706,
    n1590,
    n668,
    n1618
  );


  nor
  g2289
  (
    n2277,
    n1203,
    n1666,
    n1115,
    n1353
  );


  xor
  g2290
  (
    n1870,
    n1772,
    n1768,
    n1065,
    n1621
  );


  nand
  g2291
  (
    n1865,
    n1220,
    n1542,
    n1795,
    n1561
  );


  xnor
  g2292
  (
    n1943,
    n1650,
    n843,
    n1776,
    n1621
  );


  nand
  g2293
  (
    n1828,
    n1304,
    n1708,
    n1541,
    n1431
  );


  or
  g2294
  (
    n2416,
    n1651,
    n1652,
    n1487,
    n799
  );


  xor
  g2295
  (
    n2174,
    n971,
    n1391,
    n1785,
    n1668
  );


  nor
  g2296
  (
    n2188,
    n1543,
    n1101,
    n947,
    n1746
  );


  xnor
  g2297
  (
    n1895,
    n988,
    n1364,
    n1540,
    n912
  );


  or
  g2298
  (
    n1997,
    n1477,
    n833,
    n1537,
    n1072
  );


  or
  g2299
  (
    n1841,
    n819,
    n796,
    n1415,
    n769
  );


  nor
  g2300
  (
    n2352,
    n1745,
    n772,
    n1544,
    n1648
  );


  and
  g2301
  (
    n2378,
    n1263,
    n1689,
    n1774,
    n1600
  );


  nor
  g2302
  (
    n2295,
    n1656,
    n1530,
    n1261,
    n898
  );


  xnor
  g2303
  (
    n2267,
    n1729,
    n1672,
    n1351,
    n832
  );


  and
  g2304
  (
    n1852,
    n1124,
    n1713,
    n714,
    n1464
  );


  or
  g2305
  (
    n2328,
    n1156,
    n1479,
    n1456,
    n1777
  );


  xor
  g2306
  (
    n2403,
    n704,
    n1024,
    n1308,
    n1676
  );


  or
  g2307
  (
    n1963,
    n1051,
    n779,
    n800,
    n1043
  );


  nor
  g2308
  (
    n2025,
    n750,
    n1006,
    n903,
    n1390
  );


  nand
  g2309
  (
    n1872,
    n1801,
    n1732,
    n1267,
    n1422
  );


  xor
  g2310
  (
    n2113,
    n871,
    n1277,
    n943,
    n1809
  );


  xnor
  g2311
  (
    n2011,
    n826,
    n1156,
    n992,
    n1381
  );


  xor
  g2312
  (
    n2193,
    n1736,
    n694,
    n1325,
    n1307
  );


  nand
  g2313
  (
    n2435,
    n1174,
    n1753,
    n1335,
    n1021
  );


  and
  g2314
  (
    n2045,
    n1009,
    n939,
    n1185,
    n787
  );


  nor
  g2315
  (
    n2231,
    n1512,
    n1252,
    n899,
    n1068
  );


  nand
  g2316
  (
    n2107,
    n1777,
    n1754,
    n1784,
    n1657
  );


  and
  g2317
  (
    n2460,
    n955,
    n1529,
    n1313,
    n1730
  );


  nor
  g2318
  (
    n2436,
    n1557,
    n797,
    n1264,
    n987
  );


  and
  g2319
  (
    n1903,
    n1282,
    n848,
    n804,
    n1159
  );


  xnor
  g2320
  (
    n2309,
    n1453,
    n806,
    n1757,
    n1248
  );


  xor
  g2321
  (
    n2070,
    n1735,
    n1577,
    n1294,
    n1559
  );


  nand
  g2322
  (
    n2452,
    n1620,
    n837,
    n703,
    n1432
  );


  and
  g2323
  (
    n2208,
    n1345,
    n1748,
    n1092,
    n1580
  );


  nand
  g2324
  (
    n2440,
    n993,
    n1649,
    n1268,
    n1805
  );


  and
  g2325
  (
    n2122,
    n1744,
    n1664,
    n1075,
    n766
  );


  xnor
  g2326
  (
    n2110,
    n1551,
    n1532,
    n1200,
    n1554
  );


  xor
  g2327
  (
    n2196,
    n1205,
    n1651,
    n1286,
    n1146
  );


  nor
  g2328
  (
    n2360,
    n1377,
    n1779,
    n954,
    n978
  );


  nand
  g2329
  (
    n2441,
    n1208,
    n1120,
    n1237,
    n1322
  );


  or
  g2330
  (
    n2156,
    n1645,
    n1654,
    n769,
    n1703
  );


  nor
  g2331
  (
    n2207,
    n1500,
    n1420,
    n1665,
    n1410
  );


  nor
  g2332
  (
    n2302,
    n1045,
    n1083,
    n1397,
    n1151
  );


  nand
  g2333
  (
    n1856,
    n1184,
    n1706,
    n877,
    n894
  );


  nor
  g2334
  (
    n2381,
    n837,
    n793,
    n1350,
    n1066
  );


  xnor
  g2335
  (
    n2024,
    n1576,
    n843,
    n823,
    n1035
  );


  or
  g2336
  (
    n2008,
    n813,
    n1570,
    n1016,
    n1202
  );


  xor
  g2337
  (
    n2439,
    n1067,
    n1616,
    n995,
    n1534
  );


  or
  g2338
  (
    n1960,
    n1775,
    n1640,
    n1513,
    n1107
  );


  and
  g2339
  (
    n2218,
    n1564,
    n1709,
    n1555,
    n934
  );


  xnor
  g2340
  (
    n1922,
    n1781,
    n1627,
    n1336,
    n710
  );


  and
  g2341
  (
    n1950,
    n896,
    n1779,
    n1701,
    n834
  );


  xnor
  g2342
  (
    n1827,
    n735,
    n1686,
    n1533,
    n1688
  );


  nor
  g2343
  (
    n2410,
    n1097,
    n849,
    n1795,
    n1797
  );


  and
  g2344
  (
    n1853,
    n1535,
    n702,
    n1509,
    n1628
  );


  or
  g2345
  (
    n1961,
    n807,
    n1749,
    n988,
    n1661
  );


  nand
  g2346
  (
    n2282,
    n1738,
    n1777,
    n878,
    n1117
  );


  nand
  g2347
  (
    n2321,
    n1768,
    n1424,
    n1213,
    n1581
  );


  xor
  g2348
  (
    n2093,
    n1302,
    n1762,
    n1177,
    n1096
  );


  xor
  g2349
  (
    n2137,
    n1475,
    n1173,
    n1295,
    n743
  );


  nand
  g2350
  (
    n1947,
    n968,
    n1727,
    n1285,
    n1673
  );


  nand
  g2351
  (
    n2339,
    n685,
    n742,
    n1641,
    n1203
  );


  or
  g2352
  (
    n1908,
    n1792,
    n1061,
    n1732,
    n1465
  );


  or
  g2353
  (
    n2450,
    n1809,
    n1609,
    n1301,
    n1785
  );


  xor
  g2354
  (
    n2395,
    n701,
    n1388,
    n696,
    n1653
  );


  or
  g2355
  (
    n2141,
    n1096,
    n1729,
    n768,
    n1433
  );


  xnor
  g2356
  (
    n2135,
    n981,
    n985,
    n1692,
    n757
  );


  xnor
  g2357
  (
    n2221,
    n827,
    n1376,
    n1497,
    n788
  );


  and
  g2358
  (
    n2370,
    n1063,
    n1761,
    n1240,
    n966
  );


  nand
  g2359
  (
    n1989,
    n1251,
    n1183,
    n824,
    n705
  );


  nand
  g2360
  (
    n2240,
    n1219,
    n1716,
    n820,
    n1753
  );


  xnor
  g2361
  (
    n1949,
    n1796,
    n1309,
    n1646,
    n1125
  );


  nor
  g2362
  (
    n2185,
    n1019,
    n1577,
    n1134,
    n1275
  );


  or
  g2363
  (
    n2383,
    n1786,
    n1709,
    n1669,
    n707
  );


  nor
  g2364
  (
    n2472,
    n1687,
    n1339,
    n1022,
    n927
  );


  and
  g2365
  (
    n2152,
    n1711,
    n1471,
    n1304,
    n750
  );


  nand
  g2366
  (
    n2005,
    n1168,
    n1249,
    n1743,
    n1490
  );


  and
  g2367
  (
    n2213,
    n1158,
    n1202,
    n1808,
    n1035
  );


  or
  g2368
  (
    n2471,
    n1612,
    n835,
    n1341,
    n1675
  );


  or
  g2369
  (
    KeyWire_0_13,
    n1703,
    n1505,
    n1023,
    n1636
  );


  or
  g2370
  (
    n2242,
    n1744,
    n1628,
    n1180,
    n1460
  );


  nor
  g2371
  (
    n2057,
    n963,
    n1704,
    n1025,
    n1303
  );


  and
  g2372
  (
    n2052,
    n1689,
    n998,
    n1214,
    n753
  );


  xor
  g2373
  (
    n1993,
    n1430,
    n1217,
    n1164,
    n1499
  );


  nand
  g2374
  (
    n2173,
    n1670,
    n758,
    n1610,
    n1330
  );


  and
  g2375
  (
    n2206,
    n1071,
    n1526,
    n1562,
    n975
  );


  xnor
  g2376
  (
    n2001,
    n1087,
    n977,
    n1546,
    n1046
  );


  and
  g2377
  (
    n2256,
    n1565,
    n1015,
    n1499,
    n706
  );


  xnor
  g2378
  (
    n2296,
    n1232,
    n754,
    n1268,
    n809
  );


  nand
  g2379
  (
    n2326,
    n1429,
    n1265,
    n1730,
    n854
  );


  or
  g2380
  (
    n2424,
    n1051,
    n952,
    n1069,
    n1545
  );


  and
  g2381
  (
    n2230,
    n825,
    n1793,
    n678,
    n1372
  );


  nand
  g2382
  (
    n1906,
    n810,
    n1123,
    n1586,
    n983
  );


  or
  g2383
  (
    n2400,
    n1241,
    n1789,
    n1683,
    n1481
  );


  or
  g2384
  (
    n2239,
    n718,
    n1717,
    n1329,
    n794
  );


  nand
  g2385
  (
    n2463,
    n1690,
    n1348,
    n1359,
    n1321
  );


  or
  g2386
  (
    n2080,
    n1089,
    n782,
    n727,
    n1134
  );


  and
  g2387
  (
    n2012,
    n810,
    n1685,
    n1396,
    n1773
  );


  and
  g2388
  (
    n1897,
    n918,
    n1575,
    n1191,
    n1496
  );


  nand
  g2389
  (
    n2108,
    n839,
    n1690,
    n1803,
    n874
  );


  and
  g2390
  (
    n2148,
    n860,
    n1112,
    n1455,
    n1382
  );


  and
  g2391
  (
    n2252,
    n1766,
    n1319,
    n1744,
    n1100
  );


  nor
  g2392
  (
    n1954,
    n1273,
    n1054,
    n1658,
    n1292
  );


  xor
  g2393
  (
    n1907,
    n1043,
    n868,
    n1454,
    n930
  );


  xor
  g2394
  (
    n2083,
    n717,
    n1720,
    n933,
    n1614
  );


  nand
  g2395
  (
    n2014,
    n771,
    n1722,
    n1355,
    n1690
  );


  xor
  g2396
  (
    n2146,
    n1644,
    n1733,
    n1144,
    n1001
  );


  and
  g2397
  (
    n1972,
    n1366,
    n985,
    n1652,
    n751
  );


  nor
  g2398
  (
    n2312,
    n1206,
    n1416,
    n1395,
    n1782
  );


  and
  g2399
  (
    n2466,
    n1103,
    n1346,
    n1799,
    n1810
  );


  xnor
  g2400
  (
    n2003,
    n1405,
    n757,
    n1707,
    n1617
  );


  or
  g2401
  (
    n2341,
    n1672,
    n1467,
    n1710,
    n1150
  );


  nor
  g2402
  (
    n2202,
    n1144,
    n1755,
    n964,
    n1588
  );


  and
  g2403
  (
    n1880,
    n966,
    n960,
    n893,
    n1671
  );


  nor
  g2404
  (
    n2090,
    n1682,
    n710,
    n1718,
    n1274
  );


  nor
  g2405
  (
    n2428,
    n1373,
    n1699,
    n1443,
    n1168
  );


  and
  g2406
  (
    n2200,
    n698,
    n940,
    n1425,
    n1791
  );


  nand
  g2407
  (
    n2035,
    n1597,
    n1380,
    n1059,
    n1675
  );


  or
  g2408
  (
    n1839,
    n1728,
    n880,
    n680,
    n1102
  );


  and
  g2409
  (
    n2220,
    n1412,
    n1229,
    n755,
    n692
  );


  xor
  g2410
  (
    n1837,
    n1114,
    n1389,
    n1462,
    n873
  );


  and
  g2411
  (
    n1916,
    n744,
    n1332,
    n1236,
    n1179
  );


  or
  g2412
  (
    n2310,
    n1283,
    n713,
    n1643,
    n1525
  );


  xnor
  g2413
  (
    n1871,
    n1503,
    n1479,
    n1517,
    n1688
  );


  or
  g2414
  (
    n2357,
    n1587,
    n1783,
    n1776,
    n1482
  );


  xor
  g2415
  (
    n2315,
    n1758,
    n1404,
    n1808,
    n1769
  );


  xnor
  g2416
  (
    n2456,
    n740,
    n1686,
    n1429,
    n1190
  );


  xor
  g2417
  (
    n2431,
    n1635,
    n1374,
    n850,
    n1663
  );


  nor
  g2418
  (
    n2363,
    n1810,
    n1764,
    n1683,
    n691
  );


  and
  g2419
  (
    n2056,
    n759,
    n977,
    n1646,
    n836
  );


  xnor
  g2420
  (
    n2089,
    n793,
    n997,
    n1348,
    n1317
  );


  and
  g2421
  (
    n2191,
    n1712,
    n1756,
    n690,
    n1547
  );


  nand
  g2422
  (
    n2175,
    n734,
    n724,
    n1193,
    n1700
  );


  or
  g2423
  (
    n1921,
    n1767,
    n1340,
    n1671,
    n1684
  );


  xnor
  g2424
  (
    n2260,
    n1698,
    n1029,
    n1645,
    n909
  );


  nand
  g2425
  (
    n2109,
    n1160,
    n1556,
    n1649,
    n1225
  );


  or
  g2426
  (
    n2187,
    n1153,
    n1055,
    n1450,
    n1745
  );


  nand
  g2427
  (
    n2018,
    n897,
    n905,
    n1805,
    n912
  );


  xor
  g2428
  (
    n1914,
    n944,
    n1419,
    n1017,
    n1334
  );


  nor
  g2429
  (
    n2223,
    n1225,
    n1358,
    n1472,
    n1442
  );


  or
  g2430
  (
    n1834,
    n887,
    n1529,
    n1154,
    n1748
  );


  xor
  g2431
  (
    n2476,
    n1460,
    n1316,
    n1629,
    n1618
  );


  xor
  g2432
  (
    n2391,
    n1780,
    n1722,
    n1148,
    n1676
  );


  nor
  g2433
  (
    n2006,
    n1678,
    n761,
    n737,
    n1694
  );


  and
  g2434
  (
    n2203,
    n1310,
    n1514,
    n1209,
    n1723
  );


  xor
  g2435
  (
    n1928,
    n887,
    n1757,
    n1449,
    n714
  );


  or
  g2436
  (
    n2032,
    n1523,
    n1588,
    n1242,
    n863
  );


  nor
  g2437
  (
    n1899,
    n1804,
    n1769,
    n689,
    n955
  );


  xor
  g2438
  (
    n1956,
    n1800,
    n1667,
    n691,
    n1504
  );


  xor
  g2439
  (
    KeyWire_0_18,
    n1155,
    n1691,
    n1774,
    n1673
  );


  or
  g2440
  (
    n2384,
    n1266,
    n1771,
    n1502,
    n697
  );


  and
  g2441
  (
    n2438,
    n1787,
    n1090,
    n1659,
    n1493
  );


  or
  g2442
  (
    n1931,
    n1269,
    n1722,
    n749,
    n1131
  );


  nor
  g2443
  (
    n2337,
    n823,
    n1013,
    n1422,
    n700
  );


  nor
  g2444
  (
    n2171,
    n1365,
    n726,
    n1675,
    n1609
  );


  nand
  g2445
  (
    n2362,
    n945,
    n1768,
    n930,
    n753
  );


  nand
  g2446
  (
    n2340,
    n1658,
    n1345,
    n1327,
    n682
  );


  nor
  g2447
  (
    n2480,
    n657,
    n659
  );


  nor
  g2448
  (
    n2484,
    n1832,
    n658,
    n656,
    n660
  );


  nand
  g2449
  (
    n2482,
    n1831,
    n659,
    n656
  );


  xnor
  g2450
  (
    n2483,
    n660,
    n1825,
    n657
  );


  and
  g2451
  (
    n2481,
    n655,
    n660,
    n659
  );


  xnor
  g2452
  (
    n2486,
    n657,
    n661,
    n656,
    n658
  );


  nand
  g2453
  (
    n2485,
    n1829,
    n656,
    n658,
    n1830
  );


  nor
  g2454
  (
    n2487,
    n1828,
    n1826,
    n1827,
    n658
  );


  buf
  g2455
  (
    n2492,
    n662
  );


  buf
  g2456
  (
    n2491,
    n662
  );


  buf
  g2457
  (
    n2493,
    n2485
  );


  nor
  g2458
  (
    n2494,
    n663,
    n662,
    n2482
  );


  nand
  g2459
  (
    n2488,
    n2483,
    n2486,
    n661,
    n2484
  );


  xor
  g2460
  (
    n2490,
    n2481,
    n662,
    n2480,
    n661
  );


  xnor
  g2461
  (
    n2489,
    n661,
    n663
  );


  buf
  g2462
  (
    n2500,
    n2491
  );


  not
  g2463
  (
    n2510,
    n2490
  );


  not
  g2464
  (
    n2514,
    n2490
  );


  buf
  g2465
  (
    n2513,
    n2490
  );


  not
  g2466
  (
    n2495,
    n2491
  );


  not
  g2467
  (
    n2511,
    n2489
  );


  not
  g2468
  (
    n2501,
    n2492
  );


  not
  g2469
  (
    n2508,
    n2492
  );


  buf
  g2470
  (
    n2506,
    n2492
  );


  buf
  g2471
  (
    n2498,
    n2488
  );


  buf
  g2472
  (
    n2505,
    n2491
  );


  not
  g2473
  (
    n2502,
    n2490
  );


  buf
  g2474
  (
    n2504,
    n2489
  );


  not
  g2475
  (
    n2509,
    n2488
  );


  buf
  g2476
  (
    n2503,
    n2491
  );


  buf
  g2477
  (
    n2512,
    n2488
  );


  buf
  g2478
  (
    n2507,
    n2489
  );


  not
  g2479
  (
    n2497,
    n2489
  );


  not
  g2480
  (
    n2496,
    n2492
  );


  not
  g2481
  (
    n2499,
    n2488
  );


  xnor
  g2482
  (
    n2529,
    n1869,
    n1840
  );


  or
  g2483
  (
    n2515,
    n2497,
    n1841,
    n2496,
    n1866
  );


  and
  g2484
  (
    n2520,
    n1858,
    n1857,
    n1871,
    n2496
  );


  xnor
  g2485
  (
    n2519,
    n1843,
    n1862,
    n2495,
    n2496
  );


  and
  g2486
  (
    n2517,
    n1874,
    n2497,
    n2498,
    n1852
  );


  xnor
  g2487
  (
    n2516,
    n1872,
    n1846,
    n1854,
    n1868
  );


  nand
  g2488
  (
    n2524,
    n1839,
    n1845,
    n1856,
    n1836
  );


  xor
  g2489
  (
    n2528,
    n2495,
    n1842,
    n1838,
    n1853
  );


  nand
  g2490
  (
    n2522,
    n2496,
    n2497,
    n1847,
    n1849
  );


  and
  g2491
  (
    n2521,
    n1875,
    n1861,
    n1837,
    n1844
  );


  and
  g2492
  (
    n2518,
    n1833,
    n1870,
    n2498,
    n2497
  );


  xnor
  g2493
  (
    n2527,
    n1863,
    n1835,
    n1859,
    n2495
  );


  and
  g2494
  (
    n2526,
    n1867,
    n1855,
    n2498,
    n1873
  );


  xnor
  g2495
  (
    n2525,
    n1860,
    n1865,
    n1848,
    n1850
  );


  and
  g2496
  (
    n2523,
    n1834,
    n1851,
    n1864,
    n2495
  );


  or
  g2497
  (
    n2550,
    n1927,
    n2525,
    n1919,
    n1884
  );


  nand
  g2498
  (
    n2556,
    n1891,
    n1923,
    n2526,
    n2521
  );


  nor
  g2499
  (
    n2547,
    n1883,
    n1899,
    n1896,
    n1937
  );


  xnor
  g2500
  (
    n2548,
    n2493,
    n2493,
    n1897,
    n1902
  );


  xor
  g2501
  (
    n2535,
    n1908,
    n1885,
    n2518,
    n1913
  );


  xnor
  g2502
  (
    n2530,
    n2521,
    n1879,
    n2494,
    n2524
  );


  nand
  g2503
  (
    n2555,
    n1938,
    n2523,
    n1910,
    n1929
  );


  xor
  g2504
  (
    n2536,
    n2515,
    n2494,
    n1889,
    n2523
  );


  nand
  g2505
  (
    n2549,
    n2525,
    n1918,
    n1931,
    n2494
  );


  or
  g2506
  (
    n2543,
    n1909,
    n1921,
    n1930,
    n1912
  );


  nor
  g2507
  (
    n2551,
    n1876,
    n2520,
    n1935,
    n1936
  );


  xnor
  g2508
  (
    n2553,
    n1890,
    n1916,
    n1886,
    n1907
  );


  xnor
  g2509
  (
    n2539,
    n1941,
    n1881,
    n1926,
    n1895
  );


  nand
  g2510
  (
    n2533,
    n1915,
    n2525,
    n2516,
    n2524
  );


  or
  g2511
  (
    n2554,
    n2526,
    n2522,
    n1900,
    n2524
  );


  or
  g2512
  (
    n2531,
    n2517,
    n1878,
    n2527,
    n2493
  );


  xor
  g2513
  (
    n2546,
    n1877,
    n1924,
    n1928,
    n1925
  );


  xnor
  g2514
  (
    n2542,
    n2522,
    n2523,
    n1882,
    n2521
  );


  xnor
  g2515
  (
    n2538,
    n1940,
    n1904,
    n1892,
    n2519
  );


  xnor
  g2516
  (
    n2552,
    n1922,
    n2523,
    n1893,
    n1880
  );


  or
  g2517
  (
    n2541,
    n2521,
    n1914,
    n2522,
    n2525
  );


  xnor
  g2518
  (
    n2534,
    n1894,
    n1933,
    n1934,
    n1903
  );


  or
  g2519
  (
    n2532,
    n1911,
    n2522,
    n1901,
    n2526
  );


  or
  g2520
  (
    n2540,
    n2526,
    n2524,
    n1905,
    n1898
  );


  or
  g2521
  (
    n2537,
    n2519,
    n1917,
    n2487,
    n1939
  );


  nand
  g2522
  (
    n2544,
    n2520,
    n1920,
    n1887,
    n1888
  );


  and
  g2523
  (
    n2545,
    n1932,
    n2493,
    n2494,
    n1906
  );


  not
  g2524
  (
    n2560,
    n2544
  );


  not
  g2525
  (
    n2557,
    n2541
  );


  buf
  g2526
  (
    n2559,
    n2542
  );


  buf
  g2527
  (
    n2558,
    n2543
  );


  nand
  g2528
  (
    n2561,
    n2498,
    n2499,
    n2559
  );


  not
  g2529
  (
    n2563,
    n2561
  );


  buf
  g2530
  (
    n2562,
    n2561
  );


  not
  g2531
  (
    n2568,
    n2548
  );


  not
  g2532
  (
    n2565,
    n2562
  );


  buf
  g2533
  (
    n2564,
    n2563
  );


  not
  g2534
  (
    n2567,
    n2547
  );


  nand
  g2535
  (
    n2566,
    n2546,
    n2549,
    n2563,
    n2562
  );


  xnor
  g2536
  (
    n2569,
    n2545,
    n2550,
    n2562
  );


  not
  g2537
  (
    n2581,
    n2567
  );


  buf
  g2538
  (
    n2577,
    n1956
  );


  buf
  g2539
  (
    KeyWire_0_22,
    n2500
  );


  not
  g2540
  (
    n2579,
    n2560
  );


  and
  g2541
  (
    n2575,
    n1951,
    n2566,
    n1946,
    n2501
  );


  nor
  g2542
  (
    n2570,
    n2502,
    n2500,
    n2499,
    n2565
  );


  nor
  g2543
  (
    n2572,
    n2502,
    n1953,
    n1957,
    n2500
  );


  or
  g2544
  (
    n2580,
    n2565,
    n2502,
    n2568,
    n2501
  );


  xnor
  g2545
  (
    n2583,
    n2567,
    n2565,
    n2503,
    n1948
  );


  nor
  g2546
  (
    n2576,
    n1949,
    n2566,
    n2501
  );


  xor
  g2547
  (
    n2574,
    n1950,
    n1945,
    n1954,
    n2501
  );


  xor
  g2548
  (
    n2571,
    n2564,
    n2499,
    n2502,
    n2567
  );


  xor
  g2549
  (
    n2584,
    n1952,
    n1947,
    n2503,
    n2565
  );


  nand
  g2550
  (
    n2582,
    n1942,
    n2566,
    n2500,
    n1944
  );


  xor
  g2551
  (
    n2573,
    n1943,
    n2567,
    n1955,
    n2564
  );


  buf
  g2552
  (
    n2597,
    n2576
  );


  not
  g2553
  (
    n2603,
    n2576
  );


  not
  g2554
  (
    n2596,
    n1974
  );


  buf
  g2555
  (
    n2600,
    n2577
  );


  buf
  g2556
  (
    n2585,
    n2574
  );


  not
  g2557
  (
    n2605,
    n2570
  );


  or
  g2558
  (
    n2586,
    n1964,
    n2572
  );


  nor
  g2559
  (
    n2589,
    n1969,
    n1975,
    n2579,
    n2574
  );


  and
  g2560
  (
    n2595,
    n2571,
    n2573,
    n2575,
    n1958
  );


  and
  g2561
  (
    n2599,
    n2573,
    n2575,
    n1961,
    n2576
  );


  and
  g2562
  (
    n2591,
    n2570,
    n2577,
    n2576,
    n1972
  );


  and
  g2563
  (
    n2587,
    n1970,
    n1977,
    n2578,
    n2572
  );


  xnor
  g2564
  (
    n2594,
    n2503,
    n2575,
    n2577,
    n1976
  );


  or
  g2565
  (
    n2588,
    n2578,
    n2573,
    n1967,
    n1960
  );


  xor
  g2566
  (
    n2604,
    n2578,
    n2571,
    n2572,
    n2570
  );


  nor
  g2567
  (
    n2593,
    n1973,
    n1959,
    n1965,
    n1962
  );


  or
  g2568
  (
    n2601,
    n1980,
    n2572,
    n1979,
    n2504
  );


  or
  g2569
  (
    n2602,
    n1963,
    n1968,
    n1966,
    n2575
  );


  xnor
  g2570
  (
    n2598,
    n1971,
    n2573,
    n2578,
    n2574
  );


  or
  g2571
  (
    n2590,
    n1981,
    n2571,
    n2577
  );


  and
  g2572
  (
    n2592,
    n2574,
    n2570,
    n1978,
    n2503
  );


  xor
  g2573
  (
    n2610,
    n2586,
    n2596,
    n2593,
    n2569
  );


  and
  g2574
  (
    n2609,
    n2563,
    n2596,
    n2585,
    n2588
  );


  or
  g2575
  (
    n2617,
    n2589,
    n2568,
    n2597,
    n2585
  );


  nand
  g2576
  (
    n2619,
    n2590,
    n1987,
    n2588,
    n2595
  );


  nand
  g2577
  (
    n2607,
    n2588,
    n2589,
    n2591,
    n1982
  );


  xnor
  g2578
  (
    n2620,
    n2586,
    n2597,
    n2585,
    n2569
  );


  nor
  g2579
  (
    n2623,
    n2586,
    n2587,
    n2597,
    n2595
  );


  nor
  g2580
  (
    n2621,
    n2597,
    n2592,
    n2591
  );


  nor
  g2581
  (
    n2611,
    n2595,
    n2594,
    n2587
  );


  xnor
  g2582
  (
    n2613,
    n2568,
    n2589,
    n2596,
    n1985
  );


  xor
  g2583
  (
    n2612,
    n1988,
    n1984,
    n2563,
    n2595
  );


  xor
  g2584
  (
    n2615,
    n2598,
    n1983,
    n2585,
    n2588
  );


  and
  g2585
  (
    n2618,
    n2590,
    n2591,
    n2594,
    n2589
  );


  and
  g2586
  (
    n2616,
    n2592,
    n2587,
    n2591
  );


  xor
  g2587
  (
    n2614,
    n2599,
    n2592,
    n1986,
    n2598
  );


  nand
  g2588
  (
    n2622,
    n2598,
    n1989,
    n2593
  );


  nand
  g2589
  (
    n2608,
    n2593,
    n2596,
    n2590,
    n2586
  );


  nor
  g2590
  (
    n2606,
    n2598,
    n2590,
    n2568,
    n2594
  );


  xor
  g2591
  (
    n2624,
    n2579,
    n2569,
    n2622
  );


  not
  g2592
  (
    n2626,
    n2624
  );


  buf
  g2593
  (
    n2625,
    n2624
  );


  nand
  g2594
  (
    n2630,
    n2625,
    n2604,
    n2599,
    n2601
  );


  nand
  g2595
  (
    n2628,
    n2602,
    n2604,
    n2599,
    n2625
  );


  and
  g2596
  (
    n2634,
    n2602,
    n2602,
    n2600,
    n2625
  );


  xnor
  g2597
  (
    n2627,
    n2626,
    n2626,
    n2601,
    n2600
  );


  xnor
  g2598
  (
    n2633,
    n2602,
    n2604,
    n2600,
    n2603
  );


  xor
  g2599
  (
    n2629,
    n2601,
    n2603,
    n2605,
    n2626
  );


  and
  g2600
  (
    n2631,
    n2604,
    n2600,
    n2599,
    n2626
  );


  xnor
  g2601
  (
    n2632,
    n2625,
    n2603,
    n2601
  );


  xnor
  g2602
  (
    n2653,
    n1814,
    n1818,
    n2627,
    n2551
  );


  xnor
  g2603
  (
    n2660,
    n2630,
    n2580,
    n2581,
    n2628
  );


  nor
  g2604
  (
    n2642,
    n1817,
    n1813,
    n2529,
    n2528
  );


  nor
  g2605
  (
    n2646,
    n1811,
    n1814,
    n2631
  );


  or
  g2606
  (
    n2647,
    n1815,
    n1820,
    n2628,
    n2627
  );


  nor
  g2607
  (
    n2662,
    n2580,
    n1822,
    n1821,
    n2527
  );


  and
  g2608
  (
    n2649,
    n2527,
    n2632,
    n1991,
    n2630
  );


  xor
  g2609
  (
    n2657,
    n1811,
    n1990,
    n1814,
    n2630
  );


  nor
  g2610
  (
    n2645,
    n1820,
    n1816,
    n1824,
    n2633
  );


  xnor
  g2611
  (
    KeyWire_0_23,
    n1811,
    n1813,
    n2633,
    n2580
  );


  nand
  g2612
  (
    n2639,
    n2623,
    n1818,
    n1811
  );


  nand
  g2613
  (
    n2658,
    n1817,
    n2627,
    n2581,
    n1821
  );


  nor
  g2614
  (
    n2644,
    n2631,
    n1812,
    n2629,
    n2633
  );


  nor
  g2615
  (
    n2640,
    n2632,
    n1822,
    n2631,
    n2582
  );


  xor
  g2616
  (
    n2661,
    n1822,
    n2632,
    n2579,
    n1813
  );


  nand
  g2617
  (
    n2654,
    n1812,
    n1817,
    n1819,
    n2582
  );


  xnor
  g2618
  (
    n2648,
    n2633,
    n1820,
    n2628,
    n2581
  );


  xor
  g2619
  (
    n2652,
    n1810,
    n1823,
    n1819,
    n2529
  );


  or
  g2620
  (
    n2656,
    n1817,
    n1812,
    n1992,
    n1822
  );


  xor
  g2621
  (
    n2651,
    n1818,
    n1823,
    n2629,
    n2528
  );


  xor
  g2622
  (
    n2655,
    n1810,
    n1815,
    n2630,
    n2581
  );


  and
  g2623
  (
    n2635,
    n1819,
    n2579,
    n1816,
    n2528
  );


  xor
  g2624
  (
    n2650,
    n1994,
    n2627,
    n1820,
    n1821
  );


  xnor
  g2625
  (
    n2643,
    n2632,
    n2631,
    n2628,
    n2580
  );


  xnor
  g2626
  (
    n2638,
    n1813,
    n1815,
    n2629,
    n2582
  );


  and
  g2627
  (
    n2637,
    n1819,
    n1815,
    n1823,
    n1812
  );


  xnor
  g2628
  (
    n2659,
    n1823,
    n1816,
    n2527,
    n2629
  );


  and
  g2629
  (
    n2641,
    n2528,
    n1993,
    n1816,
    n1821
  );


  buf
  g2630
  (
    n2667,
    n2647
  );


  not
  g2631
  (
    n2675,
    n2635
  );


  buf
  g2632
  (
    n2663,
    n2646
  );


  buf
  g2633
  (
    n2670,
    n2639
  );


  buf
  g2634
  (
    n2676,
    n2637
  );


  not
  g2635
  (
    n2666,
    n2648
  );


  buf
  g2636
  (
    n2669,
    n2638
  );


  not
  g2637
  (
    n2668,
    n2645
  );


  not
  g2638
  (
    n2671,
    n2636
  );


  buf
  g2639
  (
    n2673,
    n2644
  );


  not
  g2640
  (
    n2672,
    n2642
  );


  not
  g2641
  (
    n2664,
    n2640
  );


  buf
  g2642
  (
    n2674,
    n2649
  );


  buf
  g2643
  (
    n2665,
    n2650
  );


  not
  g2644
  (
    n2677,
    n2643
  );


  buf
  g2645
  (
    n2678,
    n2641
  );


  and
  g2646
  (
    n2716,
    n2057,
    n2119,
    n2126,
    n2105
  );


  xnor
  g2647
  (
    n2708,
    n2663,
    n2068,
    n2055,
    n2018
  );


  xor
  g2648
  (
    n2687,
    n2087,
    n2665,
    n2070,
    n2663
  );


  or
  g2649
  (
    n2741,
    n2674,
    n2080,
    n2025,
    n2090
  );


  xnor
  g2650
  (
    n2737,
    n2677,
    n2083,
    n2031,
    n2058
  );


  xnor
  g2651
  (
    n2718,
    n2078,
    n2029,
    n2041,
    n2045
  );


  nand
  g2652
  (
    n2728,
    n1999,
    n2081,
    n2169,
    n2143
  );


  or
  g2653
  (
    n2726,
    n2148,
    n2634,
    n2157,
    n2674
  );


  xnor
  g2654
  (
    n2736,
    n2054,
    n2583,
    n2002,
    n2124
  );


  xnor
  g2655
  (
    n2730,
    n2065,
    n2672,
    n2127,
    n2106
  );


  nor
  g2656
  (
    n2714,
    n2060,
    n2069,
    n2678,
    n2010
  );


  xnor
  g2657
  (
    n2725,
    n2677,
    n2004,
    n2671
  );


  nand
  g2658
  (
    n2696,
    n2050,
    n2164,
    n2666,
    n2678
  );


  and
  g2659
  (
    n2734,
    n2032,
    n2158,
    n2005,
    n2059
  );


  xnor
  g2660
  (
    n2704,
    n2033,
    n2048,
    n2027,
    n2049
  );


  nand
  g2661
  (
    n2729,
    n2673,
    n2062,
    n2091,
    n2123
  );


  nand
  g2662
  (
    n2706,
    n2583,
    n664,
    n2584,
    n2103
  );


  xnor
  g2663
  (
    n2693,
    n2085,
    n2678,
    n2100,
    n2017
  );


  and
  g2664
  (
    n2692,
    n2096,
    n2012,
    n2675,
    n2672
  );


  nand
  g2665
  (
    n2723,
    n2161,
    n2584,
    n2634
  );


  nor
  g2666
  (
    n2705,
    n2044,
    n2102,
    n2142,
    n2109
  );


  or
  g2667
  (
    n2699,
    n2099,
    n2668,
    n2167,
    n2035
  );


  nand
  g2668
  (
    n2703,
    n2111,
    n2015,
    n2667,
    n2108
  );


  nor
  g2669
  (
    n2721,
    n2088,
    n2037,
    n2677,
    n2665
  );


  nor
  g2670
  (
    n2688,
    n2152,
    n2014,
    n2131,
    n2016
  );


  nor
  g2671
  (
    n2707,
    n2669,
    n2137,
    n2663,
    n2104
  );


  xnor
  g2672
  (
    n2731,
    n2664,
    n2665,
    n2671,
    n1824
  );


  or
  g2673
  (
    n2682,
    n2135,
    n2125,
    n2583,
    n2022
  );


  xnor
  g2674
  (
    n2724,
    n2666,
    n2153,
    n2084,
    n2667
  );


  xnor
  g2675
  (
    n2711,
    n2669,
    n2006,
    n2110,
    n2066
  );


  nand
  g2676
  (
    n2733,
    n2668,
    n2676,
    n2114
  );


  nor
  g2677
  (
    n2717,
    n2668,
    n2141,
    n2072,
    n2075
  );


  xor
  g2678
  (
    n2735,
    n2147,
    n2133,
    n2001,
    n2675
  );


  or
  g2679
  (
    n2694,
    n2112,
    n1824,
    n2675,
    n2140
  );


  or
  g2680
  (
    n2713,
    n2047,
    n2146,
    n2000,
    n2042
  );


  xor
  g2681
  (
    n2702,
    n2145,
    n2056,
    n2113,
    n2028
  );


  xor
  g2682
  (
    n2691,
    n2166,
    n2023,
    n2013,
    n2673
  );


  xor
  g2683
  (
    n2720,
    n2584,
    n2019,
    n2139,
    n2674
  );


  xnor
  g2684
  (
    n2740,
    n2163,
    n1824,
    n2073,
    n2064
  );


  xor
  g2685
  (
    n2697,
    n2101,
    n2021,
    n2071,
    n2007
  );


  nand
  g2686
  (
    n2712,
    n2036,
    n2030,
    n2009,
    n2043
  );


  or
  g2687
  (
    n2732,
    n2122,
    n2678,
    n2038,
    n2092
  );


  nand
  g2688
  (
    n2686,
    n2118,
    n2107,
    n2677,
    n2076
  );


  and
  g2689
  (
    n2698,
    n2159,
    n2074,
    n2168,
    n2670
  );


  nor
  g2690
  (
    n2683,
    n2117,
    n2144,
    n2095,
    n2671
  );


  nor
  g2691
  (
    n2701,
    n2666,
    n1995,
    n2155,
    n2053
  );


  or
  g2692
  (
    n2700,
    n2052,
    n2024,
    n2034,
    n2151
  );


  xnor
  g2693
  (
    n2685,
    n2067,
    n2670,
    n2136,
    n2154
  );


  xnor
  g2694
  (
    n2738,
    n2089,
    n2667,
    n2008,
    n2046
  );


  xnor
  g2695
  (
    n2727,
    n2079,
    n2675,
    n2063,
    n2132
  );


  or
  g2696
  (
    n2689,
    n2664,
    n2082,
    n2672,
    n2663
  );


  or
  g2697
  (
    KeyWire_0_6,
    n2668,
    n2003,
    n2020,
    n2674
  );


  nand
  g2698
  (
    n2715,
    n2040,
    n2666,
    n2665,
    n2634
  );


  nand
  g2699
  (
    n2709,
    n2128,
    n2094,
    n2026,
    n2150
  );


  nand
  g2700
  (
    n2690,
    n2673,
    n2664,
    n2115,
    n2130
  );


  xnor
  g2701
  (
    n2742,
    n2670,
    n2120,
    n2097,
    n2160
  );


  nand
  g2702
  (
    n2681,
    n2667,
    n2156,
    n2672,
    n2086
  );


  and
  g2703
  (
    n2695,
    n2138,
    n2077,
    n2061,
    n2093
  );


  nor
  g2704
  (
    n2679,
    n2582,
    n2149,
    n2116,
    n2129
  );


  or
  g2705
  (
    n2719,
    n2162,
    n1996,
    n2584,
    n2134
  );


  or
  g2706
  (
    n2680,
    n2039,
    n2051,
    n1998,
    n2165
  );


  nor
  g2707
  (
    n2722,
    n2098,
    n2121,
    n2673,
    n2669
  );


  and
  g2708
  (
    n2739,
    n2669,
    n2664,
    n2583,
    n2670
  );


  nand
  g2709
  (
    n2684,
    n1997,
    n2676,
    n2011
  );


  not
  g2710
  (
    n2748,
    n2679
  );


  not
  g2711
  (
    n2743,
    n2679
  );


  not
  g2712
  (
    n2749,
    n2679
  );


  buf
  g2713
  (
    n2745,
    n2679
  );


  buf
  g2714
  (
    n2746,
    n2651
  );


  buf
  g2715
  (
    n2747,
    n2680
  );


  not
  g2716
  (
    n2744,
    n2680
  );


  buf
  g2717
  (
    n2766,
    n2662
  );


  not
  g2718
  (
    n2763,
    n2747
  );


  not
  g2719
  (
    n2757,
    n2660
  );


  buf
  g2720
  (
    n2759,
    n2748
  );


  not
  g2721
  (
    n2756,
    n2747
  );


  buf
  g2722
  (
    n2754,
    n2746
  );


  not
  g2723
  (
    n2767,
    n2749
  );


  buf
  g2724
  (
    n2771,
    n2657
  );


  buf
  g2725
  (
    n2764,
    n2748
  );


  buf
  g2726
  (
    n2758,
    n2652
  );


  not
  g2727
  (
    n2768,
    n2749
  );


  buf
  g2728
  (
    n2752,
    n2745
  );


  buf
  g2729
  (
    n2762,
    n2653
  );


  buf
  g2730
  (
    n2770,
    n2654
  );


  buf
  g2731
  (
    n2773,
    n2744
  );


  buf
  g2732
  (
    n2751,
    n2749
  );


  not
  g2733
  (
    n2765,
    n2658
  );


  not
  g2734
  (
    n2772,
    n2746
  );


  buf
  g2735
  (
    n2761,
    n2744
  );


  xnor
  g2736
  (
    n2755,
    n2743,
    n2747
  );


  nand
  g2737
  (
    n2774,
    n2746,
    n2745,
    n2744
  );


  or
  g2738
  (
    n2753,
    n2659,
    n2745,
    n2743
  );


  and
  g2739
  (
    n2760,
    n2744,
    n2748,
    n2655
  );


  xnor
  g2740
  (
    n2750,
    n2748,
    n2746,
    n2661
  );


  or
  g2741
  (
    n2769,
    n2656,
    n2745,
    n2747
  );


  xnor
  g2742
  (
    n2791,
    n2686,
    n2172,
    n2700,
    n2702
  );


  and
  g2743
  (
    n2794,
    n2724,
    n2605,
    n2708,
    n2686
  );


  xnor
  g2744
  (
    n2801,
    n667,
    n2771,
    n2184,
    n2508
  );


  nor
  g2745
  (
    n2809,
    n2726,
    n2683,
    n2513,
    n2766
  );


  and
  g2746
  (
    n2821,
    n2681,
    n2759,
    n2514,
    n2707
  );


  and
  g2747
  (
    n2793,
    n2605,
    n2754,
    n2762,
    n2685
  );


  xnor
  g2748
  (
    n2781,
    n2505,
    n2509,
    n2605,
    n2702
  );


  xnor
  g2749
  (
    n2824,
    n2510,
    n2508,
    n2709,
    n2722
  );


  and
  g2750
  (
    n2787,
    n2702,
    n2707,
    n2752,
    n2717
  );


  xnor
  g2751
  (
    n2831,
    n2754,
    n2681,
    n2759,
    n2509
  );


  nor
  g2752
  (
    n2792,
    n2710,
    n2693,
    n2768,
    n2752
  );


  nand
  g2753
  (
    n2857,
    n2703,
    n2689,
    n2767,
    n2706
  );


  xnor
  g2754
  (
    n2808,
    n2754,
    n2768,
    n2710,
    n2767
  );


  xor
  g2755
  (
    n2790,
    n2750,
    n2700,
    n2755,
    n2180
  );


  xor
  g2756
  (
    n2818,
    n2719,
    n2698,
    n2699,
    n2769
  );


  xor
  g2757
  (
    n2788,
    n2683,
    n2706,
    n2766,
    n2717
  );


  and
  g2758
  (
    n2805,
    n2505,
    n2688,
    n2763,
    n2709
  );


  nand
  g2759
  (
    n2807,
    n2757,
    n2700,
    n2505,
    n2693
  );


  xnor
  g2760
  (
    n2833,
    n2716,
    n2514,
    n2723,
    n2508
  );


  nand
  g2761
  (
    n2817,
    n2716,
    n2724,
    n2699
  );


  nand
  g2762
  (
    n2853,
    n2725,
    n2718,
    n2507,
    n2719
  );


  nand
  g2763
  (
    n2826,
    n2684,
    n2688,
    n2753,
    n2687
  );


  nand
  g2764
  (
    n2778,
    n2509,
    n2181,
    n2769,
    n2755
  );


  or
  g2765
  (
    n2782,
    n2694,
    n2708,
    n664,
    n2760
  );


  nor
  g2766
  (
    n2827,
    n2753,
    n2688,
    n2715,
    n2705
  );


  xnor
  g2767
  (
    n2800,
    n2690,
    n2506,
    n2703,
    n2718
  );


  nor
  g2768
  (
    n2823,
    n2721,
    n2687,
    n2724,
    n2726
  );


  and
  g2769
  (
    n2798,
    n2751,
    n2752,
    n2696
  );


  xor
  g2770
  (
    n2775,
    n2723,
    n2763,
    n2712,
    n2770
  );


  nand
  g2771
  (
    n2848,
    n2689,
    n2715,
    n2760,
    n2505
  );


  or
  g2772
  (
    n2806,
    n2700,
    n2750,
    n2706,
    n2704
  );


  and
  g2773
  (
    n2779,
    n2718,
    n2697,
    n2720,
    n2724
  );


  nor
  g2774
  (
    n2802,
    n2715,
    n2769,
    n2514,
    n2711
  );


  xor
  g2775
  (
    n2804,
    n2712,
    n2705,
    n2685,
    n2703
  );


  xor
  g2776
  (
    n2840,
    n2506,
    n665,
    n2182,
    n2764
  );


  xor
  g2777
  (
    n2780,
    n2177,
    n2684,
    n2179,
    n2771
  );


  xor
  g2778
  (
    n2835,
    n2721,
    n2770,
    n2703,
    n2716
  );


  xnor
  g2779
  (
    n2829,
    n2715,
    n2695,
    n2693,
    n2758
  );


  or
  g2780
  (
    n2799,
    n2758,
    n2758,
    n2510,
    n2512
  );


  and
  g2781
  (
    n2836,
    n2690,
    n665,
    n2751,
    n2769
  );


  or
  g2782
  (
    n2820,
    n2510,
    n2693,
    n2756,
    n2174
  );


  nand
  g2783
  (
    n2841,
    n2725,
    n2722,
    n2756,
    n2507
  );


  xnor
  g2784
  (
    n2834,
    n665,
    n2513,
    n2504,
    n2508
  );


  or
  g2785
  (
    n2810,
    n2725,
    n2704,
    n2720,
    n2751
  );


  or
  g2786
  (
    n2851,
    n2762,
    n2767,
    n664,
    n2687
  );


  nand
  g2787
  (
    n2849,
    n2704,
    n2695,
    n2689,
    n2764
  );


  nand
  g2788
  (
    n2776,
    n2510,
    n2757,
    n2504,
    n2722
  );


  and
  g2789
  (
    n2785,
    n2764,
    n2714,
    n667
  );


  nand
  g2790
  (
    n2822,
    n2771,
    n665,
    n2756,
    n2717
  );


  xor
  g2791
  (
    n2842,
    n2767,
    n2701,
    n2712,
    n2692
  );


  xnor
  g2792
  (
    n2797,
    n2763,
    n2513,
    n2685,
    n2183
  );


  xnor
  g2793
  (
    n2845,
    n2681,
    n2717,
    n2713,
    n2685
  );


  nand
  g2794
  (
    n2847,
    n2688,
    n2682,
    n2718,
    n2711
  );


  nor
  g2795
  (
    n2814,
    n2761,
    n2723,
    n2755,
    n2708
  );


  nand
  g2796
  (
    n2828,
    n2697,
    n2694,
    n2511,
    n2765
  );


  nand
  g2797
  (
    n2844,
    n2704,
    n2170,
    n2707,
    n2691
  );


  xnor
  g2798
  (
    n2856,
    n2762,
    n2720,
    n2698,
    n2770
  );


  nand
  g2799
  (
    n2838,
    n2761,
    n2766,
    n2506,
    n2719
  );


  xnor
  g2800
  (
    n2786,
    n2175,
    n2760,
    n2708,
    n2701
  );


  and
  g2801
  (
    n2812,
    n2682,
    n2762,
    n666,
    n2723
  );


  or
  g2802
  (
    n2861,
    n2680,
    n2765,
    n2711,
    n2713
  );


  nor
  g2803
  (
    n2855,
    n2694,
    n2684,
    n2512,
    n2705
  );


  xnor
  g2804
  (
    n2813,
    n2768,
    n666,
    n2694,
    n2712
  );


  nand
  g2805
  (
    n2830,
    n2758,
    n2696,
    n2751,
    n2765
  );


  xor
  g2806
  (
    n2837,
    n2507,
    n2759,
    n2770,
    n2504
  );


  nand
  g2807
  (
    n2784,
    n2721,
    n2721,
    n2171,
    n2702
  );


  and
  g2808
  (
    n2815,
    n2710,
    n2754,
    n2691,
    n2726
  );


  xnor
  g2809
  (
    n2819,
    n2701,
    n2692,
    n2690,
    n2507
  );


  or
  g2810
  (
    n2795,
    n2750,
    n2511,
    n2753,
    n2760
  );


  nor
  g2811
  (
    n2854,
    n2698,
    n2761,
    n2719,
    n2681
  );


  nand
  g2812
  (
    n2783,
    n2756,
    n2511,
    n2695,
    n2710
  );


  nor
  g2813
  (
    n2796,
    n666,
    n2755,
    n2757
  );


  and
  g2814
  (
    n2852,
    n2697,
    n2683,
    n2178,
    n2513
  );


  nand
  g2815
  (
    n2803,
    n2682,
    n2691,
    n2720,
    n664
  );


  and
  g2816
  (
    n2816,
    n2768,
    n2701,
    n2750,
    n2711
  );


  xnor
  g2817
  (
    n2811,
    n2692,
    n2713,
    n2722,
    n2714
  );


  xnor
  g2818
  (
    n2825,
    n2686,
    n2705,
    n2697,
    n2706
  );


  nor
  g2819
  (
    n2839,
    n2691,
    n2173,
    n2512,
    n667
  );


  nand
  g2820
  (
    n2843,
    n2766,
    n2506,
    n2707,
    n2696
  );


  or
  g2821
  (
    n2859,
    n2761,
    n2725,
    n2753,
    n2687
  );


  xor
  g2822
  (
    n2777,
    n2684,
    n2763,
    n2695,
    n666
  );


  xnor
  g2823
  (
    n2789,
    n2690,
    n2699,
    n2696,
    n2682
  );


  xnor
  g2824
  (
    n2860,
    n2759,
    n2686,
    n2765,
    n2511
  );


  xnor
  g2825
  (
    n2832,
    n2726,
    n2512,
    n2709,
    n2713
  );


  nand
  g2826
  (
    n2846,
    n667,
    n2716,
    n2689,
    n2714
  );


  or
  g2827
  (
    n2858,
    n2692,
    n2683,
    n2185,
    n2709
  );


  and
  g2828
  (
    n2850,
    n2509,
    n2176,
    n2764,
    n2698
  );


  xnor
  g2829
  (
    n2981,
    n2415,
    n2314,
    n2377,
    n2352
  );


  or
  g2830
  (
    n2919,
    n2281,
    n2199,
    n2727,
    n2315
  );


  xor
  g2831
  (
    n2901,
    n2731,
    n2269,
    n2240,
    n2820
  );


  and
  g2832
  (
    n2876,
    n2740,
    n2356,
    n2851,
    n2854
  );


  xor
  g2833
  (
    n2956,
    n2749,
    n2425,
    n2738,
    n2730
  );


  nand
  g2834
  (
    n2893,
    n2358,
    n2212,
    n2220,
    n2208
  );


  and
  g2835
  (
    n2978,
    n2854,
    n2287,
    n2432,
    n2794
  );


  or
  g2836
  (
    n2977,
    n2471,
    n2254,
    n2381,
    n2291
  );


  xor
  g2837
  (
    n2914,
    n2738,
    n2393,
    n2411,
    n2379
  );


  xnor
  g2838
  (
    n2864,
    n2735,
    n2469,
    n2781,
    n2853
  );


  xor
  g2839
  (
    n2920,
    n2248,
    n2295,
    n2313,
    n2272
  );


  nand
  g2840
  (
    n2980,
    n2349,
    n2317,
    n2270,
    n2309
  );


  or
  g2841
  (
    n2868,
    n2786,
    n2728,
    n2427,
    n2221
  );


  nand
  g2842
  (
    n2930,
    n2299,
    n2331,
    n2334,
    n2328
  );


  nand
  g2843
  (
    n2950,
    n2830,
    n2729,
    n2262,
    n2337
  );


  or
  g2844
  (
    n2913,
    n2260,
    n2235,
    n2266,
    n2231
  );


  and
  g2845
  (
    n2886,
    n2843,
    n2369,
    n2232,
    n2443
  );


  nand
  g2846
  (
    n2866,
    n2456,
    n2440,
    n2330,
    n2852
  );


  and
  g2847
  (
    n2921,
    n2249,
    n2819,
    n2288,
    n2277
  );


  xnor
  g2848
  (
    n2947,
    n2853,
    n2422,
    n2735,
    n2851
  );


  nor
  g2849
  (
    n2887,
    n2441,
    n2187,
    n2308,
    n2448
  );


  and
  g2850
  (
    n2908,
    n2802,
    n2437,
    n2859,
    n2242
  );


  nor
  g2851
  (
    n2955,
    n2733,
    n2841,
    n2858,
    n2857
  );


  and
  g2852
  (
    n2940,
    n2829,
    n2850,
    n2477,
    n2849
  );


  or
  g2853
  (
    n2949,
    n2466,
    n2326,
    n2256,
    n2442
  );


  and
  g2854
  (
    n2906,
    n2435,
    n2278,
    n2738,
    n2333
  );


  nand
  g2855
  (
    n2935,
    n2261,
    n2856,
    n2206,
    n2804
  );


  or
  g2856
  (
    n2965,
    n2833,
    n2209,
    n2856,
    n2407
  );


  or
  g2857
  (
    n2896,
    n2810,
    n2338,
    n2204,
    n2391
  );


  and
  g2858
  (
    n2865,
    n2858,
    n2189,
    n2428,
    n2790
  );


  and
  g2859
  (
    n2888,
    n2324,
    n2737,
    n2801,
    n2729
  );


  nand
  g2860
  (
    n2900,
    n2263,
    n2376,
    n2461,
    n2462
  );


  and
  g2861
  (
    n2934,
    n2814,
    n2731,
    n2848,
    n2364
  );


  and
  g2862
  (
    n2915,
    n2296,
    n2234,
    n2734,
    n2342
  );


  or
  g2863
  (
    n2863,
    n2465,
    n2282,
    n2779,
    n2284
  );


  and
  g2864
  (
    n2960,
    n2417,
    n2470,
    n2405,
    n2347
  );


  xor
  g2865
  (
    n2862,
    n2449,
    n2826,
    n2741,
    n2736
  );


  nand
  g2866
  (
    n2945,
    n2401,
    n2264,
    n2849,
    n2822
  );


  and
  g2867
  (
    n2976,
    n2395,
    n2729,
    n2838,
    n2283
  );


  and
  g2868
  (
    n2875,
    n2396,
    n2265,
    n2302,
    n2807
  );


  or
  g2869
  (
    n2937,
    n2412,
    n2789,
    n2813,
    n2803
  );


  and
  g2870
  (
    n2905,
    n2384,
    n2323,
    n2365,
    n2733
  );


  xnor
  g2871
  (
    n2969,
    n2738,
    n2193,
    n2783,
    n2854
  );


  and
  g2872
  (
    n2926,
    n2355,
    n2318,
    n2293,
    n2222
  );


  or
  g2873
  (
    n2884,
    n2479,
    n2236,
    n2360,
    n2202
  );


  or
  g2874
  (
    n2871,
    n2233,
    n2230,
    n2780,
    n2275
  );


  or
  g2875
  (
    n2892,
    n2742,
    n2736,
    n2325,
    n2851
  );


  or
  g2876
  (
    n2967,
    n2430,
    n2737,
    n2856,
    n2341
  );


  nor
  g2877
  (
    n2954,
    n2292,
    n2740,
    n2808,
    n2335
  );


  and
  g2878
  (
    n2944,
    n2386,
    n2239,
    n2809,
    n2312
  );


  or
  g2879
  (
    n2973,
    n2310,
    n2739,
    n2778,
    n2827
  );


  xor
  g2880
  (
    n2979,
    n2831,
    n2359,
    n2797,
    n2823
  );


  nand
  g2881
  (
    n2961,
    n2274,
    n2363,
    n2244,
    n2343
  );


  or
  g2882
  (
    n2889,
    n2793,
    n2458,
    n2345,
    n2367
  );


  nor
  g2883
  (
    n2879,
    n2387,
    n2824,
    n2815,
    n2374
  );


  xnor
  g2884
  (
    n2877,
    n2444,
    n2431,
    n2848,
    n2728
  );


  or
  g2885
  (
    n2938,
    n2398,
    n2205,
    n2203,
    n2734
  );


  nand
  g2886
  (
    n2898,
    n2858,
    n2389,
    n2737,
    n2404
  );


  xnor
  g2887
  (
    n2941,
    n2857,
    n2741,
    n2852,
    n2201
  );


  xnor
  g2888
  (
    n2931,
    n2414,
    n2445,
    n2192,
    n2439
  );


  and
  g2889
  (
    n2948,
    n2467,
    n2733,
    n2280,
    n2854
  );


  or
  g2890
  (
    n2970,
    n2736,
    n2217,
    n2734,
    n2237
  );


  or
  g2891
  (
    n2873,
    n2421,
    n2852,
    n2730,
    n2514
  );


  nor
  g2892
  (
    n2972,
    n2846,
    n2354,
    n2303,
    n2357
  );


  xor
  g2893
  (
    n2953,
    n2373,
    n2832,
    n2739,
    n2853
  );


  nor
  g2894
  (
    n2881,
    n2859,
    n2856,
    n2416,
    n2455
  );


  xor
  g2895
  (
    n2904,
    n2216,
    n2735,
    n2474,
    n2850
  );


  nor
  g2896
  (
    n2918,
    n2798,
    n2845,
    n2740,
    n2394
  );


  nand
  g2897
  (
    n2927,
    n2268,
    n2353,
    n2464,
    n2327
  );


  and
  g2898
  (
    n2878,
    n2321,
    n2271,
    n2434,
    n2402
  );


  or
  g2899
  (
    n2963,
    n2850,
    n2227,
    n2805,
    n2849
  );


  or
  g2900
  (
    n2885,
    n2791,
    n2195,
    n2436,
    n2450
  );


  or
  g2901
  (
    n2971,
    n2733,
    n2226,
    n2800,
    n2224
  );


  xor
  g2902
  (
    n2907,
    n2255,
    n2795,
    n2285,
    n2371
  );


  xor
  g2903
  (
    n2966,
    n2346,
    n2213,
    n2191,
    n2198
  );


  nor
  g2904
  (
    n2968,
    n2273,
    n2319,
    n2378,
    n2776
  );


  or
  g2905
  (
    n2943,
    n2727,
    n2727,
    n2223,
    n2329
  );


  or
  g2906
  (
    n2917,
    n2380,
    n2848,
    n2739,
    n2459
  );


  and
  g2907
  (
    n2894,
    n2258,
    n2775,
    n2858,
    n2806
  );


  and
  g2908
  (
    n2909,
    n2457,
    n2835,
    n2452,
    n2397
  );


  nor
  g2909
  (
    n2942,
    n2253,
    n2828,
    n2408,
    n2294
  );


  xor
  g2910
  (
    n2964,
    n2251,
    n2451,
    n2855,
    n2247
  );


  xnor
  g2911
  (
    n2911,
    n2735,
    n2316,
    n2732,
    n2304
  );


  and
  g2912
  (
    n2924,
    n2736,
    n2855,
    n2739,
    n2848
  );


  nand
  g2913
  (
    n2880,
    n2850,
    n2741,
    n2228,
    n2837
  );


  and
  g2914
  (
    n2974,
    n2370,
    n2433,
    n2737,
    n2390
  );


  nand
  g2915
  (
    n2923,
    n2410,
    n2742,
    n2463,
    n2368
  );


  and
  g2916
  (
    n2925,
    n2259,
    n2816,
    n2336,
    n2728
  );


  xor
  g2917
  (
    n2929,
    n2446,
    n2241,
    n2842,
    n2290
  );


  or
  g2918
  (
    n2958,
    n2787,
    n2186,
    n2413,
    n2732
  );


  nor
  g2919
  (
    n2869,
    n2811,
    n2250,
    n2361,
    n2473
  );


  xor
  g2920
  (
    n2922,
    n2246,
    n2857,
    n2332,
    n2796
  );


  xnor
  g2921
  (
    n2951,
    n2306,
    n2799,
    n2305,
    n2219
  );


  nand
  g2922
  (
    n2902,
    n2307,
    n2478,
    n2200,
    n2286
  );


  nor
  g2923
  (
    n2867,
    n2383,
    n2818,
    n2817,
    n2252
  );


  or
  g2924
  (
    n2959,
    n2840,
    n2300,
    n2438,
    n2418
  );


  xor
  g2925
  (
    n2962,
    n2243,
    n2426,
    n2399,
    n2839
  );


  or
  g2926
  (
    n2932,
    n2188,
    n2214,
    n2403,
    n2853
  );


  xor
  g2927
  (
    n2936,
    n2740,
    n2812,
    n2406,
    n2340
  );


  or
  g2928
  (
    n2903,
    n2207,
    n2849,
    n2429,
    n2351
  );


  or
  g2929
  (
    n2890,
    n2734,
    n2821,
    n2362,
    n2460
  );


  or
  g2930
  (
    n2946,
    n2400,
    n2852,
    n2311,
    n2468
  );


  nand
  g2931
  (
    n2882,
    n2348,
    n2210,
    n2475,
    n2784
  );


  nand
  g2932
  (
    n2939,
    n2279,
    n2382,
    n2847,
    n2196
  );


  xnor
  g2933
  (
    n2912,
    n2350,
    n2190,
    n2218,
    n2855
  );


  and
  g2934
  (
    n2870,
    n2731,
    n2276,
    n2834,
    n2392
  );


  nand
  g2935
  (
    n2975,
    n2844,
    n2727,
    n2447,
    n2785
  );


  nand
  g2936
  (
    n2895,
    n2366,
    n2730,
    n2372,
    n2788
  );


  and
  g2937
  (
    n2928,
    n2741,
    n2792,
    n2825,
    n2344
  );


  or
  g2938
  (
    n2897,
    n2742,
    n2732,
    n2728,
    n2267
  );


  or
  g2939
  (
    n2952,
    n2476,
    n2424,
    n2197,
    n2215
  );


  nand
  g2940
  (
    n2899,
    n2211,
    n2301,
    n2423,
    n2731
  );


  xor
  g2941
  (
    n2916,
    n2388,
    n2229,
    n2225,
    n2729
  );


  or
  g2942
  (
    n2883,
    n2320,
    n2847,
    n2836,
    n2420
  );


  xnor
  g2943
  (
    n2874,
    n2339,
    n2238,
    n2245,
    n2851
  );


  nand
  g2944
  (
    n2872,
    n2777,
    n2857,
    n2322,
    n2742
  );


  or
  g2945
  (
    n2933,
    n2289,
    n2298,
    n2454,
    n2732
  );


  nand
  g2946
  (
    n2910,
    n2730,
    n2385,
    n2409,
    n2472
  );


  nand
  g2947
  (
    n2957,
    n2419,
    n2257,
    n2855,
    n2297
  );


  xor
  g2948
  (
    n2891,
    n2782,
    n2194,
    n2375,
    n2453
  );


  xnor
  g2949
  (
    n2983,
    n2904,
    n2866,
    n2972,
    n2953
  );


  or
  g2950
  (
    n2982,
    n2967,
    n2965,
    n2928,
    n2884
  );


  xnor
  g2951
  (
    n2996,
    n2958,
    n2864,
    n2919,
    n2966
  );


  xnor
  g2952
  (
    n2999,
    n2932,
    n2913,
    n2960,
    n2931
  );


  nor
  g2953
  (
    n3002,
    n2896,
    n2969,
    n2879,
    n2892
  );


  or
  g2954
  (
    n2985,
    n2881,
    n2954,
    n2889,
    n2915
  );


  and
  g2955
  (
    n3008,
    n2917,
    n2951,
    n2894,
    n2924
  );


  xor
  g2956
  (
    n2984,
    n2937,
    n2907,
    n2880,
    n2926
  );


  nand
  g2957
  (
    n2994,
    n2899,
    n2925,
    n2883,
    n2962
  );


  or
  g2958
  (
    n2992,
    n2968,
    n2922,
    n2959,
    n2961
  );


  xnor
  g2959
  (
    n2995,
    n2882,
    n2905,
    n2916,
    n2934
  );


  and
  g2960
  (
    n2993,
    n2940,
    n2901,
    n2971,
    n2930
  );


  nor
  g2961
  (
    n3000,
    n2888,
    n2963,
    n2955,
    n2895
  );


  and
  g2962
  (
    n3001,
    n2885,
    n2929,
    n2875,
    n2877
  );


  and
  g2963
  (
    n2987,
    n2943,
    n2903,
    n2911,
    n2949
  );


  nand
  g2964
  (
    n3006,
    n2898,
    n2910,
    n2941,
    n2908
  );


  nand
  g2965
  (
    n2988,
    n2870,
    n2876,
    n2873,
    n2869
  );


  or
  g2966
  (
    n2991,
    n2923,
    n2914,
    n2956,
    n2957
  );


  xnor
  g2967
  (
    n2998,
    n2862,
    n2947,
    n2867,
    n2933
  );


  nor
  g2968
  (
    n3007,
    n2906,
    n2891,
    n2918,
    n2921
  );


  xnor
  g2969
  (
    n3005,
    n2871,
    n2865,
    n2948,
    n2886
  );


  nand
  g2970
  (
    n3004,
    n2950,
    n2927,
    n2964,
    n2887
  );


  nand
  g2971
  (
    n2986,
    n2872,
    n2897,
    n2902,
    n2920
  );


  and
  g2972
  (
    n2997,
    n2973,
    n2938,
    n2945,
    n2946
  );


  xor
  g2973
  (
    n2990,
    n2893,
    n2909,
    n2890,
    n2935
  );


  nand
  g2974
  (
    n3003,
    n2942,
    n2900,
    n2912,
    n2939
  );


  nand
  g2975
  (
    n2989,
    n2878,
    n2874,
    n2936,
    n2868
  );


  xnor
  g2976
  (
    n3009,
    n2970,
    n2863,
    n2952,
    n2944
  );


  and
  g2977
  (
    n3024,
    n2861,
    n2861,
    n3002,
    n2992
  );


  nand
  g2978
  (
    n3016,
    n2979,
    n2774,
    n2986,
    n2773
  );


  nand
  g2979
  (
    n3019,
    n2993,
    n2772,
    n3008,
    n2984
  );


  nor
  g2980
  (
    n3017,
    n3006,
    n2999,
    n2773,
    n2860
  );


  xor
  g2981
  (
    n3014,
    n2774,
    n2998,
    n2990,
    n2996
  );


  and
  g2982
  (
    n3020,
    n2773,
    n2861,
    n2772
  );


  xor
  g2983
  (
    n3022,
    n2860,
    n2556,
    n2772,
    n3005
  );


  nor
  g2984
  (
    n3023,
    n2774,
    n2978,
    n2991,
    n3007
  );


  and
  g2985
  (
    n3021,
    n2774,
    n2529,
    n3001,
    n3000
  );


  or
  g2986
  (
    n3015,
    n2997,
    n2555,
    n2553,
    n3009
  );


  nor
  g2987
  (
    n3013,
    n2975,
    n2987,
    n2989,
    n2771
  );


  xor
  g2988
  (
    n3011,
    n3003,
    n2773,
    n2860
  );


  or
  g2989
  (
    n3012,
    n2995,
    n2859,
    n2529,
    n2552
  );


  or
  g2990
  (
    n3010,
    n2859,
    n2974,
    n2976,
    n2977
  );


  and
  g2991
  (
    n3025,
    n3004,
    n2982,
    n2985,
    n2554
  );


  xor
  g2992
  (
    n3018,
    n2772,
    n2988,
    n2994,
    n2983
  );


  not
  g2993
  (
    n3028,
    n3018
  );


  buf
  g2994
  (
    n3027,
    n3017
  );


  nor
  g2995
  (
    n3026,
    n3014,
    n3011,
    n3019,
    n3010
  );


  and
  g2996
  (
    n3029,
    n3012,
    n3015,
    n3013,
    n3016
  );


  nand
  g2997
  (
    n3030,
    n3029,
    n3020,
    n2980,
    n3024
  );


  xnor
  g2998
  (
    KeyWire_0_2,
    n3022,
    n3021,
    n3026,
    n3025
  );


  and
  g2999
  (
    n3031,
    n3028,
    n2981,
    n3027,
    n3023
  );


  xnor
  KeyGate_0_0
  (
    n286,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1525,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n3032,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n511,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1846,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1892,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n2710,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n350,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n35,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n2268,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n252,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1874,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n953,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n2338,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1729,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n2290,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1368,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n2344,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n2412,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n215,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n599,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n999,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n2578,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n2636,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n951,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n648,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n174,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n694,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1919,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1010,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n1626,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n1558,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

