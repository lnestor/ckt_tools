

module Stat_100_410
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n111,
  n106,
  n124,
  n110,
  n104,
  n132,
  n129,
  n125,
  n118,
  n119,
  n121,
  n108,
  n102,
  n109,
  n115,
  n112,
  n130,
  n123,
  n128,
  n101,
  n120,
  n131,
  n107,
  n103,
  n113,
  n117,
  n122,
  n126,
  n116,
  n105,
  n114,
  n127
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n111;output n106;output n124;output n110;output n104;output n132;output n129;output n125;output n118;output n119;output n121;output n108;output n102;output n109;output n115;output n112;output n130;output n123;output n128;output n101;output n120;output n131;output n107;output n103;output n113;output n117;output n122;output n126;output n116;output n105;output n114;output n127;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyNOTWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyWire_0_32;wire KeyNOTWire_0_32;wire KeyWire_0_33;wire KeyNOTWire_0_33;wire KeyWire_0_34;wire KeyNOTWire_0_34;wire KeyWire_0_35;wire KeyWire_0_36;wire KeyWire_0_37;wire KeyNOTWire_0_37;wire KeyWire_0_38;wire KeyWire_0_39;wire KeyNOTWire_0_39;wire KeyWire_0_40;wire KeyWire_0_41;wire KeyNOTWire_0_41;wire KeyWire_0_42;wire KeyWire_0_43;wire KeyWire_0_44;wire KeyWire_0_45;wire KeyNOTWire_0_45;wire KeyWire_0_46;wire KeyWire_0_47;wire KeyNOTWire_0_47;wire KeyWire_0_48;wire KeyWire_0_49;wire KeyNOTWire_0_49;wire KeyWire_0_50;wire KeyWire_0_51;wire KeyWire_0_52;wire KeyWire_0_53;wire KeyWire_0_54;wire KeyNOTWire_0_54;wire KeyWire_0_55;wire KeyWire_0_56;wire KeyWire_0_57;wire KeyWire_0_58;wire KeyNOTWire_0_58;wire KeyWire_0_59;wire KeyWire_0_60;wire KeyWire_0_61;wire KeyWire_0_62;wire KeyWire_0_63;wire KeyNOTWire_0_63;

  buf
  g0
  (
    KeyWire_0_45,
    n1
  );


  buf
  g1
  (
    KeyWire_0_61,
    n2
  );


  buf
  g2
  (
    KeyWire_0_7,
    n2
  );


  buf
  g3
  (
    KeyWire_0_56,
    n1
  );


  buf
  g4
  (
    n36,
    n1
  );


  buf
  g5
  (
    KeyWire_0_13,
    n34
  );


  not
  g6
  (
    KeyWire_0_29,
    n37
  );


  buf
  g7
  (
    KeyWire_0_58,
    n34
  );


  buf
  g8
  (
    n50,
    n34
  );


  buf
  g9
  (
    n53,
    n35
  );


  not
  g10
  (
    n46,
    n33
  );


  not
  g11
  (
    KeyWire_0_11,
    n36
  );


  buf
  g12
  (
    KeyWire_0_38,
    n35
  );


  not
  g13
  (
    KeyWire_0_47,
    n35
  );


  buf
  g14
  (
    KeyWire_0_36,
    n33
  );


  buf
  g15
  (
    n48,
    n37
  );


  buf
  g16
  (
    n54,
    n36
  );


  buf
  g17
  (
    KeyWire_0_43,
    n36
  );


  not
  g18
  (
    n41,
    n36
  );


  buf
  g19
  (
    n39,
    n34
  );


  not
  g20
  (
    KeyWire_0_24,
    n37
  );


  buf
  g21
  (
    KeyWire_0_52,
    n35
  );


  buf
  g22
  (
    KeyWire_0_3,
    n33
  );


  buf
  g23
  (
    KeyWire_0_14,
    n37
  );


  buf
  g24
  (
    n96,
    n54
  );


  buf
  g25
  (
    KeyWire_0_20,
    n40
  );


  not
  g26
  (
    n93,
    n54
  );


  not
  g27
  (
    KeyWire_0_19,
    n45
  );


  buf
  g28
  (
    n85,
    n9
  );


  buf
  g29
  (
    KeyWire_0_44,
    n26
  );


  xnor
  g30
  (
    KeyWire_0_53,
    n31,
    n47,
    n48
  );


  nor
  g31
  (
    KeyWire_0_22,
    n28,
    n31,
    n18,
    n4
  );


  xor
  g32
  (
    n88,
    n28,
    n38,
    n16,
    n48
  );


  xnor
  g33
  (
    n98,
    n53,
    n29,
    n14,
    n25
  );


  xor
  g34
  (
    n92,
    n16,
    n5,
    n28,
    n43
  );


  or
  g35
  (
    n82,
    n22,
    n19,
    n6,
    n21
  );


  xnor
  g36
  (
    KeyWire_0_42,
    n52,
    n10,
    n7,
    n18
  );


  xor
  g37
  (
    KeyWire_0_28,
    n22,
    n9,
    n42,
    n26
  );


  xnor
  g38
  (
    KeyWire_0_2,
    n44,
    n6,
    n32,
    n55
  );


  nor
  g39
  (
    KeyWire_0_1,
    n38,
    n25,
    n4,
    n41
  );


  xnor
  g40
  (
    n70,
    n39,
    n46,
    n49,
    n13
  );


  nor
  g41
  (
    n95,
    n27,
    n27,
    n21,
    n46
  );


  and
  g42
  (
    KeyWire_0_57,
    n25,
    n47,
    n23,
    n3
  );


  nor
  g43
  (
    KeyWire_0_26,
    n46,
    n23,
    n49,
    n19
  );


  and
  g44
  (
    KeyWire_0_59,
    n43,
    n13,
    n53,
    n2
  );


  or
  g45
  (
    KeyWire_0_16,
    n5,
    n12,
    n25,
    n56
  );


  and
  g46
  (
    KeyWire_0_60,
    n50,
    n55,
    n40,
    n29
  );


  nand
  g47
  (
    KeyWire_0_12,
    n7,
    n13,
    n39,
    n52
  );


  nand
  g48
  (
    KeyWire_0_6,
    n17,
    n32,
    n30
  );


  nor
  g49
  (
    n81,
    n18,
    n51,
    n45,
    n12
  );


  nand
  g50
  (
    KeyWire_0_15,
    n6,
    n24,
    n30,
    n28
  );


  nand
  g51
  (
    KeyWire_0_5,
    n24,
    n49,
    n27,
    n56
  );


  nand
  g52
  (
    KeyWire_0_63,
    n14,
    n11,
    n3,
    n26
  );


  and
  g53
  (
    KeyWire_0_55,
    n17,
    n27,
    n9,
    n41
  );


  nand
  g54
  (
    n59,
    n12,
    n41,
    n3,
    n8
  );


  and
  g55
  (
    KeyWire_0_30,
    n53,
    n47,
    n51,
    n44
  );


  and
  g56
  (
    KeyWire_0_8,
    n8,
    n44,
    n56,
    n24
  );


  nor
  g57
  (
    n77,
    n19,
    n17,
    n15,
    n31
  );


  and
  g58
  (
    KeyWire_0_48,
    n14,
    n15,
    n30,
    n20
  );


  xor
  g59
  (
    KeyWire_0_10,
    n23,
    n32,
    n8,
    n20
  );


  or
  g60
  (
    KeyWire_0_31,
    n31,
    n43,
    n42,
    n10
  );


  and
  g61
  (
    n74,
    n38,
    n51,
    n55,
    n11
  );


  xnor
  g62
  (
    n62,
    n29,
    n54,
    n50,
    n52
  );


  nor
  g63
  (
    KeyWire_0_18,
    n26,
    n16,
    n5,
    n15
  );


  or
  g64
  (
    n65,
    n40,
    n39,
    n7,
    n10
  );


  xnor
  g65
  (
    KeyWire_0_37,
    n32,
    n24,
    n22,
    n48
  );


  xnor
  g66
  (
    n66,
    n50,
    n21,
    n29,
    n4
  );


  nand
  g67
  (
    n97,
    n20,
    n42,
    n11,
    n45
  );


  xnor
  g68
  (
    KeyWire_0_40,
    n72,
    n78,
    n92,
    n59
  );


  nor
  g69
  (
    n117,
    n81,
    n93,
    n80,
    n85
  );


  or
  g70
  (
    KeyWire_0_27,
    n59,
    n74,
    n65,
    n93
  );


  xor
  g71
  (
    KeyWire_0_49,
    n80,
    n95,
    n67,
    n97
  );


  xor
  g72
  (
    KeyWire_0_34,
    n100,
    n84,
    n76,
    n71
  );


  nor
  g73
  (
    n124,
    n86,
    n62,
    n90,
    n59
  );


  and
  g74
  (
    KeyWire_0_39,
    n77,
    n72,
    n70,
    n63
  );


  nor
  g75
  (
    n116,
    n97,
    n83,
    n95
  );


  or
  g76
  (
    KeyWire_0_0,
    n76,
    n64,
    n80,
    n96
  );


  xnor
  g77
  (
    n103,
    n91,
    n66,
    n58,
    n98
  );


  or
  g78
  (
    n129,
    n70,
    n69,
    n62,
    n81
  );


  xnor
  g79
  (
    KeyWire_0_54,
    n98,
    n60,
    n100,
    n78
  );


  xnor
  g80
  (
    KeyWire_0_50,
    n99,
    n70,
    n85,
    n87
  );


  xnor
  g81
  (
    n121,
    n88,
    n61,
    n65,
    n77
  );


  and
  g82
  (
    KeyWire_0_46,
    n73,
    n67,
    n89,
    n63
  );


  and
  g83
  (
    KeyWire_0_4,
    n90,
    n73,
    n78,
    n72
  );


  and
  g84
  (
    KeyWire_0_21,
    n87,
    n92,
    n68,
    n79
  );


  xor
  g85
  (
    KeyWire_0_35,
    n94,
    n75,
    n74,
    n91
  );


  xor
  g86
  (
    n113,
    n87,
    n96,
    n92,
    n71
  );


  xnor
  g87
  (
    KeyWire_0_33,
    n67,
    n75,
    n94,
    n73
  );


  nor
  g88
  (
    KeyWire_0_62,
    n64,
    n71,
    n89,
    n79
  );


  or
  g89
  (
    n107,
    n63,
    n83,
    n85,
    n65
  );


  xnor
  g90
  (
    KeyWire_0_32,
    n77,
    n74,
    n88,
    n68
  );


  nor
  g91
  (
    KeyWire_0_17,
    n99,
    n60,
    n86,
    n75
  );


  nand
  g92
  (
    KeyWire_0_41,
    n99,
    n86,
    n95,
    n66
  );


  nand
  g93
  (
    n123,
    n96,
    n81,
    n57,
    n62
  );


  nor
  g94
  (
    KeyWire_0_9,
    n82,
    n84,
    n88,
    n91
  );


  xnor
  g95
  (
    n122,
    n61,
    n98,
    n90,
    n69
  );


  and
  g96
  (
    n125,
    n64,
    n61,
    n66,
    n84
  );


  xnor
  g97
  (
    KeyWire_0_23,
    n60,
    n69,
    n76,
    n68
  );


  xnor
  g98
  (
    KeyWire_0_51,
    n93,
    n79,
    n97,
    n82
  );


  xor
  g99
  (
    KeyWire_0_25,
    n89,
    n100,
    n82,
    n94
  );


  xor
  KeyGate_0_0
  (
    n105,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n64,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n63,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n43,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n111,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n86,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n80,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n35,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n100,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n132,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n90,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n55,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n89,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n40,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n47,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n67,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n87,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n120,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n73,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n72,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n94,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n127,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n79,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n130,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n51,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n108,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n78,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n115,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n71,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n56,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n84,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n91,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n112,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n110,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n118,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n119,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n42,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n75,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n44,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n131,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    n104,
    keyIn_0_40,
    KeyWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n128,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n57,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n45,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n60,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n37,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n102,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n52,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n68,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n106,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n109,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n126,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n38,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n61,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n101,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n83,
    keyIn_0_55,
    KeyWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n33,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n99,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n49,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n58,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n69,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n34,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n114,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n76,
    KeyNOTWire_0_63
  );


endmodule


