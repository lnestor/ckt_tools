

module Stat_1197_31_10
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n989,
  n996,
  n990,
  n1013,
  n1017,
  n993,
  n981,
  n1014,
  n994,
  n991,
  n1008,
  n1001,
  n999,
  n992,
  n1005,
  n987,
  n997,
  n985,
  n982,
  n1004,
  n988,
  n1028,
  n1026,
  n1031,
  n1023,
  n1029,
  n1025,
  n1022,
  n1027,
  n1181,
  n1197,
  n1220,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n989;
  output n996;
  output n990;
  output n1013;
  output n1017;
  output n993;
  output n981;
  output n1014;
  output n994;
  output n991;
  output n1008;
  output n1001;
  output n999;
  output n992;
  output n1005;
  output n987;
  output n997;
  output n985;
  output n982;
  output n1004;
  output n988;
  output n1028;
  output n1026;
  output n1031;
  output n1023;
  output n1029;
  output n1025;
  output n1022;
  output n1027;
  output n1181;
  output n1197;
  output n1220;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n983;
  wire n984;
  wire n986;
  wire n995;
  wire n998;
  wire n1000;
  wire n1002;
  wire n1003;
  wire n1006;
  wire n1007;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1015;
  wire n1016;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1024;
  wire n1030;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    n78,
    n7
  );


  buf
  g1
  (
    n82,
    n13
  );


  not
  g2
  (
    n71,
    n6
  );


  not
  g3
  (
    n36,
    n8
  );


  not
  g4
  (
    n26,
    n6
  );


  not
  g5
  (
    n113,
    n11
  );


  not
  g6
  (
    n91,
    n23
  );


  not
  g7
  (
    n114,
    n6
  );


  not
  g8
  (
    n112,
    n16
  );


  buf
  g9
  (
    n81,
    n21
  );


  buf
  g10
  (
    n84,
    n6
  );


  not
  g11
  (
    n70,
    n23
  );


  buf
  g12
  (
    n25,
    n11
  );


  not
  g13
  (
    n85,
    n18
  );


  buf
  g14
  (
    n33,
    n21
  );


  not
  g15
  (
    n34,
    n13
  );


  buf
  g16
  (
    n99,
    n18
  );


  not
  g17
  (
    n64,
    n4
  );


  not
  g18
  (
    n56,
    n8
  );


  not
  g19
  (
    n67,
    n16
  );


  buf
  g20
  (
    n59,
    n10
  );


  not
  g21
  (
    n57,
    n14
  );


  not
  g22
  (
    n51,
    n4
  );


  not
  g23
  (
    n89,
    n15
  );


  not
  g24
  (
    n100,
    n19
  );


  not
  g25
  (
    n106,
    n20
  );


  not
  g26
  (
    n76,
    n13
  );


  not
  g27
  (
    n29,
    n18
  );


  not
  g28
  (
    n44,
    n1
  );


  buf
  g29
  (
    n115,
    n20
  );


  buf
  g30
  (
    n88,
    n16
  );


  buf
  g31
  (
    n94,
    n19
  );


  buf
  g32
  (
    n48,
    n1
  );


  not
  g33
  (
    n80,
    n22
  );


  buf
  g34
  (
    n75,
    n23
  );


  not
  g35
  (
    n43,
    n19
  );


  buf
  g36
  (
    n32,
    n3
  );


  not
  g37
  (
    n60,
    n9
  );


  buf
  g38
  (
    n53,
    n9
  );


  not
  g39
  (
    n45,
    n3
  );


  buf
  g40
  (
    n95,
    n17
  );


  not
  g41
  (
    n68,
    n12
  );


  not
  g42
  (
    n27,
    n16
  );


  buf
  g43
  (
    n101,
    n2
  );


  buf
  g44
  (
    n55,
    n1
  );


  buf
  g45
  (
    n58,
    n11
  );


  buf
  g46
  (
    n105,
    n17
  );


  not
  g47
  (
    n65,
    n21
  );


  not
  g48
  (
    n49,
    n4
  );


  buf
  g49
  (
    n103,
    n15
  );


  buf
  g50
  (
    n31,
    n17
  );


  buf
  g51
  (
    n111,
    n20
  );


  not
  g52
  (
    n83,
    n12
  );


  not
  g53
  (
    n52,
    n10
  );


  buf
  g54
  (
    n73,
    n8
  );


  not
  g55
  (
    n97,
    n7
  );


  not
  g56
  (
    n28,
    n23
  );


  not
  g57
  (
    n24,
    n10
  );


  not
  g58
  (
    n61,
    n14
  );


  not
  g59
  (
    n92,
    n2
  );


  buf
  g60
  (
    n30,
    n4
  );


  buf
  g61
  (
    n47,
    n12
  );


  buf
  g62
  (
    n86,
    n15
  );


  not
  g63
  (
    n69,
    n12
  );


  not
  g64
  (
    n40,
    n9
  );


  buf
  g65
  (
    n63,
    n10
  );


  buf
  g66
  (
    n93,
    n1
  );


  not
  g67
  (
    n98,
    n3
  );


  buf
  g68
  (
    n108,
    n14
  );


  not
  g69
  (
    n109,
    n19
  );


  not
  g70
  (
    n66,
    n5
  );


  buf
  g71
  (
    n79,
    n3
  );


  not
  g72
  (
    n104,
    n15
  );


  buf
  g73
  (
    n39,
    n14
  );


  not
  g74
  (
    n107,
    n18
  );


  buf
  g75
  (
    n102,
    n21
  );


  not
  g76
  (
    n110,
    n22
  );


  buf
  g77
  (
    n90,
    n13
  );


  buf
  g78
  (
    n74,
    n7
  );


  not
  g79
  (
    n54,
    n2
  );


  not
  g80
  (
    n50,
    n22
  );


  not
  g81
  (
    n87,
    n22
  );


  not
  g82
  (
    n96,
    n5
  );


  not
  g83
  (
    n77,
    n11
  );


  not
  g84
  (
    n72,
    n17
  );


  not
  g85
  (
    n35,
    n2
  );


  not
  g86
  (
    n38,
    n5
  );


  not
  g87
  (
    n42,
    n7
  );


  buf
  g88
  (
    n62,
    n8
  );


  not
  g89
  (
    n37,
    n5
  );


  not
  g90
  (
    n41,
    n20
  );


  buf
  g91
  (
    n46,
    n9
  );


  not
  g92
  (
    n355,
    n77
  );


  buf
  g93
  (
    n343,
    n111
  );


  not
  g94
  (
    n246,
    n112
  );


  not
  g95
  (
    n414,
    n42
  );


  buf
  g96
  (
    n283,
    n31
  );


  buf
  g97
  (
    n444,
    n71
  );


  not
  g98
  (
    n135,
    n30
  );


  buf
  g99
  (
    n367,
    n25
  );


  not
  g100
  (
    KeyWire_0_30,
    n85
  );


  buf
  g101
  (
    n124,
    n38
  );


  buf
  g102
  (
    n420,
    n37
  );


  buf
  g103
  (
    n276,
    n108
  );


  not
  g104
  (
    n482,
    n57
  );


  not
  g105
  (
    n456,
    n34
  );


  not
  g106
  (
    n223,
    n45
  );


  not
  g107
  (
    n141,
    n46
  );


  buf
  g108
  (
    n221,
    n102
  );


  not
  g109
  (
    n396,
    n42
  );


  buf
  g110
  (
    n169,
    n103
  );


  buf
  g111
  (
    n303,
    n110
  );


  not
  g112
  (
    n455,
    n95
  );


  buf
  g113
  (
    n332,
    n93
  );


  not
  g114
  (
    n237,
    n47
  );


  not
  g115
  (
    n173,
    n80
  );


  buf
  g116
  (
    n277,
    n104
  );


  buf
  g117
  (
    n401,
    n40
  );


  not
  g118
  (
    n405,
    n49
  );


  buf
  g119
  (
    n447,
    n62
  );


  not
  g120
  (
    n333,
    n27
  );


  not
  g121
  (
    n361,
    n76
  );


  not
  g122
  (
    n296,
    n70
  );


  buf
  g123
  (
    n418,
    n50
  );


  not
  g124
  (
    n366,
    n54
  );


  buf
  g125
  (
    n218,
    n59
  );


  not
  g126
  (
    n119,
    n54
  );


  buf
  g127
  (
    n442,
    n67
  );


  not
  g128
  (
    n352,
    n75
  );


  not
  g129
  (
    n369,
    n97
  );


  not
  g130
  (
    n229,
    n107
  );


  buf
  g131
  (
    n335,
    n77
  );


  buf
  g132
  (
    n269,
    n69
  );


  not
  g133
  (
    n408,
    n73
  );


  buf
  g134
  (
    n323,
    n56
  );


  not
  g135
  (
    n454,
    n79
  );


  buf
  g136
  (
    n469,
    n49
  );


  buf
  g137
  (
    n285,
    n44
  );


  buf
  g138
  (
    n353,
    n98
  );


  not
  g139
  (
    n232,
    n108
  );


  buf
  g140
  (
    n429,
    n42
  );


  buf
  g141
  (
    n432,
    n102
  );


  not
  g142
  (
    n397,
    n34
  );


  not
  g143
  (
    n172,
    n85
  );


  buf
  g144
  (
    n437,
    n112
  );


  not
  g145
  (
    n165,
    n75
  );


  buf
  g146
  (
    n300,
    n110
  );


  not
  g147
  (
    n449,
    n75
  );


  buf
  g148
  (
    n242,
    n33
  );


  not
  g149
  (
    n189,
    n89
  );


  not
  g150
  (
    n194,
    n94
  );


  not
  g151
  (
    n208,
    n61
  );


  buf
  g152
  (
    n306,
    n82
  );


  buf
  g153
  (
    n328,
    n85
  );


  buf
  g154
  (
    n346,
    n27
  );


  not
  g155
  (
    n130,
    n84
  );


  not
  g156
  (
    n268,
    n82
  );


  buf
  g157
  (
    n294,
    n111
  );


  not
  g158
  (
    n251,
    n91
  );


  buf
  g159
  (
    n249,
    n101
  );


  not
  g160
  (
    n211,
    n97
  );


  not
  g161
  (
    n382,
    n41
  );


  buf
  g162
  (
    n468,
    n106
  );


  not
  g163
  (
    n471,
    n48
  );


  not
  g164
  (
    n185,
    n30
  );


  not
  g165
  (
    n458,
    n71
  );


  buf
  g166
  (
    n406,
    n99
  );


  buf
  g167
  (
    n433,
    n38
  );


  buf
  g168
  (
    n383,
    n65
  );


  not
  g169
  (
    n461,
    n92
  );


  buf
  g170
  (
    n290,
    n107
  );


  not
  g171
  (
    KeyWire_0_15,
    n46
  );


  not
  g172
  (
    n476,
    n81
  );


  not
  g173
  (
    n215,
    n48
  );


  not
  g174
  (
    n395,
    n61
  );


  not
  g175
  (
    n257,
    n104
  );


  buf
  g176
  (
    KeyWire_0_4,
    n38
  );


  buf
  g177
  (
    n180,
    n58
  );


  not
  g178
  (
    KeyWire_0_22,
    n114
  );


  not
  g179
  (
    n326,
    n68
  );


  not
  g180
  (
    n273,
    n113
  );


  buf
  g181
  (
    n117,
    n68
  );


  buf
  g182
  (
    n133,
    n28
  );


  buf
  g183
  (
    n375,
    n98
  );


  not
  g184
  (
    n402,
    n70
  );


  not
  g185
  (
    n310,
    n28
  );


  buf
  g186
  (
    n329,
    n72
  );


  not
  g187
  (
    n219,
    n68
  );


  not
  g188
  (
    n260,
    n35
  );


  not
  g189
  (
    n261,
    n51
  );


  not
  g190
  (
    n190,
    n50
  );


  buf
  g191
  (
    n132,
    n62
  );


  not
  g192
  (
    n201,
    n109
  );


  not
  g193
  (
    n336,
    n44
  );


  not
  g194
  (
    n407,
    n70
  );


  buf
  g195
  (
    n467,
    n76
  );


  not
  g196
  (
    n378,
    n46
  );


  not
  g197
  (
    n118,
    n66
  );


  buf
  g198
  (
    n143,
    n115
  );


  buf
  g199
  (
    n388,
    n52
  );


  buf
  g200
  (
    n274,
    n100
  );


  not
  g201
  (
    n216,
    n49
  );


  buf
  g202
  (
    n145,
    n109
  );


  not
  g203
  (
    n195,
    n50
  );


  not
  g204
  (
    n236,
    n75
  );


  buf
  g205
  (
    n439,
    n67
  );


  not
  g206
  (
    n428,
    n43
  );


  buf
  g207
  (
    n252,
    n57
  );


  not
  g208
  (
    n364,
    n40
  );


  not
  g209
  (
    n160,
    n100
  );


  not
  g210
  (
    n295,
    n92
  );


  buf
  g211
  (
    n142,
    n36
  );


  not
  g212
  (
    n341,
    n83
  );


  not
  g213
  (
    n234,
    n39
  );


  buf
  g214
  (
    n187,
    n71
  );


  buf
  g215
  (
    n386,
    n27
  );


  buf
  g216
  (
    n146,
    n103
  );


  not
  g217
  (
    n230,
    n84
  );


  not
  g218
  (
    n435,
    n41
  );


  buf
  g219
  (
    n253,
    n61
  );


  buf
  g220
  (
    n284,
    n101
  );


  not
  g221
  (
    n411,
    n51
  );


  not
  g222
  (
    n241,
    n91
  );


  not
  g223
  (
    n156,
    n76
  );


  not
  g224
  (
    n421,
    n53
  );


  not
  g225
  (
    n213,
    n110
  );


  buf
  g226
  (
    n379,
    n69
  );


  buf
  g227
  (
    n280,
    n47
  );


  buf
  g228
  (
    n123,
    n26
  );


  buf
  g229
  (
    n391,
    n55
  );


  buf
  g230
  (
    n116,
    n65
  );


  not
  g231
  (
    n417,
    n57
  );


  not
  g232
  (
    n462,
    n29
  );


  buf
  g233
  (
    n440,
    n51
  );


  buf
  g234
  (
    n199,
    n104
  );


  buf
  g235
  (
    n314,
    n72
  );


  not
  g236
  (
    n394,
    n69
  );


  not
  g237
  (
    n392,
    n30
  );


  not
  g238
  (
    n272,
    n76
  );


  not
  g239
  (
    n245,
    n80
  );


  buf
  g240
  (
    n321,
    n113
  );


  buf
  g241
  (
    n360,
    n32
  );


  buf
  g242
  (
    n424,
    n43
  );


  not
  g243
  (
    n288,
    n64
  );


  not
  g244
  (
    n174,
    n24
  );


  not
  g245
  (
    n316,
    n29
  );


  not
  g246
  (
    n409,
    n79
  );


  buf
  g247
  (
    n349,
    n109
  );


  not
  g248
  (
    n224,
    n100
  );


  not
  g249
  (
    n178,
    n36
  );


  not
  g250
  (
    n466,
    n24
  );


  buf
  g251
  (
    n415,
    n106
  );


  not
  g252
  (
    n176,
    n31
  );


  not
  g253
  (
    n149,
    n33
  );


  not
  g254
  (
    n450,
    n105
  );


  not
  g255
  (
    n473,
    n55
  );


  not
  g256
  (
    n151,
    n33
  );


  not
  g257
  (
    n270,
    n55
  );


  not
  g258
  (
    n319,
    n26
  );


  not
  g259
  (
    n254,
    n98
  );


  not
  g260
  (
    n400,
    n47
  );


  buf
  g261
  (
    n431,
    n68
  );


  buf
  g262
  (
    n197,
    n82
  );


  buf
  g263
  (
    n287,
    n41
  );


  buf
  g264
  (
    n203,
    n77
  );


  not
  g265
  (
    n315,
    n114
  );


  not
  g266
  (
    n330,
    n54
  );


  buf
  g267
  (
    n480,
    n113
  );


  not
  g268
  (
    n264,
    n102
  );


  buf
  g269
  (
    n479,
    n86
  );


  not
  g270
  (
    n265,
    n45
  );


  not
  g271
  (
    n168,
    n115
  );


  buf
  g272
  (
    n472,
    n43
  );


  not
  g273
  (
    n144,
    n34
  );


  buf
  g274
  (
    n183,
    n52
  );


  not
  g275
  (
    n318,
    n59
  );


  buf
  g276
  (
    n292,
    n91
  );


  buf
  g277
  (
    n210,
    n56
  );


  not
  g278
  (
    n298,
    n48
  );


  not
  g279
  (
    n281,
    n101
  );


  buf
  g280
  (
    n351,
    n93
  );


  not
  g281
  (
    n381,
    n59
  );


  not
  g282
  (
    n275,
    n83
  );


  buf
  g283
  (
    n259,
    n24
  );


  not
  g284
  (
    n419,
    n107
  );


  buf
  g285
  (
    n175,
    n53
  );


  buf
  g286
  (
    n436,
    n92
  );


  buf
  g287
  (
    n416,
    n90
  );


  buf
  g288
  (
    n475,
    n115
  );


  not
  g289
  (
    n302,
    n94
  );


  buf
  g290
  (
    n404,
    n105
  );


  buf
  g291
  (
    n164,
    n81
  );


  buf
  g292
  (
    n181,
    n67
  );


  not
  g293
  (
    n297,
    n73
  );


  buf
  g294
  (
    n425,
    n106
  );


  buf
  g295
  (
    n412,
    n59
  );


  buf
  g296
  (
    n247,
    n63
  );


  buf
  g297
  (
    n387,
    n83
  );


  not
  g298
  (
    n138,
    n72
  );


  not
  g299
  (
    n363,
    n115
  );


  not
  g300
  (
    n122,
    n53
  );


  buf
  g301
  (
    n374,
    n31
  );


  buf
  g302
  (
    n368,
    n107
  );


  not
  g303
  (
    n289,
    n24
  );


  buf
  g304
  (
    n121,
    n48
  );


  not
  g305
  (
    n293,
    n64
  );


  not
  g306
  (
    n163,
    n58
  );


  not
  g307
  (
    n186,
    n37
  );


  buf
  g308
  (
    n129,
    n96
  );


  not
  g309
  (
    n147,
    n96
  );


  buf
  g310
  (
    n354,
    n85
  );


  not
  g311
  (
    n474,
    n93
  );


  not
  g312
  (
    n206,
    n32
  );


  not
  g313
  (
    n477,
    n73
  );


  buf
  g314
  (
    n339,
    n66
  );


  not
  g315
  (
    n128,
    n78
  );


  buf
  g316
  (
    n350,
    n79
  );


  not
  g317
  (
    n157,
    n86
  );


  buf
  g318
  (
    n430,
    n65
  );


  buf
  g319
  (
    n322,
    n81
  );


  buf
  g320
  (
    n154,
    n102
  );


  buf
  g321
  (
    n403,
    n35
  );


  not
  g322
  (
    n120,
    n114
  );


  buf
  g323
  (
    n198,
    n39
  );


  not
  g324
  (
    n207,
    n97
  );


  not
  g325
  (
    n158,
    n43
  );


  buf
  g326
  (
    n214,
    n113
  );


  not
  g327
  (
    n342,
    n36
  );


  buf
  g328
  (
    n389,
    n89
  );


  buf
  g329
  (
    n271,
    n94
  );


  buf
  g330
  (
    n131,
    n90
  );


  buf
  g331
  (
    n324,
    n33
  );


  not
  g332
  (
    n347,
    n66
  );


  not
  g333
  (
    n423,
    n49
  );


  not
  g334
  (
    n313,
    n84
  );


  buf
  g335
  (
    n126,
    n82
  );


  buf
  g336
  (
    n209,
    n64
  );


  not
  g337
  (
    n483,
    n87
  );


  buf
  g338
  (
    n243,
    n103
  );


  buf
  g339
  (
    n240,
    n94
  );


  not
  g340
  (
    n202,
    n37
  );


  not
  g341
  (
    n307,
    n30
  );


  not
  g342
  (
    n309,
    n69
  );


  buf
  g343
  (
    n345,
    n112
  );


  buf
  g344
  (
    n212,
    n70
  );


  not
  g345
  (
    n365,
    n95
  );


  buf
  g346
  (
    n153,
    n88
  );


  not
  g347
  (
    n348,
    n42
  );


  not
  g348
  (
    n312,
    n109
  );


  buf
  g349
  (
    n334,
    n46
  );


  buf
  g350
  (
    n399,
    n90
  );


  buf
  g351
  (
    n279,
    n96
  );


  not
  g352
  (
    n377,
    n52
  );


  buf
  g353
  (
    n459,
    n31
  );


  not
  g354
  (
    n443,
    n78
  );


  buf
  g355
  (
    n337,
    n87
  );


  not
  g356
  (
    n311,
    n83
  );


  buf
  g357
  (
    n325,
    n60
  );


  buf
  g358
  (
    n193,
    n40
  );


  buf
  g359
  (
    n262,
    n56
  );


  buf
  g360
  (
    n255,
    n91
  );


  buf
  g361
  (
    n136,
    n105
  );


  buf
  g362
  (
    n179,
    n64
  );


  buf
  g363
  (
    KeyWire_0_11,
    n44
  );


  not
  g364
  (
    KeyWire_0_28,
    n87
  );


  buf
  g365
  (
    n463,
    n114
  );


  buf
  g366
  (
    KeyWire_0_19,
    n86
  );


  buf
  g367
  (
    n286,
    n95
  );


  buf
  g368
  (
    n384,
    n74
  );


  not
  g369
  (
    n304,
    n89
  );


  not
  g370
  (
    n267,
    n28
  );


  buf
  g371
  (
    n413,
    n101
  );


  not
  g372
  (
    n222,
    n73
  );


  buf
  g373
  (
    n427,
    n74
  );


  not
  g374
  (
    n170,
    n62
  );


  buf
  g375
  (
    n362,
    n104
  );


  not
  g376
  (
    n250,
    n99
  );


  buf
  g377
  (
    n305,
    n81
  );


  buf
  g378
  (
    n344,
    n98
  );


  buf
  g379
  (
    n438,
    n51
  );


  buf
  g380
  (
    n248,
    n87
  );


  not
  g381
  (
    n340,
    n50
  );


  buf
  g382
  (
    n227,
    n62
  );


  not
  g383
  (
    n448,
    n77
  );


  not
  g384
  (
    n191,
    n44
  );


  buf
  g385
  (
    n238,
    n108
  );


  not
  g386
  (
    n457,
    n99
  );


  buf
  g387
  (
    n148,
    n80
  );


  not
  g388
  (
    n372,
    n61
  );


  not
  g389
  (
    n239,
    n97
  );


  not
  g390
  (
    n452,
    n29
  );


  not
  g391
  (
    n139,
    n63
  );


  not
  g392
  (
    n184,
    n45
  );


  not
  g393
  (
    n226,
    n111
  );


  buf
  g394
  (
    n171,
    n78
  );


  not
  g395
  (
    n235,
    n88
  );


  buf
  g396
  (
    n233,
    n74
  );


  not
  g397
  (
    n200,
    n39
  );


  not
  g398
  (
    n451,
    n36
  );


  not
  g399
  (
    n358,
    n112
  );


  not
  g400
  (
    n478,
    n54
  );


  buf
  g401
  (
    n359,
    n92
  );


  buf
  g402
  (
    n263,
    n58
  );


  buf
  g403
  (
    n152,
    n65
  );


  buf
  g404
  (
    n140,
    n41
  );


  not
  g405
  (
    n150,
    n38
  );


  buf
  g406
  (
    n371,
    n32
  );


  buf
  g407
  (
    n162,
    n57
  );


  not
  g408
  (
    n182,
    n84
  );


  buf
  g409
  (
    n390,
    n86
  );


  not
  g410
  (
    n299,
    n89
  );


  buf
  g411
  (
    n177,
    n34
  );


  buf
  g412
  (
    n244,
    n35
  );


  not
  g413
  (
    n422,
    n37
  );


  buf
  g414
  (
    n445,
    n25
  );


  buf
  g415
  (
    n393,
    n47
  );


  buf
  g416
  (
    n446,
    n88
  );


  buf
  g417
  (
    n464,
    n111
  );


  not
  g418
  (
    n166,
    n25
  );


  buf
  g419
  (
    n385,
    n29
  );


  buf
  g420
  (
    n125,
    n103
  );


  not
  g421
  (
    n376,
    n45
  );


  not
  g422
  (
    n204,
    n110
  );


  not
  g423
  (
    n481,
    n60
  );


  not
  g424
  (
    n370,
    n105
  );


  buf
  g425
  (
    n127,
    n28
  );


  buf
  g426
  (
    n357,
    n106
  );


  not
  g427
  (
    n228,
    n60
  );


  not
  g428
  (
    n338,
    n39
  );


  buf
  g429
  (
    n137,
    n78
  );


  buf
  g430
  (
    n220,
    n80
  );


  buf
  g431
  (
    n301,
    n27
  );


  buf
  g432
  (
    n410,
    n26
  );


  buf
  g433
  (
    n161,
    n55
  );


  not
  g434
  (
    n134,
    n52
  );


  not
  g435
  (
    n317,
    n56
  );


  not
  g436
  (
    n453,
    n25
  );


  not
  g437
  (
    n398,
    n53
  );


  not
  g438
  (
    KeyWire_0_16,
    n58
  );


  buf
  g439
  (
    n441,
    n66
  );


  not
  g440
  (
    n460,
    n60
  );


  not
  g441
  (
    KeyWire_0_2,
    n40
  );


  buf
  g442
  (
    n434,
    n32
  );


  not
  g443
  (
    n291,
    n71
  );


  buf
  g444
  (
    n380,
    n99
  );


  not
  g445
  (
    n167,
    n96
  );


  not
  g446
  (
    n470,
    n93
  );


  not
  g447
  (
    n465,
    n26
  );


  buf
  g448
  (
    n192,
    n108
  );


  buf
  g449
  (
    n258,
    n74
  );


  buf
  g450
  (
    n426,
    n63
  );


  not
  g451
  (
    n217,
    n67
  );


  buf
  g452
  (
    n159,
    n72
  );


  not
  g453
  (
    n256,
    n63
  );


  buf
  g454
  (
    n331,
    n90
  );


  not
  g455
  (
    n356,
    n35
  );


  buf
  g456
  (
    n225,
    n95
  );


  not
  g457
  (
    n188,
    n79
  );


  buf
  g458
  (
    n196,
    n100
  );


  buf
  g459
  (
    n266,
    n88
  );


  nand
  g460
  (
    n671,
    n381,
    n379,
    n325,
    n332
  );


  and
  g461
  (
    n591,
    n411,
    n331,
    n281,
    n409
  );


  and
  g462
  (
    n701,
    n239,
    n331,
    n232,
    n367
  );


  nor
  g463
  (
    n533,
    n412,
    n276,
    n309,
    n248
  );


  nor
  g464
  (
    n517,
    n371,
    n420,
    n269,
    n397
  );


  nor
  g465
  (
    n546,
    n317,
    n330,
    n334,
    n400
  );


  and
  g466
  (
    n495,
    n385,
    n397,
    n434,
    n353
  );


  xnor
  g467
  (
    n624,
    n386,
    n426,
    n320,
    n409
  );


  and
  g468
  (
    n710,
    n336,
    n404,
    n291,
    n416
  );


  and
  g469
  (
    n650,
    n436,
    n357,
    n318,
    n245
  );


  nand
  g470
  (
    n513,
    n386,
    n345,
    n346,
    n348
  );


  nand
  g471
  (
    n580,
    n401,
    n199,
    n309,
    n362
  );


  nand
  g472
  (
    n519,
    n343,
    n408,
    n416,
    n310
  );


  and
  g473
  (
    n581,
    n322,
    n445,
    n382,
    n347
  );


  nand
  g474
  (
    n699,
    n315,
    n381,
    n228,
    n281
  );


  nand
  g475
  (
    n574,
    n344,
    n374,
    n417,
    n429
  );


  xor
  g476
  (
    n697,
    n447,
    n427,
    n245,
    n337
  );


  or
  g477
  (
    KeyWire_0_10,
    n272,
    n378,
    n306,
    n349
  );


  and
  g478
  (
    n622,
    n166,
    n312,
    n376,
    n165
  );


  or
  g479
  (
    n493,
    n259,
    n403,
    n424,
    n435
  );


  nor
  g480
  (
    n616,
    n424,
    n267,
    n238,
    n252
  );


  xnor
  g481
  (
    n549,
    n251,
    n418,
    n425,
    n436
  );


  xnor
  g482
  (
    n615,
    n313,
    n326,
    n442,
    n443
  );


  xnor
  g483
  (
    n526,
    n277,
    n421,
    n381,
    n375
  );


  xnor
  g484
  (
    KeyWire_0_14,
    n319,
    n301,
    n248,
    n293
  );


  xnor
  g485
  (
    n684,
    n296,
    n384,
    n441,
    n403
  );


  xnor
  g486
  (
    n536,
    n344,
    n338,
    n286,
    n194
  );


  xnor
  g487
  (
    n644,
    n361,
    n283,
    n119,
    n253
  );


  or
  g488
  (
    n523,
    n197,
    n355,
    n432,
    n363
  );


  or
  g489
  (
    n649,
    n255,
    n378,
    n148,
    n327
  );


  and
  g490
  (
    n494,
    n310,
    n279,
    n126,
    n180
  );


  xnor
  g491
  (
    n648,
    n396,
    n408,
    n325,
    n404
  );


  nor
  g492
  (
    n576,
    n379,
    n285,
    n236,
    n334
  );


  or
  g493
  (
    n658,
    n294,
    n297,
    n365,
    n332
  );


  or
  g494
  (
    n610,
    n383,
    n258,
    n213,
    n127
  );


  and
  g495
  (
    n510,
    n392,
    n273,
    n343,
    n121
  );


  xnor
  g496
  (
    n599,
    n395,
    n142,
    n431,
    n151
  );


  and
  g497
  (
    n543,
    n307,
    n370,
    n316,
    n225
  );


  xnor
  g498
  (
    n572,
    n153,
    n422,
    n313,
    n284
  );


  nor
  g499
  (
    n695,
    n304,
    n206,
    n239,
    n358
  );


  nor
  g500
  (
    n503,
    n150,
    n315,
    n221,
    n262
  );


  or
  g501
  (
    n601,
    n271,
    n441,
    n412,
    n269
  );


  xor
  g502
  (
    n652,
    n363,
    n161,
    n277,
    n359
  );


  xnor
  g503
  (
    n587,
    n227,
    n415,
    n308,
    n407
  );


  or
  g504
  (
    n609,
    n386,
    n124,
    n334,
    n341
  );


  xor
  g505
  (
    n507,
    n420,
    n278,
    n287,
    n139
  );


  or
  g506
  (
    n542,
    n144,
    n287,
    n292,
    n316
  );


  nor
  g507
  (
    n702,
    n242,
    n445,
    n177,
    n364
  );


  or
  g508
  (
    n515,
    n274,
    n303,
    n192,
    n332
  );


  and
  g509
  (
    n566,
    n274,
    n313,
    n307,
    n342
  );


  xor
  g510
  (
    n537,
    n435,
    n405,
    n446,
    n372
  );


  and
  g511
  (
    n489,
    n363,
    n339,
    n391,
    n223
  );


  nor
  g512
  (
    n682,
    n391,
    n414,
    n179,
    n247
  );


  and
  g513
  (
    n556,
    n211,
    n212,
    n130,
    n372
  );


  xor
  g514
  (
    n643,
    n438,
    n306,
    n333,
    n277
  );


  or
  g515
  (
    n598,
    n434,
    n388,
    n314,
    n353
  );


  and
  g516
  (
    n578,
    n406,
    n254,
    n277,
    n286
  );


  nand
  g517
  (
    n501,
    n422,
    n305,
    n356,
    n386
  );


  and
  g518
  (
    n540,
    n203,
    n198,
    n219,
    n325
  );


  xnor
  g519
  (
    n676,
    n351,
    n378,
    n385,
    n347
  );


  xor
  g520
  (
    n498,
    n350,
    n300,
    n327,
    n360
  );


  xor
  g521
  (
    n508,
    n355,
    n281,
    n217,
    n395
  );


  and
  g522
  (
    n618,
    n309,
    n276,
    n335,
    n387
  );


  nor
  g523
  (
    n569,
    n390,
    n176,
    n145,
    n288
  );


  nand
  g524
  (
    n612,
    n427,
    n371,
    n293
  );


  xnor
  g525
  (
    KeyWire_0_9,
    n331,
    n400,
    n357,
    n375
  );


  xor
  g526
  (
    n647,
    n275,
    n433,
    n292,
    n346
  );


  nor
  g527
  (
    n584,
    n403,
    n341,
    n417,
    n345
  );


  nand
  g528
  (
    n535,
    n364,
    n424,
    n254,
    n274
  );


  xnor
  g529
  (
    n593,
    n349,
    n437,
    n377,
    n322
  );


  nor
  g530
  (
    n573,
    n282,
    n445,
    n188,
    n131
  );


  nor
  g531
  (
    n512,
    n394,
    n430,
    n134,
    n332
  );


  or
  g532
  (
    n558,
    n258,
    n321,
    n259,
    n352
  );


  xnor
  g533
  (
    n655,
    n261,
    n380,
    n310,
    n238
  );


  xnor
  g534
  (
    n511,
    n225,
    n329,
    n439,
    n376
  );


  and
  g535
  (
    n674,
    n135,
    n421,
    n412,
    n379
  );


  xor
  g536
  (
    n588,
    n296,
    n343,
    n366,
    n270
  );


  xnor
  g537
  (
    n527,
    n383,
    n442,
    n210,
    n347
  );


  nor
  g538
  (
    n575,
    n314,
    n340,
    n370,
    n392
  );


  xnor
  g539
  (
    n504,
    n324,
    n389,
    n443,
    n339
  );


  xnor
  g540
  (
    n662,
    n302,
    n162,
    n289,
    n421
  );


  nor
  g541
  (
    n564,
    n393,
    n395,
    n381,
    n389
  );


  and
  g542
  (
    n653,
    n249,
    n222,
    n229,
    n272
  );


  and
  g543
  (
    n525,
    n326,
    n243,
    n337,
    n368
  );


  and
  g544
  (
    n611,
    n428,
    n356,
    n349,
    n233
  );


  xnor
  g545
  (
    n613,
    n444,
    n328,
    n207,
    n301
  );


  nand
  g546
  (
    n669,
    n428,
    n328,
    n402,
    n255
  );


  nor
  g547
  (
    n524,
    n307,
    n306,
    n123,
    n168
  );


  nor
  g548
  (
    n626,
    n413,
    n440,
    n367,
    n283
  );


  xor
  g549
  (
    n675,
    n435,
    n322,
    n374,
    n302
  );


  nand
  g550
  (
    n547,
    n388,
    n389,
    n440,
    n428
  );


  xor
  g551
  (
    n659,
    n402,
    n242,
    n427,
    n366
  );


  xnor
  g552
  (
    n565,
    n340,
    n415,
    n326,
    n311
  );


  xnor
  g553
  (
    n681,
    n380,
    n289,
    n337,
    n327
  );


  or
  g554
  (
    n641,
    n214,
    n323,
    n348,
    n293
  );


  nor
  g555
  (
    n585,
    n396,
    n270,
    n359,
    n330
  );


  xor
  g556
  (
    n663,
    n430,
    n411,
    n429,
    n351
  );


  xor
  g557
  (
    n545,
    n333,
    n320,
    n442,
    n291
  );


  xor
  g558
  (
    n607,
    n352,
    n424,
    n292,
    n319
  );


  nand
  g559
  (
    n531,
    n312,
    n396,
    n390,
    n374
  );


  xnor
  g560
  (
    n595,
    n404,
    n329,
    n439,
    n167
  );


  xnor
  g561
  (
    n686,
    n364,
    n300,
    n388,
    n414
  );


  nand
  g562
  (
    KeyWire_0_31,
    n299,
    n445,
    n169,
    n409
  );


  nor
  g563
  (
    n634,
    n384,
    n250,
    n183,
    n361
  );


  xor
  g564
  (
    n500,
    n260,
    n227,
    n328,
    n208
  );


  xnor
  g565
  (
    n698,
    n337,
    n361,
    n132,
    n419
  );


  and
  g566
  (
    n560,
    n354,
    n285,
    n289,
    n423
  );


  xnor
  g567
  (
    n706,
    n122,
    n283,
    n346,
    n300
  );


  nor
  g568
  (
    n561,
    n304,
    n338,
    n250,
    n195
  );


  and
  g569
  (
    n567,
    n420,
    n425,
    n307,
    n380
  );


  and
  g570
  (
    n552,
    n437,
    n251,
    n233,
    n305
  );


  nand
  g571
  (
    n705,
    n321,
    n412,
    n402,
    n365
  );


  or
  g572
  (
    n665,
    n201,
    n433,
    n368,
    n181
  );


  or
  g573
  (
    n656,
    n387,
    n432,
    n252,
    n312
  );


  nor
  g574
  (
    n538,
    n338,
    n241,
    n370,
    n284
  );


  xor
  g575
  (
    n621,
    n367,
    n247,
    n117,
    n295
  );


  nand
  g576
  (
    n497,
    n156,
    n279,
    n447,
    n370
  );


  nand
  g577
  (
    n630,
    n393,
    n446,
    n348,
    n118
  );


  xor
  g578
  (
    n603,
    n446,
    n345,
    n292,
    n191
  );


  nand
  g579
  (
    n687,
    n116,
    n322,
    n400,
    n444
  );


  and
  g580
  (
    n534,
    n387,
    n431,
    n354,
    n443
  );


  nand
  g581
  (
    n484,
    n275,
    n414,
    n383,
    n447
  );


  xnor
  g582
  (
    n492,
    n363,
    n342,
    n280,
    n244
  );


  or
  g583
  (
    n579,
    n308,
    n413,
    n320,
    n303
  );


  xor
  g584
  (
    n666,
    n407,
    n422,
    n434,
    n185
  );


  and
  g585
  (
    n677,
    n421,
    n398,
    n432,
    n265
  );


  xnor
  g586
  (
    n596,
    n289,
    n375,
    n282,
    n202
  );


  and
  g587
  (
    KeyWire_0_21,
    n266,
    n417,
    n138,
    n431
  );


  nor
  g588
  (
    n619,
    n186,
    n415,
    n273,
    n305
  );


  nor
  g589
  (
    n683,
    n297,
    n164,
    n278,
    n369
  );


  or
  g590
  (
    n532,
    n311,
    n272,
    n120,
    n315
  );


  xnor
  g591
  (
    n590,
    n246,
    n129,
    n330,
    n268
  );


  nor
  g592
  (
    n548,
    n340,
    n299,
    n403,
    n311
  );


  nor
  g593
  (
    n506,
    n405,
    n280,
    n297,
    n373
  );


  and
  g594
  (
    n638,
    n368,
    n371,
    n344,
    n352
  );


  xor
  g595
  (
    n586,
    n228,
    n359,
    n360,
    n351
  );


  nand
  g596
  (
    n680,
    n410,
    n418,
    n340,
    n444
  );


  nand
  g597
  (
    KeyWire_0_5,
    n390,
    n368,
    n365,
    n393
  );


  nand
  g598
  (
    n668,
    n323,
    n408,
    n246,
    n425
  );


  and
  g599
  (
    n505,
    n286,
    n355,
    n299,
    n205
  );


  or
  g600
  (
    n544,
    n358,
    n439,
    n318,
    n175
  );


  xnor
  g601
  (
    n516,
    n394,
    n336,
    n149,
    n288
  );


  and
  g602
  (
    n673,
    n282,
    n317,
    n434,
    n236
  );


  and
  g603
  (
    n592,
    n273,
    n290,
    n379,
    n429
  );


  xor
  g604
  (
    n707,
    n137,
    n441,
    n329,
    n360
  );


  xor
  g605
  (
    n530,
    n281,
    n172,
    n410,
    n357
  );


  nand
  g606
  (
    n559,
    n418,
    n257,
    n317,
    n350
  );


  and
  g607
  (
    n509,
    n373,
    n325,
    n282,
    n280
  );


  and
  g608
  (
    n696,
    n285,
    n304,
    n209,
    n283
  );


  nand
  g609
  (
    n642,
    n285,
    n356,
    n423,
    n157
  );


  or
  g610
  (
    n690,
    n226,
    n319,
    n298,
    n312
  );


  xor
  g611
  (
    n577,
    n290,
    n173,
    n366,
    n369
  );


  xor
  g612
  (
    n528,
    n243,
    n399,
    n384,
    n244
  );


  and
  g613
  (
    n486,
    n354,
    n399,
    n406,
    n408
  );


  or
  g614
  (
    n594,
    n398,
    n441,
    n402,
    n397
  );


  nor
  g615
  (
    n496,
    n339,
    n336,
    n367,
    n416
  );


  and
  g616
  (
    n633,
    n229,
    n348,
    n345,
    n240
  );


  nor
  g617
  (
    n488,
    n400,
    n356,
    n140,
    n411
  );


  xnor
  g618
  (
    n709,
    n392,
    n433,
    n437,
    n141
  );


  and
  g619
  (
    n554,
    n342,
    n394,
    n261,
    n335
  );


  xnor
  g620
  (
    n514,
    n216,
    n297,
    n317,
    n133
  );


  or
  g621
  (
    n667,
    n383,
    n318,
    n218,
    n329
  );


  nand
  g622
  (
    n623,
    n284,
    n387,
    n362,
    n406
  );


  nand
  g623
  (
    n637,
    n342,
    n237,
    n382,
    n302
  );


  or
  g624
  (
    n518,
    n361,
    n391,
    n235,
    n275
  );


  and
  g625
  (
    n555,
    n351,
    n313,
    n365,
    n440
  );


  nand
  g626
  (
    n678,
    n384,
    n328,
    n274,
    n419
  );


  xor
  g627
  (
    n708,
    n298,
    n350,
    n234,
    n413
  );


  and
  g628
  (
    n654,
    n136,
    n350,
    n300,
    n398
  );


  xnor
  g629
  (
    n522,
    n196,
    n291,
    n253,
    n323
  );


  and
  g630
  (
    n490,
    n318,
    n373,
    n413,
    n125
  );


  nand
  g631
  (
    n693,
    n303,
    n295,
    n237,
    n308
  );


  xnor
  g632
  (
    n632,
    n264,
    n163,
    n369,
    n260
  );


  xor
  g633
  (
    n491,
    n158,
    n366,
    n330,
    n436
  );


  nor
  g634
  (
    n664,
    n407,
    n423,
    n401,
    n428
  );


  xor
  g635
  (
    n589,
    n286,
    n439,
    n419,
    n231
  );


  xnor
  g636
  (
    n640,
    n436,
    n407,
    n257,
    n326
  );


  xnor
  g637
  (
    n600,
    n224,
    n200,
    n349,
    n397
  );


  and
  g638
  (
    n521,
    n298,
    n391,
    n429,
    n288
  );


  xor
  g639
  (
    KeyWire_0_7,
    n220,
    n288,
    n338,
    n316
  );


  nand
  g640
  (
    n606,
    n395,
    n426,
    n182,
    n343
  );


  and
  g641
  (
    n685,
    n190,
    n389,
    n392,
    n414
  );


  xor
  g642
  (
    n604,
    n334,
    n287,
    n159,
    n353
  );


  nand
  g643
  (
    n570,
    n310,
    n290,
    n422,
    n152
  );


  nand
  g644
  (
    n691,
    n360,
    n147,
    n278,
    n401
  );


  or
  g645
  (
    KeyWire_0_6,
    n438,
    n303,
    n390,
    n341
  );


  nand
  g646
  (
    n703,
    n265,
    n331,
    n426,
    n315
  );


  nand
  g647
  (
    n563,
    n278,
    n396,
    n410,
    n321
  );


  and
  g648
  (
    n539,
    n324,
    n226,
    n287,
    n430
  );


  xor
  g649
  (
    n617,
    n352,
    n170,
    n435,
    n420
  );


  nand
  g650
  (
    n704,
    n442,
    n279,
    n437,
    n362
  );


  nand
  g651
  (
    n485,
    n256,
    n333,
    n404,
    n262
  );


  xor
  g652
  (
    n614,
    n373,
    n440,
    n240,
    n146
  );


  xor
  g653
  (
    n636,
    n230,
    n358,
    n362,
    n380
  );


  and
  g654
  (
    n635,
    n372,
    n296,
    n294,
    n447
  );


  xnor
  g655
  (
    n487,
    n319,
    n143,
    n336,
    n364
  );


  xnor
  g656
  (
    n692,
    n256,
    n369,
    n446,
    n398
  );


  xnor
  g657
  (
    n550,
    n335,
    n346,
    n433,
    n423
  );


  xor
  g658
  (
    n700,
    n154,
    n430,
    n306,
    n296
  );


  nor
  g659
  (
    n639,
    n302,
    n372,
    n301,
    n275
  );


  nand
  g660
  (
    n568,
    n301,
    n241,
    n393,
    n266
  );


  and
  g661
  (
    n646,
    n432,
    n399,
    n377,
    n298
  );


  nand
  g662
  (
    n571,
    n264,
    n189,
    n410,
    n347
  );


  or
  g663
  (
    n661,
    n267,
    n359,
    n427,
    n280
  );


  xnor
  g664
  (
    n608,
    n279,
    n415,
    n378,
    n394
  );


  or
  g665
  (
    n557,
    n385,
    n294,
    n295,
    n409
  );


  or
  g666
  (
    n602,
    n295,
    n284,
    n401,
    n438
  );


  and
  g667
  (
    n597,
    n324,
    n333,
    n377,
    n271
  );


  and
  g668
  (
    n502,
    n425,
    n263,
    n234,
    n375
  );


  or
  g669
  (
    n620,
    n187,
    n128,
    n341,
    n444
  );


  nand
  g670
  (
    n541,
    n418,
    n388,
    n399,
    n323
  );


  and
  g671
  (
    n645,
    n417,
    n276,
    n155,
    n263
  );


  xor
  g672
  (
    n689,
    n204,
    n377,
    n160,
    n406
  );


  nor
  g673
  (
    n651,
    n321,
    n193,
    n405,
    n358
  );


  nor
  g674
  (
    n605,
    n316,
    n273,
    n431,
    n290
  );


  or
  g675
  (
    n499,
    n308,
    n231,
    n294,
    n299
  );


  nand
  g676
  (
    n625,
    n327,
    n215,
    n224,
    n355
  );


  nor
  g677
  (
    n629,
    n232,
    n382,
    n311,
    n374
  );


  xor
  g678
  (
    n529,
    n272,
    n304,
    n339,
    n411
  );


  or
  g679
  (
    n660,
    n353,
    n419,
    n314,
    n438
  );


  or
  g680
  (
    n583,
    n178,
    n371,
    n174,
    n249
  );


  nor
  g681
  (
    n628,
    n171,
    n268,
    n309,
    n235
  );


  and
  g682
  (
    n670,
    n184,
    n324,
    n385,
    n357
  );


  xnor
  g683
  (
    n688,
    n443,
    n405,
    n376,
    n230
  );


  xor
  g684
  (
    n679,
    n426,
    n320,
    n416,
    n376
  );


  or
  g685
  (
    n551,
    n354,
    n382,
    n314,
    n291
  );


  or
  g686
  (
    n631,
    n335,
    n305,
    n344,
    n276
  );


  not
  g687
  (
    n736,
    n513
  );


  not
  g688
  (
    n728,
    n507
  );


  not
  g689
  (
    n713,
    n497
  );


  buf
  g690
  (
    n723,
    n506
  );


  not
  g691
  (
    n739,
    n509
  );


  buf
  g692
  (
    n711,
    n511
  );


  not
  g693
  (
    n741,
    n515
  );


  not
  g694
  (
    n735,
    n505
  );


  not
  g695
  (
    n715,
    n503
  );


  buf
  g696
  (
    n731,
    n489
  );


  buf
  g697
  (
    n714,
    n514
  );


  not
  g698
  (
    n726,
    n508
  );


  not
  g699
  (
    n733,
    n491
  );


  buf
  g700
  (
    n730,
    n502
  );


  not
  g701
  (
    n721,
    n500
  );


  not
  g702
  (
    n719,
    n490
  );


  not
  g703
  (
    n724,
    n486
  );


  not
  g704
  (
    n729,
    n492
  );


  buf
  g705
  (
    n738,
    n487
  );


  buf
  g706
  (
    n712,
    n493
  );


  buf
  g707
  (
    n727,
    n501
  );


  not
  g708
  (
    n722,
    n512
  );


  buf
  g709
  (
    n717,
    n485
  );


  not
  g710
  (
    n737,
    n498
  );


  not
  g711
  (
    n716,
    n510
  );


  buf
  g712
  (
    n725,
    n494
  );


  not
  g713
  (
    n740,
    n499
  );


  not
  g714
  (
    n720,
    n484
  );


  not
  g715
  (
    n742,
    n496
  );


  not
  g716
  (
    n734,
    n488
  );


  not
  g717
  (
    n718,
    n495
  );


  not
  g718
  (
    n732,
    n504
  );


  buf
  g719
  (
    n757,
    n719
  );


  not
  g720
  (
    n762,
    n729
  );


  buf
  g721
  (
    n754,
    n713
  );


  buf
  g722
  (
    n761,
    n723
  );


  buf
  g723
  (
    n746,
    n727
  );


  buf
  g724
  (
    n750,
    n725
  );


  buf
  g725
  (
    n744,
    n730
  );


  not
  g726
  (
    n752,
    n721
  );


  buf
  g727
  (
    n743,
    n715
  );


  buf
  g728
  (
    n751,
    n717
  );


  not
  g729
  (
    n745,
    n728
  );


  not
  g730
  (
    n755,
    n716
  );


  not
  g731
  (
    n756,
    n718
  );


  not
  g732
  (
    n749,
    n722
  );


  not
  g733
  (
    n747,
    n720
  );


  not
  g734
  (
    KeyWire_0_3,
    n711
  );


  not
  g735
  (
    n759,
    n714
  );


  not
  g736
  (
    n758,
    n726
  );


  not
  g737
  (
    n753,
    n724
  );


  not
  g738
  (
    n760,
    n712
  );


  not
  g739
  (
    n801,
    n744
  );


  buf
  g740
  (
    n818,
    n538
  );


  not
  g741
  (
    KeyWire_0_8,
    n745
  );


  not
  g742
  (
    n808,
    n520
  );


  not
  g743
  (
    n814,
    n734
  );


  buf
  g744
  (
    n821,
    n756
  );


  not
  g745
  (
    n816,
    n541
  );


  buf
  g746
  (
    n786,
    n751
  );


  buf
  g747
  (
    n823,
    n548
  );


  not
  g748
  (
    n765,
    n753
  );


  not
  g749
  (
    n773,
    n745
  );


  not
  g750
  (
    n794,
    n751
  );


  not
  g751
  (
    n793,
    n750
  );


  not
  g752
  (
    n770,
    n751
  );


  buf
  g753
  (
    n817,
    n741
  );


  buf
  g754
  (
    n798,
    n543
  );


  not
  g755
  (
    n781,
    n753
  );


  not
  g756
  (
    n788,
    n741
  );


  buf
  g757
  (
    n800,
    n552
  );


  buf
  g758
  (
    n766,
    n524
  );


  not
  g759
  (
    n779,
    n523
  );


  not
  g760
  (
    n802,
    n750
  );


  not
  g761
  (
    n796,
    n742
  );


  not
  g762
  (
    n790,
    n521
  );


  buf
  g763
  (
    n769,
    n749
  );


  buf
  g764
  (
    n775,
    n747
  );


  not
  g765
  (
    n764,
    n528
  );


  not
  g766
  (
    n797,
    n540
  );


  not
  g767
  (
    n812,
    n756
  );


  not
  g768
  (
    n782,
    n745
  );


  buf
  g769
  (
    n776,
    n747
  );


  buf
  g770
  (
    n763,
    n752
  );


  not
  g771
  (
    n771,
    n743
  );


  buf
  g772
  (
    n807,
    n549
  );


  not
  g773
  (
    n813,
    n547
  );


  not
  g774
  (
    n787,
    n741
  );


  buf
  g775
  (
    n806,
    n533
  );


  not
  g776
  (
    n811,
    n530
  );


  buf
  g777
  (
    n809,
    n738
  );


  not
  g778
  (
    n767,
    n518
  );


  buf
  g779
  (
    n819,
    n516
  );


  not
  g780
  (
    n804,
    n527
  );


  and
  g781
  (
    n792,
    n746,
    n551,
    n757,
    n748
  );


  nor
  g782
  (
    n778,
    n739,
    n744,
    n748,
    n732
  );


  xor
  g783
  (
    n805,
    n537,
    n755,
    n546,
    n522
  );


  nand
  g784
  (
    n820,
    n536,
    n753,
    n757,
    n745
  );


  or
  g785
  (
    n789,
    n755,
    n735,
    n535,
    n743
  );


  nand
  g786
  (
    n783,
    n754,
    n733,
    n532,
    n517
  );


  and
  g787
  (
    n815,
    n751,
    n756,
    n746,
    n748
  );


  and
  g788
  (
    n822,
    n748,
    n553,
    n747,
    n529
  );


  xor
  g789
  (
    n774,
    n550,
    n757,
    n746,
    n754
  );


  xnor
  g790
  (
    KeyWire_0_1,
    n555,
    n525,
    n526,
    n531
  );


  xor
  g791
  (
    n780,
    n746,
    n752,
    n754,
    n554
  );


  nand
  g792
  (
    n777,
    n740,
    n545,
    n534,
    n736
  );


  or
  g793
  (
    n784,
    n756,
    n755,
    n753,
    n750
  );


  xnor
  g794
  (
    n785,
    n749,
    n749,
    n737,
    n731
  );


  nand
  g795
  (
    n795,
    n752,
    n758,
    n744,
    n743
  );


  nor
  g796
  (
    n791,
    n757,
    n519,
    n743,
    n539
  );


  nor
  g797
  (
    n803,
    n747,
    n742,
    n752,
    n542
  );


  xor
  g798
  (
    n799,
    n741,
    n744,
    n740,
    n754
  );


  xnor
  g799
  (
    n772,
    n749,
    n750,
    n544,
    n755
  );


  buf
  g800
  (
    n867,
    n570
  );


  buf
  g801
  (
    n837,
    n458
  );


  not
  g802
  (
    n858,
    n454
  );


  not
  g803
  (
    n856,
    n598
  );


  buf
  g804
  (
    n834,
    n467
  );


  not
  g805
  (
    n859,
    n473
  );


  xor
  g806
  (
    n833,
    n784,
    n592,
    n794,
    n476
  );


  xor
  g807
  (
    n826,
    n450,
    n472,
    n772,
    n580
  );


  nor
  g808
  (
    KeyWire_0_13,
    n785,
    n768,
    n808,
    n562
  );


  nor
  g809
  (
    n882,
    n449,
    n461,
    n472,
    n465
  );


  or
  g810
  (
    n852,
    n579,
    n469,
    n468
  );


  xnor
  g811
  (
    n869,
    n472,
    n587,
    n810,
    n556
  );


  and
  g812
  (
    n831,
    n822,
    n593,
    n468,
    n795
  );


  nand
  g813
  (
    n848,
    n475,
    n460,
    n456
  );


  nand
  g814
  (
    n847,
    n455,
    n458,
    n758,
    n804
  );


  and
  g815
  (
    n832,
    n459,
    n817,
    n816,
    n796
  );


  xnor
  g816
  (
    n830,
    n465,
    n459,
    n470,
    n809
  );


  xnor
  g817
  (
    n884,
    n563,
    n451,
    n813,
    n452
  );


  xor
  g818
  (
    n866,
    n814,
    n823,
    n818,
    n450
  );


  nor
  g819
  (
    n865,
    n449,
    n597,
    n461,
    n805
  );


  nand
  g820
  (
    n861,
    n448,
    n797,
    n771,
    n578
  );


  nor
  g821
  (
    n829,
    n758,
    n455,
    n470,
    n557
  );


  nor
  g822
  (
    n851,
    n450,
    n464,
    n759,
    n448
  );


  nor
  g823
  (
    n843,
    n590,
    n585,
    n467
  );


  xnor
  g824
  (
    n881,
    n476,
    n571,
    n802,
    n798
  );


  xor
  g825
  (
    n879,
    n453,
    n451,
    n474,
    n788
  );


  nor
  g826
  (
    n877,
    n470,
    n591,
    n473,
    n451
  );


  nand
  g827
  (
    n842,
    n589,
    n764,
    n453,
    n807
  );


  nand
  g828
  (
    n876,
    n779,
    n469,
    n477,
    n594
  );


  and
  g829
  (
    n840,
    n786,
    n577,
    n584,
    n462
  );


  xor
  g830
  (
    n878,
    n799,
    n778,
    n475,
    n561
  );


  and
  g831
  (
    n870,
    n811,
    n458,
    n776,
    n473
  );


  or
  g832
  (
    n874,
    n783,
    n758,
    n450,
    n567
  );


  nand
  g833
  (
    n863,
    n449,
    n466,
    n789,
    n456
  );


  nor
  g834
  (
    n827,
    n457,
    n454,
    n467,
    n560
  );


  xor
  g835
  (
    n846,
    n472,
    n466,
    n474,
    n458
  );


  nand
  g836
  (
    n845,
    n806,
    n581,
    n568,
    n462
  );


  or
  g837
  (
    n854,
    n576,
    n582,
    n463,
    n787
  );


  xor
  g838
  (
    n883,
    n466,
    n452,
    n460,
    n453
  );


  nor
  g839
  (
    n862,
    n558,
    n766,
    n469,
    n765
  );


  nor
  g840
  (
    KeyWire_0_0,
    n574,
    n453,
    n575,
    n463
  );


  and
  g841
  (
    n872,
    n572,
    n759,
    n457,
    n821
  );


  xnor
  g842
  (
    n864,
    n460,
    n763,
    n566,
    n803
  );


  and
  g843
  (
    n839,
    n464,
    n596,
    n792,
    n461
  );


  xor
  g844
  (
    n838,
    n464,
    n449,
    n473,
    n476
  );


  or
  g845
  (
    n849,
    n815,
    n455,
    n793
  );


  xnor
  g846
  (
    n825,
    n586,
    n463,
    n475,
    n460
  );


  xor
  g847
  (
    n841,
    n583,
    n565,
    n465,
    n595
  );


  nor
  g848
  (
    n873,
    n559,
    n448,
    n474,
    n465
  );


  and
  g849
  (
    n828,
    n790,
    n461,
    n454,
    n777
  );


  nand
  g850
  (
    n836,
    n463,
    n471,
    n800,
    n464
  );


  or
  g851
  (
    n835,
    n781,
    n474,
    n471,
    n564
  );


  nor
  g852
  (
    n880,
    n770,
    n791,
    n780,
    n469
  );


  xor
  g853
  (
    n853,
    n773,
    n451,
    n782,
    n452
  );


  xnor
  g854
  (
    n857,
    n819,
    n459,
    n573,
    n569
  );


  or
  g855
  (
    n871,
    n470,
    n774,
    n466,
    n459
  );


  xnor
  g856
  (
    n850,
    n769,
    n476,
    n452,
    n448
  );


  nor
  g857
  (
    KeyWire_0_20,
    n471,
    n457,
    n767,
    n462
  );


  or
  g858
  (
    n855,
    n462,
    n801,
    n454,
    n468
  );


  nand
  g859
  (
    n824,
    n471,
    n588,
    n820,
    n475
  );


  xor
  g860
  (
    n844,
    n457,
    n775,
    n456,
    n812
  );


  buf
  g861
  (
    n953,
    n610
  );


  buf
  g862
  (
    n888,
    n826
  );


  buf
  g863
  (
    n915,
    n857
  );


  buf
  g864
  (
    n949,
    n617
  );


  not
  g865
  (
    n933,
    n833
  );


  not
  g866
  (
    n889,
    n634
  );


  not
  g867
  (
    n922,
    n846
  );


  buf
  g868
  (
    n967,
    n841
  );


  buf
  g869
  (
    n886,
    n843
  );


  buf
  g870
  (
    n904,
    n850
  );


  not
  g871
  (
    n961,
    n846
  );


  buf
  g872
  (
    n979,
    n826
  );


  buf
  g873
  (
    n891,
    n833
  );


  not
  g874
  (
    n958,
    n853
  );


  buf
  g875
  (
    n962,
    n843
  );


  not
  g876
  (
    n893,
    n841
  );


  buf
  g877
  (
    n902,
    n854
  );


  buf
  g878
  (
    n931,
    n845
  );


  not
  g879
  (
    n927,
    n850
  );


  buf
  g880
  (
    n963,
    n847
  );


  not
  g881
  (
    n978,
    n852
  );


  not
  g882
  (
    n945,
    n834
  );


  buf
  g883
  (
    n950,
    n621
  );


  not
  g884
  (
    n926,
    n840
  );


  not
  g885
  (
    n914,
    n825
  );


  buf
  g886
  (
    n955,
    n632
  );


  buf
  g887
  (
    n912,
    n633
  );


  not
  g888
  (
    n906,
    n825
  );


  buf
  g889
  (
    KeyWire_0_18,
    n853
  );


  not
  g890
  (
    n939,
    n625
  );


  not
  g891
  (
    n923,
    n840
  );


  buf
  g892
  (
    n897,
    n840
  );


  not
  g893
  (
    n918,
    n836
  );


  buf
  g894
  (
    n930,
    n842
  );


  buf
  g895
  (
    n917,
    n606
  );


  not
  g896
  (
    n894,
    n603
  );


  not
  g897
  (
    n916,
    n840
  );


  buf
  g898
  (
    n934,
    n852
  );


  not
  g899
  (
    n970,
    n854
  );


  buf
  g900
  (
    n890,
    n851
  );


  not
  g901
  (
    n959,
    n824
  );


  buf
  g902
  (
    n980,
    n837
  );


  buf
  g903
  (
    n972,
    n847
  );


  not
  g904
  (
    n948,
    n612
  );


  not
  g905
  (
    n907,
    n844
  );


  buf
  g906
  (
    n947,
    n827
  );


  buf
  g907
  (
    n909,
    n848
  );


  not
  g908
  (
    n957,
    n827
  );


  not
  g909
  (
    n941,
    n834
  );


  not
  g910
  (
    n946,
    n627
  );


  not
  g911
  (
    n975,
    n849
  );


  not
  g912
  (
    n966,
    n611
  );


  not
  g913
  (
    n954,
    n858
  );


  not
  g914
  (
    n938,
    n835
  );


  not
  g915
  (
    n977,
    n830
  );


  not
  g916
  (
    n956,
    n845
  );


  not
  g917
  (
    n895,
    n623
  );


  buf
  g918
  (
    n885,
    n624
  );


  not
  g919
  (
    n965,
    n851
  );


  buf
  g920
  (
    n896,
    n619
  );


  not
  g921
  (
    n900,
    n839
  );


  not
  g922
  (
    n937,
    n857
  );


  not
  g923
  (
    n942,
    n834
  );


  buf
  g924
  (
    n932,
    n852
  );


  not
  g925
  (
    n944,
    n853
  );


  buf
  g926
  (
    n976,
    n841
  );


  buf
  g927
  (
    n943,
    n855
  );


  buf
  g928
  (
    n969,
    n836
  );


  buf
  g929
  (
    n921,
    n850
  );


  buf
  g930
  (
    n973,
    n608
  );


  xor
  g931
  (
    KeyWire_0_24,
    n832,
    n838,
    n849,
    n847
  );


  and
  g932
  (
    n892,
    n626,
    n829,
    n844,
    n848
  );


  and
  g933
  (
    n903,
    n839,
    n828,
    n629,
    n615
  );


  nand
  g934
  (
    n920,
    n857,
    n829,
    n601,
    n841
  );


  nor
  g935
  (
    n928,
    n829,
    n829,
    n852,
    n855
  );


  xor
  g936
  (
    n929,
    n837,
    n602,
    n635,
    n827
  );


  or
  g937
  (
    n887,
    n836,
    n848,
    n824,
    n856
  );


  xor
  g938
  (
    n968,
    n834,
    n599,
    n849,
    n836
  );


  or
  g939
  (
    n924,
    n830,
    n848,
    n628,
    n838
  );


  or
  g940
  (
    n901,
    n837,
    n844,
    n846,
    n616
  );


  xor
  g941
  (
    n936,
    n849,
    n855,
    n842,
    n828
  );


  nor
  g942
  (
    n899,
    n622,
    n607,
    n831,
    n609
  );


  and
  g943
  (
    n911,
    n828,
    n832,
    n855,
    n833
  );


  xnor
  g944
  (
    n964,
    n856,
    n839,
    n832,
    n631
  );


  xnor
  g945
  (
    KeyWire_0_12,
    n828,
    n856,
    n843,
    n857
  );


  nor
  g946
  (
    n925,
    n853,
    n825,
    n835,
    n854
  );


  xnor
  g947
  (
    n960,
    n605,
    n838,
    n845,
    n614
  );


  and
  g948
  (
    n974,
    n826,
    n838,
    n851,
    n831
  );


  or
  g949
  (
    n898,
    n839,
    n604,
    n835,
    n850
  );


  xnor
  g950
  (
    n940,
    n600,
    n824,
    n831,
    n613
  );


  and
  g951
  (
    n905,
    n844,
    n842,
    n830,
    n833
  );


  xor
  g952
  (
    n971,
    n826,
    n847,
    n835,
    n832
  );


  and
  g953
  (
    n919,
    n618,
    n842,
    n825,
    n831
  );


  or
  g954
  (
    n913,
    n854,
    n851,
    n824,
    n830
  );


  and
  g955
  (
    n910,
    n846,
    n843,
    n837,
    n827
  );


  xor
  g956
  (
    n908,
    n630,
    n856,
    n845,
    n620
  );


  xnor
  g957
  (
    n1012,
    n872,
    n865,
    n860,
    n893
  );


  xor
  g958
  (
    n1008,
    n933,
    n944,
    n874,
    n909
  );


  nand
  g959
  (
    n997,
    n919,
    n927,
    n876,
    n898
  );


  nand
  g960
  (
    n1003,
    n899,
    n877,
    n872,
    n878
  );


  xor
  g961
  (
    n1013,
    n861,
    n859,
    n945,
    n873
  );


  nor
  g962
  (
    n986,
    n875,
    n866,
    n938
  );


  xor
  g963
  (
    n1015,
    n871,
    n895,
    n929,
    n940
  );


  xor
  g964
  (
    n1009,
    n879,
    n874,
    n942,
    n941
  );


  xnor
  g965
  (
    n990,
    n905,
    n863,
    n930,
    n888
  );


  nand
  g966
  (
    n982,
    n932,
    n870,
    n879,
    n892
  );


  and
  g967
  (
    n995,
    n865,
    n858,
    n866,
    n876
  );


  nor
  g968
  (
    n1016,
    n939,
    n860,
    n934,
    n859
  );


  or
  g969
  (
    n981,
    n868,
    n870,
    n931,
    n860
  );


  nand
  g970
  (
    n1004,
    n928,
    n862,
    n911,
    n858
  );


  xor
  g971
  (
    n1011,
    n907,
    n863,
    n947,
    n918
  );


  xor
  g972
  (
    n993,
    n878,
    n877,
    n923,
    n912
  );


  xnor
  g973
  (
    n984,
    n894,
    n878,
    n868,
    n900
  );


  nand
  g974
  (
    n999,
    n914,
    n946,
    n876,
    n864
  );


  and
  g975
  (
    n1002,
    n902,
    n861,
    n863,
    n876
  );


  and
  g976
  (
    n988,
    n875,
    n878,
    n877,
    n915
  );


  nor
  g977
  (
    n1006,
    n867,
    n859,
    n887,
    n910
  );


  nor
  g978
  (
    n983,
    n874,
    n862,
    n864,
    n872
  );


  xnor
  g979
  (
    n998,
    n903,
    n867,
    n859
  );


  nor
  g980
  (
    n991,
    n871,
    n864,
    n913,
    n890
  );


  or
  g981
  (
    n992,
    n937,
    n858,
    n901,
    n868
  );


  nor
  g982
  (
    n985,
    n922,
    n866,
    n874,
    n873
  );


  xor
  g983
  (
    n989,
    n925,
    n935,
    n870,
    n865
  );


  nor
  g984
  (
    n1005,
    n875,
    n896,
    n865,
    n908
  );


  or
  g985
  (
    n1001,
    n861,
    n862,
    n916,
    n870
  );


  nor
  g986
  (
    n1014,
    n871,
    n943,
    n869,
    n936
  );


  or
  g987
  (
    n994,
    n906,
    n863,
    n868,
    n872
  );


  xor
  g988
  (
    KeyWire_0_29,
    n924,
    n904,
    n889,
    n886
  );


  nand
  g989
  (
    n987,
    n862,
    n917,
    n873,
    n867
  );


  nand
  g990
  (
    n996,
    n869,
    n869,
    n877,
    n920
  );


  nor
  g991
  (
    n1017,
    n875,
    n926,
    n873,
    n864
  );


  nor
  g992
  (
    n1010,
    n921,
    n885,
    n869,
    n860
  );


  xor
  g993
  (
    n1007,
    n861,
    n891,
    n897,
    n871
  );


  not
  g994
  (
    n1021,
    n1002
  );


  buf
  g995
  (
    n1018,
    n1003
  );


  buf
  g996
  (
    n1019,
    n1004
  );


  buf
  g997
  (
    n1020,
    n1005
  );


  nor
  g998
  (
    n1030,
    n644,
    n1012,
    n641,
    n646
  );


  and
  g999
  (
    n1022,
    n1018,
    n639,
    n647,
    n1013
  );


  xnor
  g1000
  (
    n1027,
    n645,
    n652,
    n648,
    n1019
  );


  nor
  g1001
  (
    KeyWire_0_26,
    n1007,
    n636,
    n1011,
    n651
  );


  nor
  g1002
  (
    n1031,
    n1020,
    n948,
    n1009,
    n642
  );


  xnor
  g1003
  (
    n1024,
    n1015,
    n649,
    n650,
    n637
  );


  xor
  g1004
  (
    n1023,
    n643,
    n1010,
    n1018,
    n1019
  );


  or
  g1005
  (
    n1026,
    n1018,
    n638,
    n1014,
    n640
  );


  and
  g1006
  (
    n1029,
    n1020,
    n1016,
    n1017,
    n1019
  );


  nand
  g1007
  (
    n1025,
    n1019,
    n1006,
    n1018,
    n1008
  );


  or
  g1008
  (
    n1032,
    n1031,
    n478,
    n1030
  );


  xnor
  g1009
  (
    n1033,
    n478,
    n477
  );


  buf
  g1010
  (
    n1039,
    n1033
  );


  buf
  g1011
  (
    n1034,
    n1033
  );


  not
  g1012
  (
    n1037,
    n1033
  );


  buf
  g1013
  (
    n1040,
    n1032
  );


  buf
  g1014
  (
    n1036,
    n1032
  );


  buf
  g1015
  (
    n1038,
    n1032
  );


  not
  g1016
  (
    n1035,
    n1032
  );


  xor
  g1017
  (
    n1041,
    n951,
    n653
  );


  xor
  g1018
  (
    n1047,
    n953,
    n655,
    n956
  );


  nor
  g1019
  (
    n1043,
    n742,
    n1037,
    n1036
  );


  nand
  g1020
  (
    n1048,
    n1038,
    n656,
    n1040
  );


  xnor
  g1021
  (
    n1042,
    n654,
    n949,
    n1039
  );


  nor
  g1022
  (
    n1046,
    n1035,
    n957,
    n1033
  );


  or
  g1023
  (
    n1049,
    n1034,
    n954,
    n958
  );


  nand
  g1024
  (
    n1045,
    n1039,
    n952,
    n1038
  );


  xor
  g1025
  (
    n1044,
    n478,
    n950,
    n955
  );


  not
  g1026
  (
    n1055,
    n479
  );


  xnor
  g1027
  (
    n1054,
    n1049,
    n961,
    n959
  );


  nand
  g1028
  (
    n1058,
    n962,
    n1049,
    n1044
  );


  or
  g1029
  (
    n1056,
    n479,
    n657,
    n1040
  );


  or
  g1030
  (
    n1052,
    n1047,
    n1040
  );


  and
  g1031
  (
    n1050,
    n1045,
    n963,
    n879
  );


  xor
  g1032
  (
    n1053,
    n965,
    n880,
    n964
  );


  xnor
  g1033
  (
    n1059,
    n1042,
    n1041,
    n1046
  );


  xnor
  g1034
  (
    n1051,
    n1048,
    n960,
    n879
  );


  nor
  g1035
  (
    n1057,
    n966,
    n479,
    n1043
  );


  not
  g1036
  (
    n1064,
    n1050
  );


  buf
  g1037
  (
    n1063,
    n1052
  );


  not
  g1038
  (
    n1061,
    n1053
  );


  buf
  g1039
  (
    n1062,
    n968
  );


  buf
  g1040
  (
    n1067,
    n1051
  );


  not
  g1041
  (
    n1066,
    n967
  );


  not
  g1042
  (
    n1060,
    n1050
  );


  and
  g1043
  (
    n1065,
    n1051,
    n1053,
    n1052
  );


  not
  g1044
  (
    n1082,
    n1056
  );


  buf
  g1045
  (
    n1076,
    n658
  );


  not
  g1046
  (
    n1084,
    n1055
  );


  not
  g1047
  (
    n1080,
    n1057
  );


  buf
  g1048
  (
    n1078,
    n481
  );


  not
  g1049
  (
    n1081,
    n659
  );


  not
  g1050
  (
    n1072,
    n1061
  );


  and
  g1051
  (
    n1069,
    n1064,
    n1063,
    n1062,
    n1061
  );


  nand
  g1052
  (
    n1083,
    n1063,
    n480,
    n1060,
    n665
  );


  and
  g1053
  (
    n1074,
    n1063,
    n668,
    n667,
    n1056
  );


  or
  g1054
  (
    n1070,
    n1062,
    n1062,
    n662,
    n661
  );


  nand
  g1055
  (
    n1079,
    n1062,
    n480,
    n1057,
    n1054
  );


  nand
  g1056
  (
    n1073,
    n1059,
    n479,
    n480,
    n1060
  );


  nand
  g1057
  (
    n1068,
    n660,
    n1064,
    n1054,
    n1058
  );


  xnor
  g1058
  (
    n1075,
    n663,
    n1059,
    n1063,
    n1061
  );


  nand
  g1059
  (
    n1071,
    n666,
    n1058,
    n664,
    n1061
  );


  xor
  g1060
  (
    n1077,
    n481,
    n1060,
    n1055,
    n480
  );


  not
  g1061
  (
    n1091,
    n1064
  );


  not
  g1062
  (
    n1096,
    n1072
  );


  buf
  g1063
  (
    n1093,
    n481
  );


  not
  g1064
  (
    n1095,
    n1070
  );


  not
  g1065
  (
    n1085,
    n669
  );


  not
  g1066
  (
    n1100,
    n1080
  );


  buf
  g1067
  (
    n1097,
    n1067
  );


  not
  g1068
  (
    n1092,
    n1066
  );


  and
  g1069
  (
    n1087,
    n1075,
    n1065
  );


  nor
  g1070
  (
    n1086,
    n1067,
    n1084,
    n1065
  );


  nand
  g1071
  (
    KeyWire_0_23,
    n1069,
    n1082,
    n670
  );


  nand
  g1072
  (
    n1094,
    n1068,
    n1065,
    n1071
  );


  nor
  g1073
  (
    n1089,
    n1079,
    n1066,
    n1078
  );


  or
  g1074
  (
    n1099,
    n1066,
    n1073,
    n1074
  );


  xor
  g1075
  (
    n1098,
    n671,
    n1064,
    n1076
  );


  or
  g1076
  (
    n1090,
    n1067,
    n1066,
    n969
  );


  and
  g1077
  (
    n1101,
    n1077,
    n1083,
    n1067,
    n1081
  );


  not
  g1078
  (
    n1104,
    n1086
  );


  buf
  g1079
  (
    n1105,
    n1088
  );


  buf
  g1080
  (
    n1103,
    n1087
  );


  buf
  g1081
  (
    n1102,
    n1085
  );


  xnor
  g1082
  (
    n1116,
    n683,
    n1102,
    n686,
    n687
  );


  nand
  g1083
  (
    n1118,
    n1095,
    n698,
    n1104,
    n695
  );


  xnor
  g1084
  (
    n1119,
    n709,
    n674,
    n676,
    n1090
  );


  nor
  g1085
  (
    n1112,
    n1094,
    n689,
    n707,
    n1104
  );


  nand
  g1086
  (
    n1117,
    n694,
    n708,
    n1105,
    n1093
  );


  nor
  g1087
  (
    n1107,
    n682,
    n1089,
    n696,
    n1103
  );


  nor
  g1088
  (
    n1115,
    n1105,
    n675,
    n1103,
    n702
  );


  xnor
  g1089
  (
    n1111,
    n692,
    n701,
    n677,
    n679
  );


  or
  g1090
  (
    n1108,
    n680,
    n681,
    n1102,
    n1105
  );


  or
  g1091
  (
    n1106,
    n699,
    n700,
    n688,
    n1105
  );


  nand
  g1092
  (
    n1121,
    n684,
    n1097,
    n691,
    n1091
  );


  xnor
  g1093
  (
    n1120,
    n1104,
    n697,
    n690,
    n1092
  );


  nor
  g1094
  (
    n1109,
    n703,
    n672,
    n693,
    n705
  );


  and
  g1095
  (
    n1113,
    n685,
    n1102,
    n1096,
    n1104
  );


  nor
  g1096
  (
    n1114,
    n1102,
    n704,
    n1098,
    n706
  );


  nand
  g1097
  (
    n1110,
    n673,
    n1103,
    n678
  );


  buf
  g1098
  (
    n1146,
    n1120
  );


  buf
  g1099
  (
    n1132,
    n1113
  );


  buf
  g1100
  (
    n1125,
    n1117
  );


  buf
  g1101
  (
    n1138,
    n1117
  );


  buf
  g1102
  (
    n1124,
    n1120
  );


  buf
  g1103
  (
    n1135,
    n1119
  );


  buf
  g1104
  (
    n1129,
    n1119
  );


  buf
  g1105
  (
    n1144,
    n1116
  );


  not
  g1106
  (
    n1128,
    n1106
  );


  buf
  g1107
  (
    n1139,
    n1118
  );


  not
  g1108
  (
    n1133,
    n1108
  );


  not
  g1109
  (
    KeyWire_0_17,
    n1119
  );


  not
  g1110
  (
    n1131,
    n1117
  );


  buf
  g1111
  (
    n1151,
    n1109
  );


  buf
  g1112
  (
    n1123,
    n1118
  );


  not
  g1113
  (
    n1147,
    n1120
  );


  not
  g1114
  (
    n1141,
    n1118
  );


  buf
  g1115
  (
    n1140,
    n1117
  );


  not
  g1116
  (
    n1136,
    n1121
  );


  not
  g1117
  (
    n1126,
    n1121
  );


  buf
  g1118
  (
    n1145,
    n1118
  );


  buf
  g1119
  (
    n1149,
    n1119
  );


  not
  g1120
  (
    n1134,
    n1114
  );


  buf
  g1121
  (
    n1122,
    n1121
  );


  not
  g1122
  (
    n1137,
    n1111
  );


  not
  g1123
  (
    n1127,
    n1120
  );


  not
  g1124
  (
    n1130,
    n1115
  );


  buf
  g1125
  (
    n1143,
    n1107
  );


  buf
  g1126
  (
    n1148,
    n1112
  );


  buf
  g1127
  (
    n1150,
    n1110
  );


  not
  g1128
  (
    n1152,
    n1122
  );


  not
  g1129
  (
    n1153,
    n1123
  );


  buf
  g1130
  (
    n1156,
    n1153
  );


  xor
  g1131
  (
    n1160,
    n1153,
    n1126,
    n1129
  );


  and
  g1132
  (
    n1154,
    n1152,
    n1133,
    n1128,
    n1134
  );


  nand
  g1133
  (
    n1157,
    n1135,
    n1141,
    n1132,
    n1130
  );


  nor
  g1134
  (
    n1155,
    n1139,
    n1143,
    n1138,
    n1153
  );


  xor
  g1135
  (
    n1158,
    n1152,
    n1131,
    n1136,
    n1127
  );


  nor
  g1136
  (
    n1159,
    n1124,
    n1137,
    n1152
  );


  nor
  g1137
  (
    n1161,
    n1125,
    n1142,
    n1140,
    n1153
  );


  and
  g1138
  (
    n1164,
    n482,
    n482,
    n1155,
    n483
  );


  or
  g1139
  (
    n1163,
    n1154,
    n482,
    n483
  );


  and
  g1140
  (
    n1162,
    n481,
    n1154,
    n483
  );


  and
  g1141
  (
    n1169,
    n1164,
    n1163,
    n1158,
    n1155
  );


  or
  g1142
  (
    n1167,
    n1158,
    n972,
    n1159,
    n1163
  );


  xor
  g1143
  (
    n1166,
    n1156,
    n970,
    n973,
    n1160
  );


  or
  g1144
  (
    n1168,
    n971,
    n1156,
    n1164,
    n1162
  );


  nand
  g1145
  (
    n1165,
    n1159,
    n1157,
    n974
  );


  not
  g1146
  (
    n1173,
    n1166
  );


  not
  g1147
  (
    n1176,
    n1165
  );


  buf
  g1148
  (
    n1172,
    n1166
  );


  not
  g1149
  (
    n1174,
    n1165
  );


  buf
  g1150
  (
    n1170,
    n1165
  );


  not
  g1151
  (
    n1171,
    n1166
  );


  not
  g1152
  (
    n1175,
    n1165
  );


  nand
  g1153
  (
    n1197,
    n1020,
    n1168,
    n1172
  );


  and
  g1154
  (
    n1186,
    n975,
    n977,
    n1176,
    n761
  );


  or
  g1155
  (
    n1183,
    n1172,
    n1161,
    n762,
    n1167
  );


  nor
  g1156
  (
    n1195,
    n1021,
    n1161,
    n1175,
    n1160
  );


  xor
  g1157
  (
    KeyWire_0_25,
    n1170,
    n759,
    n1166,
    n760
  );


  nor
  g1158
  (
    n1187,
    n1173,
    n978,
    n1167
  );


  nor
  g1159
  (
    KeyWire_0_27,
    n1168,
    n882,
    n1171,
    n1173
  );


  and
  g1160
  (
    n1196,
    n761,
    n1021,
    n1175,
    n1169
  );


  nand
  g1161
  (
    n1188,
    n1175,
    n1169,
    n1168,
    n1176
  );


  and
  g1162
  (
    n1191,
    n976,
    n880,
    n760
  );


  and
  g1163
  (
    n1189,
    n1101,
    n1021,
    n762,
    n1100
  );


  xnor
  g1164
  (
    n1182,
    n1172,
    n1174,
    n1169,
    n1170
  );


  xor
  g1165
  (
    n1178,
    n761,
    n759,
    n1170
  );


  and
  g1166
  (
    n1193,
    n881,
    n1099,
    n1171,
    n762
  );


  xor
  g1167
  (
    n1184,
    n1174,
    n1121,
    n881
  );


  xnor
  g1168
  (
    n1185,
    n1176,
    n742,
    n1100,
    n979
  );


  xnor
  g1169
  (
    n1190,
    n1169,
    n762,
    n1172,
    n1171
  );


  or
  g1170
  (
    n1181,
    n1173,
    n881,
    n1171,
    n761
  );


  or
  g1171
  (
    n1194,
    n1176,
    n1101,
    n1173,
    n1021
  );


  or
  g1172
  (
    n1179,
    n880,
    n1174,
    n760,
    n1020
  );


  nor
  g1173
  (
    n1192,
    n1167,
    n880,
    n1174,
    n1175
  );


  buf
  g1174
  (
    n1198,
    n1179
  );


  buf
  g1175
  (
    n1202,
    n1181
  );


  buf
  g1176
  (
    n1201,
    n1180
  );


  buf
  g1177
  (
    n1199,
    n1182
  );


  not
  g1178
  (
    n1200,
    n1183
  );


  nor
  g1179
  (
    n1213,
    n883,
    n980,
    n882,
    n1201
  );


  nand
  g1180
  (
    n1204,
    n1191,
    n882,
    n1199,
    n710
  );


  and
  g1181
  (
    n1203,
    n1201,
    n1190,
    n1146,
    n1150
  );


  xor
  g1182
  (
    n1206,
    n1200,
    n883
  );


  and
  g1183
  (
    n1211,
    n1193,
    n1200,
    n1201,
    n1198
  );


  xnor
  g1184
  (
    n1210,
    n1147,
    n1148,
    n884,
    n1201
  );


  xnor
  g1185
  (
    n1209,
    n1145,
    n1149,
    n1198,
    n882
  );


  xnor
  g1186
  (
    n1205,
    n1199,
    n1198,
    n1188,
    n1189
  );


  xor
  g1187
  (
    n1214,
    n1192,
    n884,
    n1202,
    n1199
  );


  or
  g1188
  (
    n1208,
    n884,
    n1194,
    n1197,
    n1198
  );


  xnor
  g1189
  (
    n1212,
    n1185,
    n884,
    n1199,
    n1184
  );


  nor
  g1190
  (
    n1215,
    n1187,
    n1196,
    n883,
    n1186
  );


  or
  g1191
  (
    n1207,
    n1200,
    n1195,
    n1144,
    n1151
  );


  xnor
  g1192
  (
    n1219,
    n1215,
    n1212,
    n1202
  );


  or
  g1193
  (
    n1217,
    n1210,
    n1208,
    n1207,
    n1214
  );


  xor
  g1194
  (
    n1216,
    n1211,
    n1213,
    n1205,
    n1203
  );


  and
  g1195
  (
    n1218,
    n1204,
    n1202,
    n1206,
    n1209
  );


  xnor
  g1196
  (
    n1220,
    n1219,
    n1218,
    n1217,
    n1216
  );


  xor
  KeyGate_0_0
  (
    n875,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n768,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n231,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n748,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n373,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n694,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n672,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n627,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n810,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n657,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n582,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n205,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n951,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n868,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n562,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n282,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n308,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1142,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n952,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n278,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n860,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n553,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n327,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1088,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n935,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1177,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n1028,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1180,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n320,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1000,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n155,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n520,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

