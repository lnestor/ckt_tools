// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_203 written by SynthGen on 2021/04/05 11:08:35
module Stat_1000_203( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n550, n622, n656, n640, n637, n620, n616, n638,
 n652, n641, n643, n621, n615, n624, n626, n639,
 n631, n979, n1008, n1000, n1006, n1013, n1025, n1016,
 n1022, n1024, n1011, n1021, n1012, n1032, n1031, n1030);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n550, n622, n656, n640, n637, n620, n616, n638,
 n652, n641, n643, n621, n615, n624, n626, n639,
 n631, n979, n1008, n1000, n1006, n1013, n1025, n1016,
 n1022, n1024, n1011, n1021, n1012, n1032, n1031, n1030;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n617, n618, n619,
 n623, n625, n627, n628, n629, n630, n632, n633,
 n634, n635, n636, n642, n644, n645, n646, n647,
 n648, n649, n650, n651, n653, n654, n655, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1001, n1002, n1003,
 n1004, n1005, n1007, n1009, n1010, n1014, n1015, n1017,
 n1018, n1019, n1020, n1023, n1026, n1027, n1028, n1029;

not  g0 (n41, n14);
buf  g1 (n91, n9);
buf  g2 (n40, n15);
not  g3 (n83, n19);
not  g4 (n68, n19);
not  g5 (n62, n16);
not  g6 (n48, n5);
buf  g7 (n102, n11);
buf  g8 (n38, n17);
buf  g9 (n101, n20);
buf  g10 (n100, n16);
buf  g11 (n37, n6);
not  g12 (n35, n12);
buf  g13 (n36, n9);
buf  g14 (n34, n19);
not  g15 (n33, n21);
not  g16 (n65, n20);
not  g17 (n58, n17);
not  g18 (n80, n8);
buf  g19 (n39, n8);
not  g20 (n97, n5);
not  g21 (n77, n8);
buf  g22 (n44, n11);
buf  g23 (n94, n11);
buf  g24 (n50, n21);
buf  g25 (n89, n22);
buf  g26 (n54, n17);
not  g27 (n76, n4);
not  g28 (n43, n7);
buf  g29 (n99, n14);
not  g30 (n66, n7);
not  g31 (n86, n4);
buf  g32 (n84, n10);
buf  g33 (n90, n7);
not  g34 (n63, n5);
not  g35 (n64, n13);
buf  g36 (n42, n17);
buf  g37 (n46, n20);
not  g38 (n98, n16);
not  g39 (n78, n6);
buf  g40 (n69, n2);
buf  g41 (n71, n5);
not  g42 (n74, n16);
not  g43 (n67, n8);
not  g44 (n45, n6);
not  g45 (n49, n15);
not  g46 (n47, n19);
not  g47 (n85, n6);
buf  g48 (n72, n12);
not  g49 (n73, n22);
buf  g50 (n51, n13);
not  g51 (n53, n13);
not  g52 (n95, n18);
not  g53 (n82, n3);
buf  g54 (n81, n20);
not  g55 (n87, n14);
not  g56 (n70, n4);
buf  g57 (n59, n13);
not  g58 (n104, n10);
not  g59 (n56, n14);
buf  g60 (n61, n12);
buf  g61 (n103, n18);
not  g62 (n96, n10);
not  g63 (n57, n15);
not  g64 (n93, n1);
not  g65 (n55, n11);
not  g66 (n79, n21);
buf  g67 (n75, n9);
not  g68 (n88, n15);
buf  g69 (n52, n22);
xnor g70 (n60, n18, n18, n10, n9);
xor  g71 (n92, n4, n12, n21, n7);
buf  g72 (n196, n54);
buf  g73 (n223, n63);
not  g74 (n140, n49);
buf  g75 (n216, n64);
not  g76 (n284, n38);
buf  g77 (n229, n34);
buf  g78 (n277, n75);
buf  g79 (n181, n38);
buf  g80 (n156, n75);
not  g81 (n226, n72);
buf  g82 (n250, n46);
buf  g83 (n221, n67);
buf  g84 (n153, n63);
not  g85 (n213, n63);
buf  g86 (n279, n65);
buf  g87 (n139, n59);
not  g88 (n272, n73);
not  g89 (n105, n70);
not  g90 (n182, n56);
not  g91 (n234, n71);
buf  g92 (n138, n66);
not  g93 (n188, n53);
not  g94 (n168, n40);
buf  g95 (n290, n37);
not  g96 (n256, n48);
buf  g97 (n253, n64);
buf  g98 (n283, n35);
not  g99 (n200, n65);
buf  g100 (n254, n41);
not  g101 (n113, n40);
not  g102 (n195, n58);
buf  g103 (n151, n39);
not  g104 (n165, n47);
not  g105 (n117, n73);
buf  g106 (n269, n62);
buf  g107 (n133, n50);
not  g108 (n162, n68);
buf  g109 (n131, n47);
buf  g110 (n237, n78);
not  g111 (n172, n62);
not  g112 (n194, n59);
buf  g113 (n235, n60);
not  g114 (n210, n58);
not  g115 (n218, n71);
buf  g116 (n144, n68);
buf  g117 (n110, n70);
not  g118 (n289, n65);
buf  g119 (n288, n71);
buf  g120 (n246, n52);
not  g121 (n108, n68);
not  g122 (n219, n70);
not  g123 (n189, n66);
not  g124 (n285, n36);
not  g125 (n228, n61);
not  g126 (n201, n75);
not  g127 (n206, n35);
buf  g128 (n192, n51);
not  g129 (n255, n37);
buf  g130 (n114, n54);
buf  g131 (n119, n76);
not  g132 (n115, n50);
not  g133 (n152, n41);
buf  g134 (n247, n46);
not  g135 (n170, n34);
not  g136 (n106, n43);
not  g137 (n273, n52);
not  g138 (n262, n35);
buf  g139 (n186, n66);
not  g140 (n251, n62);
not  g141 (n123, n62);
buf  g142 (n267, n42);
buf  g143 (n160, n33);
buf  g144 (n190, n78);
buf  g145 (n124, n40);
not  g146 (n177, n67);
not  g147 (n281, n79);
buf  g148 (n149, n70);
buf  g149 (n161, n64);
not  g150 (n159, n77);
buf  g151 (n282, n40);
not  g152 (n164, n46);
not  g153 (n230, n69);
buf  g154 (n180, n37);
not  g155 (n276, n36);
buf  g156 (n122, n61);
buf  g157 (n265, n59);
buf  g158 (n109, n39);
not  g159 (n154, n42);
buf  g160 (n174, n55);
buf  g161 (n214, n57);
buf  g162 (n249, n44);
not  g163 (n286, n56);
not  g164 (n155, n57);
buf  g165 (n121, n33);
buf  g166 (n111, n69);
buf  g167 (n143, n54);
buf  g168 (n204, n48);
not  g169 (n227, n74);
not  g170 (n130, n56);
not  g171 (n199, n58);
not  g172 (n175, n41);
not  g173 (n239, n58);
buf  g174 (n211, n65);
buf  g175 (n191, n78);
buf  g176 (n187, n64);
not  g177 (n112, n74);
buf  g178 (n148, n45);
buf  g179 (n236, n50);
buf  g180 (n241, n56);
buf  g181 (n163, n61);
not  g182 (n193, n34);
not  g183 (n127, n39);
not  g184 (n268, n72);
buf  g185 (n185, n59);
buf  g186 (n260, n72);
not  g187 (n135, n60);
not  g188 (n176, n69);
buf  g189 (n280, n77);
buf  g190 (n274, n76);
not  g191 (n134, n73);
buf  g192 (n287, n75);
buf  g193 (n157, n39);
buf  g194 (n198, n55);
buf  g195 (n118, n38);
buf  g196 (n258, n73);
not  g197 (n261, n36);
not  g198 (n263, n42);
not  g199 (n166, n55);
buf  g200 (n145, n76);
buf  g201 (n242, n35);
not  g202 (n212, n63);
buf  g203 (n183, n71);
not  g204 (n184, n47);
not  g205 (n128, n34);
not  g206 (n203, n79);
buf  g207 (n208, n78);
buf  g208 (n142, n60);
not  g209 (n270, n49);
not  g210 (n120, n33);
not  g211 (n179, n51);
buf  g212 (n146, n61);
not  g213 (n158, n53);
buf  g214 (n173, n44);
not  g215 (n126, n48);
not  g216 (n107, n57);
not  g217 (n264, n74);
not  g218 (n178, n53);
buf  g219 (n220, n77);
buf  g220 (n125, n36);
not  g221 (n243, n37);
buf  g222 (n252, n66);
buf  g223 (n238, n69);
buf  g224 (n171, n76);
buf  g225 (n244, n60);
buf  g226 (n136, n38);
not  g227 (n129, n41);
not  g228 (n225, n74);
not  g229 (n150, n43);
not  g230 (n257, n47);
not  g231 (n224, n72);
not  g232 (n222, n48);
buf  g233 (n275, n53);
buf  g234 (n245, n45);
not  g235 (n266, n33);
not  g236 (n215, n43);
not  g237 (n232, n67);
buf  g238 (n132, n49);
buf  g239 (n209, n49);
buf  g240 (n248, n54);
not  g241 (n207, n77);
buf  g242 (n233, n46);
buf  g243 (n231, n50);
not  g244 (n205, n68);
buf  g245 (n271, n67);
not  g246 (n147, n51);
not  g247 (n137, n57);
not  g248 (n202, n52);
not  g249 (n217, n51);
not  g250 (n240, n44);
buf  g251 (n259, n45);
not  g252 (n197, n52);
buf  g253 (n141, n45);
buf  g254 (n278, n42);
buf  g255 (n167, n44);
buf  g256 (n116, n55);
buf  g257 (n169, n43);
buf  g258 (n338, n272);
not  g259 (n349, n207);
buf  g260 (n454, n98);
not  g261 (n490, n80);
not  g262 (n325, n105);
not  g263 (n361, n189);
buf  g264 (n434, n121);
buf  g265 (n386, n164);
buf  g266 (n462, n209);
not  g267 (n380, n268);
not  g268 (n491, n149);
buf  g269 (n368, n194);
buf  g270 (n427, n164);
buf  g271 (n296, n144);
not  g272 (n464, n272);
not  g273 (n308, n171);
not  g274 (n298, n239);
buf  g275 (n399, n128);
buf  g276 (n517, n229);
buf  g277 (n457, n224);
not  g278 (n404, n85);
not  g279 (n449, n211);
not  g280 (n385, n288);
buf  g281 (n421, n175);
buf  g282 (n416, n264);
buf  g283 (n415, n170);
buf  g284 (n396, n264);
not  g285 (n480, n105);
xor  g286 (n329, n117, n135, n150, n268);
or   g287 (n374, n166, n118, n254, n240);
or   g288 (n514, n185, n83, n285, n216);
xnor g289 (n486, n213, n263, n220, n212);
xor  g290 (n458, n157, n168, n273, n281);
xor  g291 (n388, n92, n275, n267, n274);
nor  g292 (n472, n120, n286, n222, n202);
xor  g293 (n412, n211, n261, n270, n93);
nand g294 (n419, n225, n165, n212, n248);
nor  g295 (n305, n200, n282, n231, n111);
and  g296 (n381, n171, n206, n179, n152);
nor  g297 (n377, n232, n154, n220, n186);
nor  g298 (n451, n132, n130, n180, n262);
nand g299 (n442, n191, n209, n178, n221);
or   g300 (n471, n225, n192, n114, n91);
xnor g301 (n301, n113, n134, n287, n85);
xor  g302 (n468, n285, n198, n194, n163);
or   g303 (n474, n196, n152, n167, n226);
xnor g304 (n467, n116, n288, n139, n236);
nand g305 (n352, n216, n231, n154, n241);
or   g306 (n379, n227, n186, n125, n163);
nand g307 (n513, n273, n180, n107, n199);
nand g308 (n369, n251, n218, n147, n124);
nand g309 (n346, n220, n217, n219, n157);
xor  g310 (n433, n145, n134, n215, n148);
xnor g311 (n481, n258, n227, n214, n156);
or   g312 (n351, n230, n184, n108, n208);
and  g313 (n402, n121, n171, n149);
xor  g314 (n477, n108, n218, n89, n169);
nor  g315 (n487, n190, n162, n133, n112);
and  g316 (n340, n247, n251, n266, n155);
or   g317 (n339, n249, n90, n206, n137);
or   g318 (n297, n178, n258, n105, n123);
and  g319 (n398, n126, n110, n225);
xnor g320 (n510, n282, n258, n135, n259);
and  g321 (n341, n247, n130, n174, n279);
nand g322 (n494, n140, n256, n187, n181);
xor  g323 (n364, n245, n258, n242, n170);
xor  g324 (n366, n269, n167, n82, n286);
or   g325 (n470, n109, n252, n106, n84);
nand g326 (n327, n131, n275, n181, n215);
nand g327 (n429, n99, n82, n111, n184);
xnor g328 (n485, n200, n90, n158, n252);
xor  g329 (n445, n127, n238, n138, n212);
xor  g330 (n293, n254, n172, n263, n214);
nand g331 (n420, n264, n250, n184, n203);
nor  g332 (n303, n148, n137, n142, n160);
and  g333 (n432, n273, n153, n186, n84);
xnor g334 (n370, n198, n240, n280, n284);
nand g335 (n418, n143, n87, n129, n280);
xnor g336 (n410, n150, n83, n94, n114);
nor  g337 (n446, n159, n199, n140, n182);
or   g338 (n373, n119, n234, n225, n249);
and  g339 (n306, n155, n245, n233, n195);
or   g340 (n359, n133, n207, n289, n161);
xnor g341 (n372, n159, n120, n243, n228);
and  g342 (n392, n281, n196, n213, n243);
nand g343 (n356, n276, n88, n132, n123);
xnor g344 (n319, n173, n250, n281, n120);
and  g345 (n318, n213, n121, n232, n277);
nand g346 (n406, n118, n137, n90, n132);
nand g347 (n466, n205, n80, n237, n261);
and  g348 (n507, n261, n217, n229, n277);
nor  g349 (n300, n265, n274, n281, n257);
xor  g350 (n417, n242, n264, n219, n216);
xor  g351 (n328, n202, n189, n150, n149);
or   g352 (n413, n214, n112, n176, n204);
nand g353 (n501, n223, n97, n252, n128);
or   g354 (n342, n130, n157, n238, n197);
or   g355 (n394, n126, n154, n249, n149);
nand g356 (n314, n106, n94, n211, n125);
xor  g357 (n294, n110, n98, n164, n82);
xor  g358 (n322, n245, n271, n199);
and  g359 (n292, n266, n108, n253, n129);
xnor g360 (n358, n80, n93, n280, n250);
nand g361 (n335, n269, n96, n92, n197);
xor  g362 (n321, n205, n165, n204, n162);
or   g363 (n515, n162, n113, n129, n145);
xor  g364 (n334, n263, n172, n202, n242);
and  g365 (n407, n167, n141, n117, n289);
or   g366 (n307, n254, n156, n183, n142);
xor  g367 (n426, n95, n262, n176, n89);
nor  g368 (n483, n236, n127, n224, n215);
nand g369 (n409, n231, n210, n271, n246);
nor  g370 (n475, n205, n157, n244, n235);
or   g371 (n465, n277, n211, n253, n250);
xnor g372 (n291, n134, n177, n228, n181);
nor  g373 (n405, n213, n176, n147, n83);
and  g374 (n367, n232, n216, n270);
nand g375 (n389, n161, n166, n153, n123);
xnor g376 (n363, n181, n151, n133, n201);
nand g377 (n503, n159, n139, n91, n146);
or   g378 (n493, n219, n239, n185, n283);
nand g379 (n347, n136, n207, n197, n252);
xor  g380 (n295, n284, n247, n248, n173);
and  g381 (n443, n255, n151, n91, n210);
nor  g382 (n505, n128, n248, n273, n203);
xnor g383 (n425, n162, n97, n239, n210);
and  g384 (n344, n268, n166, n109, n283);
xor  g385 (n400, n175, n197, n87, n231);
xnor g386 (n343, n266, n138, n272, n148);
xnor g387 (n489, n173, n90, n253, n230);
xor  g388 (n492, n166, n165, n175, n170);
nand g389 (n350, n289, n190, n240, n127);
nor  g390 (n383, n182, n283, n191, n256);
xnor g391 (n313, n188, n251, n164, n98);
and  g392 (n357, n285, n265, n195, n95);
xnor g393 (n508, n269, n140, n236, n125);
nand g394 (n509, n112, n262, n278, n122);
and  g395 (n378, n119, n218, n222, n247);
xor  g396 (n430, n106, n260, n145, n238);
xnor g397 (n309, n208, n195, n259, n152);
or   g398 (n436, n141, n208, n88, n260);
or   g399 (n460, n141, n159, n185, n94);
nand g400 (n316, n99, n155, n108, n86);
xnor g401 (n362, n119, n86, n111, n263);
and  g402 (n326, n278, n160, n212, n163);
xnor g403 (n497, n287, n168, n260, n232);
nand g404 (n384, n85, n81, n189, n287);
xnor g405 (n516, n142, n114, n185, n175);
and  g406 (n302, n229, n98, n118, n122);
or   g407 (n453, n131, n153, n201, n272);
and  g408 (n304, n158, n173, n99, n182);
xor  g409 (n376, n92, n126, n191, n113);
xnor g410 (n310, n81, n84, n223, n174);
xnor g411 (n439, n97, n100, n275, n143);
xor  g412 (n324, n190, n84, n139, n244);
and  g413 (n437, n158, n282, n136, n246);
nor  g414 (n484, n246, n80, n187, n186);
xnor g415 (n375, n161, n177, n183, n286);
xor  g416 (n441, n260, n183, n136, n178);
and  g417 (n469, n191, n203, n178, n276);
nor  g418 (n428, n163, n116, n93, n82);
xnor g419 (n431, n205, n248, n122, n237);
xor  g420 (n337, n112, n274, n176, n168);
or   g421 (n512, n198, n279, n244, n223);
xor  g422 (n411, n141, n193, n243, n192);
xnor g423 (n479, n119, n276, n115, n184);
nand g424 (n482, n196, n135, n218, n131);
xor  g425 (n456, n246, n96, n174, n160);
nand g426 (n511, n196, n288, n245, n267);
nand g427 (n382, n132, n138, n255, n267);
and  g428 (n391, n279, n237, n137, n189);
or   g429 (n390, n279, n148, n115, n128);
or   g430 (n414, n187, n194, n215, n124);
xnor g431 (n403, n95, n204, n221, n188);
and  g432 (n395, n249, n282, n115, n79);
nand g433 (n447, n156, n257, n129, n174);
and  g434 (n498, n97, n105, n123, n136);
or   g435 (n488, n193, n242, n114, n217);
and  g436 (n435, n117, n224, n111, n251);
nor  g437 (n355, n235, n190, n86, n152);
or   g438 (n463, n241, n130, n228, n193);
xnor g439 (n299, n221, n262, n126, n256);
nor  g440 (n478, n161, n131, n83, n203);
xnor g441 (n336, n88, n287, n169, n210);
xor  g442 (n353, n233, n187, n86, n115);
nand g443 (n320, n100, n234, n142, n94);
or   g444 (n504, n261, n234, n107, n116);
nor  g445 (n459, n278, n202, n155, n228);
nand g446 (n444, n95, n199, n200, n234);
and  g447 (n499, n284, n217, n167, n214);
and  g448 (n496, n285, n280, n172, n222);
xor  g449 (n330, n233, n198, n237, n206);
nor  g450 (n397, n256, n150, n269, n177);
or   g451 (n424, n89, n89, n156, n192);
nand g452 (n365, n99, n233, n107, n146);
nand g453 (n495, n183, n268, n227, n220);
nor  g454 (n438, n201, n79, n92, n134);
nand g455 (n311, n81, n91, n139, n209);
or   g456 (n371, n219, n271, n201, n179);
xor  g457 (n450, n170, n172, n124, n188);
nand g458 (n333, n200, n106, n182, n226);
nor  g459 (n440, n127, n276, n153, n259);
xor  g460 (n401, n288, n122, n154, n87);
nand g461 (n452, n208, n144, n88, n147);
nor  g462 (n354, n240, n143, n151);
xnor g463 (n506, n267, n124, n275, n144);
or   g464 (n502, n116, n146, n235, n110);
nor  g465 (n423, n206, n180, n169);
or   g466 (n345, n192, n207, n179, n257);
nor  g467 (n473, n257, n265, n284, n146);
or   g468 (n387, n144, n277, n270, n117);
or   g469 (n348, n243, n125, n235, n188);
nor  g470 (n461, n209, n147, n239, n135);
xnor g471 (n323, n236, n118, n87, n81);
nand g472 (n331, n145, n244, n107, n113);
and  g473 (n455, n238, n230, n177);
and  g474 (n315, n93, n254, n195, n241);
or   g475 (n500, n255, n283, n158, n168);
nor  g476 (n448, n227, n194, n109, n133);
or   g477 (n360, n179, n140, n169, n253);
xor  g478 (n408, n241, n151, n286, n229);
nand g479 (n422, n266, n278, n121, n138);
xnor g480 (n317, n221, n96, n120, n274);
xor  g481 (n476, n109, n193, n224, n222);
xnor g482 (n393, n259, n226, n160, n289);
nor  g483 (n332, n265, n226, n255, n204);
or   g484 (n312, n165, n85, n223, n96);
buf  g485 (n547, n401);
buf  g486 (n570, n295);
not  g487 (n557, n292);
not  g488 (n554, n485);
nor  g489 (n533, n405, n406);
xnor g490 (n548, n344, n354, n316, n440);
or   g491 (n528, n395, n412, n392, n384);
nor  g492 (n560, n341, n375, n351, n389);
nand g493 (n546, n333, n298, n476, n414);
xnor g494 (n563, n457, n486, n449, n346);
or   g495 (n550, n381, n368, n408, n294);
xnor g496 (n524, n312, n443, n420, n332);
nand g497 (n536, n437, n371, n398, n442);
and  g498 (n559, n452, n355, n338, n369);
and  g499 (n545, n478, n313, n309, n471);
nand g500 (n539, n446, n393, n422, n303);
nand g501 (n519, n315, n453, n349, n366);
xnor g502 (n543, n376, n320, n402, n424);
nand g503 (n525, n328, n467, n327, n466);
nor  g504 (n555, n307, n318, n365, n324);
nand g505 (n542, n461, n435, n407, n374);
nor  g506 (n556, n394, n329, n445, n396);
xor  g507 (n562, n474, n441, n444, n310);
nand g508 (n537, n317, n464, n410, n431);
xor  g509 (n531, n390, n308, n319, n339);
nor  g510 (n569, n411, n475, n345, n304);
xnor g511 (n532, n300, n306, n387, n483);
nand g512 (n549, n469, n359, n334, n382);
nand g513 (n526, n472, n314, n348, n323);
xor  g514 (n544, n372, n343, n330, n385);
and  g515 (n566, n399, n347, n380, n409);
nor  g516 (n538, n463, n311, n462, n356);
xnor g517 (n520, n415, n439, n326, n297);
xnor g518 (n567, n488, n425, n373, n379);
xnor g519 (n553, n403, n305, n477, n454);
xnor g520 (n568, n448, n352, n481, n299);
xor  g521 (n530, n378, n342, n465, n426);
or   g522 (n534, n337, n386, n302, n447);
nand g523 (n518, n450, n391, n357, n322);
xor  g524 (n552, n388, n459, n423, n456);
and  g525 (n541, n331, n336, n404, n479);
xnor g526 (n521, n416, n436, n480, n487);
nand g527 (n523, n360, n421, n484, n430);
nor  g528 (n540, n301, n350, n361, n428);
xor  g529 (n551, n468, n335, n353, n400);
xnor g530 (n564, n418, n362, n427, n417);
and  g531 (n565, n434, n460, n429, n458);
nor  g532 (n561, n364, n433, n291, n367);
nand g533 (n535, n482, n419, n293, n438);
xor  g534 (n527, n377, n296, n432, n363);
xor  g535 (n529, n451, n321, n325, n383);
or   g536 (n558, n455, n397, n470, n358);
xor  g537 (n522, n473, n370, n340, n413);
buf  g538 (n579, n525);
not  g539 (n594, n528);
not  g540 (n595, n520);
not  g541 (n576, n529);
not  g542 (n572, n521);
buf  g543 (n574, n530);
not  g544 (n600, n523);
not  g545 (n597, n522);
not  g546 (n580, n522);
not  g547 (n591, n527);
buf  g548 (n577, n520);
not  g549 (n585, n530);
buf  g550 (n582, n527);
not  g551 (n587, n530);
not  g552 (n599, n518);
buf  g553 (n584, n529);
not  g554 (n601, n521);
not  g555 (n596, n528);
buf  g556 (n589, n529);
not  g557 (n588, n524);
buf  g558 (n598, n519);
buf  g559 (n583, n525);
buf  g560 (n581, n523);
buf  g561 (n593, n526);
buf  g562 (n590, n526);
and  g563 (n592, n519, n529, n524);
xnor g564 (n578, n528, n521, n527, n530);
nand g565 (n573, n518, n520, n523, n526);
and  g566 (n571, n525, n520, n524, n528);
and  g567 (n586, n524, n527, n522, n525);
nand g568 (n575, n523, n526, n521, n522);
not  g569 (n605, n535);
not  g570 (n603, n533);
buf  g571 (n608, n571);
buf  g572 (n604, n532);
buf  g573 (n607, n532);
buf  g574 (n602, n535);
nand g575 (n610, n574, n533);
xor  g576 (n613, n573, n535, n533, n574);
xor  g577 (n612, n572, n571, n534, n531);
xor  g578 (n606, n574, n532, n531);
xnor g579 (n609, n533, n572, n534);
xnor g580 (n614, n532, n573, n572);
nor  g581 (n611, n534, n531, n572, n573);
or   g582 (n623, n588, n602, n612, n540);
nand g583 (n648, n610, n538, n585, n595);
xor  g584 (n634, n598, n603, n542, n594);
xor  g585 (n619, n579, n610, n585, n611);
and  g586 (n631, n594, n578, n577);
nor  g587 (n620, n539, n578, n541, n612);
xnor g588 (n615, n595, n587, n609, n604);
xor  g589 (n617, n606, n609, n593, n586);
and  g590 (n650, n593, n606, n541, n598);
and  g591 (n624, n536, n582, n580, n606);
or   g592 (n638, n598, n607, n583);
or   g593 (n645, n598, n597, n605, n586);
nand g594 (n651, n593, n540, n577, n590);
xor  g595 (n642, n575, n576, n581, n542);
nand g596 (n641, n539, n590, n608, n537);
nor  g597 (n654, n587, n597, n581, n589);
and  g598 (n630, n542, n612, n538, n611);
xor  g599 (n621, n605, n588, n591, n595);
xnor g600 (n639, n593, n595, n604, n585);
xnor g601 (n632, n586, n536, n607, n603);
nand g602 (n633, n609, n592, n605, n604);
xnor g603 (n628, n608, n539, n579, n580);
nor  g604 (n656, n596, n537, n592, n540);
xor  g605 (n640, n589, n579, n584, n582);
or   g606 (n625, n582, n603, n611, n538);
or   g607 (n635, n604, n596, n581, n590);
and  g608 (n637, n586, n591, n608, n540);
nand g609 (n644, n613, n575, n584, n576);
nor  g610 (n616, n579, n603, n537, n612);
xnor g611 (n652, n587, n589, n577, n581);
nand g612 (n629, n541, n596, n542);
nor  g613 (n653, n610, n541, n574, n577);
xnor g614 (n636, n607, n576, n592, n538);
or   g615 (n646, n597, n588, n594, n606);
nor  g616 (n618, n608, n537, n591, n578);
nor  g617 (n647, n611, n535, n536, n594);
xor  g618 (n627, n584, n575, n605, n607);
and  g619 (n655, n589, n592, n597, n583);
xor  g620 (n649, n582, n536, n591, n580);
and  g621 (n626, n576, n583, n590, n580);
nor  g622 (n643, n539, n587, n610, n575);
or   g623 (n622, n585, n584, n588, n609);
buf  g624 (n661, n643);
buf  g625 (n664, n544);
and  g626 (n659, n640, n544);
nor  g627 (n663, n637, n645, n648);
xor  g628 (n670, n543, n546, n544);
and  g629 (n672, n614, n613, n543);
and  g630 (n657, n651, n601, n599);
xnor g631 (n662, n546, n634, n545);
nor  g632 (n674, n631, n546, n649);
xnor g633 (n660, n632, n543, n635);
or   g634 (n673, n646, n642, n599);
xnor g635 (n669, n613, n600);
nand g636 (n668, n641, n601, n639);
or   g637 (n667, n650, n638, n644);
nand g638 (n666, n636, n633, n599);
nor  g639 (n665, n545, n543, n601);
nor  g640 (n676, n600, n545);
xor  g641 (n658, n546, n614, n600);
nand g642 (n671, n614, n647, n601);
nand g643 (n675, n613, n599, n614);
or   g644 (n678, n663, n676);
xor  g645 (n681, n659, n548, n100, n658);
and  g646 (n680, n657, n490, n547, n658);
xor  g647 (n690, n502, n663, n666, n662);
nor  g648 (n684, n23, n661, n547, n492);
nor  g649 (n704, n25, n669, n26, n654);
and  g650 (n691, n670, n667, n661, n550);
and  g651 (n708, n499, n672, n673, n494);
and  g652 (n687, n25, n676, n496, n668);
nand g653 (n700, n663, n101, n500, n497);
nor  g654 (n689, n662, n549, n674, n658);
nor  g655 (n703, n103, n24, n673, n671);
or   g656 (n713, n24, n670, n669, n22);
xnor g657 (n697, n666, n655, n550);
and  g658 (n706, n23, n101, n668, n659);
xnor g659 (n696, n550, n661, n676, n675);
xor  g660 (n695, n24, n661, n664);
and  g661 (n711, n657, n665, n101, n674);
or   g662 (n685, n674, n101, n548);
xnor g663 (n677, n26, n659, n504, n102);
and  g664 (n688, n549, n652, n100, n23);
or   g665 (n683, n666, n547, n676, n658);
and  g666 (n702, n665, n489, n548, n503);
and  g667 (n710, n671, n660, n495, n664);
xnor g668 (n679, n674, n549, n665, n671);
and  g669 (n699, n26, n675, n670, n657);
and  g670 (n701, n23, n491, n660, n673);
nand g671 (n692, n662, n672);
xor  g672 (n705, n666, n663, n25, n669);
or   g673 (n698, n24, n672, n656, n675);
nor  g674 (n693, n102, n657, n653, n25);
or   g675 (n694, n660, n670, n103, n668);
or   g676 (n686, n660, n659, n501, n665);
xor  g677 (n707, n549, n675, n102, n498);
or   g678 (n682, n667, n547, n673, n103);
and  g679 (n709, n102, n664, n667);
nor  g680 (n712, n493, n668, n669, n671);
buf  g681 (n718, n688);
not  g682 (n747, n694);
buf  g683 (n731, n686);
buf  g684 (n735, n695);
buf  g685 (n726, n682);
buf  g686 (n716, n692);
not  g687 (n715, n683);
not  g688 (n737, n690);
not  g689 (n740, n690);
buf  g690 (n714, n684);
buf  g691 (n725, n694);
not  g692 (n732, n679);
buf  g693 (n736, n679);
not  g694 (n745, n680);
not  g695 (n741, n691);
buf  g696 (n748, n686);
buf  g697 (n742, n677);
not  g698 (n730, n678);
buf  g699 (n743, n685);
not  g700 (n746, n683);
buf  g701 (n723, n681);
buf  g702 (n717, n684);
buf  g703 (n727, n689);
buf  g704 (n721, n685);
buf  g705 (n738, n693);
buf  g706 (n733, n691);
buf  g707 (n729, n687);
not  g708 (n720, n680);
not  g709 (n722, n687);
not  g710 (n744, n682);
buf  g711 (n728, n692);
not  g712 (n749, n689);
not  g713 (n734, n693);
not  g714 (n739, n681);
buf  g715 (n719, n688);
not  g716 (n724, n678);
nor  g717 (n753, n723, n708, n728);
or   g718 (n784, n707, n746, n729, n559);
or   g719 (n757, n710, n735, n704, n552);
nand g720 (n789, n712, n745, n735, n741);
nand g721 (n773, n734, n725, n556, n737);
xor  g722 (n762, n554, n742, n719, n732);
or   g723 (n794, n716, n698, n725, n746);
or   g724 (n763, n731, n558, n709, n739);
or   g725 (n801, n725, n740, n732, n743);
xnor g726 (n752, n560, n560, n742, n555);
or   g727 (n797, n741, n718, n559, n748);
xor  g728 (n769, n702, n730, n554, n700);
nor  g729 (n798, n728, n711, n745, n727);
xor  g730 (n778, n557, n551, n731, n727);
and  g731 (n779, n747, n723, n749, n702);
nor  g732 (n785, n714, n558, n715, n744);
or   g733 (n782, n720, n749, n552, n719);
nor  g734 (n800, n737, n700, n716, n710);
xnor g735 (n772, n728, n734, n557, n743);
nand g736 (n787, n727, n722, n555, n720);
xor  g737 (n796, n738, n747, n708, n733);
xnor g738 (n765, n713, n747, n722, n736);
xnor g739 (n764, n723, n719, n714, n737);
xnor g740 (n771, n557, n727, n720, n705);
and  g741 (n776, n722, n729, n740, n747);
xnor g742 (n802, n735, n714, n701, n712);
xor  g743 (n760, n703, n715, n558, n722);
xnor g744 (n759, n733, n724, n706, n697);
xor  g745 (n790, n699, n726, n555, n748);
or   g746 (n770, n730, n743, n721, n749);
xnor g747 (n799, n717, n744, n552, n725);
nand g748 (n767, n717, n717, n704, n696);
xor  g749 (n750, n729, n744, n558, n748);
xor  g750 (n775, n744, n716, n717);
or   g751 (n783, n554, n739, n553, n697);
or   g752 (n792, n556, n742, n738, n731);
xnor g753 (n804, n559, n554, n557, n741);
or   g754 (n803, n719, n748, n726, n745);
nand g755 (n755, n551, n721, n701, n740);
xor  g756 (n788, n729, n706, n715, n734);
and  g757 (n761, n738, n555, n724, n707);
xnor g758 (n756, n723, n734, n721, n735);
nand g759 (n795, n713, n741, n556, n718);
nand g760 (n786, n705, n721, n736, n738);
xor  g761 (n780, n709, n740, n699, n718);
xor  g762 (n766, n732, n746, n726, n724);
nor  g763 (n768, n736, n746, n743, n726);
and  g764 (n781, n715, n730, n737, n714);
nand g765 (n777, n736, n553, n731, n551);
xnor g766 (n791, n718, n698, n745, n739);
nor  g767 (n793, n552, n553, n559, n711);
nand g768 (n758, n730, n695, n703, n733);
and  g769 (n751, n553, n696, n733, n739);
nor  g770 (n774, n720, n551, n728, n749);
and  g771 (n754, n742, n556, n732, n724);
not  g772 (n859, n797);
not  g773 (n824, n790);
not  g774 (n855, n795);
not  g775 (n845, n791);
buf  g776 (n808, n789);
not  g777 (n850, n776);
not  g778 (n838, n786);
buf  g779 (n836, n793);
buf  g780 (n854, n789);
buf  g781 (n831, n804);
not  g782 (n858, n802);
not  g783 (n809, n797);
not  g784 (n819, n765);
not  g785 (n813, n789);
buf  g786 (n844, n760);
buf  g787 (n835, n770);
buf  g788 (n846, n766);
not  g789 (n842, n752);
buf  g790 (n852, n795);
not  g791 (n867, n787);
not  g792 (n848, n782);
not  g793 (n865, n799);
not  g794 (n869, n751);
buf  g795 (n832, n791);
buf  g796 (n810, n788);
buf  g797 (n833, n794);
not  g798 (n805, n759);
not  g799 (n834, n756);
not  g800 (n823, n791);
not  g801 (n806, n778);
not  g802 (n829, n787);
not  g803 (n821, n804);
not  g804 (n856, n787);
not  g805 (n870, n753);
buf  g806 (n817, n802);
not  g807 (n843, n803);
buf  g808 (n847, n797);
buf  g809 (n818, n773);
not  g810 (n828, n803);
buf  g811 (n820, n795);
not  g812 (n851, n757);
not  g813 (n866, n780);
buf  g814 (n822, n771);
buf  g815 (n830, n772);
buf  g816 (n827, n799);
buf  g817 (n807, n801);
and  g818 (n853, n796, n804);
xnor g819 (n826, n800, n796, n783);
nor  g820 (n814, n801, n798, n775);
nor  g821 (n868, n785, n796, n800);
or   g822 (n812, n763, n799, n769);
nand g823 (n825, n794, n801, n790);
and  g824 (n839, n798, n794, n800);
nor  g825 (n840, n802, n789, n755);
nor  g826 (n863, n787, n801, n781);
and  g827 (n849, n799, n790, n792);
xnor g828 (n864, n788, n777, n784);
nor  g829 (n862, n758, n792, n795);
xor  g830 (n815, n774, n792, n788);
xor  g831 (n860, n767, n761, n792);
and  g832 (n857, n794, n788, n798);
xnor g833 (n811, n754, n803, n796);
nor  g834 (n837, n798, n793);
xor  g835 (n861, n803, n802, n779);
and  g836 (n871, n797, n800, n793);
nand g837 (n841, n791, n762, n764);
or   g838 (n816, n790, n768, n804);
buf  g839 (n887, n811);
buf  g840 (n877, n813);
buf  g841 (n875, n812);
buf  g842 (n872, n811);
not  g843 (n884, n807);
not  g844 (n885, n805);
not  g845 (n888, n808);
buf  g846 (n890, n810);
buf  g847 (n882, n808);
buf  g848 (n876, n814);
not  g849 (n891, n807);
buf  g850 (n881, n809);
not  g851 (n883, n808);
not  g852 (n874, n806);
or   g853 (n889, n807, n806, n805, n812);
xor  g854 (n886, n810, n810, n811, n806);
xor  g855 (n873, n807, n806, n812, n805);
xnor g856 (n879, n810, n813, n809);
xor  g857 (n880, n813, n814, n811, n809);
xor  g858 (n878, n812, n813, n805, n808);
or   g859 (n971, n859, n818);
xor  g860 (n918, n880, n888, n863, n846);
and  g861 (n904, n847, n839, n816, n832);
nor  g862 (n969, n838, n876, n883, n817);
nand g863 (n911, n814, n876, n840, n824);
nor  g864 (n899, n883, n842, n853, n854);
nor  g865 (n945, n837, n833, n850, n891);
and  g866 (n928, n850, n890, n824, n836);
nor  g867 (n946, n823, n882, n868, n855);
and  g868 (n953, n819, n857, n861, n871);
xnor g869 (n898, n867, n857, n828, n849);
or   g870 (n968, n858, n873, n881, n854);
nor  g871 (n967, n863, n855, n833, n879);
nor  g872 (n938, n848, n830, n815, n863);
xor  g873 (n935, n835, n891, n877, n882);
or   g874 (n936, n839, n821, n827, n814);
or   g875 (n919, n875, n857, n852, n863);
or   g876 (n939, n884, n845, n834, n829);
xnor g877 (n917, n820, n888, n827, n831);
or   g878 (n940, n835, n846, n870, n887);
xnor g879 (n920, n837, n859, n832, n857);
nor  g880 (n965, n862, n878, n821, n888);
nor  g881 (n896, n841, n865, n844, n883);
xnor g882 (n970, n849, n844, n866, n840);
xnor g883 (n925, n824, n824, n855, n817);
nor  g884 (n951, n861, n881, n828, n825);
or   g885 (n895, n885, n831, n839, n891);
nand g886 (n916, n871, n836, n875, n822);
or   g887 (n947, n871, n837, n846, n856);
or   g888 (n892, n817, n831, n561, n877);
xnor g889 (n927, n822, n877, n886);
nor  g890 (n963, n816, n860, n828, n858);
nor  g891 (n921, n837, n832, n879);
xnor g892 (n934, n887, n889, n838, n848);
xnor g893 (n893, n838, n831, n834, n866);
xnor g894 (n931, n884, n889, n859, n870);
xnor g895 (n957, n873, n864, n880, n823);
and  g896 (n933, n561, n890, n887, n816);
nor  g897 (n960, n816, n886, n858, n855);
and  g898 (n955, n841, n835, n843, n842);
xnor g899 (n948, n870, n820, n562, n832);
nor  g900 (n929, n853, n826, n873, n877);
xnor g901 (n966, n885, n842, n852, n817);
nor  g902 (n924, n838, n883, n833, n867);
xnor g903 (n894, n830, n875, n862, n815);
or   g904 (n897, n849, n875, n818, n847);
xor  g905 (n932, n872, n844, n876, n829);
xnor g906 (n942, n866, n836, n865, n864);
xnor g907 (n910, n868, n871, n872, n820);
nor  g908 (n941, n818, n884, n890, n825);
xnor g909 (n937, n562, n851, n865, n849);
and  g910 (n923, n826, n836, n835, n861);
nand g911 (n912, n868, n858, n840, n827);
nand g912 (n914, n820, n854, n822, n846);
nand g913 (n949, n815, n880, n827, n560);
and  g914 (n913, n842, n885, n860, n847);
xnor g915 (n900, n865, n830, n822, n845);
xnor g916 (n902, n862, n825, n867);
xnor g917 (n952, n874, n874, n869, n882);
xnor g918 (n901, n885, n841, n850, n881);
nand g919 (n903, n869, n853, n889, n851);
and  g920 (n950, n860, n828, n829, n834);
xnor g921 (n909, n826, n834, n853, n860);
or   g922 (n905, n866, n845, n879, n561);
nor  g923 (n962, n874, n862, n856, n864);
xnor g924 (n922, n874, n856, n888, n819);
nand g925 (n956, n852, n843, n818, n819);
xnor g926 (n944, n867, n560, n878, n861);
nand g927 (n958, n850, n876, n841, n823);
or   g928 (n959, n848, n884, n881, n859);
xnor g929 (n915, n869, n856, n819, n891);
and  g930 (n907, n873, n839, n840, n869);
nor  g931 (n954, n844, n851, n829, n821);
nand g932 (n906, n826, n848, n886, n843);
xor  g933 (n964, n889, n821, n854, n890);
nor  g934 (n926, n878, n864, n872, n847);
xnor g935 (n930, n882, n830, n823, n845);
nor  g936 (n961, n868, n878, n815, n870);
xnor g937 (n943, n851, n880, n872, n833);
xor  g938 (n908, n561, n887, n843, n852);
and  g939 (n984, n956, n562, n955);
xnor g940 (n973, n936, n919, n932, n940);
xor  g941 (n991, n931, n908, n963, n926);
xnor g942 (n990, n944, n902, n918, n898);
nand g943 (n989, n943, n900, n892, n894);
nor  g944 (n974, n962, n960, n964, n947);
and  g945 (n985, n925, n895, n953, n945);
nor  g946 (n977, n912, n927, n921, n924);
and  g947 (n983, n933, n911, n958, n910);
nand g948 (n992, n906, n916, n913, n920);
nor  g949 (n981, n960, n951, n939, n930);
and  g950 (n975, n952, n923, n935, n962);
xnor g951 (n986, n948, n903, n961, n942);
and  g952 (n982, n914, n962, n922, n949);
nor  g953 (n976, n961, n907, n963, n959);
xor  g954 (n972, n937, n899, n964, n901);
xor  g955 (n988, n893, n904, n929, n946);
or   g956 (n978, n928, n905, n962, n950);
and  g957 (n979, n917, n896, n957, n963);
and  g958 (n987, n909, n941, n938, n954);
nand g959 (n980, n897, n963, n934, n915);
xor  g960 (n1010, n564, n968, n565, n103);
xor  g961 (n1000, n983, n991, n565, n964);
and  g962 (n1004, n990, n567, n976, n566);
and  g963 (n1003, n967, n975, n992, n565);
xnor g964 (n996, n104, n971, n977, n979);
and  g965 (n993, n563, n970, n985, n964);
or   g966 (n1006, n104, n971, n965, n966);
and  g967 (n1009, n970, n968, n563, n965);
nand g968 (n997, n987, n563, n970);
or   g969 (n1008, n104, n967, n969, n968);
nor  g970 (n999, n968, n988, n566, n981);
xnor g971 (n998, n966, n967, n566, n565);
nor  g972 (n1001, n563, n965, n986, n564);
xnor g973 (n995, n967, n969, n971, n564);
nor  g974 (n1007, n989, n980, n104, n973);
and  g975 (n994, n971, n965, n982, n966);
nand g976 (n1005, n969, n966, n974, n978);
nand g977 (n1002, n564, n984, n969, n566);
or   g978 (n1024, n511, n29, n31, n30);
xnor g979 (n1017, n569, n26, n31, n514);
nand g980 (n1012, n998, n32, n567, n1008);
nand g981 (n1023, n513, n30, n508);
xnor g982 (n1018, n27, n1006, n31, n28);
nand g983 (n1016, n515, n509, n997, n32);
nor  g984 (n1015, n568, n27, n1004, n569);
and  g985 (n1013, n568, n1001, n507, n1010);
xor  g986 (n1022, n568, n1007, n28, n32);
xnor g987 (n1011, n512, n28, n999, n567);
xnor g988 (n1019, n31, n29, n32, n27);
xnor g989 (n1021, n1009, n1005, n996, n1003);
nor  g990 (n1025, n506, n568, n1002, n29);
nor  g991 (n1014, n28, n567, n505, n29);
xor  g992 (n1020, n1000, n30, n510, n27);
xnor g993 (n1026, n569, n1024, n1022);
and  g994 (n1027, n1020, n570, n1021);
xnor g995 (n1028, n569, n1019, n1023, n1025);
nor  g996 (n1029, n1026, n570);
or   g997 (n1031, n1027, n1029, n516, n1028);
xnor g998 (n1032, n517, n1029, n290);
or   g999 (n1030, n1029, n290);
endmodule
