

module Stat_2000_223
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n731,
  n741,
  n737,
  n736,
  n739,
  n740,
  n738,
  n733,
  n730,
  n748,
  n747,
  n729,
  n746,
  n745,
  n742,
  n734,
  n744,
  n743,
  n2019,
  n2021,
  n2025,
  n2023,
  n2026,
  n2032,
  n2031,
  n2030,
  n2024,
  n2022,
  n2028,
  n2029,
  n2020,
  n2027
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n731;output n741;output n737;output n736;output n739;output n740;output n738;output n733;output n730;output n748;output n747;output n729;output n746;output n745;output n742;output n734;output n744;output n743;output n2019;output n2021;output n2025;output n2023;output n2026;output n2032;output n2031;output n2030;output n2024;output n2022;output n2028;output n2029;output n2020;output n2027;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n732;wire n735;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  buf
  g0
  (
    n43,
    n22
  );


  buf
  g1
  (
    n90,
    n29
  );


  buf
  g2
  (
    n114,
    n7
  );


  buf
  g3
  (
    n104,
    n28
  );


  buf
  g4
  (
    n100,
    n11
  );


  buf
  g5
  (
    n136,
    n4
  );


  buf
  g6
  (
    n141,
    n7
  );


  buf
  g7
  (
    n96,
    n26
  );


  not
  g8
  (
    n93,
    n29
  );


  buf
  g9
  (
    n95,
    n13
  );


  buf
  g10
  (
    n72,
    n16
  );


  buf
  g11
  (
    n53,
    n9
  );


  buf
  g12
  (
    n110,
    n4
  );


  buf
  g13
  (
    n92,
    n5
  );


  buf
  g14
  (
    n121,
    n21
  );


  not
  g15
  (
    n148,
    n9
  );


  buf
  g16
  (
    n40,
    n19
  );


  buf
  g17
  (
    n76,
    n10
  );


  buf
  g18
  (
    n140,
    n8
  );


  not
  g19
  (
    n78,
    n12
  );


  not
  g20
  (
    n49,
    n3
  );


  not
  g21
  (
    n108,
    n2
  );


  buf
  g22
  (
    n87,
    n30
  );


  not
  g23
  (
    n97,
    n10
  );


  buf
  g24
  (
    n130,
    n21
  );


  not
  g25
  (
    n55,
    n24
  );


  not
  g26
  (
    n57,
    n27
  );


  buf
  g27
  (
    n41,
    n15
  );


  not
  g28
  (
    n42,
    n1
  );


  not
  g29
  (
    n81,
    n18
  );


  not
  g30
  (
    n124,
    n11
  );


  not
  g31
  (
    n37,
    n25
  );


  not
  g32
  (
    n139,
    n6
  );


  buf
  g33
  (
    n132,
    n12
  );


  not
  g34
  (
    n88,
    n14
  );


  not
  g35
  (
    n61,
    n17
  );


  buf
  g36
  (
    n51,
    n20
  );


  buf
  g37
  (
    n116,
    n4
  );


  not
  g38
  (
    n71,
    n16
  );


  not
  g39
  (
    KeyWire_0_2,
    n10
  );


  buf
  g40
  (
    n79,
    n14
  );


  buf
  g41
  (
    n33,
    n1
  );


  buf
  g42
  (
    n120,
    n7
  );


  not
  g43
  (
    n138,
    n13
  );


  not
  g44
  (
    n115,
    n28
  );


  not
  g45
  (
    n119,
    n7
  );


  not
  g46
  (
    n128,
    n18
  );


  buf
  g47
  (
    n137,
    n23
  );


  buf
  g48
  (
    n39,
    n24
  );


  not
  g49
  (
    n46,
    n12
  );


  buf
  g50
  (
    n60,
    n20
  );


  not
  g51
  (
    n58,
    n26
  );


  buf
  g52
  (
    n36,
    n2
  );


  not
  g53
  (
    n99,
    n30
  );


  buf
  g54
  (
    n82,
    n8
  );


  buf
  g55
  (
    n52,
    n29
  );


  buf
  g56
  (
    n68,
    n23
  );


  buf
  g57
  (
    n133,
    n22
  );


  not
  g58
  (
    n131,
    n27
  );


  buf
  g59
  (
    n50,
    n8
  );


  buf
  g60
  (
    n69,
    n29
  );


  buf
  g61
  (
    n149,
    n28
  );


  buf
  g62
  (
    n45,
    n3
  );


  buf
  g63
  (
    n70,
    n4
  );


  buf
  g64
  (
    n47,
    n24
  );


  not
  g65
  (
    n105,
    n22
  );


  not
  g66
  (
    n56,
    n18
  );


  not
  g67
  (
    n80,
    n9
  );


  buf
  g68
  (
    n38,
    n20
  );


  not
  g69
  (
    n123,
    n15
  );


  not
  g70
  (
    n129,
    n13
  );


  not
  g71
  (
    n135,
    n17
  );


  not
  g72
  (
    n59,
    n13
  );


  not
  g73
  (
    n94,
    n6
  );


  not
  g74
  (
    n83,
    n24
  );


  buf
  g75
  (
    n64,
    n5
  );


  buf
  g76
  (
    n134,
    n3
  );


  buf
  g77
  (
    n34,
    n26
  );


  not
  g78
  (
    n84,
    n23
  );


  not
  g79
  (
    KeyWire_0_12,
    n12
  );


  not
  g80
  (
    n127,
    n2
  );


  not
  g81
  (
    n86,
    n20
  );


  buf
  g82
  (
    n143,
    n25
  );


  buf
  g83
  (
    n62,
    n19
  );


  not
  g84
  (
    n89,
    n17
  );


  buf
  g85
  (
    n117,
    n21
  );


  not
  g86
  (
    n101,
    n1
  );


  not
  g87
  (
    n65,
    n14
  );


  buf
  g88
  (
    n113,
    n23
  );


  buf
  g89
  (
    n122,
    n19
  );


  buf
  g90
  (
    n142,
    n25
  );


  not
  g91
  (
    n112,
    n8
  );


  buf
  g92
  (
    n54,
    n22
  );


  not
  g93
  (
    n151,
    n15
  );


  buf
  g94
  (
    n125,
    n25
  );


  not
  g95
  (
    n106,
    n11
  );


  buf
  g96
  (
    n85,
    n16
  );


  not
  g97
  (
    n126,
    n30
  );


  buf
  g98
  (
    n102,
    n14
  );


  not
  g99
  (
    n147,
    n18
  );


  not
  g100
  (
    n44,
    n27
  );


  not
  g101
  (
    n66,
    n10
  );


  buf
  g102
  (
    n75,
    n27
  );


  not
  g103
  (
    n77,
    n17
  );


  buf
  g104
  (
    n111,
    n15
  );


  not
  g105
  (
    n91,
    n21
  );


  buf
  g106
  (
    n98,
    n28
  );


  not
  g107
  (
    n150,
    n1
  );


  not
  g108
  (
    n146,
    n19
  );


  not
  g109
  (
    n74,
    n9
  );


  buf
  g110
  (
    n35,
    n16
  );


  buf
  g111
  (
    n144,
    n5
  );


  not
  g112
  (
    n48,
    n11
  );


  buf
  g113
  (
    n63,
    n2
  );


  not
  g114
  (
    n145,
    n5
  );


  not
  g115
  (
    n103,
    n3
  );


  buf
  g116
  (
    n67,
    n6
  );


  buf
  g117
  (
    n73,
    n26
  );


  buf
  g118
  (
    n118,
    n6
  );


  not
  g119
  (
    n335,
    n140
  );


  buf
  g120
  (
    n551,
    n111
  );


  buf
  g121
  (
    n349,
    n75
  );


  not
  g122
  (
    n322,
    n55
  );


  not
  g123
  (
    n540,
    n50
  );


  buf
  g124
  (
    n352,
    n36
  );


  buf
  g125
  (
    n171,
    n37
  );


  not
  g126
  (
    n556,
    n95
  );


  not
  g127
  (
    n180,
    n97
  );


  not
  g128
  (
    n497,
    n35
  );


  buf
  g129
  (
    n324,
    n38
  );


  buf
  g130
  (
    n248,
    n128
  );


  not
  g131
  (
    n523,
    n71
  );


  buf
  g132
  (
    n474,
    n51
  );


  not
  g133
  (
    n371,
    n85
  );


  not
  g134
  (
    n276,
    n90
  );


  buf
  g135
  (
    n513,
    n53
  );


  not
  g136
  (
    n301,
    n115
  );


  buf
  g137
  (
    n380,
    n114
  );


  buf
  g138
  (
    n220,
    n90
  );


  not
  g139
  (
    n168,
    n139
  );


  not
  g140
  (
    n234,
    n40
  );


  buf
  g141
  (
    n267,
    n58
  );


  not
  g142
  (
    n297,
    n107
  );


  not
  g143
  (
    n264,
    n131
  );


  not
  g144
  (
    n161,
    n127
  );


  not
  g145
  (
    n461,
    n141
  );


  not
  g146
  (
    n366,
    n108
  );


  not
  g147
  (
    n369,
    n56
  );


  not
  g148
  (
    n411,
    n112
  );


  buf
  g149
  (
    n299,
    n98
  );


  not
  g150
  (
    n412,
    n74
  );


  buf
  g151
  (
    n339,
    n106
  );


  buf
  g152
  (
    n174,
    n89
  );


  not
  g153
  (
    n280,
    n86
  );


  not
  g154
  (
    n244,
    n89
  );


  not
  g155
  (
    n166,
    n42
  );


  buf
  g156
  (
    n320,
    n135
  );


  buf
  g157
  (
    n392,
    n63
  );


  not
  g158
  (
    n178,
    n136
  );


  not
  g159
  (
    n545,
    n108
  );


  not
  g160
  (
    n510,
    n128
  );


  buf
  g161
  (
    n293,
    n95
  );


  buf
  g162
  (
    n365,
    n73
  );


  not
  g163
  (
    n268,
    n48
  );


  buf
  g164
  (
    n478,
    n118
  );


  not
  g165
  (
    n585,
    n137
  );


  not
  g166
  (
    n323,
    n116
  );


  not
  g167
  (
    n194,
    n62
  );


  not
  g168
  (
    n399,
    n60
  );


  not
  g169
  (
    n457,
    n113
  );


  not
  g170
  (
    n415,
    n43
  );


  buf
  g171
  (
    n527,
    n108
  );


  not
  g172
  (
    n203,
    n119
  );


  not
  g173
  (
    n406,
    n42
  );


  buf
  g174
  (
    n395,
    n78
  );


  not
  g175
  (
    n390,
    n72
  );


  not
  g176
  (
    n259,
    n117
  );


  not
  g177
  (
    n218,
    n45
  );


  not
  g178
  (
    n193,
    n48
  );


  buf
  g179
  (
    n153,
    n134
  );


  buf
  g180
  (
    n524,
    n38
  );


  not
  g181
  (
    n489,
    n133
  );


  buf
  g182
  (
    n450,
    n60
  );


  not
  g183
  (
    n331,
    n84
  );


  buf
  g184
  (
    n182,
    n140
  );


  buf
  g185
  (
    n359,
    n98
  );


  buf
  g186
  (
    n566,
    n53
  );


  buf
  g187
  (
    n375,
    n54
  );


  not
  g188
  (
    n228,
    n105
  );


  buf
  g189
  (
    n177,
    n113
  );


  not
  g190
  (
    n291,
    n67
  );


  not
  g191
  (
    n424,
    n56
  );


  not
  g192
  (
    n295,
    n101
  );


  buf
  g193
  (
    n572,
    n107
  );


  buf
  g194
  (
    n567,
    n62
  );


  buf
  g195
  (
    n209,
    n46
  );


  buf
  g196
  (
    n360,
    n107
  );


  buf
  g197
  (
    n443,
    n115
  );


  buf
  g198
  (
    n515,
    n121
  );


  buf
  g199
  (
    n285,
    n110
  );


  not
  g200
  (
    n441,
    n81
  );


  buf
  g201
  (
    n482,
    n67
  );


  not
  g202
  (
    n238,
    n36
  );


  buf
  g203
  (
    n310,
    n90
  );


  not
  g204
  (
    n314,
    n34
  );


  not
  g205
  (
    n184,
    n37
  );


  not
  g206
  (
    n189,
    n38
  );


  buf
  g207
  (
    n356,
    n104
  );


  buf
  g208
  (
    n451,
    n132
  );


  buf
  g209
  (
    n565,
    n127
  );


  buf
  g210
  (
    n345,
    n130
  );


  not
  g211
  (
    n281,
    n103
  );


  not
  g212
  (
    n553,
    n92
  );


  buf
  g213
  (
    n508,
    n72
  );


  not
  g214
  (
    n517,
    n134
  );


  buf
  g215
  (
    n577,
    n66
  );


  buf
  g216
  (
    n408,
    n121
  );


  buf
  g217
  (
    n200,
    n68
  );


  buf
  g218
  (
    n219,
    n123
  );


  buf
  g219
  (
    n284,
    n89
  );


  buf
  g220
  (
    n279,
    n75
  );


  buf
  g221
  (
    n377,
    n52
  );


  buf
  g222
  (
    n463,
    n82
  );


  buf
  g223
  (
    n422,
    n81
  );


  not
  g224
  (
    n444,
    n33
  );


  not
  g225
  (
    n420,
    n51
  );


  buf
  g226
  (
    n315,
    n54
  );


  not
  g227
  (
    n470,
    n137
  );


  buf
  g228
  (
    n459,
    n137
  );


  buf
  g229
  (
    n409,
    n130
  );


  not
  g230
  (
    n475,
    n77
  );


  buf
  g231
  (
    n430,
    n132
  );


  buf
  g232
  (
    n346,
    n141
  );


  buf
  g233
  (
    n538,
    n66
  );


  buf
  g234
  (
    n312,
    n122
  );


  buf
  g235
  (
    n247,
    n125
  );


  buf
  g236
  (
    n340,
    n132
  );


  buf
  g237
  (
    n266,
    n41
  );


  not
  g238
  (
    n256,
    n66
  );


  buf
  g239
  (
    n319,
    n53
  );


  buf
  g240
  (
    n574,
    n129
  );


  not
  g241
  (
    n531,
    n33
  );


  not
  g242
  (
    n535,
    n129
  );


  buf
  g243
  (
    n169,
    n139
  );


  buf
  g244
  (
    n428,
    n94
  );


  buf
  g245
  (
    n313,
    n126
  );


  buf
  g246
  (
    n418,
    n36
  );


  not
  g247
  (
    n544,
    n73
  );


  buf
  g248
  (
    n208,
    n101
  );


  buf
  g249
  (
    n271,
    n125
  );


  buf
  g250
  (
    n576,
    n100
  );


  buf
  g251
  (
    n241,
    n111
  );


  buf
  g252
  (
    n274,
    n71
  );


  not
  g253
  (
    n192,
    n49
  );


  buf
  g254
  (
    n170,
    n136
  );


  buf
  g255
  (
    n385,
    n46
  );


  not
  g256
  (
    n373,
    n76
  );


  not
  g257
  (
    n158,
    n48
  );


  not
  g258
  (
    n221,
    n94
  );


  buf
  g259
  (
    n325,
    n96
  );


  buf
  g260
  (
    n536,
    n64
  );


  buf
  g261
  (
    n202,
    n74
  );


  not
  g262
  (
    n476,
    n51
  );


  buf
  g263
  (
    n442,
    n114
  );


  not
  g264
  (
    n492,
    n99
  );


  not
  g265
  (
    n229,
    n76
  );


  buf
  g266
  (
    n456,
    n122
  );


  buf
  g267
  (
    n296,
    n98
  );


  not
  g268
  (
    n254,
    n33
  );


  not
  g269
  (
    n507,
    n82
  );


  buf
  g270
  (
    n403,
    n121
  );


  buf
  g271
  (
    n439,
    n99
  );


  buf
  g272
  (
    n205,
    n58
  );


  buf
  g273
  (
    n197,
    n62
  );


  buf
  g274
  (
    n288,
    n91
  );


  buf
  g275
  (
    n199,
    n50
  );


  buf
  g276
  (
    n386,
    n61
  );


  not
  g277
  (
    n462,
    n56
  );


  not
  g278
  (
    n374,
    n58
  );


  not
  g279
  (
    n488,
    n122
  );


  buf
  g280
  (
    n250,
    n80
  );


  not
  g281
  (
    n258,
    n92
  );


  not
  g282
  (
    n173,
    n55
  );


  not
  g283
  (
    n491,
    n46
  );


  not
  g284
  (
    n486,
    n113
  );


  not
  g285
  (
    n216,
    n108
  );


  not
  g286
  (
    n519,
    n60
  );


  not
  g287
  (
    n330,
    n78
  );


  not
  g288
  (
    n448,
    n109
  );


  buf
  g289
  (
    n563,
    n40
  );


  buf
  g290
  (
    n179,
    n103
  );


  buf
  g291
  (
    n480,
    n72
  );


  not
  g292
  (
    n225,
    n104
  );


  not
  g293
  (
    n546,
    n44
  );


  buf
  g294
  (
    n263,
    n100
  );


  buf
  g295
  (
    n298,
    n64
  );


  not
  g296
  (
    n530,
    n129
  );


  not
  g297
  (
    n466,
    n95
  );


  not
  g298
  (
    n525,
    n84
  );


  buf
  g299
  (
    n217,
    n87
  );


  buf
  g300
  (
    n398,
    n86
  );


  buf
  g301
  (
    n223,
    n90
  );


  not
  g302
  (
    n410,
    n122
  );


  buf
  g303
  (
    n554,
    n119
  );


  not
  g304
  (
    n210,
    n52
  );


  not
  g305
  (
    n469,
    n118
  );


  buf
  g306
  (
    n505,
    n93
  );


  buf
  g307
  (
    n164,
    n116
  );


  not
  g308
  (
    n240,
    n39
  );


  buf
  g309
  (
    n560,
    n80
  );


  buf
  g310
  (
    n532,
    n119
  );


  not
  g311
  (
    n342,
    n100
  );


  not
  g312
  (
    n309,
    n47
  );


  buf
  g313
  (
    n394,
    n95
  );


  buf
  g314
  (
    n245,
    n79
  );


  buf
  g315
  (
    n372,
    n116
  );


  buf
  g316
  (
    n440,
    n49
  );


  buf
  g317
  (
    n494,
    n43
  );


  buf
  g318
  (
    n431,
    n94
  );


  buf
  g319
  (
    n575,
    n65
  );


  buf
  g320
  (
    n472,
    n36
  );


  not
  g321
  (
    n239,
    n137
  );


  buf
  g322
  (
    n578,
    n127
  );


  buf
  g323
  (
    n433,
    n106
  );


  buf
  g324
  (
    n368,
    n117
  );


  buf
  g325
  (
    n351,
    n65
  );


  not
  g326
  (
    n286,
    n99
  );


  buf
  g327
  (
    n396,
    n59
  );


  buf
  g328
  (
    n304,
    n97
  );


  buf
  g329
  (
    n569,
    n34
  );


  not
  g330
  (
    n224,
    n135
  );


  buf
  g331
  (
    n552,
    n93
  );


  buf
  g332
  (
    n300,
    n126
  );


  buf
  g333
  (
    n485,
    n105
  );


  buf
  g334
  (
    n159,
    n39
  );


  not
  g335
  (
    n405,
    n44
  );


  buf
  g336
  (
    n487,
    n43
  );


  buf
  g337
  (
    n232,
    n73
  );


  not
  g338
  (
    n452,
    n61
  );


  not
  g339
  (
    n435,
    n66
  );


  not
  g340
  (
    n465,
    n128
  );


  buf
  g341
  (
    n432,
    n105
  );


  buf
  g342
  (
    n337,
    n110
  );


  buf
  g343
  (
    n358,
    n123
  );


  buf
  g344
  (
    n512,
    n91
  );


  buf
  g345
  (
    KeyWire_0_0,
    n102
  );


  buf
  g346
  (
    n383,
    n48
  );


  buf
  g347
  (
    n287,
    n138
  );


  buf
  g348
  (
    n260,
    n127
  );


  buf
  g349
  (
    n413,
    n85
  );


  not
  g350
  (
    n581,
    n125
  );


  buf
  g351
  (
    n355,
    n49
  );


  buf
  g352
  (
    n455,
    n37
  );


  not
  g353
  (
    n548,
    n49
  );


  not
  g354
  (
    n270,
    n57
  );


  buf
  g355
  (
    n167,
    n67
  );


  not
  g356
  (
    n363,
    n138
  );


  not
  g357
  (
    n155,
    n71
  );


  not
  g358
  (
    n176,
    n115
  );


  not
  g359
  (
    n561,
    n80
  );


  buf
  g360
  (
    n496,
    n72
  );


  not
  g361
  (
    n437,
    n101
  );


  buf
  g362
  (
    n318,
    n109
  );


  not
  g363
  (
    n294,
    n124
  );


  not
  g364
  (
    n391,
    n77
  );


  buf
  g365
  (
    n357,
    n104
  );


  buf
  g366
  (
    KeyWire_0_3,
    n91
  );


  not
  g367
  (
    n490,
    n35
  );


  not
  g368
  (
    n367,
    n126
  );


  buf
  g369
  (
    n378,
    n98
  );


  not
  g370
  (
    n427,
    n123
  );


  buf
  g371
  (
    n233,
    n104
  );


  buf
  g372
  (
    n582,
    n70
  );


  buf
  g373
  (
    n332,
    n80
  );


  buf
  g374
  (
    n506,
    n77
  );


  not
  g375
  (
    n446,
    n78
  );


  buf
  g376
  (
    KeyWire_0_4,
    n97
  );


  buf
  g377
  (
    n157,
    n71
  );


  buf
  g378
  (
    n269,
    n69
  );


  buf
  g379
  (
    n160,
    n106
  );


  not
  g380
  (
    n550,
    n40
  );


  buf
  g381
  (
    n213,
    n76
  );


  not
  g382
  (
    n206,
    n76
  );


  not
  g383
  (
    n384,
    n46
  );


  buf
  g384
  (
    n328,
    n105
  );


  not
  g385
  (
    n484,
    n120
  );


  not
  g386
  (
    n252,
    n83
  );


  not
  g387
  (
    n400,
    n33
  );


  buf
  g388
  (
    n542,
    n140
  );


  buf
  g389
  (
    n343,
    n65
  );


  buf
  g390
  (
    n231,
    n87
  );


  not
  g391
  (
    n584,
    n68
  );


  not
  g392
  (
    n334,
    n56
  );


  buf
  g393
  (
    n483,
    n57
  );


  not
  g394
  (
    n501,
    n92
  );


  buf
  g395
  (
    n235,
    n103
  );


  not
  g396
  (
    n547,
    n64
  );


  not
  g397
  (
    n500,
    n124
  );


  not
  g398
  (
    n562,
    n59
  );


  not
  g399
  (
    n163,
    n42
  );


  buf
  g400
  (
    n308,
    n132
  );


  not
  g401
  (
    n201,
    n83
  );


  buf
  g402
  (
    n282,
    n126
  );


  buf
  g403
  (
    n471,
    n39
  );


  buf
  g404
  (
    n212,
    n78
  );


  not
  g405
  (
    n207,
    n79
  );


  buf
  g406
  (
    n481,
    n55
  );


  not
  g407
  (
    n555,
    n118
  );


  not
  g408
  (
    n521,
    n84
  );


  buf
  g409
  (
    n283,
    n138
  );


  buf
  g410
  (
    n196,
    n111
  );


  buf
  g411
  (
    n255,
    n52
  );


  not
  g412
  (
    n573,
    n100
  );


  buf
  g413
  (
    n479,
    n59
  );


  buf
  g414
  (
    n579,
    n89
  );


  not
  g415
  (
    n539,
    n118
  );


  not
  g416
  (
    n460,
    n69
  );


  not
  g417
  (
    n425,
    n77
  );


  not
  g418
  (
    n195,
    n131
  );


  not
  g419
  (
    n382,
    n124
  );


  buf
  g420
  (
    n407,
    n96
  );


  buf
  g421
  (
    n502,
    n51
  );


  not
  g422
  (
    n516,
    n88
  );


  not
  g423
  (
    n580,
    n74
  );


  not
  g424
  (
    n388,
    n120
  );


  not
  g425
  (
    n570,
    n37
  );


  not
  g426
  (
    n447,
    n34
  );


  buf
  g427
  (
    n421,
    n61
  );


  buf
  g428
  (
    n243,
    n140
  );


  not
  g429
  (
    n272,
    n120
  );


  not
  g430
  (
    n185,
    n53
  );


  buf
  g431
  (
    n237,
    n74
  );


  buf
  g432
  (
    n341,
    n130
  );


  buf
  g433
  (
    n426,
    n133
  );


  not
  g434
  (
    n503,
    n45
  );


  buf
  g435
  (
    n215,
    n41
  );


  not
  g436
  (
    n242,
    n134
  );


  buf
  g437
  (
    n273,
    n93
  );


  buf
  g438
  (
    n533,
    n68
  );


  not
  g439
  (
    n321,
    n87
  );


  buf
  g440
  (
    n190,
    n44
  );


  not
  g441
  (
    n175,
    n120
  );


  not
  g442
  (
    n156,
    n110
  );


  buf
  g443
  (
    n226,
    n54
  );


  not
  g444
  (
    n379,
    n114
  );


  buf
  g445
  (
    n541,
    n61
  );


  not
  g446
  (
    n528,
    n42
  );


  buf
  g447
  (
    n333,
    n65
  );


  buf
  g448
  (
    n227,
    n55
  );


  buf
  g449
  (
    n558,
    n85
  );


  buf
  g450
  (
    n236,
    n133
  );


  not
  g451
  (
    n204,
    n59
  );


  buf
  g452
  (
    n376,
    n107
  );


  not
  g453
  (
    n514,
    n102
  );


  buf
  g454
  (
    n289,
    n63
  );


  buf
  g455
  (
    n222,
    n70
  );


  buf
  g456
  (
    n152,
    n121
  );


  not
  g457
  (
    n518,
    n45
  );


  buf
  g458
  (
    n436,
    n45
  );


  not
  g459
  (
    n559,
    n63
  );


  buf
  g460
  (
    n181,
    n79
  );


  buf
  g461
  (
    n529,
    n35
  );


  buf
  g462
  (
    n162,
    n115
  );


  buf
  g463
  (
    n564,
    n112
  );


  buf
  g464
  (
    n526,
    n81
  );


  not
  g465
  (
    n230,
    n75
  );


  buf
  g466
  (
    n557,
    n113
  );


  not
  g467
  (
    n419,
    n47
  );


  not
  g468
  (
    n262,
    n112
  );


  not
  g469
  (
    n265,
    n79
  );


  not
  g470
  (
    n317,
    n96
  );


  not
  g471
  (
    n417,
    n106
  );


  not
  g472
  (
    n416,
    n136
  );


  buf
  g473
  (
    n292,
    n62
  );


  buf
  g474
  (
    n543,
    n47
  );


  not
  g475
  (
    n348,
    n123
  );


  buf
  g476
  (
    n172,
    n96
  );


  buf
  g477
  (
    n571,
    n124
  );


  buf
  g478
  (
    n290,
    n117
  );


  not
  g479
  (
    n303,
    n101
  );


  not
  g480
  (
    n338,
    n60
  );


  not
  g481
  (
    n336,
    n97
  );


  not
  g482
  (
    n249,
    n88
  );


  not
  g483
  (
    n458,
    n58
  );


  not
  g484
  (
    n520,
    n88
  );


  not
  g485
  (
    n381,
    n82
  );


  buf
  g486
  (
    n568,
    n99
  );


  not
  g487
  (
    n393,
    n133
  );


  buf
  g488
  (
    n493,
    n129
  );


  not
  g489
  (
    n198,
    n131
  );


  not
  g490
  (
    n498,
    n102
  );


  buf
  g491
  (
    n454,
    n110
  );


  not
  g492
  (
    n404,
    n57
  );


  buf
  g493
  (
    n509,
    n109
  );


  not
  g494
  (
    n347,
    n69
  );


  not
  g495
  (
    n350,
    n92
  );


  buf
  g496
  (
    n522,
    n86
  );


  buf
  g497
  (
    n246,
    n70
  );


  buf
  g498
  (
    n537,
    n130
  );


  buf
  g499
  (
    n495,
    n52
  );


  buf
  g500
  (
    n473,
    n41
  );


  not
  g501
  (
    n401,
    n85
  );


  buf
  g502
  (
    n499,
    n82
  );


  buf
  g503
  (
    n468,
    n114
  );


  not
  g504
  (
    n534,
    n134
  );


  buf
  g505
  (
    n504,
    n54
  );


  buf
  g506
  (
    n397,
    n83
  );


  not
  g507
  (
    n186,
    n69
  );


  not
  g508
  (
    n353,
    n109
  );


  buf
  g509
  (
    n211,
    n70
  );


  buf
  g510
  (
    n305,
    n50
  );


  not
  g511
  (
    n307,
    n64
  );


  not
  g512
  (
    n361,
    n41
  );


  not
  g513
  (
    n275,
    n84
  );


  not
  g514
  (
    n438,
    n103
  );


  buf
  g515
  (
    n434,
    n35
  );


  not
  g516
  (
    n326,
    n102
  );


  not
  g517
  (
    n154,
    n93
  );


  buf
  g518
  (
    n445,
    n63
  );


  buf
  g519
  (
    n278,
    n86
  );


  not
  g520
  (
    n467,
    n34
  );


  not
  g521
  (
    n302,
    n111
  );


  not
  g522
  (
    n370,
    n83
  );


  buf
  g523
  (
    n453,
    n125
  );


  buf
  g524
  (
    n165,
    n40
  );


  not
  g525
  (
    n261,
    n47
  );


  not
  g526
  (
    n316,
    n38
  );


  buf
  g527
  (
    n414,
    n57
  );


  not
  g528
  (
    n257,
    n88
  );


  not
  g529
  (
    n344,
    n75
  );


  buf
  g530
  (
    n387,
    n139
  );


  not
  g531
  (
    n389,
    n81
  );


  not
  g532
  (
    n253,
    n139
  );


  not
  g533
  (
    n429,
    n43
  );


  not
  g534
  (
    n188,
    n44
  );


  not
  g535
  (
    n362,
    n68
  );


  not
  g536
  (
    n464,
    n136
  );


  not
  g537
  (
    n306,
    n135
  );


  not
  g538
  (
    n511,
    n116
  );


  not
  g539
  (
    n354,
    n128
  );


  not
  g540
  (
    n423,
    n112
  );


  buf
  g541
  (
    n311,
    n87
  );


  buf
  g542
  (
    n277,
    n73
  );


  not
  g543
  (
    n329,
    n135
  );


  buf
  g544
  (
    n449,
    n94
  );


  buf
  g545
  (
    n183,
    n39
  );


  not
  g546
  (
    n549,
    n138
  );


  not
  g547
  (
    n251,
    n91
  );


  not
  g548
  (
    n364,
    n50
  );


  not
  g549
  (
    n214,
    n67
  );


  not
  g550
  (
    n477,
    n119
  );


  buf
  g551
  (
    n327,
    n117
  );


  buf
  g552
  (
    n402,
    n131
  );


  xor
  g553
  (
    n600,
    n222,
    n162,
    n186,
    n160
  );


  or
  g554
  (
    n596,
    n169,
    n212,
    n223,
    n185
  );


  nand
  g555
  (
    n595,
    n167,
    n220,
    n164,
    n166
  );


  xor
  g556
  (
    n597,
    n156,
    n179,
    n210,
    n218
  );


  nand
  g557
  (
    n601,
    n201,
    n174,
    n182,
    n171
  );


  and
  g558
  (
    n593,
    n202,
    n177,
    n193,
    n163
  );


  or
  g559
  (
    n589,
    n197,
    n189,
    n204,
    n213
  );


  or
  g560
  (
    n598,
    n184,
    n208,
    n195,
    n209
  );


  nor
  g561
  (
    n594,
    n217,
    n176,
    n173,
    n219
  );


  xnor
  g562
  (
    n590,
    n194,
    n191,
    n157,
    n198
  );


  xnor
  g563
  (
    n587,
    n158,
    n206,
    n196,
    n161
  );


  and
  g564
  (
    n592,
    n155,
    n200,
    n203,
    n153
  );


  nand
  g565
  (
    n602,
    n221,
    n211,
    n183,
    n159
  );


  xor
  g566
  (
    n586,
    n165,
    n154,
    n188,
    n168
  );


  nor
  g567
  (
    n588,
    n199,
    n205,
    n181,
    n216
  );


  xnor
  g568
  (
    n599,
    n170,
    n172,
    n180,
    n187
  );


  and
  g569
  (
    n603,
    n207,
    n190,
    n214,
    n215
  );


  or
  g570
  (
    n591,
    n175,
    n178,
    n152,
    n192
  );


  or
  g571
  (
    n604,
    n592,
    n141,
    n143
  );


  nor
  g572
  (
    n609,
    n146,
    n586,
    n142,
    n144
  );


  nand
  g573
  (
    n605,
    n142,
    n588,
    n143
  );


  or
  g574
  (
    n611,
    n596,
    n595,
    n589,
    n144
  );


  or
  g575
  (
    n607,
    n143,
    n146,
    n142,
    n594
  );


  nand
  g576
  (
    n606,
    n591,
    n593,
    n145,
    n144
  );


  nor
  g577
  (
    n610,
    n590,
    n142,
    n146,
    n144
  );


  nand
  g578
  (
    n608,
    n587,
    n145
  );


  not
  g579
  (
    n612,
    n605
  );


  not
  g580
  (
    n613,
    n604
  );


  not
  g581
  (
    n616,
    n612
  );


  not
  g582
  (
    n614,
    n613
  );


  buf
  g583
  (
    n615,
    n613
  );


  not
  g584
  (
    n621,
    n612
  );


  buf
  g585
  (
    n618,
    n612
  );


  not
  g586
  (
    n617,
    n612
  );


  buf
  g587
  (
    n619,
    n613
  );


  buf
  g588
  (
    n620,
    n613
  );


  buf
  g589
  (
    n627,
    n619
  );


  not
  g590
  (
    n634,
    n148
  );


  not
  g591
  (
    n637,
    n32
  );


  buf
  g592
  (
    n624,
    n30
  );


  buf
  g593
  (
    n632,
    n614
  );


  buf
  g594
  (
    n639,
    n621
  );


  not
  g595
  (
    n649,
    n225
  );


  not
  g596
  (
    n622,
    n226
  );


  not
  g597
  (
    n623,
    n150
  );


  buf
  g598
  (
    n628,
    n618
  );


  not
  g599
  (
    n652,
    n614
  );


  buf
  g600
  (
    n631,
    n617
  );


  not
  g601
  (
    n650,
    n147
  );


  buf
  g602
  (
    n629,
    n615
  );


  buf
  g603
  (
    n641,
    n615
  );


  buf
  g604
  (
    n625,
    n227
  );


  buf
  g605
  (
    n644,
    n148
  );


  buf
  g606
  (
    n646,
    n620
  );


  nand
  g607
  (
    n638,
    n31,
    n32,
    n618
  );


  xnor
  g608
  (
    n647,
    n607,
    n620,
    n610,
    n614
  );


  or
  g609
  (
    n651,
    n147,
    n619,
    n32
  );


  and
  g610
  (
    n640,
    n619,
    n617,
    n31,
    n148
  );


  xnor
  g611
  (
    n643,
    n609,
    n224,
    n150,
    n228
  );


  xnor
  g612
  (
    n645,
    n597,
    n147,
    n618,
    n232
  );


  nor
  g613
  (
    n633,
    n31,
    n148,
    n615
  );


  nand
  g614
  (
    n648,
    n617,
    n617,
    n620,
    n149
  );


  xor
  g615
  (
    n635,
    n231,
    n611,
    n620,
    n621
  );


  and
  g616
  (
    n642,
    n233,
    n606,
    n616,
    n150
  );


  xor
  g617
  (
    n630,
    n31,
    n149,
    n146,
    n147
  );


  nor
  g618
  (
    n626,
    n621,
    n614,
    n616,
    n149
  );


  nand
  g619
  (
    n636,
    n618,
    n229,
    n608,
    n230
  );


  nand
  g620
  (
    n653,
    n621,
    n149,
    n616
  );


  not
  g621
  (
    n669,
    n650
  );


  not
  g622
  (
    n654,
    n629
  );


  buf
  g623
  (
    n679,
    n640
  );


  buf
  g624
  (
    n673,
    n635
  );


  not
  g625
  (
    n697,
    n622
  );


  buf
  g626
  (
    n683,
    n643
  );


  buf
  g627
  (
    n662,
    n649
  );


  not
  g628
  (
    n698,
    n625
  );


  not
  g629
  (
    n708,
    n634
  );


  not
  g630
  (
    n699,
    n643
  );


  buf
  g631
  (
    n688,
    n624
  );


  buf
  g632
  (
    n684,
    n636
  );


  not
  g633
  (
    n674,
    n644
  );


  buf
  g634
  (
    n657,
    n624
  );


  not
  g635
  (
    n676,
    n641
  );


  buf
  g636
  (
    n691,
    n640
  );


  not
  g637
  (
    n671,
    n647
  );


  not
  g638
  (
    n686,
    n628
  );


  not
  g639
  (
    n678,
    n648
  );


  buf
  g640
  (
    n656,
    n622
  );


  not
  g641
  (
    n682,
    n647
  );


  not
  g642
  (
    n705,
    n642
  );


  nand
  g643
  (
    n670,
    n622,
    n646
  );


  xnor
  g644
  (
    KeyWire_0_11,
    n642,
    n639,
    n649
  );


  xor
  g645
  (
    n681,
    n625,
    n638,
    n623
  );


  and
  g646
  (
    n692,
    n645,
    n630
  );


  nor
  g647
  (
    n696,
    n631,
    n622,
    n623
  );


  xnor
  g648
  (
    n703,
    n650,
    n647,
    n632
  );


  xnor
  g649
  (
    n664,
    n627,
    n629,
    n637
  );


  xnor
  g650
  (
    n693,
    n625,
    n645,
    n639
  );


  nor
  g651
  (
    n701,
    n646,
    n641,
    n647
  );


  nand
  g652
  (
    n680,
    n626,
    n645,
    n634
  );


  xor
  g653
  (
    n702,
    n627,
    n630,
    n631
  );


  nand
  g654
  (
    n706,
    n627,
    n646,
    n649
  );


  xor
  g655
  (
    n685,
    n648,
    n643,
    n651
  );


  or
  g656
  (
    n660,
    n633,
    n627,
    n630
  );


  nor
  g657
  (
    n694,
    n623,
    n641,
    n637
  );


  nor
  g658
  (
    n668,
    n640,
    n631,
    n646
  );


  nand
  g659
  (
    n690,
    n640,
    n650,
    n624
  );


  or
  g660
  (
    n689,
    n642,
    n626,
    n636
  );


  xnor
  g661
  (
    n655,
    n638,
    n633
  );


  xor
  g662
  (
    n707,
    n635,
    n644,
    n651
  );


  and
  g663
  (
    n663,
    n624,
    n626,
    n638
  );


  nand
  g664
  (
    n677,
    n644,
    n634,
    n651
  );


  xor
  g665
  (
    n672,
    n629,
    n636,
    n635
  );


  and
  g666
  (
    KeyWire_0_10,
    n639,
    n628
  );


  and
  g667
  (
    n665,
    n629,
    n634,
    n648
  );


  nand
  g668
  (
    n700,
    n642,
    n639,
    n631
  );


  or
  g669
  (
    n658,
    n633,
    n632,
    n644
  );


  and
  g670
  (
    n695,
    n637,
    n649,
    n632
  );


  or
  g671
  (
    n659,
    n638,
    n623,
    n628
  );


  nor
  g672
  (
    n704,
    n650,
    n635,
    n641
  );


  xor
  g673
  (
    n687,
    n626,
    n643,
    n636
  );


  xor
  g674
  (
    n667,
    n632,
    n637,
    n645
  );


  or
  g675
  (
    n675,
    n648,
    n625,
    n651
  );


  buf
  g676
  (
    n709,
    n656
  );


  not
  g677
  (
    n711,
    n654
  );


  not
  g678
  (
    n710,
    n657
  );


  buf
  g679
  (
    n712,
    n655
  );


  not
  g680
  (
    n723,
    n709
  );


  buf
  g681
  (
    n716,
    n709
  );


  buf
  g682
  (
    n728,
    n711
  );


  buf
  g683
  (
    n721,
    n709
  );


  not
  g684
  (
    n714,
    n709
  );


  buf
  g685
  (
    n719,
    n711
  );


  buf
  g686
  (
    n722,
    n712
  );


  not
  g687
  (
    n727,
    n710
  );


  not
  g688
  (
    n717,
    n712
  );


  buf
  g689
  (
    n718,
    n712
  );


  buf
  g690
  (
    n715,
    n710
  );


  not
  g691
  (
    n726,
    n711
  );


  not
  g692
  (
    n720,
    n710
  );


  buf
  g693
  (
    n713,
    n711
  );


  buf
  g694
  (
    n724,
    n712
  );


  buf
  g695
  (
    n725,
    n710
  );


  or
  g696
  (
    n735,
    n675,
    n727,
    n714,
    n245
  );


  and
  g697
  (
    n737,
    n686,
    n664,
    n720,
    n728
  );


  nor
  g698
  (
    n741,
    n728,
    n684,
    n683,
    n249
  );


  xor
  g699
  (
    n744,
    n723,
    n676,
    n695,
    n693
  );


  xor
  g700
  (
    n734,
    n724,
    n680,
    n725,
    n238
  );


  xnor
  g701
  (
    n739,
    n726,
    n678,
    n719,
    n660
  );


  nor
  g702
  (
    n743,
    n679,
    n718,
    n244,
    n671
  );


  nand
  g703
  (
    n731,
    n692,
    n722,
    n235,
    n728
  );


  nor
  g704
  (
    n736,
    n674,
    n243,
    n687,
    n236
  );


  and
  g705
  (
    n748,
    n682,
    n728,
    n713,
    n669
  );


  xnor
  g706
  (
    n738,
    n662,
    n688,
    n670,
    n239
  );


  xnor
  g707
  (
    n733,
    n667,
    n247,
    n241,
    n237
  );


  and
  g708
  (
    n729,
    n727,
    n727,
    n663,
    n673
  );


  and
  g709
  (
    n730,
    n716,
    n248,
    n726,
    n721
  );


  and
  g710
  (
    n745,
    n725,
    n668,
    n661,
    n658
  );


  xor
  g711
  (
    n742,
    n234,
    n694,
    n685,
    n691
  );


  xnor
  g712
  (
    n740,
    n677,
    n242,
    n666,
    n681
  );


  nand
  g713
  (
    n732,
    n727,
    n696,
    n690,
    n697
  );


  and
  g714
  (
    n746,
    n659,
    n689,
    n715,
    n717
  );


  xor
  g715
  (
    n747,
    n246,
    n240,
    n665,
    n672
  );


  not
  g716
  (
    n750,
    n747
  );


  not
  g717
  (
    n749,
    n748
  );


  buf
  g718
  (
    n755,
    n749
  );


  not
  g719
  (
    n754,
    n749
  );


  not
  g720
  (
    n753,
    n750
  );


  buf
  g721
  (
    n752,
    n250
  );


  buf
  g722
  (
    n751,
    n749
  );


  not
  g723
  (
    n758,
    n751
  );


  buf
  g724
  (
    n757,
    n752
  );


  buf
  g725
  (
    n756,
    n753
  );


  not
  g726
  (
    n759,
    n752
  );


  not
  g727
  (
    n766,
    n262
  );


  not
  g728
  (
    n772,
    n756
  );


  xor
  g729
  (
    n760,
    n255,
    n750
  );


  or
  g730
  (
    n769,
    n757,
    n702,
    n603,
    n267
  );


  nand
  g731
  (
    KeyWire_0_14,
    n759,
    n600,
    n251,
    n252
  );


  and
  g732
  (
    n771,
    n264,
    n759,
    n256,
    n758
  );


  xor
  g733
  (
    n770,
    n258,
    n757,
    n759,
    n652
  );


  nand
  g734
  (
    n767,
    n700,
    n652,
    n750,
    n261
  );


  xor
  g735
  (
    n773,
    n704,
    n756,
    n758
  );


  or
  g736
  (
    n768,
    n703,
    n759,
    n652,
    n599
  );


  and
  g737
  (
    n761,
    n653,
    n259,
    n601,
    n699
  );


  xor
  g738
  (
    n775,
    n263,
    n698,
    n757,
    n602
  );


  nand
  g739
  (
    n774,
    n652,
    n653,
    n253,
    n750
  );


  or
  g740
  (
    n765,
    n266,
    n757,
    n257,
    n701
  );


  xor
  g741
  (
    n763,
    n653,
    n758,
    n260,
    n756
  );


  or
  g742
  (
    n764,
    n598,
    n758,
    n265,
    n254
  );


  buf
  g743
  (
    n791,
    n773
  );


  buf
  g744
  (
    n789,
    n754
  );


  not
  g745
  (
    n831,
    n772
  );


  not
  g746
  (
    n832,
    n275
  );


  not
  g747
  (
    n827,
    n771
  );


  not
  g748
  (
    n784,
    n774
  );


  not
  g749
  (
    n787,
    n761
  );


  not
  g750
  (
    n814,
    n764
  );


  buf
  g751
  (
    n810,
    n771
  );


  buf
  g752
  (
    n822,
    n766
  );


  buf
  g753
  (
    n786,
    n281
  );


  not
  g754
  (
    n777,
    n273
  );


  not
  g755
  (
    n798,
    n774
  );


  buf
  g756
  (
    n819,
    n764
  );


  buf
  g757
  (
    n839,
    n770
  );


  not
  g758
  (
    n817,
    n755
  );


  not
  g759
  (
    n779,
    n768
  );


  not
  g760
  (
    n824,
    n283
  );


  buf
  g761
  (
    n776,
    n765
  );


  not
  g762
  (
    n838,
    n754
  );


  not
  g763
  (
    n793,
    n774
  );


  not
  g764
  (
    n830,
    n753
  );


  buf
  g765
  (
    n836,
    n286
  );


  buf
  g766
  (
    n804,
    n769
  );


  buf
  g767
  (
    n781,
    n754
  );


  not
  g768
  (
    n790,
    n770
  );


  not
  g769
  (
    n807,
    n767
  );


  buf
  g770
  (
    n828,
    n768
  );


  not
  g771
  (
    n783,
    n274
  );


  not
  g772
  (
    n809,
    n770
  );


  not
  g773
  (
    n801,
    n280
  );


  not
  g774
  (
    n820,
    n768
  );


  buf
  g775
  (
    n797,
    n767
  );


  not
  g776
  (
    n825,
    n285
  );


  buf
  g777
  (
    n813,
    n769
  );


  buf
  g778
  (
    n803,
    n271
  );


  not
  g779
  (
    n834,
    n765
  );


  buf
  g780
  (
    n808,
    n772
  );


  buf
  g781
  (
    n835,
    n753
  );


  buf
  g782
  (
    n821,
    n282
  );


  buf
  g783
  (
    n785,
    n761
  );


  not
  g784
  (
    n826,
    n284
  );


  buf
  g785
  (
    n833,
    n269
  );


  not
  g786
  (
    n823,
    n763
  );


  buf
  g787
  (
    n815,
    n763
  );


  buf
  g788
  (
    n837,
    n766
  );


  buf
  g789
  (
    n799,
    n288
  );


  buf
  g790
  (
    n816,
    n762
  );


  not
  g791
  (
    n794,
    n773
  );


  buf
  g792
  (
    n818,
    n763
  );


  not
  g793
  (
    n795,
    n764
  );


  not
  g794
  (
    n800,
    n772
  );


  not
  g795
  (
    n805,
    n771
  );


  nand
  g796
  (
    n806,
    n774,
    n773,
    n775
  );


  nand
  g797
  (
    n802,
    n766,
    n763,
    n761,
    n771
  );


  nand
  g798
  (
    n780,
    n279,
    n760,
    n755,
    n268
  );


  nor
  g799
  (
    n782,
    n769,
    n760,
    n775,
    n762
  );


  nand
  g800
  (
    n811,
    n767,
    n762,
    n270,
    n769
  );


  xor
  g801
  (
    n788,
    n765,
    n755,
    n773,
    n277
  );


  and
  g802
  (
    n796,
    n760,
    n772,
    n761,
    n753
  );


  xor
  g803
  (
    n829,
    n768,
    n775,
    n272,
    n278
  );


  or
  g804
  (
    n792,
    n762,
    n760,
    n767,
    n765
  );


  nand
  g805
  (
    n812,
    n287,
    n764,
    n755,
    n766
  );


  xor
  g806
  (
    n778,
    n754,
    n770,
    n775,
    n276
  );


  buf
  g807
  (
    n879,
    n787
  );


  not
  g808
  (
    n850,
    n793
  );


  buf
  g809
  (
    n842,
    n788
  );


  not
  g810
  (
    n889,
    n791
  );


  not
  g811
  (
    n863,
    n784
  );


  not
  g812
  (
    n853,
    n786
  );


  not
  g813
  (
    n887,
    n793
  );


  not
  g814
  (
    n877,
    n784
  );


  buf
  g815
  (
    n880,
    n783
  );


  not
  g816
  (
    n847,
    n785
  );


  buf
  g817
  (
    n876,
    n789
  );


  not
  g818
  (
    n845,
    n790
  );


  not
  g819
  (
    n854,
    n782
  );


  buf
  g820
  (
    n872,
    n776
  );


  buf
  g821
  (
    n884,
    n782
  );


  not
  g822
  (
    n883,
    n791
  );


  buf
  g823
  (
    n897,
    n786
  );


  not
  g824
  (
    n893,
    n780
  );


  not
  g825
  (
    n894,
    n782
  );


  buf
  g826
  (
    n873,
    n784
  );


  not
  g827
  (
    n857,
    n784
  );


  buf
  g828
  (
    n866,
    n792
  );


  buf
  g829
  (
    n888,
    n787
  );


  buf
  g830
  (
    n844,
    n785
  );


  not
  g831
  (
    n890,
    n783
  );


  not
  g832
  (
    n849,
    n781
  );


  not
  g833
  (
    n869,
    n790
  );


  not
  g834
  (
    n841,
    n782
  );


  buf
  g835
  (
    n867,
    n789
  );


  buf
  g836
  (
    n899,
    n792
  );


  not
  g837
  (
    n871,
    n790
  );


  not
  g838
  (
    n862,
    n787
  );


  not
  g839
  (
    n852,
    n780
  );


  buf
  g840
  (
    n878,
    n792
  );


  buf
  g841
  (
    n840,
    n789
  );


  not
  g842
  (
    n875,
    n781
  );


  buf
  g843
  (
    n856,
    n791
  );


  not
  g844
  (
    n865,
    n783
  );


  not
  g845
  (
    KeyWire_0_8,
    n793
  );


  buf
  g846
  (
    n851,
    n790
  );


  not
  g847
  (
    n860,
    n793
  );


  buf
  g848
  (
    n859,
    n786
  );


  not
  g849
  (
    n896,
    n788
  );


  not
  g850
  (
    n895,
    n778
  );


  buf
  g851
  (
    n846,
    n780
  );


  buf
  g852
  (
    n885,
    n792
  );


  buf
  g853
  (
    n858,
    n783
  );


  buf
  g854
  (
    n891,
    n779
  );


  not
  g855
  (
    n843,
    n785
  );


  buf
  g856
  (
    n882,
    n787
  );


  not
  g857
  (
    n864,
    n791
  );


  buf
  g858
  (
    n881,
    n785
  );


  not
  g859
  (
    n886,
    n780
  );


  not
  g860
  (
    n868,
    n788
  );


  not
  g861
  (
    n870,
    n781
  );


  buf
  g862
  (
    n848,
    n786
  );


  buf
  g863
  (
    n898,
    n781
  );


  not
  g864
  (
    n861,
    n788
  );


  buf
  g865
  (
    n855,
    n777
  );


  not
  g866
  (
    n874,
    n789
  );


  not
  g867
  (
    n1125,
    n895
  );


  not
  g868
  (
    n1070,
    n882
  );


  buf
  g869
  (
    n942,
    n853
  );


  buf
  g870
  (
    n1049,
    n871
  );


  not
  g871
  (
    n1055,
    n862
  );


  not
  g872
  (
    n975,
    n874
  );


  buf
  g873
  (
    n956,
    n847
  );


  not
  g874
  (
    n977,
    n841
  );


  not
  g875
  (
    n900,
    n855
  );


  not
  g876
  (
    n976,
    n840
  );


  buf
  g877
  (
    n1040,
    n851
  );


  buf
  g878
  (
    n924,
    n873
  );


  buf
  g879
  (
    n1091,
    n887
  );


  buf
  g880
  (
    n967,
    n865
  );


  not
  g881
  (
    n1024,
    n875
  );


  not
  g882
  (
    n991,
    n862
  );


  buf
  g883
  (
    n911,
    n878
  );


  not
  g884
  (
    n1135,
    n886
  );


  buf
  g885
  (
    n902,
    n872
  );


  buf
  g886
  (
    n1058,
    n855
  );


  buf
  g887
  (
    n1011,
    n868
  );


  not
  g888
  (
    n1128,
    n881
  );


  buf
  g889
  (
    n901,
    n875
  );


  not
  g890
  (
    n1065,
    n868
  );


  not
  g891
  (
    n908,
    n874
  );


  not
  g892
  (
    n1073,
    n857
  );


  buf
  g893
  (
    n1068,
    n858
  );


  not
  g894
  (
    n928,
    n881
  );


  not
  g895
  (
    n912,
    n898
  );


  not
  g896
  (
    n966,
    n858
  );


  buf
  g897
  (
    n962,
    n846
  );


  buf
  g898
  (
    n1111,
    n883
  );


  buf
  g899
  (
    n907,
    n891
  );


  buf
  g900
  (
    n1021,
    n893
  );


  buf
  g901
  (
    n1114,
    n861
  );


  buf
  g902
  (
    n1094,
    n856
  );


  not
  g903
  (
    n1134,
    n895
  );


  not
  g904
  (
    n1052,
    n883
  );


  not
  g905
  (
    n1069,
    n865
  );


  buf
  g906
  (
    n1085,
    n890
  );


  buf
  g907
  (
    n905,
    n849
  );


  not
  g908
  (
    n981,
    n896
  );


  not
  g909
  (
    n936,
    n854
  );


  not
  g910
  (
    n1139,
    n878
  );


  buf
  g911
  (
    n1131,
    n851
  );


  not
  g912
  (
    n973,
    n854
  );


  not
  g913
  (
    n910,
    n880
  );


  not
  g914
  (
    n937,
    n860
  );


  buf
  g915
  (
    n1014,
    n897
  );


  not
  g916
  (
    n1121,
    n899
  );


  buf
  g917
  (
    n1099,
    n846
  );


  not
  g918
  (
    n1130,
    n880
  );


  not
  g919
  (
    n1109,
    n874
  );


  not
  g920
  (
    n1071,
    n875
  );


  not
  g921
  (
    n926,
    n885
  );


  not
  g922
  (
    n1084,
    n882
  );


  buf
  g923
  (
    n959,
    n856
  );


  buf
  g924
  (
    n1115,
    n849
  );


  buf
  g925
  (
    n1098,
    n840
  );


  buf
  g926
  (
    n1132,
    n891
  );


  not
  g927
  (
    n1087,
    n884
  );


  buf
  g928
  (
    n1063,
    n897
  );


  not
  g929
  (
    n992,
    n855
  );


  not
  g930
  (
    n1056,
    n863
  );


  not
  g931
  (
    n927,
    n877
  );


  not
  g932
  (
    n929,
    n883
  );


  buf
  g933
  (
    n906,
    n869
  );


  buf
  g934
  (
    n1017,
    n850
  );


  not
  g935
  (
    n1015,
    n846
  );


  buf
  g936
  (
    n1077,
    n888
  );


  not
  g937
  (
    n1076,
    n874
  );


  buf
  g938
  (
    n957,
    n844
  );


  buf
  g939
  (
    n918,
    n892
  );


  buf
  g940
  (
    n999,
    n878
  );


  buf
  g941
  (
    n1127,
    n894
  );


  not
  g942
  (
    n1036,
    n871
  );


  buf
  g943
  (
    n1006,
    n867
  );


  buf
  g944
  (
    n913,
    n888
  );


  buf
  g945
  (
    n1054,
    n842
  );


  not
  g946
  (
    n1030,
    n871
  );


  buf
  g947
  (
    n1074,
    n859
  );


  buf
  g948
  (
    n1003,
    n858
  );


  buf
  g949
  (
    n1051,
    n843
  );


  not
  g950
  (
    n1007,
    n853
  );


  buf
  g951
  (
    n909,
    n292
  );


  not
  g952
  (
    n1045,
    n886
  );


  not
  g953
  (
    n1105,
    n867
  );


  not
  g954
  (
    n994,
    n853
  );


  not
  g955
  (
    n948,
    n867
  );


  buf
  g956
  (
    n1062,
    n842
  );


  buf
  g957
  (
    n1061,
    n842
  );


  buf
  g958
  (
    n922,
    n290
  );


  not
  g959
  (
    n1082,
    n861
  );


  not
  g960
  (
    n1057,
    n846
  );


  buf
  g961
  (
    n1008,
    n863
  );


  not
  g962
  (
    n1079,
    n847
  );


  not
  g963
  (
    n982,
    n896
  );


  not
  g964
  (
    n960,
    n847
  );


  buf
  g965
  (
    n938,
    n879
  );


  not
  g966
  (
    n1112,
    n877
  );


  buf
  g967
  (
    n947,
    n877
  );


  not
  g968
  (
    n904,
    n891
  );


  buf
  g969
  (
    n955,
    n879
  );


  not
  g970
  (
    n1039,
    n864
  );


  buf
  g971
  (
    n958,
    n857
  );


  not
  g972
  (
    n1103,
    n860
  );


  buf
  g973
  (
    n1089,
    n894
  );


  buf
  g974
  (
    n1022,
    n872
  );


  not
  g975
  (
    n1119,
    n876
  );


  buf
  g976
  (
    n1026,
    n875
  );


  not
  g977
  (
    n954,
    n893
  );


  not
  g978
  (
    n1032,
    n873
  );


  not
  g979
  (
    n1004,
    n885
  );


  buf
  g980
  (
    n985,
    n868
  );


  buf
  g981
  (
    n1047,
    n843
  );


  not
  g982
  (
    n978,
    n889
  );


  buf
  g983
  (
    n1104,
    n841
  );


  not
  g984
  (
    n1133,
    n890
  );


  not
  g985
  (
    n1137,
    n870
  );


  not
  g986
  (
    n1031,
    n856
  );


  buf
  g987
  (
    n1050,
    n849
  );


  buf
  g988
  (
    n1023,
    n848
  );


  not
  g989
  (
    n1046,
    n848
  );


  buf
  g990
  (
    n903,
    n289
  );


  buf
  g991
  (
    n965,
    n852
  );


  buf
  g992
  (
    n1092,
    n854
  );


  buf
  g993
  (
    n1126,
    n887
  );


  not
  g994
  (
    n1093,
    n880
  );


  buf
  g995
  (
    n915,
    n866
  );


  buf
  g996
  (
    n939,
    n892
  );


  not
  g997
  (
    n963,
    n850
  );


  not
  g998
  (
    n1038,
    n843
  );


  not
  g999
  (
    n933,
    n845
  );


  not
  g1000
  (
    n1122,
    n881
  );


  not
  g1001
  (
    n1083,
    n879
  );


  buf
  g1002
  (
    n993,
    n879
  );


  buf
  g1003
  (
    n951,
    n864
  );


  not
  g1004
  (
    n1095,
    n293
  );


  not
  g1005
  (
    n974,
    n860
  );


  not
  g1006
  (
    n1113,
    n887
  );


  not
  g1007
  (
    n1090,
    n889
  );


  not
  g1008
  (
    n997,
    n892
  );


  not
  g1009
  (
    n1086,
    n882
  );


  buf
  g1010
  (
    n1066,
    n876
  );


  not
  g1011
  (
    n931,
    n851
  );


  not
  g1012
  (
    n1000,
    n841
  );


  buf
  g1013
  (
    n1012,
    n876
  );


  buf
  g1014
  (
    n1059,
    n852
  );


  buf
  g1015
  (
    n972,
    n854
  );


  buf
  g1016
  (
    n1097,
    n890
  );


  not
  g1017
  (
    n920,
    n863
  );


  not
  g1018
  (
    n1019,
    n878
  );


  buf
  g1019
  (
    n968,
    n882
  );


  not
  g1020
  (
    n953,
    n899
  );


  not
  g1021
  (
    n914,
    n841
  );


  buf
  g1022
  (
    n916,
    n898
  );


  buf
  g1023
  (
    n950,
    n859
  );


  buf
  g1024
  (
    n1108,
    n873
  );


  buf
  g1025
  (
    n1088,
    n862
  );


  buf
  g1026
  (
    n1067,
    n899
  );


  not
  g1027
  (
    n945,
    n845
  );


  buf
  g1028
  (
    n1118,
    n857
  );


  not
  g1029
  (
    n1060,
    n867
  );


  not
  g1030
  (
    n1025,
    n844
  );


  not
  g1031
  (
    n1009,
    n894
  );


  buf
  g1032
  (
    n1001,
    n893
  );


  not
  g1033
  (
    n961,
    n843
  );


  buf
  g1034
  (
    n1064,
    n852
  );


  not
  g1035
  (
    n946,
    n848
  );


  buf
  g1036
  (
    n1081,
    n291
  );


  buf
  g1037
  (
    n935,
    n899
  );


  not
  g1038
  (
    n1107,
    n884
  );


  not
  g1039
  (
    n1029,
    n872
  );


  buf
  g1040
  (
    n984,
    n840
  );


  not
  g1041
  (
    n995,
    n844
  );


  not
  g1042
  (
    n1037,
    n892
  );


  buf
  g1043
  (
    n990,
    n898
  );


  buf
  g1044
  (
    n1048,
    n866
  );


  not
  g1045
  (
    n941,
    n853
  );


  not
  g1046
  (
    n998,
    n884
  );


  buf
  g1047
  (
    n1106,
    n849
  );


  buf
  g1048
  (
    n971,
    n888
  );


  buf
  g1049
  (
    n923,
    n860
  );


  buf
  g1050
  (
    n952,
    n866
  );


  buf
  g1051
  (
    n1080,
    n861
  );


  buf
  g1052
  (
    n1041,
    n859
  );


  buf
  g1053
  (
    n940,
    n856
  );


  not
  g1054
  (
    n979,
    n872
  );


  not
  g1055
  (
    n930,
    n898
  );


  buf
  g1056
  (
    n921,
    n895
  );


  buf
  g1057
  (
    n1005,
    n869
  );


  not
  g1058
  (
    n1124,
    n868
  );


  not
  g1059
  (
    n1075,
    n897
  );


  buf
  g1060
  (
    n943,
    n894
  );


  not
  g1061
  (
    n919,
    n889
  );


  buf
  g1062
  (
    n964,
    n865
  );


  not
  g1063
  (
    n1078,
    n869
  );


  buf
  g1064
  (
    n986,
    n895
  );


  not
  g1065
  (
    n1013,
    n870
  );


  not
  g1066
  (
    n980,
    n885
  );


  not
  g1067
  (
    n1018,
    n847
  );


  buf
  g1068
  (
    n949,
    n851
  );


  buf
  g1069
  (
    n1123,
    n850
  );


  not
  g1070
  (
    n1096,
    n864
  );


  not
  g1071
  (
    n1110,
    n884
  );


  not
  g1072
  (
    n1034,
    n896
  );


  buf
  g1073
  (
    n1129,
    n896
  );


  not
  g1074
  (
    n944,
    n871
  );


  buf
  g1075
  (
    n983,
    n840
  );


  buf
  g1076
  (
    n970,
    n865
  );


  buf
  g1077
  (
    n1027,
    n880
  );


  buf
  g1078
  (
    n1116,
    n862
  );


  buf
  g1079
  (
    n1042,
    n881
  );


  not
  g1080
  (
    n1136,
    n864
  );


  buf
  g1081
  (
    n934,
    n889
  );


  not
  g1082
  (
    n987,
    n869
  );


  buf
  g1083
  (
    n1044,
    n842
  );


  buf
  g1084
  (
    n932,
    n850
  );


  buf
  g1085
  (
    n917,
    n885
  );


  not
  g1086
  (
    n1020,
    n858
  );


  not
  g1087
  (
    n1138,
    n857
  );


  buf
  g1088
  (
    n1043,
    n852
  );


  buf
  g1089
  (
    n988,
    n863
  );


  buf
  g1090
  (
    n1102,
    n845
  );


  buf
  g1091
  (
    n925,
    n890
  );


  buf
  g1092
  (
    n989,
    n861
  );


  buf
  g1093
  (
    n1117,
    n876
  );


  buf
  g1094
  (
    n1101,
    n883
  );


  buf
  g1095
  (
    n1035,
    n870
  );


  buf
  g1096
  (
    n1053,
    n866
  );


  not
  g1097
  (
    n1033,
    n893
  );


  buf
  g1098
  (
    n1120,
    n886
  );


  buf
  g1099
  (
    n1028,
    n859
  );


  not
  g1100
  (
    n1016,
    n886
  );


  buf
  g1101
  (
    n1100,
    n891
  );


  not
  g1102
  (
    n1072,
    n848
  );


  not
  g1103
  (
    n969,
    n870
  );


  not
  g1104
  (
    n996,
    n855
  );


  and
  g1105
  (
    n1002,
    n877,
    n845,
    n887
  );


  nor
  g1106
  (
    n1010,
    n873,
    n897,
    n844,
    n888
  );


  not
  g1107
  (
    n1695,
    n1096
  );


  not
  g1108
  (
    n1517,
    n1091
  );


  buf
  g1109
  (
    n1722,
    n921
  );


  buf
  g1110
  (
    n1373,
    n817
  );


  buf
  g1111
  (
    n1582,
    n814
  );


  buf
  g1112
  (
    n1151,
    n1035
  );


  buf
  g1113
  (
    n1554,
    n931
  );


  buf
  g1114
  (
    n1666,
    n1025
  );


  buf
  g1115
  (
    n1306,
    n1032
  );


  not
  g1116
  (
    n1661,
    n1011
  );


  not
  g1117
  (
    n1431,
    n929
  );


  buf
  g1118
  (
    n1522,
    n834
  );


  buf
  g1119
  (
    n1273,
    n1002
  );


  buf
  g1120
  (
    n1312,
    n1048
  );


  buf
  g1121
  (
    n1544,
    n960
  );


  not
  g1122
  (
    n1552,
    n969
  );


  buf
  g1123
  (
    n1725,
    n1111
  );


  not
  g1124
  (
    n1732,
    n1008
  );


  not
  g1125
  (
    n1399,
    n1015
  );


  buf
  g1126
  (
    n1527,
    n978
  );


  buf
  g1127
  (
    n1147,
    n1027
  );


  buf
  g1128
  (
    n1228,
    n296
  );


  buf
  g1129
  (
    n1409,
    n799
  );


  not
  g1130
  (
    n1202,
    n794
  );


  buf
  g1131
  (
    n1503,
    n801
  );


  buf
  g1132
  (
    n1618,
    n813
  );


  buf
  g1133
  (
    n1420,
    n1080
  );


  not
  g1134
  (
    n1516,
    n1104
  );


  not
  g1135
  (
    n1324,
    n1133
  );


  not
  g1136
  (
    n1304,
    n1006
  );


  not
  g1137
  (
    n1419,
    n1031
  );


  buf
  g1138
  (
    n1177,
    n1057
  );


  buf
  g1139
  (
    n1737,
    n1064
  );


  buf
  g1140
  (
    n1193,
    n1100
  );


  not
  g1141
  (
    n1238,
    n1012
  );


  buf
  g1142
  (
    n1677,
    n1087
  );


  buf
  g1143
  (
    n1691,
    n1083
  );


  buf
  g1144
  (
    n1640,
    n1063
  );


  not
  g1145
  (
    n1162,
    n985
  );


  not
  g1146
  (
    n1268,
    n1094
  );


  buf
  g1147
  (
    n1621,
    n1040
  );


  not
  g1148
  (
    n1693,
    n963
  );


  buf
  g1149
  (
    n1458,
    n1042
  );


  not
  g1150
  (
    n1510,
    n1120
  );


  not
  g1151
  (
    n1519,
    n1097
  );


  not
  g1152
  (
    n1371,
    n834
  );


  buf
  g1153
  (
    n1543,
    n1109
  );


  buf
  g1154
  (
    n1298,
    n1022
  );


  not
  g1155
  (
    n1674,
    n1044
  );


  not
  g1156
  (
    n1495,
    n1040
  );


  buf
  g1157
  (
    n1612,
    n1026
  );


  buf
  g1158
  (
    n1616,
    n1130
  );


  not
  g1159
  (
    n1351,
    n968
  );


  not
  g1160
  (
    n1140,
    n1007
  );


  buf
  g1161
  (
    n1289,
    n1045
  );


  not
  g1162
  (
    n1319,
    n837
  );


  not
  g1163
  (
    KeyWire_0_5,
    n1096
  );


  not
  g1164
  (
    n1609,
    n833
  );


  not
  g1165
  (
    n1288,
    n1015
  );


  not
  g1166
  (
    n1689,
    n815
  );


  buf
  g1167
  (
    n1217,
    n939
  );


  buf
  g1168
  (
    n1209,
    n821
  );


  not
  g1169
  (
    n1507,
    n1064
  );


  not
  g1170
  (
    n1641,
    n1033
  );


  not
  g1171
  (
    n1300,
    n817
  );


  not
  g1172
  (
    n1179,
    n833
  );


  not
  g1173
  (
    n1508,
    n911
  );


  not
  g1174
  (
    n1276,
    n942
  );


  buf
  g1175
  (
    n1343,
    n1023
  );


  buf
  g1176
  (
    n1190,
    n1081
  );


  not
  g1177
  (
    n1599,
    n1050
  );


  not
  g1178
  (
    n1412,
    n798
  );


  not
  g1179
  (
    n1484,
    n1000
  );


  buf
  g1180
  (
    n1559,
    n1108
  );


  buf
  g1181
  (
    n1729,
    n1107
  );


  buf
  g1182
  (
    n1272,
    n827
  );


  not
  g1183
  (
    n1704,
    n1081
  );


  not
  g1184
  (
    n1296,
    n823
  );


  not
  g1185
  (
    n1428,
    n1126
  );


  not
  g1186
  (
    n1470,
    n907
  );


  buf
  g1187
  (
    n1212,
    n1007
  );


  not
  g1188
  (
    n1713,
    n1020
  );


  buf
  g1189
  (
    n1648,
    n1122
  );


  not
  g1190
  (
    n1628,
    n1028
  );


  not
  g1191
  (
    n1500,
    n983
  );


  buf
  g1192
  (
    n1701,
    n1021
  );


  not
  g1193
  (
    n1197,
    n1030
  );


  buf
  g1194
  (
    n1252,
    n1053
  );


  buf
  g1195
  (
    n1392,
    n1076
  );


  buf
  g1196
  (
    n1482,
    n1123
  );


  buf
  g1197
  (
    n1264,
    n1023
  );


  buf
  g1198
  (
    n1480,
    n923
  );


  not
  g1199
  (
    n1328,
    n1089
  );


  buf
  g1200
  (
    n1655,
    n915
  );


  buf
  g1201
  (
    n1174,
    n1001
  );


  not
  g1202
  (
    n1381,
    n823
  );


  buf
  g1203
  (
    n1301,
    n996
  );


  not
  g1204
  (
    n1646,
    n969
  );


  buf
  g1205
  (
    n1625,
    n816
  );


  buf
  g1206
  (
    n1259,
    n1008
  );


  buf
  g1207
  (
    n1368,
    n805
  );


  not
  g1208
  (
    n1358,
    n1098
  );


  not
  g1209
  (
    n1489,
    n1043
  );


  not
  g1210
  (
    n1660,
    n1061
  );


  buf
  g1211
  (
    n1388,
    n1102
  );


  buf
  g1212
  (
    n1529,
    n988
  );


  buf
  g1213
  (
    n1430,
    n1079
  );


  buf
  g1214
  (
    n1709,
    n1010
  );


  buf
  g1215
  (
    n1587,
    n826
  );


  not
  g1216
  (
    n1687,
    n1004
  );


  buf
  g1217
  (
    n1583,
    n830
  );


  not
  g1218
  (
    n1553,
    n1115
  );


  buf
  g1219
  (
    n1734,
    n1046
  );


  buf
  g1220
  (
    n1490,
    n806
  );


  buf
  g1221
  (
    n1332,
    n1024
  );


  not
  g1222
  (
    n1464,
    n837
  );


  buf
  g1223
  (
    n1326,
    n1002
  );


  not
  g1224
  (
    n1230,
    n1082
  );


  buf
  g1225
  (
    n1683,
    n1094
  );


  not
  g1226
  (
    n1270,
    n797
  );


  not
  g1227
  (
    n1176,
    n1040
  );


  not
  g1228
  (
    n1261,
    n819
  );


  buf
  g1229
  (
    n1218,
    n1118
  );


  not
  g1230
  (
    n1665,
    n821
  );


  buf
  g1231
  (
    n1535,
    n1137
  );


  not
  g1232
  (
    n1188,
    n1019
  );


  not
  g1233
  (
    n1654,
    n1037
  );


  buf
  g1234
  (
    n1606,
    n1048
  );


  not
  g1235
  (
    n1619,
    n987
  );


  not
  g1236
  (
    KeyWire_0_1,
    n811
  );


  not
  g1237
  (
    n1717,
    n1092
  );


  buf
  g1238
  (
    n1251,
    n1067
  );


  not
  g1239
  (
    n1205,
    n1138
  );


  not
  g1240
  (
    n1608,
    n914
  );


  buf
  g1241
  (
    n1295,
    n1066
  );


  not
  g1242
  (
    n1465,
    n1106
  );


  not
  g1243
  (
    n1233,
    n1062
  );


  buf
  g1244
  (
    n1334,
    n812
  );


  buf
  g1245
  (
    n1438,
    n916
  );


  buf
  g1246
  (
    n1148,
    n828
  );


  buf
  g1247
  (
    n1345,
    n1095
  );


  buf
  g1248
  (
    n1727,
    n1068
  );


  not
  g1249
  (
    n1410,
    n810
  );


  buf
  g1250
  (
    n1342,
    n806
  );


  buf
  g1251
  (
    n1242,
    n1106
  );


  not
  g1252
  (
    n1168,
    n1071
  );


  buf
  g1253
  (
    n1391,
    n1058
  );


  buf
  g1254
  (
    n1322,
    n1036
  );


  buf
  g1255
  (
    n1413,
    n1135
  );


  not
  g1256
  (
    n1467,
    n984
  );


  buf
  g1257
  (
    n1243,
    n822
  );


  buf
  g1258
  (
    n1537,
    n812
  );


  not
  g1259
  (
    n1222,
    n1036
  );


  buf
  g1260
  (
    n1283,
    n973
  );


  not
  g1261
  (
    n1633,
    n1059
  );


  buf
  g1262
  (
    n1325,
    n805
  );


  buf
  g1263
  (
    n1688,
    n1106
  );


  not
  g1264
  (
    n1627,
    n804
  );


  not
  g1265
  (
    n1454,
    n1047
  );


  not
  g1266
  (
    n1207,
    n1056
  );


  buf
  g1267
  (
    n1153,
    n1087
  );


  buf
  g1268
  (
    n1313,
    n1066
  );


  buf
  g1269
  (
    n1199,
    n1073
  );


  not
  g1270
  (
    n1398,
    n1061
  );


  buf
  g1271
  (
    n1707,
    n1056
  );


  buf
  g1272
  (
    n1323,
    n1068
  );


  not
  g1273
  (
    n1443,
    n1088
  );


  not
  g1274
  (
    n1602,
    n1128
  );


  buf
  g1275
  (
    n1163,
    n934
  );


  buf
  g1276
  (
    n1378,
    n812
  );


  buf
  g1277
  (
    n1662,
    n1020
  );


  not
  g1278
  (
    n1210,
    n830
  );


  not
  g1279
  (
    n1652,
    n1039
  );


  buf
  g1280
  (
    n1387,
    n1127
  );


  not
  g1281
  (
    n1672,
    n1115
  );


  buf
  g1282
  (
    n1172,
    n1026
  );


  not
  g1283
  (
    n1285,
    n966
  );


  buf
  g1284
  (
    n1634,
    n1071
  );


  buf
  g1285
  (
    n1329,
    n1009
  );


  buf
  g1286
  (
    n1679,
    n811
  );


  not
  g1287
  (
    n1303,
    n1046
  );


  buf
  g1288
  (
    n1198,
    n1022
  );


  not
  g1289
  (
    n1447,
    n1010
  );


  not
  g1290
  (
    n1630,
    n1057
  );


  not
  g1291
  (
    n1597,
    n794
  );


  not
  g1292
  (
    n1485,
    n987
  );


  buf
  g1293
  (
    n1206,
    n1096
  );


  not
  g1294
  (
    n1684,
    n1124
  );


  buf
  g1295
  (
    n1194,
    n904
  );


  not
  g1296
  (
    n1244,
    n1110
  );


  buf
  g1297
  (
    n1639,
    n1053
  );


  not
  g1298
  (
    n1248,
    n836
  );


  not
  g1299
  (
    n1340,
    n815
  );


  not
  g1300
  (
    n1397,
    n992
  );


  buf
  g1301
  (
    n1711,
    n950
  );


  not
  g1302
  (
    n1269,
    n1117
  );


  not
  g1303
  (
    n1415,
    n818
  );


  not
  g1304
  (
    n1445,
    n1105
  );


  buf
  g1305
  (
    n1542,
    n1120
  );


  not
  g1306
  (
    n1635,
    n1130
  );


  not
  g1307
  (
    n1545,
    n1099
  );


  not
  g1308
  (
    n1676,
    n832
  );


  not
  g1309
  (
    n1521,
    n1112
  );


  not
  g1310
  (
    n1383,
    n1072
  );


  not
  g1311
  (
    n1372,
    n1055
  );


  not
  g1312
  (
    n1700,
    n933
  );


  buf
  g1313
  (
    n1560,
    n1069
  );


  not
  g1314
  (
    n1638,
    n1128
  );


  not
  g1315
  (
    n1338,
    n1045
  );


  not
  g1316
  (
    n1149,
    n1052
  );


  buf
  g1317
  (
    n1308,
    n1067
  );


  buf
  g1318
  (
    n1367,
    n1138
  );


  buf
  g1319
  (
    n1647,
    n826
  );


  buf
  g1320
  (
    n1571,
    n815
  );


  not
  g1321
  (
    n1407,
    n819
  );


  not
  g1322
  (
    n1310,
    n925
  );


  not
  g1323
  (
    n1728,
    n1114
  );


  not
  g1324
  (
    n1551,
    n1013
  );


  buf
  g1325
  (
    n1169,
    n1136
  );


  not
  g1326
  (
    n1255,
    n1010
  );


  buf
  g1327
  (
    n1708,
    n924
  );


  buf
  g1328
  (
    n1363,
    n1088
  );


  not
  g1329
  (
    n1370,
    n802
  );


  not
  g1330
  (
    n1339,
    n1069
  );


  buf
  g1331
  (
    n1366,
    n803
  );


  not
  g1332
  (
    n1333,
    n920
  );


  not
  g1333
  (
    n1331,
    n1025
  );


  buf
  g1334
  (
    n1196,
    n1014
  );


  buf
  g1335
  (
    n1389,
    n1090
  );


  not
  g1336
  (
    n1686,
    n905
  );


  buf
  g1337
  (
    n1473,
    n1040
  );


  buf
  g1338
  (
    n1416,
    n1105
  );


  buf
  g1339
  (
    n1515,
    n1108
  );


  buf
  g1340
  (
    n1337,
    n825
  );


  buf
  g1341
  (
    n1187,
    n1119
  );


  not
  g1342
  (
    n1265,
    n806
  );


  buf
  g1343
  (
    n1309,
    n1097
  );


  buf
  g1344
  (
    n1352,
    n813
  );


  buf
  g1345
  (
    n1594,
    n1127
  );


  not
  g1346
  (
    n1578,
    n1065
  );


  not
  g1347
  (
    n1236,
    n1011
  );


  not
  g1348
  (
    n1615,
    n1114
  );


  not
  g1349
  (
    n1267,
    n1052
  );


  not
  g1350
  (
    n1315,
    n1016
  );


  buf
  g1351
  (
    n1286,
    n1112
  );


  buf
  g1352
  (
    n1692,
    n961
  );


  buf
  g1353
  (
    n1254,
    n1090
  );


  not
  g1354
  (
    n1155,
    n1099
  );


  not
  g1355
  (
    n1493,
    n1103
  );


  buf
  g1356
  (
    n1565,
    n1028
  );


  not
  g1357
  (
    n1492,
    n1119
  );


  not
  g1358
  (
    n1318,
    n1086
  );


  not
  g1359
  (
    n1282,
    n1053
  );


  buf
  g1360
  (
    n1241,
    n802
  );


  not
  g1361
  (
    n1327,
    n1005
  );


  not
  g1362
  (
    n1466,
    n981
  );


  buf
  g1363
  (
    n1414,
    n1028
  );


  buf
  g1364
  (
    n1611,
    n1075
  );


  buf
  g1365
  (
    n1595,
    n965
  );


  not
  g1366
  (
    n1716,
    n1134
  );


  buf
  g1367
  (
    n1463,
    n1093
  );


  not
  g1368
  (
    n1402,
    n1054
  );


  buf
  g1369
  (
    n1703,
    n1035
  );


  not
  g1370
  (
    n1150,
    n802
  );


  not
  g1371
  (
    n1569,
    n294
  );


  buf
  g1372
  (
    n1256,
    n1013
  );


  not
  g1373
  (
    n1305,
    n1138
  );


  not
  g1374
  (
    n1441,
    n971
  );


  not
  g1375
  (
    n1546,
    n1121
  );


  buf
  g1376
  (
    n1723,
    n1029
  );


  buf
  g1377
  (
    n1245,
    n1034
  );


  buf
  g1378
  (
    n1253,
    n1111
  );


  buf
  g1379
  (
    n1557,
    n1116
  );


  not
  g1380
  (
    KeyWire_0_9,
    n813
  );


  not
  g1381
  (
    n1164,
    n828
  );


  buf
  g1382
  (
    n1731,
    n1135
  );


  buf
  g1383
  (
    n1453,
    n1132
  );


  not
  g1384
  (
    n1705,
    n1048
  );


  buf
  g1385
  (
    n1685,
    n985
  );


  not
  g1386
  (
    n1446,
    n1116
  );


  buf
  g1387
  (
    n1681,
    n1021
  );


  not
  g1388
  (
    n1375,
    n1029
  );


  not
  g1389
  (
    n1513,
    n1037
  );


  not
  g1390
  (
    n1673,
    n1111
  );


  not
  g1391
  (
    n1505,
    n809
  );


  not
  g1392
  (
    n1299,
    n1054
  );


  not
  g1393
  (
    n1620,
    n1086
  );


  buf
  g1394
  (
    n1219,
    n1124
  );


  buf
  g1395
  (
    n1180,
    n1080
  );


  not
  g1396
  (
    n1733,
    n836
  );


  not
  g1397
  (
    n1525,
    n901
  );


  buf
  g1398
  (
    n1246,
    n948
  );


  buf
  g1399
  (
    n1487,
    n831
  );


  not
  g1400
  (
    n1393,
    n1054
  );


  buf
  g1401
  (
    n1539,
    n1089
  );


  not
  g1402
  (
    n1321,
    n1130
  );


  buf
  g1403
  (
    n1214,
    n1025
  );


  buf
  g1404
  (
    n1523,
    n919
  );


  not
  g1405
  (
    n1498,
    n816
  );


  not
  g1406
  (
    n1534,
    n1035
  );


  buf
  g1407
  (
    n1511,
    n1133
  );


  buf
  g1408
  (
    n1478,
    n1046
  );


  buf
  g1409
  (
    n1541,
    n1038
  );


  buf
  g1410
  (
    n1592,
    n1025
  );


  not
  g1411
  (
    n1408,
    n1004
  );


  not
  g1412
  (
    n1675,
    n972
  );


  not
  g1413
  (
    n1223,
    n977
  );


  buf
  g1414
  (
    n1422,
    n1077
  );


  buf
  g1415
  (
    n1405,
    n1135
  );


  not
  g1416
  (
    n1653,
    n807
  );


  buf
  g1417
  (
    n1668,
    n839
  );


  buf
  g1418
  (
    n1341,
    n1063
  );


  buf
  g1419
  (
    n1650,
    n1123
  );


  not
  g1420
  (
    n1144,
    n1051
  );


  not
  g1421
  (
    n1158,
    n821
  );


  buf
  g1422
  (
    n1528,
    n810
  );


  not
  g1423
  (
    n1614,
    n1113
  );


  buf
  g1424
  (
    n1694,
    n1041
  );


  buf
  g1425
  (
    n1400,
    n829
  );


  not
  g1426
  (
    n1266,
    n1030
  );


  not
  g1427
  (
    n1292,
    n1109
  );


  buf
  g1428
  (
    n1294,
    n834
  );


  not
  g1429
  (
    n1433,
    n1091
  );


  not
  g1430
  (
    n1221,
    n838
  );


  not
  g1431
  (
    n1736,
    n981
  );


  buf
  g1432
  (
    n1538,
    n795
  );


  buf
  g1433
  (
    n1649,
    n810
  );


  not
  g1434
  (
    n1718,
    n800
  );


  buf
  g1435
  (
    n1380,
    n1012
  );


  buf
  g1436
  (
    n1555,
    n983
  );


  buf
  g1437
  (
    n1536,
    n1084
  );


  buf
  g1438
  (
    n1533,
    n903
  );


  buf
  g1439
  (
    n1146,
    n968
  );


  not
  g1440
  (
    n1591,
    n1092
  );


  not
  g1441
  (
    n1213,
    n804
  );


  not
  g1442
  (
    n1509,
    n1108
  );


  buf
  g1443
  (
    n1330,
    n1070
  );


  buf
  g1444
  (
    n1237,
    n1019
  );


  not
  g1445
  (
    n1706,
    n1112
  );


  not
  g1446
  (
    n1586,
    n900
  );


  buf
  g1447
  (
    n1354,
    n1049
  );


  buf
  g1448
  (
    n1497,
    n1032
  );


  buf
  g1449
  (
    n1488,
    n1113
  );


  buf
  g1450
  (
    n1145,
    n1070
  );


  not
  g1451
  (
    n1362,
    n1052
  );


  buf
  g1452
  (
    n1426,
    n1059
  );


  buf
  g1453
  (
    n1152,
    n1132
  );


  buf
  g1454
  (
    n1316,
    n1073
  );


  buf
  g1455
  (
    n1235,
    n1119
  );


  buf
  g1456
  (
    n1526,
    n817
  );


  buf
  g1457
  (
    n1624,
    n1099
  );


  not
  g1458
  (
    n1156,
    n1033
  );


  not
  g1459
  (
    n1494,
    n1076
  );


  buf
  g1460
  (
    n1631,
    n1033
  );


  not
  g1461
  (
    n1171,
    n1065
  );


  not
  g1462
  (
    n1448,
    n1034
  );


  not
  g1463
  (
    n1610,
    n1138
  );


  buf
  g1464
  (
    n1643,
    n1107
  );


  not
  g1465
  (
    n1384,
    n1139
  );


  buf
  g1466
  (
    n1590,
    n1044
  );


  buf
  g1467
  (
    n1604,
    n803
  );


  buf
  g1468
  (
    n1735,
    n1007
  );


  buf
  g1469
  (
    n1434,
    n1128
  );


  buf
  g1470
  (
    n1281,
    n1060
  );


  not
  g1471
  (
    n1437,
    n994
  );


  not
  g1472
  (
    n1585,
    n1090
  );


  buf
  g1473
  (
    n1506,
    n1018
  );


  buf
  g1474
  (
    n1249,
    n941
  );


  buf
  g1475
  (
    n1215,
    n824
  );


  buf
  g1476
  (
    n1182,
    n808
  );


  buf
  g1477
  (
    n1239,
    n1060
  );


  not
  g1478
  (
    n1664,
    n823
  );


  not
  g1479
  (
    n1603,
    n1032
  );


  not
  g1480
  (
    n1574,
    n1014
  );


  not
  g1481
  (
    n1667,
    n990
  );


  not
  g1482
  (
    n1678,
    n1016
  );


  not
  g1483
  (
    n1257,
    n1022
  );


  not
  g1484
  (
    n1178,
    n993
  );


  not
  g1485
  (
    n1486,
    n839
  );


  not
  g1486
  (
    n1165,
    n1017
  );


  not
  g1487
  (
    n1721,
    n824
  );


  buf
  g1488
  (
    n1429,
    n1071
  );


  not
  g1489
  (
    n1471,
    n1136
  );


  not
  g1490
  (
    n1696,
    n980
  );


  buf
  g1491
  (
    n1593,
    n1137
  );


  buf
  g1492
  (
    n1403,
    n1115
  );


  not
  g1493
  (
    n1154,
    n1077
  );


  not
  g1494
  (
    n1385,
    n796
  );


  not
  g1495
  (
    n1232,
    n1011
  );


  not
  g1496
  (
    n1702,
    n1103
  );


  not
  g1497
  (
    n1451,
    n839
  );


  not
  g1498
  (
    KeyWire_0_6,
    n1082
  );


  not
  g1499
  (
    n1186,
    n940
  );


  not
  g1500
  (
    n1382,
    n1023
  );


  buf
  g1501
  (
    n1314,
    n1055
  );


  buf
  g1502
  (
    n1663,
    n1065
  );


  not
  g1503
  (
    n1469,
    n818
  );


  buf
  g1504
  (
    n1141,
    n1086
  );


  buf
  g1505
  (
    n1435,
    n814
  );


  not
  g1506
  (
    n1262,
    n1114
  );


  not
  g1507
  (
    n1573,
    n1117
  );


  buf
  g1508
  (
    n1561,
    n918
  );


  not
  g1509
  (
    n1360,
    n935
  );


  not
  g1510
  (
    n1353,
    n1075
  );


  buf
  g1511
  (
    n1658,
    n1075
  );


  not
  g1512
  (
    n1290,
    n1062
  );


  not
  g1513
  (
    n1417,
    n815
  );


  buf
  g1514
  (
    n1607,
    n1132
  );


  buf
  g1515
  (
    n1195,
    n1088
  );


  not
  g1516
  (
    n1726,
    n827
  );


  buf
  g1517
  (
    n1183,
    n989
  );


  not
  g1518
  (
    n1657,
    n955
  );


  not
  g1519
  (
    n1320,
    n1059
  );


  not
  g1520
  (
    n1359,
    n817
  );


  buf
  g1521
  (
    n1659,
    n986
  );


  buf
  g1522
  (
    n1203,
    n1139
  );


  not
  g1523
  (
    n1496,
    n988
  );


  buf
  g1524
  (
    n1715,
    n1078
  );


  not
  g1525
  (
    n1349,
    n796
  );


  not
  g1526
  (
    n1530,
    n1005
  );


  buf
  g1527
  (
    n1344,
    n1088
  );


  not
  g1528
  (
    n1297,
    n1087
  );


  buf
  g1529
  (
    n1626,
    n936
  );


  buf
  g1530
  (
    n1394,
    n1072
  );


  not
  g1531
  (
    n1142,
    n1126
  );


  not
  g1532
  (
    n1450,
    n833
  );


  buf
  g1533
  (
    n1302,
    n932
  );


  buf
  g1534
  (
    n1364,
    n1039
  );


  not
  g1535
  (
    n1184,
    n1019
  );


  not
  g1536
  (
    n1424,
    n1067
  );


  buf
  g1537
  (
    n1632,
    n1006
  );


  buf
  g1538
  (
    n1481,
    n1099
  );


  buf
  g1539
  (
    n1670,
    n1006
  );


  not
  g1540
  (
    n1280,
    n795
  );


  buf
  g1541
  (
    n1396,
    n909
  );


  not
  g1542
  (
    n1201,
    n1083
  );


  not
  g1543
  (
    n1629,
    n824
  );


  not
  g1544
  (
    n1432,
    n653
  );


  buf
  g1545
  (
    n1556,
    n1066
  );


  not
  g1546
  (
    n1401,
    n964
  );


  not
  g1547
  (
    n1226,
    n794
  );


  not
  g1548
  (
    n1348,
    n930
  );


  buf
  g1549
  (
    n1477,
    n1074
  );


  buf
  g1550
  (
    n1287,
    n1058
  );


  buf
  g1551
  (
    n1143,
    n1104
  );


  buf
  g1552
  (
    n1291,
    n800
  );


  buf
  g1553
  (
    n1449,
    n976
  );


  not
  g1554
  (
    n1577,
    n1120
  );


  buf
  g1555
  (
    n1271,
    n818
  );


  not
  g1556
  (
    n1564,
    n820
  );


  buf
  g1557
  (
    n1229,
    n945
  );


  not
  g1558
  (
    n1220,
    n839
  );


  not
  g1559
  (
    n1547,
    n1137
  );


  not
  g1560
  (
    n1699,
    n1118
  );


  not
  g1561
  (
    n1514,
    n1072
  );


  buf
  g1562
  (
    n1697,
    n1063
  );


  buf
  g1563
  (
    n1379,
    n967
  );


  not
  g1564
  (
    n1680,
    n1029
  );


  not
  g1565
  (
    n1258,
    n952
  );


  buf
  g1566
  (
    n1293,
    n991
  );


  not
  g1567
  (
    n1311,
    n1034
  );


  not
  g1568
  (
    n1562,
    n996
  );


  buf
  g1569
  (
    n1170,
    n825
  );


  buf
  g1570
  (
    n1548,
    n1085
  );


  buf
  g1571
  (
    n1211,
    n1102
  );


  buf
  g1572
  (
    n1192,
    n830
  );


  not
  g1573
  (
    n1600,
    n1073
  );


  buf
  g1574
  (
    n1710,
    n1094
  );


  buf
  g1575
  (
    n1622,
    n1136
  );


  not
  g1576
  (
    n1275,
    n1057
  );


  buf
  g1577
  (
    n1277,
    n1026
  );


  not
  g1578
  (
    n1440,
    n803
  );


  buf
  g1579
  (
    n1642,
    n1124
  );


  not
  g1580
  (
    n1455,
    n1037
  );


  not
  g1581
  (
    KeyWire_0_15,
    n1086
  );


  not
  g1582
  (
    n1346,
    n1065
  );


  buf
  g1583
  (
    n1475,
    n1115
  );


  not
  g1584
  (
    n1365,
    n943
  );


  not
  g1585
  (
    n1637,
    n975
  );


  buf
  g1586
  (
    n1225,
    n1097
  );


  buf
  g1587
  (
    n1566,
    n1020
  );


  buf
  g1588
  (
    n1231,
    n827
  );


  buf
  g1589
  (
    n1436,
    n799
  );


  not
  g1590
  (
    n1439,
    n1058
  );


  buf
  g1591
  (
    n1570,
    n831
  );


  not
  g1592
  (
    n1524,
    n1023
  );


  not
  g1593
  (
    n1518,
    n819
  );


  buf
  g1594
  (
    n1549,
    n1050
  );


  not
  g1595
  (
    n1427,
    n1070
  );


  buf
  g1596
  (
    n1200,
    n837
  );


  buf
  g1597
  (
    n1656,
    n832
  );


  not
  g1598
  (
    n1605,
    n807
  );


  not
  g1599
  (
    n1719,
    n1050
  );


  buf
  g1600
  (
    n1645,
    n998
  );


  not
  g1601
  (
    n1350,
    n1016
  );


  not
  g1602
  (
    n1730,
    n1081
  );


  not
  g1603
  (
    n1563,
    n1055
  );


  not
  g1604
  (
    n1386,
    n838
  );


  not
  g1605
  (
    n1532,
    n1104
  );


  not
  g1606
  (
    n1234,
    n1095
  );


  not
  g1607
  (
    n1457,
    n1130
  );


  not
  g1608
  (
    n1390,
    n1019
  );


  buf
  g1609
  (
    n1374,
    n838
  );


  not
  g1610
  (
    n1317,
    n1066
  );


  buf
  g1611
  (
    n1491,
    n829
  );


  not
  g1612
  (
    n1617,
    n927
  );


  buf
  g1613
  (
    n1307,
    n956
  );


  buf
  g1614
  (
    n1460,
    n832
  );


  and
  g1615
  (
    n1501,
    n1122,
    n804,
    n962,
    n705
  );


  nand
  g1616
  (
    n1227,
    n997,
    n1042,
    n1044,
    n1123
  );


  xor
  g1617
  (
    n1444,
    n1103,
    n820,
    n1133,
    n974
  );


  nor
  g1618
  (
    n1166,
    n971,
    n1074,
    n1045,
    n1129
  );


  nand
  g1619
  (
    n1483,
    n824,
    n1021,
    n825,
    n1084
  );


  nand
  g1620
  (
    n1216,
    n797,
    n958,
    n1079,
    n812
  );


  or
  g1621
  (
    n1567,
    n795,
    n975,
    n928,
    n1051
  );


  xnor
  g1622
  (
    n1191,
    n1131,
    n1024,
    n1117,
    n1041
  );


  and
  g1623
  (
    n1160,
    n1084,
    n1125,
    n978,
    n822
  );


  xor
  g1624
  (
    n1596,
    n1005,
    n1054,
    n1121,
    n1092
  );


  and
  g1625
  (
    n1499,
    n1081,
    n798,
    n801,
    n1085
  );


  xor
  g1626
  (
    n1568,
    n1075,
    n926,
    n1134,
    n1098
  );


  xor
  g1627
  (
    n1462,
    n1029,
    n1098,
    n819,
    n1047
  );


  nor
  g1628
  (
    n1623,
    n1059,
    n1007,
    n1015,
    n1073
  );


  xnor
  g1629
  (
    n1167,
    n1017,
    n822,
    n917,
    n1036
  );


  xnor
  g1630
  (
    n1274,
    n1060,
    n1064,
    n1026,
    n1043
  );


  nor
  g1631
  (
    n1452,
    n1126,
    n1009,
    n1001,
    n990
  );


  and
  g1632
  (
    n1550,
    n1083,
    n982,
    n989,
    n1125
  );


  xnor
  g1633
  (
    n1336,
    n1033,
    n1098,
    n828,
    n798
  );


  or
  g1634
  (
    n1159,
    n1027,
    n1102,
    n831,
    n954
  );


  and
  g1635
  (
    n1411,
    n1043,
    n1121,
    n1106,
    n1079
  );


  xor
  g1636
  (
    n1279,
    n1100,
    n836,
    n797,
    n796
  );


  nor
  g1637
  (
    n1502,
    n1101,
    n1003,
    n1129,
    n1131
  );


  or
  g1638
  (
    n1263,
    n980,
    n837,
    n1129,
    n993
  );


  xnor
  g1639
  (
    n1669,
    n1076,
    n1125,
    n822,
    n836
  );


  nor
  g1640
  (
    n1558,
    n1006,
    n1078,
    n833,
    n829
  );


  xor
  g1641
  (
    n1601,
    n913,
    n995,
    n1091,
    n1070
  );


  nor
  g1642
  (
    n1738,
    n1016,
    n1123,
    n795,
    n1083
  );


  xor
  g1643
  (
    n1208,
    n1017,
    n801,
    n1121,
    n1038
  );


  nand
  g1644
  (
    n1584,
    n1022,
    n1042,
    n809,
    n1131
  );


  or
  g1645
  (
    n1442,
    n1087,
    n1063,
    n1012,
    n1103
  );


  nor
  g1646
  (
    n1278,
    n827,
    n1038,
    n1110,
    n1111
  );


  or
  g1647
  (
    n1355,
    n910,
    n1049,
    n813,
    n800
  );


  and
  g1648
  (
    n1474,
    n994,
    n1032,
    n1095,
    n1076
  );


  xnor
  g1649
  (
    n1504,
    n1105,
    n830,
    n1010,
    n1107
  );


  nand
  g1650
  (
    n1406,
    n1048,
    n800,
    n951,
    n1045
  );


  xnor
  g1651
  (
    n1575,
    n816,
    n1041,
    n1078
  );


  and
  g1652
  (
    n1540,
    n1136,
    n1102,
    n1061,
    n992
  );


  nand
  g1653
  (
    n1161,
    n998,
    n1003,
    n801,
    n1028
  );


  xor
  g1654
  (
    n1720,
    n1039,
    n1122,
    n829,
    n1085
  );


  nor
  g1655
  (
    n1335,
    n1133,
    n1056,
    n1127,
    n1047
  );


  xnor
  g1656
  (
    n1712,
    n959,
    n834,
    n906,
    n1052
  );


  or
  g1657
  (
    n1724,
    n825,
    n1053,
    n970,
    n1009
  );


  nand
  g1658
  (
    n1189,
    n1101,
    n1060,
    n1109,
    n979
  );


  xor
  g1659
  (
    n1459,
    n1080,
    n1093,
    n814,
    n949
  );


  or
  g1660
  (
    n1423,
    n1018,
    n1092,
    n835,
    n809
  );


  xor
  g1661
  (
    n1250,
    n1100,
    n808,
    n1129,
    n1082
  );


  or
  g1662
  (
    n1247,
    n1126,
    n1071,
    n972,
    n973
  );


  nand
  g1663
  (
    n1356,
    n797,
    n946,
    n823,
    n1038
  );


  nor
  g1664
  (
    n1240,
    n1134,
    n1089,
    n1062,
    n1043
  );


  or
  g1665
  (
    n1425,
    n295,
    n1015,
    n810,
    n1112
  );


  xor
  g1666
  (
    n1671,
    n1108,
    n1122,
    n1080,
    n938
  );


  or
  g1667
  (
    n1613,
    n999,
    n1008,
    n1031,
    n807
  );


  nand
  g1668
  (
    n1204,
    n1035,
    n1068,
    n1005,
    n1109
  );


  nand
  g1669
  (
    n1644,
    n799,
    n912,
    n1116,
    n1094
  );


  or
  g1670
  (
    n1347,
    n1135,
    n1012,
    n1046,
    n1049
  );


  and
  g1671
  (
    n1260,
    n820,
    n799,
    n808,
    n1030
  );


  xor
  g1672
  (
    n1376,
    n1009,
    n1134,
    n804,
    n1064
  );


  xor
  g1673
  (
    n1520,
    n984,
    n1120,
    n828,
    n1084
  );


  nor
  g1674
  (
    n1479,
    n1137,
    n1014,
    n1082,
    n838
  );


  and
  g1675
  (
    n1175,
    n1077,
    n1051,
    n1101,
    n794
  );


  xor
  g1676
  (
    n1636,
    n967,
    n806,
    n1050,
    n1062
  );


  or
  g1677
  (
    n1690,
    n1008,
    n1024,
    n1055,
    n1072
  );


  nor
  g1678
  (
    n1181,
    n974,
    n816,
    n1091,
    n811
  );


  xnor
  g1679
  (
    n1461,
    n1117,
    n1027,
    n944,
    n1118
  );


  xnor
  g1680
  (
    n1580,
    n1018,
    n953,
    n1047,
    n1042
  );


  and
  g1681
  (
    n1369,
    n1132,
    n805,
    n1058,
    n826
  );


  or
  g1682
  (
    n1589,
    n835,
    n1079,
    n1031,
    n947
  );


  xor
  g1683
  (
    n1581,
    n999,
    n796,
    n1014,
    n1074
  );


  xnor
  g1684
  (
    n1418,
    n1017,
    n805,
    n832,
    n826
  );


  xor
  g1685
  (
    n1173,
    n902,
    n1089,
    n1051,
    n1107
  );


  xnor
  g1686
  (
    n1395,
    n1127,
    n1105,
    n802,
    n1119
  );


  xor
  g1687
  (
    n1576,
    n1093,
    n1027,
    n1131,
    n1039
  );


  xor
  g1688
  (
    n1714,
    n1021,
    n1077,
    n970,
    n1128
  );


  and
  g1689
  (
    n1698,
    n977,
    n808,
    n1100,
    n1139
  );


  or
  g1690
  (
    n1598,
    n991,
    n1104,
    n1139,
    n803
  );


  xnor
  g1691
  (
    n1512,
    n995,
    n1020,
    n1113,
    n820
  );


  nor
  g1692
  (
    n1284,
    n1013,
    n1030,
    n908,
    n1011
  );


  nor
  g1693
  (
    n1456,
    n1018,
    n807,
    n1069,
    n1024
  );


  nor
  g1694
  (
    n1361,
    n1101,
    n979,
    n1093,
    n997
  );


  xor
  g1695
  (
    n1572,
    n1044,
    n821,
    n831,
    n1124
  );


  or
  g1696
  (
    n1157,
    n1067,
    n1013,
    n957,
    n986
  );


  and
  g1697
  (
    n1531,
    n1069,
    n1097,
    n1125,
    n1049
  );


  and
  g1698
  (
    n1357,
    n1096,
    n1085,
    n1116,
    n811
  );


  xor
  g1699
  (
    n1421,
    n1061,
    n1074,
    n1036,
    n1037
  );


  and
  g1700
  (
    n1404,
    n1000,
    n818,
    n982,
    n1090
  );


  xnor
  g1701
  (
    n1476,
    n976,
    n1118,
    n814,
    n835
  );


  nand
  g1702
  (
    n1224,
    n1078,
    n1114,
    n937,
    n798
  );


  xnor
  g1703
  (
    n1468,
    n922,
    n1110,
    n835,
    n1057
  );


  xnor
  g1704
  (
    n1651,
    n809,
    n1110,
    n1113,
    n1068
  );


  xor
  g1705
  (
    n1377,
    n1034,
    n1095,
    n1031,
    n1056
  );


  nor
  g1706
  (
    n1881,
    n1211,
    n1620,
    n1356,
    n1489
  );


  or
  g1707
  (
    n1834,
    n373,
    n1616,
    n1680,
    n1215
  );


  xor
  g1708
  (
    n1905,
    n383,
    n1160,
    n503,
    n512
  );


  xnor
  g1709
  (
    n1828,
    n1173,
    n1263,
    n298,
    n1608
  );


  or
  g1710
  (
    n1786,
    n1538,
    n377,
    n1380,
    n1695
  );


  nand
  g1711
  (
    n1929,
    n547,
    n1705,
    n1479,
    n1732
  );


  or
  g1712
  (
    n1760,
    n1627,
    n441,
    n1504,
    n1443
  );


  xor
  g1713
  (
    n1936,
    n539,
    n1687,
    n1487,
    n1614
  );


  nand
  g1714
  (
    n1769,
    n1283,
    n1244,
    n1654,
    n359
  );


  or
  g1715
  (
    n1831,
    n1426,
    n1152,
    n1253,
    n1631
  );


  xnor
  g1716
  (
    n1867,
    n1256,
    n341,
    n1451,
    n1255
  );


  nand
  g1717
  (
    n1773,
    n1606,
    n1516,
    n1526,
    n1600
  );


  nor
  g1718
  (
    n1808,
    n1327,
    n1488,
    n1722,
    n1247
  );


  nor
  g1719
  (
    n1857,
    n1517,
    n345,
    n360,
    n1394
  );


  xor
  g1720
  (
    n1942,
    n1469,
    n335,
    n1532,
    n1601
  );


  or
  g1721
  (
    n1849,
    n1636,
    n394,
    n1369,
    n1200
  );


  or
  g1722
  (
    n1959,
    n1448,
    n482,
    n1351,
    n1509
  );


  nor
  g1723
  (
    n1815,
    n1581,
    n336,
    n1447,
    n1389
  );


  nand
  g1724
  (
    n1889,
    n1424,
    n1164,
    n1667,
    n1465
  );


  nand
  g1725
  (
    n1770,
    n1251,
    n574,
    n303,
    n1148
  );


  or
  g1726
  (
    n1824,
    n1725,
    n1198,
    n1219,
    n1652
  );


  xor
  g1727
  (
    n1844,
    n1734,
    n542,
    n1460,
    n1243
  );


  nor
  g1728
  (
    n1860,
    n342,
    n520,
    n1578,
    n317
  );


  nand
  g1729
  (
    n1894,
    n1323,
    n444,
    n1359,
    n1186
  );


  xor
  g1730
  (
    n1757,
    n1337,
    n1298,
    n1728,
    n1252
  );


  and
  g1731
  (
    n1741,
    n399,
    n308,
    n1669,
    n384
  );


  nand
  g1732
  (
    n1768,
    n1299,
    n1378,
    n416,
    n1333
  );


  nor
  g1733
  (
    n1906,
    n1681,
    n1672,
    n1473,
    n1557
  );


  nor
  g1734
  (
    n1863,
    n1153,
    n1408,
    n1724,
    n1403
  );


  xor
  g1735
  (
    n1784,
    n1259,
    n1726,
    n1582,
    n1268
  );


  and
  g1736
  (
    n1838,
    n374,
    n1735,
    n1275,
    n391
  );


  xor
  g1737
  (
    n1961,
    n1611,
    n1413,
    n1657,
    n1206
  );


  xor
  g1738
  (
    n1861,
    n1232,
    n1587,
    n1257,
    n521
  );


  nor
  g1739
  (
    n1954,
    n1676,
    n1315,
    n1508,
    n1157
  );


  and
  g1740
  (
    n1941,
    n1446,
    n544,
    n1317,
    n1635
  );


  xnor
  g1741
  (
    n1858,
    n389,
    n418,
    n1521,
    n1466
  );


  nor
  g1742
  (
    n1928,
    n1320,
    n579,
    n1233,
    n463
  );


  nand
  g1743
  (
    n1866,
    n1518,
    n1150,
    n1593,
    n1549
  );


  nand
  g1744
  (
    n1829,
    n1352,
    n1335,
    n1273,
    n1503
  );


  or
  g1745
  (
    n1744,
    n363,
    n518,
    n1617,
    n504
  );


  and
  g1746
  (
    n1767,
    n306,
    n1267,
    n1213,
    n1332
  );


  xor
  g1747
  (
    n1746,
    n1632,
    n307,
    n526,
    n1621
  );


  xor
  g1748
  (
    n1806,
    n1397,
    n1499,
    n1300,
    n1190
  );


  nor
  g1749
  (
    n1917,
    n1541,
    n456,
    n1468,
    n1625
  );


  and
  g1750
  (
    n1750,
    n1575,
    n1607,
    n1368,
    n509
  );


  and
  g1751
  (
    n1899,
    n1195,
    n1280,
    n405,
    n465
  );


  or
  g1752
  (
    n1765,
    n1348,
    n385,
    n550,
    n572
  );


  and
  g1753
  (
    n1926,
    n1573,
    n1714,
    n1441,
    n1360
  );


  nand
  g1754
  (
    n1912,
    n583,
    n1506,
    n1480,
    n489
  );


  or
  g1755
  (
    n1803,
    n1427,
    n496,
    n1421,
    n1192
  );


  xor
  g1756
  (
    n1877,
    n375,
    n1502,
    n1203,
    n1530
  );


  nor
  g1757
  (
    n1782,
    n1303,
    n437,
    n479,
    n1553
  );


  nor
  g1758
  (
    n1810,
    n1277,
    n338,
    n1535,
    n573
  );


  xnor
  g1759
  (
    n1921,
    n423,
    n1143,
    n1241,
    n1453
  );


  xor
  g1760
  (
    n1843,
    n1703,
    n1240,
    n1286,
    n1640
  );


  xnor
  g1761
  (
    n1895,
    n1476,
    n321,
    n528,
    n1189
  );


  xor
  g1762
  (
    n1809,
    n1289,
    n1710,
    n1520,
    n1534
  );


  nor
  g1763
  (
    n1891,
    n443,
    n1296,
    n1694,
    n366
  );


  nor
  g1764
  (
    n1790,
    n1653,
    n1603,
    n1391,
    n315
  );


  or
  g1765
  (
    n1864,
    n1628,
    n1347,
    n1513,
    n1589
  );


  nand
  g1766
  (
    n1915,
    n1527,
    n1341,
    n1224,
    n708
  );


  nor
  g1767
  (
    n1900,
    n1629,
    n316,
    n1444,
    n1647
  );


  and
  g1768
  (
    n1886,
    n1254,
    n1339,
    n1295,
    n580
  );


  and
  g1769
  (
    n1903,
    n1477,
    n1210,
    n1586,
    n707
  );


  nor
  g1770
  (
    n1871,
    n1715,
    n1602,
    n1528,
    n468
  );


  xor
  g1771
  (
    n1837,
    n535,
    n1434,
    n464,
    n1677
  );


  nand
  g1772
  (
    n1931,
    n1161,
    n415,
    n372,
    n1439
  );


  or
  g1773
  (
    n1911,
    n368,
    n1462,
    n1623,
    n540
  );


  nor
  g1774
  (
    n1953,
    n1155,
    n1709,
    n1361,
    n1498
  );


  or
  g1775
  (
    n1874,
    n1472,
    n1235,
    n1459,
    n1718
  );


  and
  g1776
  (
    n1885,
    n1605,
    n1495,
    n1552,
    n1383
  );


  xnor
  g1777
  (
    n1848,
    n1505,
    n461,
    n1220,
    n1171
  );


  nor
  g1778
  (
    n1934,
    n553,
    n404,
    n421,
    n1696
  );


  nand
  g1779
  (
    n1797,
    n538,
    n537,
    n1218,
    n1551
  );


  xnor
  g1780
  (
    n1949,
    n523,
    n1234,
    n1562,
    n1682
  );


  nand
  g1781
  (
    n1745,
    n1537,
    n1305,
    n1306,
    n1212
  );


  and
  g1782
  (
    n1827,
    n1656,
    n493,
    n1387,
    n1436
  );


  or
  g1783
  (
    n1791,
    n1420,
    n1674,
    n408,
    n1363
  );


  nor
  g1784
  (
    n1920,
    n151,
    n1491,
    n566,
    n330
  );


  or
  g1785
  (
    n1778,
    n1440,
    n1338,
    n1556,
    n1358
  );


  xnor
  g1786
  (
    n1839,
    n1633,
    n393,
    n525,
    n561
  );


  nand
  g1787
  (
    n1960,
    n1577,
    n1272,
    n376,
    n1438
  );


  nor
  g1788
  (
    n1887,
    n1641,
    n483,
    n1177,
    n1683
  );


  and
  g1789
  (
    n1814,
    n1217,
    n1730,
    n472,
    n1490
  );


  or
  g1790
  (
    n1851,
    n1425,
    n478,
    n551,
    n406
  );


  nand
  g1791
  (
    n1804,
    n1242,
    n490,
    n1342,
    n1159
  );


  xnor
  g1792
  (
    n1742,
    n1384,
    n451,
    n318,
    n1227
  );


  xor
  g1793
  (
    n1854,
    n1284,
    n488,
    n1619,
    n499
  );


  xor
  g1794
  (
    n1937,
    n1416,
    n1548,
    n1555,
    n1291
  );


  xnor
  g1795
  (
    n1842,
    n438,
    n1308,
    n519,
    n1501
  );


  nand
  g1796
  (
    n1811,
    n1313,
    n1258,
    n1184,
    n1178
  );


  xor
  g1797
  (
    n1780,
    n1409,
    n365,
    n1692,
    n151
  );


  xor
  g1798
  (
    n1792,
    n1497,
    n1209,
    n1561,
    n1467
  );


  or
  g1799
  (
    n1904,
    n1165,
    n300,
    n581,
    n1319
  );


  xor
  g1800
  (
    n1832,
    n1330,
    n382,
    n1376,
    n1454
  );


  xor
  g1801
  (
    n1759,
    n1464,
    n1547,
    n299,
    n1329
  );


  xor
  g1802
  (
    n1787,
    n350,
    n1156,
    n541,
    n388
  );


  xor
  g1803
  (
    n1749,
    n344,
    n1545,
    n434,
    n452
  );


  xor
  g1804
  (
    n1840,
    n1510,
    n390,
    n1716,
    n1570
  );


  or
  g1805
  (
    n1907,
    n1226,
    n407,
    n1388,
    n348
  );


  and
  g1806
  (
    n1743,
    n1287,
    n304,
    n1540,
    n1365
  );


  nand
  g1807
  (
    n1785,
    n1452,
    n430,
    n322,
    n449
  );


  or
  g1808
  (
    n1764,
    n536,
    n1585,
    n325,
    n1396
  );


  xnor
  g1809
  (
    n1927,
    n1326,
    n1613,
    n455,
    n427
  );


  xnor
  g1810
  (
    n1795,
    n1316,
    n558,
    n1717,
    n1412
  );


  xor
  g1811
  (
    n1836,
    n1288,
    n530,
    n1314,
    n1353
  );


  and
  g1812
  (
    n1799,
    n1398,
    n369,
    n474,
    n1366
  );


  nor
  g1813
  (
    n1932,
    n1248,
    n347,
    n386,
    n1738
  );


  nor
  g1814
  (
    n1916,
    n1673,
    n436,
    n1646,
    n1598
  );


  xnor
  g1815
  (
    n1957,
    n313,
    n1515,
    n1546,
    n1324
  );


  nand
  g1816
  (
    n1908,
    n1223,
    n1230,
    n1225,
    n445
  );


  xor
  g1817
  (
    n1870,
    n1590,
    n571,
    n334,
    n1231
  );


  xor
  g1818
  (
    n1865,
    n1712,
    n1370,
    n1174,
    n356
  );


  nand
  g1819
  (
    n1852,
    n312,
    n1665,
    n1643,
    n1594
  );


  nor
  g1820
  (
    n1846,
    n398,
    n1310,
    n1554,
    n457
  );


  nand
  g1821
  (
    n1758,
    n314,
    n1279,
    n1325,
    n1658
  );


  xor
  g1822
  (
    n1747,
    n1381,
    n151,
    n1482,
    n469
  );


  or
  g1823
  (
    n1879,
    n1334,
    n1307,
    n1612,
    n1437
  );


  nand
  g1824
  (
    n1800,
    n1393,
    n1512,
    n1292,
    n1731
  );


  nand
  g1825
  (
    n1962,
    n527,
    n1733,
    n1265,
    n1450
  );


  or
  g1826
  (
    n1862,
    n397,
    n1697,
    n1592,
    n510
  );


  xor
  g1827
  (
    n1873,
    n1470,
    n554,
    n1345,
    n565
  );


  or
  g1828
  (
    n1869,
    n1474,
    n1367,
    n569,
    n1390
  );


  xor
  g1829
  (
    n1816,
    n1168,
    n1167,
    n1346,
    n706
  );


  and
  g1830
  (
    n1924,
    n400,
    n1689,
    n1566,
    n320
  );


  and
  g1831
  (
    n1913,
    n476,
    n1456,
    n301,
    n1662
  );


  and
  g1832
  (
    n1756,
    n1216,
    n302,
    n428,
    n502
  );


  nor
  g1833
  (
    n1868,
    n1221,
    n508,
    n1290,
    n1264
  );


  nand
  g1834
  (
    n1830,
    n559,
    n339,
    n576,
    n506
  );


  nor
  g1835
  (
    n1948,
    n1442,
    n1236,
    n1691,
    n151
  );


  xor
  g1836
  (
    n1823,
    n584,
    n1648,
    n433,
    n1642
  );


  and
  g1837
  (
    n1763,
    n454,
    n531,
    n1180,
    n522
  );


  and
  g1838
  (
    n1918,
    n450,
    n435,
    n1418,
    n413
  );


  nand
  g1839
  (
    n1923,
    n578,
    n1321,
    n432,
    n1344
  );


  nand
  g1840
  (
    n1950,
    n1430,
    n473,
    n1663,
    n420
  );


  nor
  g1841
  (
    n1820,
    n1395,
    n1559,
    n1407,
    n353
  );


  xnor
  g1842
  (
    n1940,
    n1169,
    n1163,
    n1525,
    n1331
  );


  xnor
  g1843
  (
    n1855,
    n524,
    n1250,
    n1149,
    n392
  );


  nor
  g1844
  (
    n1896,
    n460,
    n1141,
    n1194,
    n1514
  );


  and
  g1845
  (
    n1914,
    n1507,
    n501,
    n1630,
    n563
  );


  or
  g1846
  (
    n1783,
    n1208,
    n1609,
    n453,
    n1357
  );


  nand
  g1847
  (
    n1955,
    n1706,
    n1435,
    n1649,
    n1187
  );


  xor
  g1848
  (
    n1802,
    n1661,
    n1659,
    n500,
    n1579
  );


  and
  g1849
  (
    n1788,
    n1519,
    n1563,
    n549,
    n1588
  );


  or
  g1850
  (
    n1892,
    n1493,
    n568,
    n1297,
    n410
  );


  nor
  g1851
  (
    n1938,
    n354,
    n1622,
    n1644,
    n1246
  );


  or
  g1852
  (
    n1777,
    n1151,
    n1140,
    n1322,
    n1340
  );


  xnor
  g1853
  (
    n1902,
    n1543,
    n1639,
    n466,
    n297
  );


  or
  g1854
  (
    n1951,
    n1404,
    n358,
    n409,
    n1522
  );


  or
  g1855
  (
    n1835,
    n1276,
    n1261,
    n1281,
    n1432
  );


  nand
  g1856
  (
    n1952,
    n387,
    n1637,
    n332,
    n349
  );


  nor
  g1857
  (
    n1825,
    n331,
    n492,
    n1567,
    n355
  );


  or
  g1858
  (
    n1909,
    n1471,
    n1170,
    n380,
    n1433
  );


  and
  g1859
  (
    n1751,
    n1604,
    n1597,
    n477,
    n343
  );


  xor
  g1860
  (
    n1922,
    n1486,
    n1707,
    n1599,
    n1670
  );


  nand
  g1861
  (
    n1805,
    n442,
    n1671,
    n1708,
    n1615
  );


  or
  g1862
  (
    n1925,
    n1626,
    n333,
    n396,
    n505
  );


  nand
  g1863
  (
    n1933,
    n1529,
    n1729,
    n319,
    n516
  );


  nand
  g1864
  (
    n1775,
    n494,
    n1191,
    n1354,
    n517
  );


  xnor
  g1865
  (
    n1818,
    n1318,
    n1595,
    n1572,
    n1197
  );


  nand
  g1866
  (
    n1878,
    n1249,
    n486,
    n311,
    n1428
  );


  xor
  g1867
  (
    n1772,
    n529,
    n513,
    n487,
    n1349
  );


  xnor
  g1868
  (
    n1946,
    n426,
    n1182,
    n1270,
    n1569
  );


  nand
  g1869
  (
    n1753,
    n1539,
    n1302,
    n1309,
    n1524
  );


  xnor
  g1870
  (
    n1893,
    n1202,
    n1343,
    n425,
    n1172
  );


  nor
  g1871
  (
    n1819,
    n1142,
    n412,
    n1458,
    n1401
  );


  xnor
  g1872
  (
    n1781,
    n1415,
    n1723,
    n1229,
    n1701
  );


  xnor
  g1873
  (
    n1813,
    n485,
    n1584,
    n1147,
    n1544
  );


  nor
  g1874
  (
    n1793,
    n381,
    n1145,
    n422,
    n1580
  );


  or
  g1875
  (
    n1817,
    n395,
    n1274,
    n1410,
    n1311
  );


  nand
  g1876
  (
    n1947,
    n1711,
    n326,
    n491,
    n1419
  );


  nor
  g1877
  (
    n1740,
    n1542,
    n1721,
    n1238,
    n577
  );


  xor
  g1878
  (
    n1748,
    n1684,
    n1176,
    n1699,
    n1624
  );


  xor
  g1879
  (
    n1919,
    n1583,
    n1727,
    n1162,
    n1523
  );


  nor
  g1880
  (
    n1821,
    n1196,
    n429,
    n1500,
    n1461
  );


  nor
  g1881
  (
    n1880,
    n1445,
    n401,
    n324,
    n439
  );


  or
  g1882
  (
    KeyWire_0_13,
    n1400,
    n351,
    n564,
    n557
  );


  and
  g1883
  (
    n1771,
    n1237,
    n1478,
    n495,
    n364
  );


  nor
  g1884
  (
    n1956,
    n431,
    n1576,
    n1457,
    n533
  );


  xnor
  g1885
  (
    n1875,
    n340,
    n309,
    n480,
    n1417
  );


  nand
  g1886
  (
    n1807,
    n1713,
    n150,
    n567,
    n328
  );


  nor
  g1887
  (
    n1761,
    n1423,
    n1328,
    n1199,
    n1431
  );


  or
  g1888
  (
    n1888,
    n1245,
    n560,
    n470,
    n414
  );


  nor
  g1889
  (
    n1901,
    n1350,
    n1618,
    n1278,
    n1154
  );


  xor
  g1890
  (
    n1930,
    n1638,
    n1411,
    n1405,
    n582
  );


  xor
  g1891
  (
    n1845,
    n402,
    n585,
    n1429,
    n1651
  );


  nor
  g1892
  (
    n1798,
    n1193,
    n411,
    n1678,
    n327
  );


  and
  g1893
  (
    n1833,
    n1406,
    n346,
    n1449,
    n357
  );


  nor
  g1894
  (
    n1897,
    n1650,
    n462,
    n1704,
    n1285
  );


  nor
  g1895
  (
    n1789,
    n1664,
    n1266,
    n1166,
    n562
  );


  nor
  g1896
  (
    n1762,
    n1269,
    n1565,
    n1558,
    n1571
  );


  nand
  g1897
  (
    n1774,
    n305,
    n1550,
    n1693,
    n1355
  );


  nand
  g1898
  (
    n1841,
    n379,
    n548,
    n511,
    n1228
  );


  or
  g1899
  (
    n1776,
    n1201,
    n1492,
    n507,
    n362
  );


  nor
  g1900
  (
    n1794,
    n371,
    n1371,
    n1205,
    n1312
  );


  xnor
  g1901
  (
    n1856,
    n1481,
    n1214,
    n1146,
    n440
  );


  xnor
  g1902
  (
    n1883,
    n403,
    n1183,
    n1685,
    n1700
  );


  nor
  g1903
  (
    n1859,
    n1294,
    n1690,
    n1375,
    n424
  );


  nand
  g1904
  (
    n1890,
    n448,
    n1282,
    n497,
    n484
  );


  or
  g1905
  (
    n1822,
    n1144,
    n1645,
    n1702,
    n1239
  );


  nor
  g1906
  (
    n1801,
    n1610,
    n1719,
    n1362,
    n570
  );


  or
  g1907
  (
    n1826,
    n1373,
    n467,
    n1222,
    n310
  );


  xnor
  g1908
  (
    n1779,
    n1686,
    n1660,
    n475,
    n1260
  );


  nand
  g1909
  (
    n1796,
    n1207,
    n1591,
    n329,
    n1392
  );


  or
  g1910
  (
    n1945,
    n1364,
    n1737,
    n1181,
    n498
  );


  nand
  g1911
  (
    n1935,
    n545,
    n1385,
    n1655,
    n459
  );


  xor
  g1912
  (
    n1910,
    n361,
    n556,
    n1399,
    n1455
  );


  xnor
  g1913
  (
    n1847,
    n575,
    n1188,
    n1574,
    n1386
  );


  or
  g1914
  (
    n1766,
    n534,
    n1511,
    n1531,
    n1271
  );


  nor
  g1915
  (
    n1898,
    n1596,
    n1736,
    n1679,
    n552
  );


  or
  g1916
  (
    n1958,
    n323,
    n1301,
    n1675,
    n419
  );


  nor
  g1917
  (
    n1939,
    n1668,
    n1377,
    n1564,
    n1204
  );


  nor
  g1918
  (
    n1876,
    n1568,
    n1475,
    n378,
    n1536
  );


  or
  g1919
  (
    n1943,
    n1175,
    n1533,
    n1185,
    n1634
  );


  xor
  g1920
  (
    n1944,
    n543,
    n1463,
    n1422,
    n532
  );


  nand
  g1921
  (
    n1754,
    n555,
    n446,
    n370,
    n1666
  );


  and
  g1922
  (
    n1884,
    n515,
    n1496,
    n1698,
    n1374
  );


  and
  g1923
  (
    n1755,
    n1382,
    n1179,
    n1485,
    n447
  );


  or
  g1924
  (
    n1739,
    n458,
    n1494,
    n367,
    n546
  );


  nor
  g1925
  (
    n1850,
    n471,
    n1720,
    n352,
    n1379
  );


  and
  g1926
  (
    n1853,
    n1336,
    n514,
    n1158,
    n1262
  );


  nor
  g1927
  (
    n1882,
    n1483,
    n1402,
    n1372,
    n481
  );


  or
  g1928
  (
    n1812,
    n337,
    n1560,
    n1414,
    n1293
  );


  nor
  g1929
  (
    n1872,
    n1484,
    n417,
    n1304,
    n1688
  );


  nor
  g1930
  (
    n2014,
    n1802,
    n1892,
    n1913,
    n1849
  );


  nand
  g1931
  (
    n1978,
    n1767,
    n1805,
    n1751,
    n1877
  );


  and
  g1932
  (
    n2016,
    n1899,
    n1939,
    n1782,
    n1831
  );


  nand
  g1933
  (
    n2015,
    n1862,
    n1911,
    n1932,
    n1827
  );


  and
  g1934
  (
    n2012,
    n1817,
    n1902,
    n1914,
    n1785
  );


  nor
  g1935
  (
    n2009,
    n1920,
    n1840,
    n1953,
    n1949
  );


  nand
  g1936
  (
    n2017,
    n1850,
    n1740,
    n1834,
    n1815
  );


  or
  g1937
  (
    n1998,
    n1837,
    n1762,
    n1739,
    n1886
  );


  nor
  g1938
  (
    n1970,
    n1833,
    n1763,
    n1760,
    n1947
  );


  xnor
  g1939
  (
    n1984,
    n1957,
    n1803,
    n1883,
    n1746
  );


  xnor
  g1940
  (
    n1976,
    n1839,
    n1942,
    n1761,
    n1934
  );


  xnor
  g1941
  (
    n2007,
    n1943,
    n1797,
    n1859,
    n1874
  );


  nand
  g1942
  (
    n2008,
    n1770,
    n1845,
    n1878,
    n1853
  );


  xor
  g1943
  (
    n1972,
    n1756,
    n1855,
    n1945,
    n1844
  );


  xnor
  g1944
  (
    n1996,
    n1961,
    n1933,
    n1868,
    n1959
  );


  xnor
  g1945
  (
    n1988,
    n1876,
    n1822,
    n1880,
    n1752
  );


  or
  g1946
  (
    n2010,
    n1848,
    n1935,
    n1937,
    n1944
  );


  xor
  g1947
  (
    n2011,
    n1956,
    n1888,
    n1931,
    n1808
  );


  nor
  g1948
  (
    n1989,
    n1893,
    n1768,
    n1936,
    n1904
  );


  and
  g1949
  (
    n2013,
    n1789,
    n1940,
    n1794,
    n1783
  );


  nor
  g1950
  (
    n2000,
    n1766,
    n1791,
    n1869,
    n1809
  );


  xnor
  g1951
  (
    n1999,
    n1830,
    n1912,
    n1918,
    n1922
  );


  nor
  g1952
  (
    n1975,
    n1753,
    n1865,
    n1744,
    n1851
  );


  xnor
  g1953
  (
    n1991,
    n1901,
    n1941,
    n1796,
    n1842
  );


  nor
  g1954
  (
    n1971,
    n1800,
    n1798,
    n1925,
    n1905
  );


  nor
  g1955
  (
    n1993,
    n1758,
    n1906,
    n1929,
    n1769
  );


  or
  g1956
  (
    n1981,
    n1743,
    n1780,
    n1872,
    n1801
  );


  xnor
  g1957
  (
    n1967,
    n1856,
    n1776,
    n1821,
    n1793
  );


  nand
  g1958
  (
    KeyWire_0_7,
    n1788,
    n1861,
    n1806,
    n1835
  );


  nor
  g1959
  (
    n2004,
    n1896,
    n1747,
    n1928,
    n1773
  );


  xor
  g1960
  (
    n1966,
    n1887,
    n1813,
    n1759,
    n1807
  );


  and
  g1961
  (
    n2018,
    n1749,
    n1757,
    n1907,
    n1946
  );


  nand
  g1962
  (
    n1980,
    n1960,
    n1819,
    n1777,
    n1864
  );


  xnor
  g1963
  (
    n2005,
    n1814,
    n1921,
    n1854,
    n1919
  );


  or
  g1964
  (
    n1986,
    n1898,
    n1951,
    n1950,
    n1910
  );


  nor
  g1965
  (
    n1995,
    n1870,
    n1952,
    n1741,
    n1779
  );


  or
  g1966
  (
    n1994,
    n1897,
    n1875,
    n1765,
    n1908
  );


  nor
  g1967
  (
    n1964,
    n1867,
    n1841,
    n1786,
    n1812
  );


  or
  g1968
  (
    n2003,
    n1852,
    n1954,
    n1818,
    n1863
  );


  xor
  g1969
  (
    n1985,
    n1778,
    n1832,
    n1771,
    n1894
  );


  xnor
  g1970
  (
    n1982,
    n1775,
    n1926,
    n1847,
    n1917
  );


  xor
  g1971
  (
    n1990,
    n1909,
    n1900,
    n1804,
    n1890
  );


  and
  g1972
  (
    n2006,
    n1916,
    n1774,
    n1858,
    n1781
  );


  xnor
  g1973
  (
    n1973,
    n1799,
    n1879,
    n1784,
    n1824
  );


  nor
  g1974
  (
    n1963,
    n1825,
    n1857,
    n1930,
    n1871
  );


  nand
  g1975
  (
    n1992,
    n1792,
    n1828,
    n1955,
    n1829
  );


  and
  g1976
  (
    n1983,
    n1843,
    n1866,
    n1795,
    n1754
  );


  or
  g1977
  (
    n1979,
    n1895,
    n1903,
    n1924,
    n1881
  );


  and
  g1978
  (
    n1974,
    n1742,
    n1823,
    n1772,
    n1826
  );


  xor
  g1979
  (
    n2001,
    n1873,
    n1836,
    n1889,
    n1820
  );


  xnor
  g1980
  (
    n1987,
    n1927,
    n1962,
    n1846,
    n1764
  );


  xor
  g1981
  (
    n1965,
    n1882,
    n1787,
    n1938,
    n1958
  );


  xor
  g1982
  (
    n1968,
    n1810,
    n1755,
    n1885,
    n1790
  );


  or
  g1983
  (
    n1997,
    n1811,
    n1915,
    n1860,
    n1838
  );


  or
  g1984
  (
    n1977,
    n1923,
    n1748,
    n1750,
    n1884
  );


  nor
  g1985
  (
    n2002,
    n1891,
    n1816,
    n1745,
    n1948
  );


  nor
  g1986
  (
    n2020,
    n2016,
    n2014,
    n1983,
    n1974
  );


  xnor
  g1987
  (
    n2022,
    n2003,
    n1992,
    n1995,
    n1998
  );


  nor
  g1988
  (
    n2021,
    n1963,
    n2013,
    n1999,
    n1981
  );


  and
  g1989
  (
    n2024,
    n1982,
    n2010,
    n1969,
    n1965
  );


  or
  g1990
  (
    n2028,
    n1977,
    n1964,
    n1987,
    n1985
  );


  xnor
  g1991
  (
    n2026,
    n1997,
    n2004,
    n2008,
    n1973
  );


  nor
  g1992
  (
    n2025,
    n1968,
    n1978,
    n1988,
    n1986
  );


  nor
  g1993
  (
    n2029,
    n1972,
    n1990,
    n2005,
    n1993
  );


  or
  g1994
  (
    n2019,
    n2006,
    n2012,
    n1967,
    n1970
  );


  xor
  g1995
  (
    n2027,
    n1966,
    n1991,
    n1994,
    n1989
  );


  and
  g1996
  (
    n2031,
    n2009,
    n1975,
    n2015,
    n2017
  );


  and
  g1997
  (
    n2023,
    n1984,
    n1979,
    n2000,
    n1996
  );


  xor
  g1998
  (
    n2032,
    n1980,
    n2007,
    n2018,
    n2001
  );


  or
  g1999
  (
    n2030,
    n1971,
    n1976,
    n2011,
    n2002
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n191,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1682,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n107,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n187,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n583,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1472,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1579,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1969,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n892,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n1588,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n661,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n666,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n109,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1752,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n762,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1185,
    KeyNOTWire_0_15
  );


endmodule


