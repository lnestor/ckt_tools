

module Stat_3000_434
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1316,
  n2048,
  n2051,
  n2065,
  n2071,
  n2075,
  n2074,
  n2081,
  n2080,
  n2892,
  n2895,
  n2896,
  n2894,
  n3030,
  n3029,
  n3024,
  n3023,
  n3022,
  n3015,
  n3031,
  n3027,
  n3021,
  n3032,
  n3018,
  n3020,
  n3026,
  n3019,
  n3014,
  n3016,
  n3025,
  n3017,
  n3028,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n1316;
  output n2048;
  output n2051;
  output n2065;
  output n2071;
  output n2075;
  output n2074;
  output n2081;
  output n2080;
  output n2892;
  output n2895;
  output n2896;
  output n2894;
  output n3030;
  output n3029;
  output n3024;
  output n3023;
  output n3022;
  output n3015;
  output n3031;
  output n3027;
  output n3021;
  output n3032;
  output n3018;
  output n3020;
  output n3026;
  output n3019;
  output n3014;
  output n3016;
  output n3025;
  output n3017;
  output n3028;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2049;
  wire n2050;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2072;
  wire n2073;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2893;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  buf
  g0
  (
    n149,
    n30
  );


  buf
  g1
  (
    n40,
    n21
  );


  buf
  g2
  (
    n134,
    n10
  );


  not
  g3
  (
    n142,
    n3
  );


  buf
  g4
  (
    n53,
    n15
  );


  buf
  g5
  (
    n54,
    n19
  );


  not
  g6
  (
    n60,
    n15
  );


  not
  g7
  (
    n58,
    n6
  );


  buf
  g8
  (
    n153,
    n25
  );


  buf
  g9
  (
    n104,
    n5
  );


  not
  g10
  (
    n110,
    n20
  );


  buf
  g11
  (
    n70,
    n4
  );


  not
  g12
  (
    n85,
    n8
  );


  buf
  g13
  (
    n99,
    n7
  );


  buf
  g14
  (
    n97,
    n20
  );


  not
  g15
  (
    n79,
    n3
  );


  buf
  g16
  (
    n124,
    n13
  );


  buf
  g17
  (
    n117,
    n13
  );


  not
  g18
  (
    n74,
    n2
  );


  buf
  g19
  (
    n137,
    n21
  );


  buf
  g20
  (
    n90,
    n22
  );


  not
  g21
  (
    n62,
    n10
  );


  not
  g22
  (
    n100,
    n5
  );


  buf
  g23
  (
    n86,
    n7
  );


  not
  g24
  (
    n92,
    n10
  );


  buf
  g25
  (
    n47,
    n32
  );


  not
  g26
  (
    n82,
    n9
  );


  not
  g27
  (
    n154,
    n27
  );


  not
  g28
  (
    n71,
    n2
  );


  buf
  g29
  (
    n157,
    n25
  );


  buf
  g30
  (
    n101,
    n1
  );


  not
  g31
  (
    n135,
    n26
  );


  not
  g32
  (
    n93,
    n28
  );


  not
  g33
  (
    n141,
    n21
  );


  not
  g34
  (
    n108,
    n13
  );


  buf
  g35
  (
    n75,
    n12
  );


  not
  g36
  (
    n143,
    n23
  );


  buf
  g37
  (
    n42,
    n29
  );


  buf
  g38
  (
    n50,
    n27
  );


  buf
  g39
  (
    n35,
    n22
  );


  not
  g40
  (
    n129,
    n2
  );


  not
  g41
  (
    n45,
    n7
  );


  not
  g42
  (
    n144,
    n31
  );


  buf
  g43
  (
    n120,
    n14
  );


  buf
  g44
  (
    n147,
    n15
  );


  buf
  g45
  (
    n111,
    n17
  );


  not
  g46
  (
    n106,
    n11
  );


  buf
  g47
  (
    n160,
    n14
  );


  not
  g48
  (
    n132,
    n16
  );


  buf
  g49
  (
    n72,
    n31
  );


  buf
  g50
  (
    n145,
    n10
  );


  buf
  g51
  (
    n121,
    n29
  );


  buf
  g52
  (
    n33,
    n24
  );


  not
  g53
  (
    n68,
    n8
  );


  buf
  g54
  (
    n76,
    n16
  );


  buf
  g55
  (
    n119,
    n18
  );


  not
  g56
  (
    n150,
    n17
  );


  buf
  g57
  (
    n64,
    n11
  );


  buf
  g58
  (
    n146,
    n19
  );


  buf
  g59
  (
    n34,
    n3
  );


  buf
  g60
  (
    n148,
    n24
  );


  not
  g61
  (
    n98,
    n17
  );


  not
  g62
  (
    n39,
    n28
  );


  buf
  g63
  (
    n122,
    n9
  );


  buf
  g64
  (
    n123,
    n32
  );


  buf
  g65
  (
    n112,
    n22
  );


  buf
  g66
  (
    n115,
    n23
  );


  not
  g67
  (
    n52,
    n32
  );


  buf
  g68
  (
    n140,
    n13
  );


  buf
  g69
  (
    n125,
    n15
  );


  buf
  g70
  (
    n65,
    n5
  );


  not
  g71
  (
    n38,
    n26
  );


  buf
  g72
  (
    n114,
    n19
  );


  not
  g73
  (
    n77,
    n27
  );


  not
  g74
  (
    n84,
    n5
  );


  buf
  g75
  (
    n118,
    n28
  );


  not
  g76
  (
    n113,
    n6
  );


  not
  g77
  (
    n44,
    n6
  );


  buf
  g78
  (
    n67,
    n8
  );


  not
  g79
  (
    n158,
    n22
  );


  not
  g80
  (
    n51,
    n1
  );


  buf
  g81
  (
    n151,
    n21
  );


  buf
  g82
  (
    n49,
    n4
  );


  buf
  g83
  (
    n152,
    n26
  );


  not
  g84
  (
    n87,
    n31
  );


  not
  g85
  (
    n109,
    n11
  );


  not
  g86
  (
    n37,
    n18
  );


  not
  g87
  (
    n46,
    n16
  );


  not
  g88
  (
    n116,
    n4
  );


  buf
  g89
  (
    n131,
    n20
  );


  buf
  g90
  (
    n127,
    n18
  );


  not
  g91
  (
    n103,
    n25
  );


  not
  g92
  (
    n126,
    n2
  );


  buf
  g93
  (
    n94,
    n9
  );


  buf
  g94
  (
    n83,
    n9
  );


  not
  g95
  (
    n59,
    n30
  );


  buf
  g96
  (
    n155,
    n29
  );


  not
  g97
  (
    n81,
    n29
  );


  not
  g98
  (
    n57,
    n23
  );


  not
  g99
  (
    n69,
    n3
  );


  buf
  g100
  (
    n156,
    n1
  );


  buf
  g101
  (
    n78,
    n7
  );


  not
  g102
  (
    n89,
    n14
  );


  not
  g103
  (
    n43,
    n12
  );


  buf
  g104
  (
    n80,
    n28
  );


  buf
  g105
  (
    n105,
    n32
  );


  not
  g106
  (
    n130,
    n26
  );


  not
  g107
  (
    n63,
    n18
  );


  not
  g108
  (
    KeyWire_0_11,
    n31
  );


  buf
  g109
  (
    n41,
    n23
  );


  not
  g110
  (
    n138,
    n4
  );


  not
  g111
  (
    n133,
    n14
  );


  buf
  g112
  (
    n55,
    n11
  );


  not
  g113
  (
    n66,
    n27
  );


  not
  g114
  (
    n48,
    n30
  );


  buf
  g115
  (
    n61,
    n1
  );


  not
  g116
  (
    n96,
    n6
  );


  buf
  g117
  (
    n107,
    n16
  );


  buf
  g118
  (
    n102,
    n12
  );


  buf
  g119
  (
    n73,
    n24
  );


  buf
  g120
  (
    n36,
    n30
  );


  buf
  g121
  (
    n128,
    n25
  );


  not
  g122
  (
    n95,
    n8
  );


  not
  g123
  (
    n56,
    n20
  );


  buf
  g124
  (
    n136,
    n24
  );


  not
  g125
  (
    n159,
    n17
  );


  buf
  g126
  (
    n91,
    n12
  );


  not
  g127
  (
    n139,
    n19
  );


  not
  g128
  (
    n389,
    n41
  );


  buf
  g129
  (
    n445,
    n140
  );


  not
  g130
  (
    n503,
    n138
  );


  not
  g131
  (
    n330,
    n52
  );


  buf
  g132
  (
    n638,
    n71
  );


  buf
  g133
  (
    n277,
    n49
  );


  buf
  g134
  (
    n343,
    n71
  );


  buf
  g135
  (
    n496,
    n142
  );


  not
  g136
  (
    n208,
    n100
  );


  not
  g137
  (
    n339,
    n110
  );


  buf
  g138
  (
    n164,
    n101
  );


  buf
  g139
  (
    n593,
    n136
  );


  not
  g140
  (
    n667,
    n130
  );


  not
  g141
  (
    n415,
    n152
  );


  buf
  g142
  (
    n669,
    n53
  );


  buf
  g143
  (
    n295,
    n125
  );


  not
  g144
  (
    n449,
    n145
  );


  buf
  g145
  (
    n641,
    n48
  );


  buf
  g146
  (
    n314,
    n77
  );


  not
  g147
  (
    n434,
    n153
  );


  buf
  g148
  (
    n554,
    n42
  );


  buf
  g149
  (
    n644,
    n53
  );


  buf
  g150
  (
    n300,
    n103
  );


  not
  g151
  (
    n358,
    n152
  );


  buf
  g152
  (
    n285,
    n68
  );


  buf
  g153
  (
    n359,
    n90
  );


  buf
  g154
  (
    n211,
    n99
  );


  buf
  g155
  (
    n301,
    n50
  );


  buf
  g156
  (
    n501,
    n35
  );


  not
  g157
  (
    n258,
    n112
  );


  not
  g158
  (
    n469,
    n117
  );


  not
  g159
  (
    n625,
    n158
  );


  not
  g160
  (
    n651,
    n124
  );


  buf
  g161
  (
    n630,
    n127
  );


  not
  g162
  (
    n443,
    n124
  );


  buf
  g163
  (
    n601,
    n85
  );


  not
  g164
  (
    n409,
    n149
  );


  not
  g165
  (
    n391,
    n94
  );


  buf
  g166
  (
    n255,
    n90
  );


  not
  g167
  (
    n612,
    n127
  );


  buf
  g168
  (
    n354,
    n88
  );


  buf
  g169
  (
    n231,
    n74
  );


  not
  g170
  (
    n329,
    n91
  );


  buf
  g171
  (
    n193,
    n35
  );


  buf
  g172
  (
    n517,
    n61
  );


  buf
  g173
  (
    n221,
    n105
  );


  buf
  g174
  (
    n397,
    n159
  );


  buf
  g175
  (
    n390,
    n92
  );


  buf
  g176
  (
    n523,
    n62
  );


  buf
  g177
  (
    n542,
    n85
  );


  not
  g178
  (
    n332,
    n146
  );


  not
  g179
  (
    n637,
    n57
  );


  buf
  g180
  (
    n666,
    n156
  );


  buf
  g181
  (
    n439,
    n136
  );


  not
  g182
  (
    n514,
    n71
  );


  buf
  g183
  (
    n513,
    n65
  );


  not
  g184
  (
    n336,
    n127
  );


  buf
  g185
  (
    n305,
    n142
  );


  buf
  g186
  (
    n217,
    n141
  );


  not
  g187
  (
    n273,
    n36
  );


  buf
  g188
  (
    n200,
    n76
  );


  buf
  g189
  (
    n440,
    n57
  );


  not
  g190
  (
    n356,
    n50
  );


  not
  g191
  (
    n189,
    n64
  );


  not
  g192
  (
    n518,
    n81
  );


  not
  g193
  (
    n649,
    n115
  );


  not
  g194
  (
    n392,
    n88
  );


  buf
  g195
  (
    n214,
    n73
  );


  buf
  g196
  (
    n576,
    n89
  );


  not
  g197
  (
    n377,
    n140
  );


  not
  g198
  (
    n302,
    n85
  );


  buf
  g199
  (
    n408,
    n128
  );


  buf
  g200
  (
    n410,
    n120
  );


  not
  g201
  (
    n290,
    n108
  );


  not
  g202
  (
    n372,
    n145
  );


  buf
  g203
  (
    n490,
    n52
  );


  not
  g204
  (
    n228,
    n84
  );


  not
  g205
  (
    n163,
    n75
  );


  buf
  g206
  (
    n642,
    n139
  );


  not
  g207
  (
    n448,
    n78
  );


  buf
  g208
  (
    n286,
    n116
  );


  not
  g209
  (
    n324,
    n60
  );


  not
  g210
  (
    n592,
    n44
  );


  buf
  g211
  (
    n253,
    n104
  );


  buf
  g212
  (
    n657,
    n120
  );


  buf
  g213
  (
    n478,
    n39
  );


  buf
  g214
  (
    n369,
    n157
  );


  buf
  g215
  (
    n316,
    n111
  );


  buf
  g216
  (
    n287,
    n47
  );


  not
  g217
  (
    n450,
    n105
  );


  not
  g218
  (
    n639,
    n86
  );


  buf
  g219
  (
    n348,
    n61
  );


  not
  g220
  (
    n432,
    n36
  );


  buf
  g221
  (
    n522,
    n152
  );


  buf
  g222
  (
    n446,
    n65
  );


  buf
  g223
  (
    n237,
    n53
  );


  buf
  g224
  (
    n232,
    n160
  );


  not
  g225
  (
    n325,
    n136
  );


  not
  g226
  (
    n559,
    n131
  );


  not
  g227
  (
    n395,
    n107
  );


  not
  g228
  (
    n210,
    n159
  );


  buf
  g229
  (
    n613,
    n52
  );


  buf
  g230
  (
    n241,
    n143
  );


  buf
  g231
  (
    n321,
    n103
  );


  not
  g232
  (
    n583,
    n66
  );


  not
  g233
  (
    n480,
    n94
  );


  not
  g234
  (
    n174,
    n45
  );


  not
  g235
  (
    n235,
    n70
  );


  not
  g236
  (
    n615,
    n101
  );


  not
  g237
  (
    n203,
    n56
  );


  buf
  g238
  (
    n239,
    n51
  );


  not
  g239
  (
    n291,
    n95
  );


  buf
  g240
  (
    n540,
    n57
  );


  not
  g241
  (
    n247,
    n114
  );


  not
  g242
  (
    n484,
    n76
  );


  not
  g243
  (
    n352,
    n155
  );


  not
  g244
  (
    n606,
    n75
  );


  buf
  g245
  (
    n201,
    n67
  );


  buf
  g246
  (
    n378,
    n75
  );


  not
  g247
  (
    n547,
    n154
  );


  not
  g248
  (
    n624,
    n48
  );


  buf
  g249
  (
    n328,
    n145
  );


  not
  g250
  (
    n527,
    n54
  );


  buf
  g251
  (
    n627,
    n41
  );


  buf
  g252
  (
    n310,
    n116
  );


  buf
  g253
  (
    n257,
    n38
  );


  buf
  g254
  (
    n368,
    n141
  );


  buf
  g255
  (
    n187,
    n69
  );


  buf
  g256
  (
    n171,
    n61
  );


  buf
  g257
  (
    n278,
    n111
  );


  buf
  g258
  (
    n620,
    n153
  );


  not
  g259
  (
    n653,
    n44
  );


  buf
  g260
  (
    n526,
    n46
  );


  not
  g261
  (
    n505,
    n151
  );


  buf
  g262
  (
    n441,
    n119
  );


  buf
  g263
  (
    n197,
    n38
  );


  buf
  g264
  (
    n182,
    n126
  );


  not
  g265
  (
    n584,
    n33
  );


  buf
  g266
  (
    n281,
    n55
  );


  not
  g267
  (
    n212,
    n144
  );


  buf
  g268
  (
    n388,
    n115
  );


  not
  g269
  (
    n347,
    n34
  );


  not
  g270
  (
    n455,
    n82
  );


  not
  g271
  (
    n580,
    n78
  );


  buf
  g272
  (
    n616,
    n141
  );


  buf
  g273
  (
    n313,
    n137
  );


  buf
  g274
  (
    n312,
    n134
  );


  buf
  g275
  (
    n532,
    n148
  );


  not
  g276
  (
    n230,
    n83
  );


  buf
  g277
  (
    n426,
    n36
  );


  not
  g278
  (
    n456,
    n61
  );


  buf
  g279
  (
    n355,
    n88
  );


  not
  g280
  (
    n509,
    n45
  );


  not
  g281
  (
    n394,
    n64
  );


  not
  g282
  (
    n166,
    n83
  );


  buf
  g283
  (
    n553,
    n68
  );


  buf
  g284
  (
    n393,
    n123
  );


  buf
  g285
  (
    n462,
    n101
  );


  buf
  g286
  (
    n672,
    n97
  );


  buf
  g287
  (
    n351,
    n46
  );


  not
  g288
  (
    n419,
    n117
  );


  buf
  g289
  (
    n631,
    n59
  );


  not
  g290
  (
    n566,
    n85
  );


  not
  g291
  (
    n585,
    n117
  );


  not
  g292
  (
    n447,
    n49
  );


  buf
  g293
  (
    n563,
    n94
  );


  buf
  g294
  (
    n402,
    n146
  );


  not
  g295
  (
    n550,
    n95
  );


  not
  g296
  (
    n371,
    n122
  );


  not
  g297
  (
    n383,
    n129
  );


  buf
  g298
  (
    n524,
    n55
  );


  not
  g299
  (
    n646,
    n100
  );


  buf
  g300
  (
    n635,
    n156
  );


  buf
  g301
  (
    n519,
    n68
  );


  not
  g302
  (
    n628,
    n110
  );


  not
  g303
  (
    n299,
    n97
  );


  not
  g304
  (
    n401,
    n91
  );


  not
  g305
  (
    n579,
    n134
  );


  not
  g306
  (
    n474,
    n51
  );


  not
  g307
  (
    n564,
    n104
  );


  buf
  g308
  (
    n655,
    n107
  );


  not
  g309
  (
    n209,
    n103
  );


  buf
  g310
  (
    n417,
    n86
  );


  buf
  g311
  (
    n364,
    n160
  );


  not
  g312
  (
    n233,
    n137
  );


  not
  g313
  (
    n574,
    n144
  );


  not
  g314
  (
    n254,
    n149
  );


  not
  g315
  (
    n226,
    n157
  );


  buf
  g316
  (
    n412,
    n92
  );


  not
  g317
  (
    n340,
    n35
  );


  buf
  g318
  (
    n353,
    n109
  );


  not
  g319
  (
    n413,
    n144
  );


  buf
  g320
  (
    n326,
    n102
  );


  not
  g321
  (
    n650,
    n86
  );


  not
  g322
  (
    n227,
    n108
  );


  buf
  g323
  (
    n344,
    n80
  );


  not
  g324
  (
    n387,
    n66
  );


  not
  g325
  (
    n508,
    n125
  );


  buf
  g326
  (
    n528,
    n66
  );


  buf
  g327
  (
    n497,
    n56
  );


  not
  g328
  (
    n400,
    n120
  );


  not
  g329
  (
    n246,
    n122
  );


  not
  g330
  (
    n327,
    n154
  );


  not
  g331
  (
    n216,
    n87
  );


  not
  g332
  (
    n261,
    n54
  );


  not
  g333
  (
    n489,
    n129
  );


  not
  g334
  (
    n555,
    n131
  );


  not
  g335
  (
    n619,
    n121
  );


  not
  g336
  (
    n640,
    n69
  );


  not
  g337
  (
    n575,
    n73
  );


  buf
  g338
  (
    n168,
    n69
  );


  buf
  g339
  (
    n453,
    n78
  );


  buf
  g340
  (
    n596,
    n49
  );


  not
  g341
  (
    n424,
    n47
  );


  buf
  g342
  (
    n173,
    n139
  );


  not
  g343
  (
    n486,
    n146
  );


  not
  g344
  (
    n176,
    n65
  );


  not
  g345
  (
    n269,
    n113
  );


  not
  g346
  (
    n205,
    n89
  );


  buf
  g347
  (
    n498,
    n67
  );


  buf
  g348
  (
    n483,
    n128
  );


  not
  g349
  (
    n457,
    n123
  );


  buf
  g350
  (
    n403,
    n118
  );


  buf
  g351
  (
    n184,
    n46
  );


  buf
  g352
  (
    n659,
    n109
  );


  not
  g353
  (
    n303,
    n143
  );


  buf
  g354
  (
    n647,
    n56
  );


  not
  g355
  (
    n552,
    n62
  );


  buf
  g356
  (
    n181,
    n47
  );


  not
  g357
  (
    n557,
    n81
  );


  buf
  g358
  (
    n609,
    n113
  );


  not
  g359
  (
    n185,
    n45
  );


  buf
  g360
  (
    n218,
    n79
  );


  buf
  g361
  (
    n495,
    n135
  );


  buf
  g362
  (
    n488,
    n110
  );


  not
  g363
  (
    n538,
    n134
  );


  not
  g364
  (
    n506,
    n126
  );


  buf
  g365
  (
    n345,
    n46
  );


  buf
  g366
  (
    n643,
    n74
  );


  buf
  g367
  (
    n418,
    n72
  );


  not
  g368
  (
    n262,
    n48
  );


  not
  g369
  (
    n591,
    n112
  );


  not
  g370
  (
    n379,
    n89
  );


  not
  g371
  (
    n267,
    n143
  );


  not
  g372
  (
    n454,
    n140
  );


  buf
  g373
  (
    n452,
    n150
  );


  buf
  g374
  (
    n536,
    n87
  );


  buf
  g375
  (
    n420,
    n151
  );


  not
  g376
  (
    n236,
    n69
  );


  not
  g377
  (
    n222,
    n128
  );


  buf
  g378
  (
    n323,
    n146
  );


  buf
  g379
  (
    n274,
    n96
  );


  not
  g380
  (
    n560,
    n90
  );


  not
  g381
  (
    n487,
    n49
  );


  buf
  g382
  (
    n570,
    n129
  );


  buf
  g383
  (
    n341,
    n58
  );


  not
  g384
  (
    n665,
    n94
  );


  buf
  g385
  (
    n265,
    n156
  );


  not
  g386
  (
    n479,
    n82
  );


  buf
  g387
  (
    n468,
    n60
  );


  buf
  g388
  (
    n520,
    n159
  );


  buf
  g389
  (
    n477,
    n105
  );


  buf
  g390
  (
    n636,
    n110
  );


  not
  g391
  (
    n461,
    n98
  );


  buf
  g392
  (
    n442,
    n56
  );


  not
  g393
  (
    n533,
    n152
  );


  buf
  g394
  (
    n319,
    n101
  );


  not
  g395
  (
    n198,
    n109
  );


  not
  g396
  (
    n539,
    n77
  );


  buf
  g397
  (
    n617,
    n102
  );


  buf
  g398
  (
    n296,
    n83
  );


  not
  g399
  (
    n428,
    n65
  );


  not
  g400
  (
    n618,
    n59
  );


  buf
  g401
  (
    n350,
    n107
  );


  buf
  g402
  (
    n365,
    n135
  );


  not
  g403
  (
    n435,
    n128
  );


  not
  g404
  (
    n458,
    n63
  );


  buf
  g405
  (
    n167,
    n40
  );


  not
  g406
  (
    n525,
    n57
  );


  not
  g407
  (
    n362,
    n34
  );


  buf
  g408
  (
    n219,
    n91
  );


  buf
  g409
  (
    n234,
    n64
  );


  not
  g410
  (
    n662,
    n40
  );


  buf
  g411
  (
    n175,
    n99
  );


  not
  g412
  (
    n334,
    n84
  );


  buf
  g413
  (
    n648,
    n70
  );


  not
  g414
  (
    n404,
    n40
  );


  not
  g415
  (
    n475,
    n36
  );


  buf
  g416
  (
    n600,
    n62
  );


  buf
  g417
  (
    n634,
    n119
  );


  not
  g418
  (
    n282,
    n140
  );


  not
  g419
  (
    n521,
    n100
  );


  buf
  g420
  (
    n623,
    n93
  );


  buf
  g421
  (
    n590,
    n134
  );


  not
  g422
  (
    n562,
    n124
  );


  not
  g423
  (
    n614,
    n88
  );


  buf
  g424
  (
    n582,
    n124
  );


  not
  g425
  (
    n386,
    n139
  );


  buf
  g426
  (
    n473,
    n149
  );


  not
  g427
  (
    n658,
    n104
  );


  buf
  g428
  (
    n331,
    n81
  );


  not
  g429
  (
    n206,
    n108
  );


  buf
  g430
  (
    n367,
    n150
  );


  not
  g431
  (
    n288,
    n105
  );


  not
  g432
  (
    n602,
    n102
  );


  buf
  g433
  (
    n491,
    n52
  );


  buf
  g434
  (
    n633,
    n100
  );


  buf
  g435
  (
    n224,
    n41
  );


  buf
  g436
  (
    n169,
    n74
  );


  not
  g437
  (
    n304,
    n72
  );


  buf
  g438
  (
    n283,
    n60
  );


  buf
  g439
  (
    n587,
    n64
  );


  buf
  g440
  (
    n357,
    n153
  );


  buf
  g441
  (
    n306,
    n148
  );


  not
  g442
  (
    n500,
    n129
  );


  buf
  g443
  (
    n346,
    n147
  );


  buf
  g444
  (
    n199,
    n93
  );


  not
  g445
  (
    n380,
    n116
  );


  buf
  g446
  (
    n433,
    n79
  );


  buf
  g447
  (
    n349,
    n108
  );


  buf
  g448
  (
    n406,
    n67
  );


  not
  g449
  (
    n411,
    n132
  );


  not
  g450
  (
    n292,
    n38
  );


  buf
  g451
  (
    n541,
    n34
  );


  buf
  g452
  (
    n178,
    n37
  );


  buf
  g453
  (
    n422,
    n76
  );


  not
  g454
  (
    n196,
    n42
  );


  buf
  g455
  (
    n668,
    n133
  );


  buf
  g456
  (
    n546,
    n45
  );


  not
  g457
  (
    n240,
    n37
  );


  buf
  g458
  (
    n431,
    n66
  );


  buf
  g459
  (
    n252,
    n137
  );


  not
  g460
  (
    n376,
    n43
  );


  buf
  g461
  (
    n573,
    n113
  );


  not
  g462
  (
    n337,
    n135
  );


  not
  g463
  (
    n405,
    n99
  );


  not
  g464
  (
    n317,
    n127
  );


  not
  g465
  (
    n229,
    n147
  );


  buf
  g466
  (
    n511,
    n83
  );


  not
  g467
  (
    n248,
    n153
  );


  buf
  g468
  (
    n581,
    n147
  );


  not
  g469
  (
    n268,
    n121
  );


  not
  g470
  (
    n249,
    n120
  );


  not
  g471
  (
    n507,
    n115
  );


  buf
  g472
  (
    n276,
    n53
  );


  not
  g473
  (
    n482,
    n158
  );


  not
  g474
  (
    n537,
    n115
  );


  buf
  g475
  (
    n543,
    n60
  );


  not
  g476
  (
    n190,
    n59
  );


  buf
  g477
  (
    n396,
    n38
  );


  buf
  g478
  (
    n204,
    n39
  );


  buf
  g479
  (
    n556,
    n119
  );


  buf
  g480
  (
    n607,
    n155
  );


  buf
  g481
  (
    n451,
    n106
  );


  not
  g482
  (
    n597,
    n119
  );


  buf
  g483
  (
    n465,
    n104
  );


  buf
  g484
  (
    n366,
    n54
  );


  buf
  g485
  (
    n629,
    n132
  );


  buf
  g486
  (
    n568,
    n73
  );


  buf
  g487
  (
    n605,
    n125
  );


  buf
  g488
  (
    n586,
    n84
  );


  not
  g489
  (
    n549,
    n81
  );


  not
  g490
  (
    n626,
    n43
  );


  not
  g491
  (
    n567,
    n155
  );


  not
  g492
  (
    n294,
    n138
  );


  not
  g493
  (
    n264,
    n97
  );


  not
  g494
  (
    n476,
    n122
  );


  buf
  g495
  (
    n467,
    n106
  );


  not
  g496
  (
    n162,
    n33
  );


  not
  g497
  (
    n333,
    n130
  );


  buf
  g498
  (
    n244,
    n43
  );


  not
  g499
  (
    n194,
    n126
  );


  buf
  g500
  (
    n275,
    n112
  );


  not
  g501
  (
    n170,
    n82
  );


  buf
  g502
  (
    n611,
    n63
  );


  buf
  g503
  (
    n569,
    n93
  );


  not
  g504
  (
    n338,
    n87
  );


  buf
  g505
  (
    n308,
    n138
  );


  not
  g506
  (
    n280,
    n158
  );


  not
  g507
  (
    n595,
    n71
  );


  not
  g508
  (
    n172,
    n67
  );


  not
  g509
  (
    n385,
    n51
  );


  not
  g510
  (
    n504,
    n150
  );


  buf
  g511
  (
    n608,
    n156
  );


  buf
  g512
  (
    n284,
    n106
  );


  not
  g513
  (
    n438,
    n63
  );


  buf
  g514
  (
    n515,
    n149
  );


  not
  g515
  (
    n481,
    n112
  );


  not
  g516
  (
    n256,
    n54
  );


  buf
  g517
  (
    n179,
    n58
  );


  not
  g518
  (
    n494,
    n50
  );


  buf
  g519
  (
    n460,
    n95
  );


  not
  g520
  (
    n664,
    n98
  );


  not
  g521
  (
    n363,
    n58
  );


  not
  g522
  (
    n360,
    n75
  );


  not
  g523
  (
    n670,
    n84
  );


  not
  g524
  (
    n444,
    n151
  );


  not
  g525
  (
    n561,
    n35
  );


  not
  g526
  (
    KeyWire_0_12,
    n42
  );


  buf
  g527
  (
    n421,
    n58
  );


  not
  g528
  (
    n407,
    n33
  );


  not
  g529
  (
    n430,
    n126
  );


  buf
  g530
  (
    n272,
    n131
  );


  not
  g531
  (
    n213,
    n70
  );


  buf
  g532
  (
    n263,
    n147
  );


  not
  g533
  (
    n381,
    n138
  );


  not
  g534
  (
    n361,
    n150
  );


  not
  g535
  (
    n289,
    n143
  );


  buf
  g536
  (
    n466,
    n103
  );


  not
  g537
  (
    n250,
    n98
  );


  not
  g538
  (
    n207,
    n109
  );


  buf
  g539
  (
    n621,
    n160
  );


  not
  g540
  (
    n502,
    n68
  );


  not
  g541
  (
    n186,
    n33
  );


  not
  g542
  (
    n335,
    n78
  );


  buf
  g543
  (
    n188,
    n50
  );


  buf
  g544
  (
    n297,
    n80
  );


  not
  g545
  (
    n373,
    n118
  );


  buf
  g546
  (
    n622,
    n123
  );


  buf
  g547
  (
    n251,
    n121
  );


  not
  g548
  (
    n656,
    n132
  );


  buf
  g549
  (
    n598,
    n114
  );


  not
  g550
  (
    n183,
    n96
  );


  buf
  g551
  (
    n177,
    n91
  );


  not
  g552
  (
    n558,
    n96
  );


  buf
  g553
  (
    n245,
    n142
  );


  buf
  g554
  (
    n382,
    n130
  );


  buf
  g555
  (
    n423,
    n160
  );


  buf
  g556
  (
    n548,
    n121
  );


  buf
  g557
  (
    n493,
    n90
  );


  not
  g558
  (
    n499,
    n102
  );


  not
  g559
  (
    n534,
    n73
  );


  not
  g560
  (
    n399,
    n155
  );


  not
  g561
  (
    n603,
    n63
  );


  not
  g562
  (
    n671,
    n142
  );


  buf
  g563
  (
    n565,
    n89
  );


  not
  g564
  (
    n242,
    n114
  );


  buf
  g565
  (
    n293,
    n72
  );


  buf
  g566
  (
    n663,
    n107
  );


  not
  g567
  (
    n374,
    n51
  );


  not
  g568
  (
    n271,
    n79
  );


  buf
  g569
  (
    n191,
    n158
  );


  buf
  g570
  (
    n654,
    n113
  );


  buf
  g571
  (
    n238,
    n70
  );


  not
  g572
  (
    n315,
    n37
  );


  not
  g573
  (
    n578,
    n48
  );


  buf
  g574
  (
    n425,
    n72
  );


  not
  g575
  (
    n298,
    n80
  );


  buf
  g576
  (
    n551,
    n98
  );


  buf
  g577
  (
    n599,
    n154
  );


  buf
  g578
  (
    n279,
    n117
  );


  not
  g579
  (
    n572,
    n44
  );


  not
  g580
  (
    n309,
    n137
  );


  buf
  g581
  (
    n223,
    n118
  );


  buf
  g582
  (
    n320,
    n44
  );


  buf
  g583
  (
    n588,
    n154
  );


  not
  g584
  (
    n195,
    n41
  );


  not
  g585
  (
    n516,
    n34
  );


  not
  g586
  (
    n202,
    n136
  );


  not
  g587
  (
    n660,
    n77
  );


  not
  g588
  (
    n311,
    n148
  );


  not
  g589
  (
    n370,
    n122
  );


  not
  g590
  (
    n318,
    n59
  );


  buf
  g591
  (
    n436,
    n80
  );


  buf
  g592
  (
    n571,
    n77
  );


  buf
  g593
  (
    n270,
    n55
  );


  buf
  g594
  (
    n463,
    n157
  );


  buf
  g595
  (
    n645,
    n96
  );


  buf
  g596
  (
    n604,
    n42
  );


  buf
  g597
  (
    n471,
    n111
  );


  not
  g598
  (
    n165,
    n106
  );


  not
  g599
  (
    n225,
    n92
  );


  buf
  g600
  (
    n414,
    n118
  );


  buf
  g601
  (
    n531,
    n40
  );


  not
  g602
  (
    n342,
    n82
  );


  buf
  g603
  (
    n510,
    n74
  );


  not
  g604
  (
    n259,
    n79
  );


  not
  g605
  (
    n161,
    n135
  );


  not
  g606
  (
    n464,
    n133
  );


  buf
  g607
  (
    n416,
    n55
  );


  not
  g608
  (
    n215,
    n62
  );


  not
  g609
  (
    n459,
    n133
  );


  buf
  g610
  (
    n485,
    n141
  );


  buf
  g611
  (
    n180,
    n47
  );


  buf
  g612
  (
    n307,
    n99
  );


  buf
  g613
  (
    n632,
    n97
  );


  not
  g614
  (
    n529,
    n39
  );


  buf
  g615
  (
    n472,
    n132
  );


  buf
  g616
  (
    n266,
    n87
  );


  not
  g617
  (
    n594,
    n130
  );


  not
  g618
  (
    n652,
    n43
  );


  not
  g619
  (
    n470,
    n114
  );


  not
  g620
  (
    n437,
    n131
  );


  buf
  g621
  (
    n384,
    n39
  );


  buf
  g622
  (
    n398,
    n37
  );


  not
  g623
  (
    n429,
    n133
  );


  not
  g624
  (
    n322,
    n93
  );


  not
  g625
  (
    n544,
    n144
  );


  buf
  g626
  (
    n220,
    n116
  );


  buf
  g627
  (
    n243,
    n95
  );


  not
  g628
  (
    n530,
    n123
  );


  buf
  g629
  (
    n492,
    n125
  );


  not
  g630
  (
    n577,
    n151
  );


  buf
  g631
  (
    n610,
    n145
  );


  not
  g632
  (
    n375,
    n111
  );


  buf
  g633
  (
    n535,
    n76
  );


  buf
  g634
  (
    n589,
    n148
  );


  buf
  g635
  (
    n427,
    n86
  );


  buf
  g636
  (
    n260,
    n159
  );


  buf
  g637
  (
    n545,
    n157
  );


  buf
  g638
  (
    n512,
    n139
  );


  buf
  g639
  (
    n661,
    n92
  );


  not
  g640
  (
    n900,
    n363
  );


  not
  g641
  (
    n948,
    n488
  );


  buf
  g642
  (
    n1408,
    n269
  );


  buf
  g643
  (
    n1624,
    n321
  );


  not
  g644
  (
    n1229,
    n223
  );


  not
  g645
  (
    n1015,
    n186
  );


  not
  g646
  (
    n1199,
    n313
  );


  not
  g647
  (
    n1145,
    n234
  );


  not
  g648
  (
    n1717,
    n372
  );


  not
  g649
  (
    n1122,
    n418
  );


  buf
  g650
  (
    n1186,
    n300
  );


  not
  g651
  (
    n1604,
    n398
  );


  not
  g652
  (
    n896,
    n440
  );


  buf
  g653
  (
    n904,
    n282
  );


  not
  g654
  (
    n882,
    n164
  );


  not
  g655
  (
    n1739,
    n519
  );


  buf
  g656
  (
    n1582,
    n237
  );


  buf
  g657
  (
    n1388,
    n344
  );


  buf
  g658
  (
    n1305,
    n408
  );


  not
  g659
  (
    n1528,
    n617
  );


  buf
  g660
  (
    n1072,
    n272
  );


  buf
  g661
  (
    n914,
    n437
  );


  buf
  g662
  (
    n1236,
    n373
  );


  buf
  g663
  (
    n1602,
    n622
  );


  buf
  g664
  (
    n814,
    n188
  );


  buf
  g665
  (
    n1466,
    n252
  );


  not
  g666
  (
    n1175,
    n537
  );


  buf
  g667
  (
    n738,
    n543
  );


  buf
  g668
  (
    n1482,
    n182
  );


  buf
  g669
  (
    n1000,
    n618
  );


  not
  g670
  (
    n1143,
    n628
  );


  not
  g671
  (
    n1415,
    n362
  );


  buf
  g672
  (
    n834,
    n593
  );


  not
  g673
  (
    n1046,
    n620
  );


  buf
  g674
  (
    n1068,
    n636
  );


  not
  g675
  (
    n805,
    n466
  );


  buf
  g676
  (
    n1210,
    n511
  );


  buf
  g677
  (
    n1427,
    n392
  );


  buf
  g678
  (
    n1029,
    n628
  );


  buf
  g679
  (
    n1665,
    n204
  );


  not
  g680
  (
    n1153,
    n342
  );


  not
  g681
  (
    n1403,
    n353
  );


  buf
  g682
  (
    n930,
    n625
  );


  buf
  g683
  (
    n815,
    n331
  );


  not
  g684
  (
    n787,
    n605
  );


  buf
  g685
  (
    n1189,
    n263
  );


  not
  g686
  (
    n1348,
    n433
  );


  buf
  g687
  (
    n680,
    n469
  );


  buf
  g688
  (
    n1018,
    n567
  );


  not
  g689
  (
    n1090,
    n184
  );


  buf
  g690
  (
    n843,
    n612
  );


  buf
  g691
  (
    n1457,
    n270
  );


  buf
  g692
  (
    n1276,
    n558
  );


  not
  g693
  (
    n978,
    n443
  );


  not
  g694
  (
    n1540,
    n612
  );


  buf
  g695
  (
    n1643,
    n290
  );


  buf
  g696
  (
    n1462,
    n439
  );


  buf
  g697
  (
    n1592,
    n375
  );


  buf
  g698
  (
    n694,
    n217
  );


  buf
  g699
  (
    n1649,
    n348
  );


  not
  g700
  (
    n869,
    n560
  );


  buf
  g701
  (
    n1343,
    n361
  );


  not
  g702
  (
    n1323,
    n314
  );


  buf
  g703
  (
    n830,
    n640
  );


  buf
  g704
  (
    n1197,
    n214
  );


  buf
  g705
  (
    n1254,
    n255
  );


  not
  g706
  (
    n944,
    n571
  );


  not
  g707
  (
    n1487,
    n467
  );


  buf
  g708
  (
    n731,
    n496
  );


  buf
  g709
  (
    n689,
    n566
  );


  not
  g710
  (
    n1455,
    n338
  );


  buf
  g711
  (
    n1715,
    n201
  );


  buf
  g712
  (
    n730,
    n498
  );


  not
  g713
  (
    n823,
    n239
  );


  buf
  g714
  (
    n1438,
    n278
  );


  not
  g715
  (
    n1631,
    n262
  );


  not
  g716
  (
    n1125,
    n210
  );


  buf
  g717
  (
    n1079,
    n393
  );


  not
  g718
  (
    n1483,
    n227
  );


  buf
  g719
  (
    n1237,
    n431
  );


  buf
  g720
  (
    n1579,
    n363
  );


  not
  g721
  (
    n1746,
    n340
  );


  not
  g722
  (
    n887,
    n288
  );


  buf
  g723
  (
    n691,
    n533
  );


  buf
  g724
  (
    n1431,
    n290
  );


  buf
  g725
  (
    n1569,
    n427
  );


  not
  g726
  (
    n1622,
    n564
  );


  not
  g727
  (
    n1373,
    n595
  );


  buf
  g728
  (
    n746,
    n635
  );


  buf
  g729
  (
    n1545,
    n608
  );


  buf
  g730
  (
    n1283,
    n226
  );


  buf
  g731
  (
    n886,
    n213
  );


  not
  g732
  (
    n862,
    n265
  );


  not
  g733
  (
    n932,
    n592
  );


  not
  g734
  (
    n1391,
    n590
  );


  not
  g735
  (
    n1190,
    n216
  );


  buf
  g736
  (
    n1620,
    n515
  );


  buf
  g737
  (
    n802,
    n457
  );


  not
  g738
  (
    n1084,
    n512
  );


  buf
  g739
  (
    n1508,
    n393
  );


  buf
  g740
  (
    n683,
    n538
  );


  buf
  g741
  (
    n1671,
    n621
  );


  not
  g742
  (
    n1270,
    n214
  );


  not
  g743
  (
    n1085,
    n341
  );


  buf
  g744
  (
    n1273,
    n332
  );


  not
  g745
  (
    n1014,
    n244
  );


  not
  g746
  (
    n1727,
    n228
  );


  buf
  g747
  (
    n1736,
    n502
  );


  not
  g748
  (
    n1365,
    n549
  );


  not
  g749
  (
    n1110,
    n205
  );


  buf
  g750
  (
    n1382,
    n358
  );


  buf
  g751
  (
    n723,
    n592
  );


  not
  g752
  (
    n1439,
    n629
  );


  buf
  g753
  (
    n1633,
    n325
  );


  not
  g754
  (
    n1251,
    n304
  );


  not
  g755
  (
    n1499,
    n518
  );


  not
  g756
  (
    n1514,
    n389
  );


  buf
  g757
  (
    n1241,
    n390
  );


  not
  g758
  (
    n1688,
    n322
  );


  not
  g759
  (
    n1109,
    n232
  );


  not
  g760
  (
    n1686,
    n504
  );


  not
  g761
  (
    n1493,
    n635
  );


  buf
  g762
  (
    n1362,
    n306
  );


  not
  g763
  (
    n726,
    n188
  );


  not
  g764
  (
    n1726,
    n224
  );


  not
  g765
  (
    n1045,
    n544
  );


  not
  g766
  (
    n1676,
    n204
  );


  buf
  g767
  (
    n875,
    n359
  );


  not
  g768
  (
    n724,
    n610
  );


  buf
  g769
  (
    n1291,
    n397
  );


  not
  g770
  (
    n1692,
    n603
  );


  buf
  g771
  (
    n852,
    n579
  );


  not
  g772
  (
    n1004,
    n540
  );


  buf
  g773
  (
    n826,
    n509
  );


  buf
  g774
  (
    n1345,
    n162
  );


  buf
  g775
  (
    n850,
    n446
  );


  buf
  g776
  (
    n1720,
    n550
  );


  buf
  g777
  (
    n854,
    n188
  );


  buf
  g778
  (
    n877,
    n242
  );


  not
  g779
  (
    n808,
    n283
  );


  not
  g780
  (
    n1734,
    n590
  );


  not
  g781
  (
    n1207,
    n616
  );


  buf
  g782
  (
    n1171,
    n166
  );


  not
  g783
  (
    n1695,
    n456
  );


  not
  g784
  (
    n1553,
    n609
  );


  not
  g785
  (
    n903,
    n608
  );


  not
  g786
  (
    n873,
    n200
  );


  not
  g787
  (
    n1627,
    n447
  );


  not
  g788
  (
    n1418,
    n212
  );


  buf
  g789
  (
    n1435,
    n435
  );


  buf
  g790
  (
    n1394,
    n504
  );


  not
  g791
  (
    n1521,
    n585
  );


  buf
  g792
  (
    n1637,
    n234
  );


  not
  g793
  (
    n1541,
    n220
  );


  buf
  g794
  (
    n728,
    n369
  );


  buf
  g795
  (
    n937,
    n588
  );


  buf
  g796
  (
    n1663,
    n484
  );


  buf
  g797
  (
    n1678,
    n510
  );


  not
  g798
  (
    n1269,
    n268
  );


  buf
  g799
  (
    n1081,
    n405
  );


  not
  g800
  (
    n1687,
    n470
  );


  buf
  g801
  (
    n1028,
    n395
  );


  buf
  g802
  (
    n960,
    n453
  );


  not
  g803
  (
    n784,
    n164
  );


  buf
  g804
  (
    n1589,
    n561
  );


  buf
  g805
  (
    n870,
    n417
  );


  buf
  g806
  (
    n1129,
    n199
  );


  buf
  g807
  (
    n1214,
    n667
  );


  buf
  g808
  (
    n1076,
    n602
  );


  not
  g809
  (
    n1165,
    n284
  );


  buf
  g810
  (
    n801,
    n234
  );


  buf
  g811
  (
    n1581,
    n606
  );


  buf
  g812
  (
    n1167,
    n407
  );


  not
  g813
  (
    n1013,
    n633
  );


  buf
  g814
  (
    n1070,
    n565
  );


  not
  g815
  (
    n686,
    n530
  );


  not
  g816
  (
    n758,
    n321
  );


  buf
  g817
  (
    n890,
    n581
  );


  not
  g818
  (
    n1689,
    n363
  );


  buf
  g819
  (
    n773,
    n340
  );


  buf
  g820
  (
    n1211,
    n223
  );


  not
  g821
  (
    n1098,
    n314
  );


  not
  g822
  (
    KeyWire_0_4,
    n598
  );


  not
  g823
  (
    n1096,
    n419
  );


  buf
  g824
  (
    n1326,
    n383
  );


  not
  g825
  (
    n1445,
    n455
  );


  not
  g826
  (
    n1538,
    n225
  );


  not
  g827
  (
    n881,
    n292
  );


  not
  g828
  (
    n1547,
    n213
  );


  not
  g829
  (
    n766,
    n576
  );


  not
  g830
  (
    n1234,
    n310
  );


  buf
  g831
  (
    n1037,
    n283
  );


  buf
  g832
  (
    n692,
    n639
  );


  buf
  g833
  (
    n1747,
    n189
  );


  buf
  g834
  (
    n856,
    n258
  );


  buf
  g835
  (
    n1127,
    n540
  );


  buf
  g836
  (
    n798,
    n667
  );


  buf
  g837
  (
    n969,
    n243
  );


  buf
  g838
  (
    n1477,
    n634
  );


  buf
  g839
  (
    n1616,
    n647
  );


  buf
  g840
  (
    n1465,
    n637
  );


  not
  g841
  (
    n1169,
    n343
  );


  not
  g842
  (
    n1527,
    n258
  );


  not
  g843
  (
    n684,
    n671
  );


  buf
  g844
  (
    n1142,
    n196
  );


  not
  g845
  (
    n866,
    n505
  );


  not
  g846
  (
    n1510,
    n277
  );


  not
  g847
  (
    n1126,
    n410
  );


  buf
  g848
  (
    n1651,
    n387
  );


  buf
  g849
  (
    n1668,
    n582
  );


  not
  g850
  (
    n927,
    n660
  );


  buf
  g851
  (
    n1414,
    n484
  );


  buf
  g852
  (
    n1262,
    n421
  );


  not
  g853
  (
    n999,
    n385
  );


  not
  g854
  (
    n1550,
    n370
  );


  buf
  g855
  (
    n1063,
    n365
  );


  buf
  g856
  (
    n682,
    n601
  );


  buf
  g857
  (
    n1201,
    n275
  );


  buf
  g858
  (
    n1750,
    n286
  );


  buf
  g859
  (
    n1137,
    n438
  );


  not
  g860
  (
    n1342,
    n352
  );


  buf
  g861
  (
    n712,
    n568
  );


  not
  g862
  (
    n1312,
    n197
  );


  buf
  g863
  (
    n1131,
    n231
  );


  not
  g864
  (
    n996,
    n436
  );


  buf
  g865
  (
    n1044,
    n429
  );


  buf
  g866
  (
    n1259,
    n274
  );


  buf
  g867
  (
    n1032,
    n571
  );


  not
  g868
  (
    n1255,
    n582
  );


  not
  g869
  (
    n673,
    n487
  );


  buf
  g870
  (
    n1371,
    n442
  );


  buf
  g871
  (
    n1516,
    n453
  );


  not
  g872
  (
    n1378,
    n207
  );


  buf
  g873
  (
    n983,
    n163
  );


  not
  g874
  (
    KeyWire_0_8,
    n656
  );


  not
  g875
  (
    n1456,
    n493
  );


  buf
  g876
  (
    n1601,
    n555
  );


  buf
  g877
  (
    n1213,
    n331
  );


  not
  g878
  (
    n1011,
    n581
  );


  not
  g879
  (
    n1712,
    n411
  );


  buf
  g880
  (
    n1181,
    n326
  );


  not
  g881
  (
    n1570,
    n600
  );


  not
  g882
  (
    n806,
    n597
  );


  buf
  g883
  (
    n1558,
    n374
  );


  not
  g884
  (
    n1536,
    n556
  );


  buf
  g885
  (
    n1648,
    n524
  );


  not
  g886
  (
    n735,
    n334
  );


  not
  g887
  (
    n1699,
    n542
  );


  buf
  g888
  (
    n1156,
    n171
  );


  buf
  g889
  (
    n1708,
    n238
  );


  not
  g890
  (
    n1603,
    n239
  );


  not
  g891
  (
    n1352,
    n343
  );


  not
  g892
  (
    n1574,
    n480
  );


  buf
  g893
  (
    n1433,
    n248
  );


  buf
  g894
  (
    n1194,
    n226
  );


  buf
  g895
  (
    n1192,
    n241
  );


  not
  g896
  (
    n1467,
    n653
  );


  buf
  g897
  (
    n1621,
    n523
  );


  buf
  g898
  (
    n1667,
    n553
  );


  buf
  g899
  (
    n911,
    n562
  );


  not
  g900
  (
    n816,
    n603
  );


  buf
  g901
  (
    n1200,
    n168
  );


  buf
  g902
  (
    n1022,
    n565
  );


  buf
  g903
  (
    n1390,
    n486
  );


  buf
  g904
  (
    n845,
    n618
  );


  buf
  g905
  (
    n1705,
    n540
  );


  not
  g906
  (
    n1218,
    n654
  );


  not
  g907
  (
    n751,
    n525
  );


  buf
  g908
  (
    n1202,
    n670
  );


  not
  g909
  (
    n936,
    n453
  );


  not
  g910
  (
    n1405,
    n636
  );


  buf
  g911
  (
    n1203,
    n208
  );


  not
  g912
  (
    n1740,
    n395
  );


  not
  g913
  (
    n1025,
    n340
  );


  buf
  g914
  (
    n1718,
    n238
  );


  buf
  g915
  (
    n1074,
    n460
  );


  not
  g916
  (
    n961,
    n231
  );


  buf
  g917
  (
    n1755,
    n282
  );


  not
  g918
  (
    n1010,
    n552
  );


  not
  g919
  (
    n1421,
    n320
  );


  buf
  g920
  (
    n1048,
    n537
  );


  not
  g921
  (
    n1635,
    n423
  );


  buf
  g922
  (
    n1132,
    n557
  );


  not
  g923
  (
    n1441,
    n245
  );


  not
  g924
  (
    n1480,
    n469
  );


  buf
  g925
  (
    n1675,
    n668
  );


  not
  g926
  (
    n796,
    n204
  );


  buf
  g927
  (
    n1400,
    n293
  );


  not
  g928
  (
    n1134,
    n191
  );


  buf
  g929
  (
    n1031,
    n592
  );


  buf
  g930
  (
    n1094,
    n523
  );


  buf
  g931
  (
    n1702,
    n406
  );


  buf
  g932
  (
    n864,
    n358
  );


  buf
  g933
  (
    n1662,
    n483
  );


  buf
  g934
  (
    n1056,
    n599
  );


  buf
  g935
  (
    n1555,
    n591
  );


  buf
  g936
  (
    n1017,
    n343
  );


  not
  g937
  (
    n1092,
    n330
  );


  buf
  g938
  (
    n1488,
    n631
  );


  buf
  g939
  (
    n1151,
    n550
  );


  buf
  g940
  (
    n965,
    n400
  );


  not
  g941
  (
    n963,
    n349
  );


  buf
  g942
  (
    n1425,
    n188
  );


  not
  g943
  (
    n839,
    n326
  );


  buf
  g944
  (
    n1474,
    n505
  );


  buf
  g945
  (
    n1083,
    n658
  );


  buf
  g946
  (
    n788,
    n549
  );


  buf
  g947
  (
    n1544,
    n497
  );


  buf
  g948
  (
    n1288,
    n199
  );


  buf
  g949
  (
    n708,
    n402
  );


  buf
  g950
  (
    n1412,
    n194
  );


  not
  g951
  (
    n702,
    n175
  );


  not
  g952
  (
    n1614,
    n322
  );


  not
  g953
  (
    n1231,
    n167
  );


  not
  g954
  (
    n1120,
    n320
  );


  not
  g955
  (
    n1650,
    n613
  );


  not
  g956
  (
    n1308,
    n405
  );


  not
  g957
  (
    n987,
    n256
  );


  not
  g958
  (
    n1337,
    n318
  );


  not
  g959
  (
    n1006,
    n659
  );


  buf
  g960
  (
    n1728,
    n461
  );


  buf
  g961
  (
    n1461,
    n332
  );


  not
  g962
  (
    n1193,
    n629
  );


  buf
  g963
  (
    n1335,
    n169
  );


  not
  g964
  (
    n1419,
    n533
  );


  not
  g965
  (
    n951,
    n508
  );


  not
  g966
  (
    n1113,
    n326
  );


  buf
  g967
  (
    n1626,
    n470
  );


  not
  g968
  (
    n804,
    n650
  );


  buf
  g969
  (
    n1166,
    n174
  );


  buf
  g970
  (
    n1407,
    n546
  );


  not
  g971
  (
    n1674,
    n478
  );


  buf
  g972
  (
    n1257,
    n517
  );


  not
  g973
  (
    n1500,
    n517
  );


  not
  g974
  (
    n696,
    n568
  );


  buf
  g975
  (
    n827,
    n162
  );


  buf
  g976
  (
    n1443,
    n409
  );


  buf
  g977
  (
    n872,
    n445
  );


  not
  g978
  (
    n1517,
    n567
  );


  buf
  g979
  (
    n1454,
    n594
  );


  not
  g980
  (
    n1141,
    n666
  );


  not
  g981
  (
    KeyWire_0_5,
    n373
  );


  not
  g982
  (
    n1606,
    n179
  );


  buf
  g983
  (
    n835,
    n165
  );


  not
  g984
  (
    n1226,
    n387
  );


  not
  g985
  (
    n876,
    n296
  );


  buf
  g986
  (
    n720,
    n335
  );


  not
  g987
  (
    n952,
    n426
  );


  buf
  g988
  (
    n1178,
    n508
  );


  not
  g989
  (
    n1372,
    n483
  );


  buf
  g990
  (
    n1248,
    n171
  );


  buf
  g991
  (
    n1318,
    n471
  );


  not
  g992
  (
    n1387,
    n482
  );


  buf
  g993
  (
    n1356,
    n515
  );


  buf
  g994
  (
    n1330,
    n359
  );


  not
  g995
  (
    n1507,
    n272
  );


  buf
  g996
  (
    n943,
    n315
  );


  buf
  g997
  (
    n1227,
    n654
  );


  not
  g998
  (
    n1656,
    n530
  );


  buf
  g999
  (
    n1422,
    n190
  );


  buf
  g1000
  (
    n1331,
    n491
  );


  buf
  g1001
  (
    n956,
    n346
  );


  not
  g1002
  (
    n1157,
    n636
  );


  not
  g1003
  (
    n1118,
    n323
  );


  not
  g1004
  (
    n1173,
    n665
  );


  buf
  g1005
  (
    n1685,
    n516
  );


  not
  g1006
  (
    n849,
    n268
  );


  not
  g1007
  (
    n1080,
    n222
  );


  not
  g1008
  (
    n1353,
    n304
  );


  not
  g1009
  (
    n759,
    n304
  );


  not
  g1010
  (
    n878,
    n521
  );


  not
  g1011
  (
    n837,
    n589
  );


  buf
  g1012
  (
    n942,
    n480
  );


  buf
  g1013
  (
    n754,
    n279
  );


  buf
  g1014
  (
    n1473,
    n405
  );


  not
  g1015
  (
    n1180,
    n520
  );


  not
  g1016
  (
    n842,
    n613
  );


  buf
  g1017
  (
    n1583,
    n655
  );


  buf
  g1018
  (
    n1424,
    n412
  );


  buf
  g1019
  (
    n981,
    n230
  );


  not
  g1020
  (
    n1495,
    n210
  );


  buf
  g1021
  (
    n1311,
    n198
  );


  not
  g1022
  (
    n953,
    n652
  );


  not
  g1023
  (
    n1355,
    n406
  );


  buf
  g1024
  (
    n789,
    n383
  );


  not
  g1025
  (
    n1358,
    n658
  );


  buf
  g1026
  (
    n1672,
    n351
  );


  buf
  g1027
  (
    n777,
    n348
  );


  not
  g1028
  (
    n690,
    n215
  );


  not
  g1029
  (
    n1016,
    n252
  );


  not
  g1030
  (
    n1485,
    n534
  );


  buf
  g1031
  (
    n1534,
    n474
  );


  buf
  g1032
  (
    n1069,
    n502
  );


  buf
  g1033
  (
    n1591,
    n350
  );


  not
  g1034
  (
    n1059,
    n260
  );


  buf
  g1035
  (
    n863,
    n589
  );


  buf
  g1036
  (
    n976,
    n424
  );


  buf
  g1037
  (
    n1600,
    n548
  );


  buf
  g1038
  (
    n1677,
    n166
  );


  not
  g1039
  (
    n1148,
    n172
  );


  not
  g1040
  (
    n1138,
    n660
  );


  buf
  g1041
  (
    n1494,
    n324
  );


  buf
  g1042
  (
    n1344,
    n587
  );


  not
  g1043
  (
    n1754,
    n604
  );


  buf
  g1044
  (
    n1082,
    n572
  );


  buf
  g1045
  (
    n1741,
    n325
  );


  buf
  g1046
  (
    n855,
    n465
  );


  not
  g1047
  (
    n1710,
    n664
  );


  not
  g1048
  (
    n1459,
    n507
  );


  buf
  g1049
  (
    n1266,
    n416
  );


  not
  g1050
  (
    n1304,
    n283
  );


  buf
  g1051
  (
    n1701,
    n605
  );


  not
  g1052
  (
    n1347,
    n347
  );


  not
  g1053
  (
    n1205,
    n503
  );


  buf
  g1054
  (
    n1047,
    n666
  );


  buf
  g1055
  (
    n1641,
    n627
  );


  buf
  g1056
  (
    n1263,
    n665
  );


  not
  g1057
  (
    n1449,
    n327
  );


  buf
  g1058
  (
    n1130,
    n434
  );


  buf
  g1059
  (
    n1289,
    n301
  );


  buf
  g1060
  (
    n1529,
    n259
  );


  buf
  g1061
  (
    n1376,
    n551
  );


  not
  g1062
  (
    n844,
    n452
  );


  buf
  g1063
  (
    n714,
    n219
  );


  not
  g1064
  (
    n1489,
    n330
  );


  not
  g1065
  (
    n1168,
    n353
  );


  buf
  g1066
  (
    n1379,
    n215
  );


  buf
  g1067
  (
    n915,
    n209
  );


  buf
  g1068
  (
    n1155,
    n473
  );


  buf
  g1069
  (
    n707,
    n462
  );


  not
  g1070
  (
    n966,
    n385
  );


  buf
  g1071
  (
    n1426,
    n631
  );


  not
  g1072
  (
    n1357,
    n665
  );


  not
  g1073
  (
    n1543,
    n449
  );


  buf
  g1074
  (
    n1265,
    n461
  );


  buf
  g1075
  (
    n909,
    n543
  );


  not
  g1076
  (
    n1354,
    n440
  );


  not
  g1077
  (
    n954,
    n183
  );


  not
  g1078
  (
    n1417,
    n389
  );


  buf
  g1079
  (
    n1531,
    n197
  );


  buf
  g1080
  (
    n1292,
    n246
  );


  buf
  g1081
  (
    n770,
    n211
  );


  not
  g1082
  (
    n711,
    n484
  );


  buf
  g1083
  (
    n1282,
    n168
  );


  buf
  g1084
  (
    n832,
    n302
  );


  not
  g1085
  (
    n1632,
    n420
  );


  buf
  g1086
  (
    n1560,
    n409
  );


  buf
  g1087
  (
    n1654,
    n418
  );


  not
  g1088
  (
    n737,
    n345
  );


  not
  g1089
  (
    n1097,
    n346
  );


  buf
  g1090
  (
    n1406,
    n389
  );


  not
  g1091
  (
    n946,
    n615
  );


  buf
  g1092
  (
    n1723,
    n585
  );


  not
  g1093
  (
    n973,
    n481
  );


  buf
  g1094
  (
    n970,
    n426
  );


  not
  g1095
  (
    n1216,
    n356
  );


  buf
  g1096
  (
    n955,
    n377
  );


  buf
  g1097
  (
    n744,
    n363
  );


  buf
  g1098
  (
    n1468,
    n174
  );


  not
  g1099
  (
    n775,
    n625
  );


  buf
  g1100
  (
    n1209,
    n180
  );


  not
  g1101
  (
    n1470,
    n329
  );


  buf
  g1102
  (
    n889,
    n220
  );


  not
  g1103
  (
    n1617,
    n630
  );


  not
  g1104
  (
    n1206,
    n556
  );


  buf
  g1105
  (
    n957,
    n475
  );


  not
  g1106
  (
    n1522,
    n266
  );


  not
  g1107
  (
    n1170,
    n191
  );


  buf
  g1108
  (
    n1172,
    n367
  );


  not
  g1109
  (
    n879,
    n585
  );


  buf
  g1110
  (
    n1611,
    n337
  );


  not
  g1111
  (
    n908,
    n342
  );


  buf
  g1112
  (
    n1307,
    n353
  );


  buf
  g1113
  (
    n1586,
    n601
  );


  not
  g1114
  (
    n1511,
    n421
  );


  not
  g1115
  (
    n985,
    n307
  );


  not
  g1116
  (
    n913,
    n284
  );


  not
  g1117
  (
    n1112,
    n627
  );


  buf
  g1118
  (
    n1146,
    n247
  );


  not
  g1119
  (
    n779,
    n282
  );


  buf
  g1120
  (
    n1232,
    n593
  );


  buf
  g1121
  (
    n1562,
    n285
  );


  not
  g1122
  (
    n1735,
    n267
  );


  not
  g1123
  (
    n1525,
    n528
  );


  not
  g1124
  (
    n1339,
    n416
  );


  not
  g1125
  (
    n1472,
    n247
  );


  not
  g1126
  (
    n1370,
    n339
  );


  buf
  g1127
  (
    n964,
    n615
  );


  buf
  g1128
  (
    n1077,
    n514
  );


  not
  g1129
  (
    n782,
    n583
  );


  buf
  g1130
  (
    n1316,
    n263
  );


  buf
  g1131
  (
    n1060,
    n291
  );


  not
  g1132
  (
    n1154,
    n639
  );


  buf
  g1133
  (
    n1277,
    n602
  );


  buf
  g1134
  (
    n1588,
    n211
  );


  not
  g1135
  (
    n1233,
    n260
  );


  buf
  g1136
  (
    n764,
    n513
  );


  buf
  g1137
  (
    n681,
    n350
  );


  not
  g1138
  (
    n1149,
    n596
  );


  buf
  g1139
  (
    n742,
    n475
  );


  not
  g1140
  (
    n1225,
    n515
  );


  buf
  g1141
  (
    n1578,
    n470
  );


  buf
  g1142
  (
    n945,
    n564
  );


  not
  g1143
  (
    n828,
    n270
  );


  not
  g1144
  (
    n819,
    n601
  );


  buf
  g1145
  (
    n1286,
    n384
  );


  not
  g1146
  (
    n971,
    n420
  );


  not
  g1147
  (
    n1250,
    n482
  );


  buf
  g1148
  (
    n1103,
    n388
  );


  not
  g1149
  (
    n1369,
    n428
  );


  buf
  g1150
  (
    n757,
    n345
  );


  buf
  g1151
  (
    n1599,
    n503
  );


  buf
  g1152
  (
    n891,
    n347
  );


  buf
  g1153
  (
    n1374,
    n391
  );


  buf
  g1154
  (
    n1402,
    n203
  );


  not
  g1155
  (
    n1324,
    n296
  );


  not
  g1156
  (
    n949,
    n284
  );


  buf
  g1157
  (
    n1551,
    n197
  );


  not
  g1158
  (
    n1359,
    n579
  );


  not
  g1159
  (
    n1515,
    n666
  );


  buf
  g1160
  (
    n717,
    n495
  );


  not
  g1161
  (
    n1646,
    n255
  );


  buf
  g1162
  (
    n885,
    n315
  );


  buf
  g1163
  (
    n1036,
    n534
  );


  buf
  g1164
  (
    n1666,
    n198
  );


  buf
  g1165
  (
    n678,
    n341
  );


  buf
  g1166
  (
    n979,
    n397
  );


  not
  g1167
  (
    n1630,
    n322
  );


  buf
  g1168
  (
    n821,
    n558
  );


  buf
  g1169
  (
    n1301,
    n462
  );


  buf
  g1170
  (
    n749,
    n435
  );


  not
  g1171
  (
    n1101,
    n439
  );


  not
  g1172
  (
    KeyWire_0_3,
    n275
  );


  not
  g1173
  (
    n1733,
    n186
  );


  buf
  g1174
  (
    n1243,
    n324
  );


  buf
  g1175
  (
    n933,
    n324
  );


  not
  g1176
  (
    n926,
    n669
  );


  buf
  g1177
  (
    n1571,
    n448
  );


  buf
  g1178
  (
    n1722,
    n265
  );


  buf
  g1179
  (
    n1049,
    n440
  );


  buf
  g1180
  (
    n1590,
    n456
  );


  buf
  g1181
  (
    n1296,
    n551
  );


  not
  g1182
  (
    n1327,
    n581
  );


  not
  g1183
  (
    n1664,
    n476
  );


  not
  g1184
  (
    n1451,
    n439
  );


  not
  g1185
  (
    n703,
    n442
  );


  buf
  g1186
  (
    n1160,
    n307
  );


  buf
  g1187
  (
    n1554,
    n194
  );


  not
  g1188
  (
    n1546,
    n267
  );


  not
  g1189
  (
    n1052,
    n220
  );


  not
  g1190
  (
    n790,
    n657
  );


  not
  g1191
  (
    n1444,
    n492
  );


  not
  g1192
  (
    n1751,
    n662
  );


  buf
  g1193
  (
    n786,
    n638
  );


  not
  g1194
  (
    n1598,
    n596
  );


  buf
  g1195
  (
    n1033,
    n538
  );


  not
  g1196
  (
    n1279,
    n212
  );


  not
  g1197
  (
    n1410,
    n336
  );


  buf
  g1198
  (
    n1274,
    n536
  );


  buf
  g1199
  (
    n825,
    n167
  );


  not
  g1200
  (
    n1158,
    n615
  );


  buf
  g1201
  (
    n1386,
    n349
  );


  not
  g1202
  (
    n1310,
    n260
  );


  buf
  g1203
  (
    n1220,
    n382
  );


  buf
  g1204
  (
    n1752,
    n478
  );


  not
  g1205
  (
    n1690,
    n512
  );


  not
  g1206
  (
    n1224,
    n496
  );


  buf
  g1207
  (
    n1434,
    n367
  );


  not
  g1208
  (
    n1346,
    n355
  );


  buf
  g1209
  (
    n1089,
    n361
  );


  buf
  g1210
  (
    n990,
    n417
  );


  not
  g1211
  (
    n1389,
    n589
  );


  buf
  g1212
  (
    n1008,
    n608
  );


  not
  g1213
  (
    n1636,
    n518
  );


  buf
  g1214
  (
    n1593,
    n190
  );


  buf
  g1215
  (
    n1567,
    n475
  );


  not
  g1216
  (
    KeyWire_0_14,
    n627
  );


  not
  g1217
  (
    n793,
    n392
  );


  not
  g1218
  (
    n1246,
    n328
  );


  buf
  g1219
  (
    n928,
    n364
  );


  buf
  g1220
  (
    n739,
    n542
  );


  buf
  g1221
  (
    n1164,
    n499
  );


  buf
  g1222
  (
    n1518,
    n174
  );


  buf
  g1223
  (
    n1298,
    n212
  );


  buf
  g1224
  (
    n1564,
    n396
  );


  not
  g1225
  (
    n1613,
    n226
  );


  not
  g1226
  (
    n1469,
    n652
  );


  buf
  g1227
  (
    n1235,
    n251
  );


  buf
  g1228
  (
    n986,
    n218
  );


  not
  g1229
  (
    n1284,
    n610
  );


  not
  g1230
  (
    n1644,
    n451
  );


  buf
  g1231
  (
    n829,
    n228
  );


  not
  g1232
  (
    n1245,
    n327
  );


  buf
  g1233
  (
    n1716,
    n447
  );


  not
  g1234
  (
    n1071,
    n459
  );


  buf
  g1235
  (
    n1306,
    n279
  );


  buf
  g1236
  (
    n1260,
    n354
  );


  not
  g1237
  (
    n721,
    n366
  );


  buf
  g1238
  (
    n1340,
    n651
  );


  not
  g1239
  (
    n699,
    n647
  );


  buf
  g1240
  (
    n781,
    n418
  );


  not
  g1241
  (
    n962,
    n399
  );


  buf
  g1242
  (
    n1395,
    n391
  );


  buf
  g1243
  (
    n760,
    n457
  );


  not
  g1244
  (
    n1612,
    n396
  );


  buf
  g1245
  (
    n1729,
    n360
  );


  not
  g1246
  (
    n705,
    n624
  );


  buf
  g1247
  (
    n1272,
    n572
  );


  buf
  g1248
  (
    n1416,
    n392
  );


  buf
  g1249
  (
    n818,
    n189
  );


  buf
  g1250
  (
    n734,
    n371
  );


  not
  g1251
  (
    KeyWire_0_0,
    n612
  );


  not
  g1252
  (
    n1490,
    n597
  );


  not
  g1253
  (
    n824,
    n558
  );


  buf
  g1254
  (
    n1639,
    n295
  );


  not
  g1255
  (
    n1238,
    n399
  );


  buf
  g1256
  (
    n1524,
    n670
  );


  buf
  g1257
  (
    n894,
    n381
  );


  buf
  g1258
  (
    n1577,
    n531
  );


  not
  g1259
  (
    n1714,
    n662
  );


  buf
  g1260
  (
    n1385,
    n582
  );


  buf
  g1261
  (
    n1038,
    n362
  );


  buf
  g1262
  (
    n884,
    n342
  );


  not
  g1263
  (
    n1580,
    n174
  );


  not
  g1264
  (
    n1315,
    n594
  );


  buf
  g1265
  (
    n1280,
    n465
  );


  buf
  g1266
  (
    n675,
    n438
  );


  not
  g1267
  (
    n1698,
    n491
  );


  not
  g1268
  (
    n1302,
    n373
  );


  not
  g1269
  (
    n1001,
    n476
  );


  not
  g1270
  (
    n1043,
    n317
  );


  buf
  g1271
  (
    n685,
    n627
  );


  buf
  g1272
  (
    n1432,
    n326
  );


  not
  g1273
  (
    n677,
    n235
  );


  buf
  g1274
  (
    n1065,
    n346
  );


  buf
  g1275
  (
    n939,
    n547
  );


  not
  g1276
  (
    KeyWire_0_6,
    n574
  );


  not
  g1277
  (
    n1509,
    n652
  );


  buf
  g1278
  (
    n1478,
    n365
  );


  not
  g1279
  (
    n995,
    n214
  );


  buf
  g1280
  (
    n1064,
    n631
  );


  not
  g1281
  (
    n1659,
    n339
  );


  not
  g1282
  (
    n1607,
    n522
  );


  buf
  g1283
  (
    n1737,
    n262
  );


  not
  g1284
  (
    n1573,
    n380
  );


  not
  g1285
  (
    n1268,
    n512
  );


  not
  g1286
  (
    n1703,
    n519
  );


  not
  g1287
  (
    n1121,
    n525
  );


  not
  g1288
  (
    n1332,
    n194
  );


  not
  g1289
  (
    n1303,
    n264
  );


  not
  g1290
  (
    n1563,
    n235
  );


  buf
  g1291
  (
    n809,
    n280
  );


  buf
  g1292
  (
    n1486,
    n618
  );


  not
  g1293
  (
    n695,
    n433
  );


  buf
  g1294
  (
    n1670,
    n425
  );


  not
  g1295
  (
    n867,
    n236
  );


  not
  g1296
  (
    n732,
    n619
  );


  not
  g1297
  (
    n1709,
    n661
  );


  buf
  g1298
  (
    n1661,
    n477
  );


  not
  g1299
  (
    n1730,
    n498
  );


  not
  g1300
  (
    n719,
    n161
  );


  buf
  g1301
  (
    n1351,
    n355
  );


  not
  g1302
  (
    n1123,
    n472
  );


  buf
  g1303
  (
    n1360,
    n565
  );


  buf
  g1304
  (
    n1035,
    n330
  );


  not
  g1305
  (
    n1680,
    n466
  );


  not
  g1306
  (
    n1293,
    n532
  );


  buf
  g1307
  (
    n1334,
    n467
  );


  not
  g1308
  (
    n1116,
    n423
  );


  buf
  g1309
  (
    n977,
    n502
  );


  not
  g1310
  (
    n1423,
    n643
  );


  not
  g1311
  (
    n1396,
    n432
  );


  not
  g1312
  (
    n984,
    n542
  );


  buf
  g1313
  (
    n1204,
    n424
  );


  buf
  g1314
  (
    n1683,
    n621
  );


  not
  g1315
  (
    n994,
    n382
  );


  not
  g1316
  (
    n706,
    n338
  );


  buf
  g1317
  (
    n1230,
    n624
  );


  not
  g1318
  (
    n1256,
    n339
  );


  buf
  g1319
  (
    n772,
    n560
  );


  buf
  g1320
  (
    n1475,
    n463
  );


  buf
  g1321
  (
    n1102,
    n467
  );


  buf
  g1322
  (
    n769,
    n555
  );


  not
  g1323
  (
    n1411,
    n423
  );


  buf
  g1324
  (
    n799,
    n233
  );


  not
  g1325
  (
    n688,
    n341
  );


  not
  g1326
  (
    n1139,
    n429
  );


  not
  g1327
  (
    n778,
    n580
  );


  not
  g1328
  (
    n831,
    n294
  );


  buf
  g1329
  (
    n820,
    n195
  );


  not
  g1330
  (
    n972,
    n452
  );


  not
  g1331
  (
    n1278,
    n297
  );


  buf
  g1332
  (
    n1329,
    n345
  );


  not
  g1333
  (
    n727,
    n422
  );


  not
  g1334
  (
    n807,
    n469
  );


  not
  g1335
  (
    n910,
    n525
  );


  not
  g1336
  (
    n1152,
    n311
  );


  not
  g1337
  (
    n1561,
    n445
  );


  buf
  g1338
  (
    n833,
    n214
  );


  buf
  g1339
  (
    n1542,
    n561
  );


  not
  g1340
  (
    n1240,
    n464
  );


  buf
  g1341
  (
    n1399,
    n472
  );


  not
  g1342
  (
    n935,
    n404
  );


  not
  g1343
  (
    n761,
    n177
  );


  not
  g1344
  (
    n947,
    n198
  );


  not
  g1345
  (
    n1497,
    n497
  );


  buf
  g1346
  (
    n1183,
    n274
  );


  buf
  g1347
  (
    n1691,
    n276
  );


  not
  g1348
  (
    n1219,
    n195
  );


  not
  g1349
  (
    n1450,
    n306
  );


  not
  g1350
  (
    n917,
    n184
  );


  buf
  g1351
  (
    n1392,
    n544
  );


  not
  g1352
  (
    n1088,
    n289
  );


  buf
  g1353
  (
    n1533,
    n274
  );


  buf
  g1354
  (
    n1140,
    n583
  );


  not
  g1355
  (
    n1610,
    n526
  );


  not
  g1356
  (
    n1187,
    n167
  );


  buf
  g1357
  (
    n1095,
    n312
  );


  buf
  g1358
  (
    n701,
    n309
  );


  buf
  g1359
  (
    n1679,
    n635
  );


  buf
  g1360
  (
    n1322,
    n527
  );


  not
  g1361
  (
    n1707,
    n276
  );


  buf
  g1362
  (
    n1212,
    n621
  );


  buf
  g1363
  (
    n1012,
    n243
  );


  not
  g1364
  (
    n1681,
    n463
  );


  not
  g1365
  (
    n921,
    n331
  );


  buf
  g1366
  (
    n958,
    n539
  );


  not
  g1367
  (
    n1496,
    n316
  );


  not
  g1368
  (
    n1361,
    n210
  );


  buf
  g1369
  (
    n1520,
    n280
  );


  buf
  g1370
  (
    n902,
    n329
  );


  buf
  g1371
  (
    n1453,
    n374
  );


  not
  g1372
  (
    n1328,
    n567
  );


  buf
  g1373
  (
    n1195,
    n598
  );


  buf
  g1374
  (
    n676,
    n181
  );


  buf
  g1375
  (
    n741,
    n292
  );


  buf
  g1376
  (
    n974,
    n599
  );


  buf
  g1377
  (
    n857,
    n209
  );


  not
  g1378
  (
    n1696,
    n431
  );


  buf
  g1379
  (
    n975,
    n624
  );


  buf
  g1380
  (
    n763,
    n473
  );


  buf
  g1381
  (
    n1003,
    n372
  );


  not
  g1382
  (
    n861,
    n637
  );


  not
  g1383
  (
    n1397,
    n602
  );


  not
  g1384
  (
    n733,
    n613
  );


  not
  g1385
  (
    n771,
    n658
  );


  not
  g1386
  (
    n1448,
    n438
  );


  not
  g1387
  (
    n988,
    n401
  );


  not
  g1388
  (
    n1176,
    n450
  );


  not
  g1389
  (
    n700,
    n432
  );


  not
  g1390
  (
    n800,
    n255
  );


  buf
  g1391
  (
    n1549,
    n404
  );


  not
  g1392
  (
    n1697,
    n228
  );


  not
  g1393
  (
    n853,
    n479
  );


  buf
  g1394
  (
    n1684,
    n370
  );


  not
  g1395
  (
    n1073,
    n209
  );


  not
  g1396
  (
    n745,
    n287
  );


  not
  g1397
  (
    n1242,
    n585
  );


  not
  g1398
  (
    n747,
    n193
  );


  not
  g1399
  (
    n1673,
    n614
  );


  not
  g1400
  (
    n1133,
    n271
  );


  not
  g1401
  (
    n1026,
    n481
  );


  nand
  g1402
  (
    n1128,
    n485,
    n429
  );


  nand
  g1403
  (
    n1314,
    n301,
    n318,
    n218,
    n308
  );


  xor
  g1404
  (
    n1258,
    n376,
    n437,
    n538,
    n477
  );


  nor
  g1405
  (
    n1104,
    n233,
    n332,
    n410,
    n556
  );


  or
  g1406
  (
    n1252,
    n568,
    n638,
    n574,
    n357
  );


  nor
  g1407
  (
    n1460,
    n439,
    n470,
    n370,
    n407
  );


  or
  g1408
  (
    n1748,
    n350,
    n201,
    n667,
    n540
  );


  nor
  g1409
  (
    n1535,
    n435,
    n413,
    n402,
    n494
  );


  nor
  g1410
  (
    n1290,
    n206,
    n664,
    n413,
    n403
  );


  nor
  g1411
  (
    n1264,
    n445,
    n530,
    n570,
    n463
  );


  nor
  g1412
  (
    n918,
    n223,
    n503,
    n414,
    n386
  );


  or
  g1413
  (
    n1669,
    n222,
    n254,
    n452,
    n238
  );


  and
  g1414
  (
    n1117,
    n431,
    n451,
    n281,
    n654
  );


  nand
  g1415
  (
    n1163,
    n251,
    n441,
    n514,
    n259
  );


  and
  g1416
  (
    n895,
    n169,
    n241,
    n305,
    n552
  );


  nand
  g1417
  (
    n1498,
    n207,
    n212,
    n341,
    n318
  );


  xnor
  g1418
  (
    n1594,
    n557,
    n300,
    n648,
    n569
  );


  nand
  g1419
  (
    n1309,
    n413,
    n267,
    n408,
    n301
  );


  xor
  g1420
  (
    n1584,
    n529,
    n600,
    n582,
    n535
  );


  and
  g1421
  (
    n1285,
    n655,
    n370,
    n610,
    n646
  );


  and
  g1422
  (
    n1253,
    n332,
    n449,
    n310,
    n594
  );


  xor
  g1423
  (
    n1576,
    n328,
    n596,
    n502,
    n671
  );


  nand
  g1424
  (
    n1215,
    n213,
    n319,
    n415,
    n270
  );


  nand
  g1425
  (
    n892,
    n649,
    n279,
    n389,
    n262
  );


  and
  g1426
  (
    n848,
    n551,
    n173,
    n281,
    n327
  );


  and
  g1427
  (
    n1519,
    n544,
    n264,
    n289,
    n624
  );


  xnor
  g1428
  (
    n1317,
    n362,
    n431,
    n426,
    n290
  );


  xnor
  g1429
  (
    n1009,
    n444,
    n485,
    n619,
    n489
  );


  xnor
  g1430
  (
    n1368,
    n471,
    n252,
    n283,
    n463
  );


  xor
  g1431
  (
    n1384,
    n545,
    n656,
    n280,
    n526
  );


  and
  g1432
  (
    n880,
    n361,
    n653,
    n495,
    n202
  );


  xor
  g1433
  (
    n1724,
    n187,
    n593,
    n524,
    n337
  );


  xnor
  g1434
  (
    n967,
    n218,
    n535,
    n541,
    n514
  );


  or
  g1435
  (
    n1021,
    n498,
    n573,
    n381,
    n250
  );


  xor
  g1436
  (
    n1053,
    n622,
    n219,
    n471,
    n246
  );


  nand
  g1437
  (
    n1609,
    n601,
    n307,
    n632,
    n287
  );


  xnor
  g1438
  (
    n1704,
    n368,
    n497,
    n526
  );


  xor
  g1439
  (
    n1513,
    n176,
    n344,
    n245,
    n205
  );


  nand
  g1440
  (
    n1271,
    n482,
    n464,
    n456,
    n488
  );


  xor
  g1441
  (
    n1377,
    n516,
    n428,
    n298,
    n184
  );


  xnor
  g1442
  (
    n1144,
    n368,
    n253,
    n220,
    n554
  );


  xnor
  g1443
  (
    n1481,
    n185,
    n380,
    n507,
    n464
  );


  xor
  g1444
  (
    n1501,
    n244,
    n360,
    n479,
    n516
  );


  xor
  g1445
  (
    n1066,
    n251,
    n505,
    n357,
    n483
  );


  and
  g1446
  (
    n1420,
    n371,
    n460,
    n280,
    n587
  );


  xnor
  g1447
  (
    n1363,
    n641,
    n565,
    n564,
    n450
  );


  nand
  g1448
  (
    n1642,
    n287,
    n183,
    n654,
    n489
  );


  and
  g1449
  (
    n1476,
    n206,
    n491,
    n193,
    n625
  );


  nor
  g1450
  (
    n1364,
    n417,
    n511,
    n257,
    n545
  );


  xor
  g1451
  (
    n1711,
    n264,
    n506,
    n448,
    n238
  );


  xor
  g1452
  (
    n1512,
    n273,
    n460,
    n205,
    n490
  );


  xor
  g1453
  (
    n1523,
    n237,
    n577,
    n561,
    n367
  );


  xor
  g1454
  (
    n1198,
    n305,
    n426,
    n620,
    n671
  );


  nor
  g1455
  (
    n1294,
    n529,
    n180,
    n430,
    n216
  );


  nand
  g1456
  (
    n1099,
    n421,
    n267,
    n414,
    n411
  );


  and
  g1457
  (
    n1655,
    n634,
    n452,
    n172,
    n586
  );


  xnor
  g1458
  (
    n992,
    n602,
    n513,
    n261,
    n610
  );


  nand
  g1459
  (
    n1267,
    n400,
    n390,
    n248,
    n387
  );


  or
  g1460
  (
    n1557,
    n614,
    n613,
    n236,
    n162
  );


  xnor
  g1461
  (
    n1559,
    n166,
    n317,
    n480,
    n455
  );


  xor
  g1462
  (
    n718,
    n285,
    n655,
    n378,
    n529
  );


  nor
  g1463
  (
    n1484,
    n479,
    n383,
    n482,
    n577
  );


  xnor
  g1464
  (
    n1657,
    n517,
    n450,
    n434,
    n244
  );


  and
  g1465
  (
    n941,
    n659,
    n201,
    n523,
    n391
  );


  nor
  g1466
  (
    n1297,
    n534,
    n412,
    n400,
    n199
  );


  nor
  g1467
  (
    n795,
    n401,
    n367,
    n356,
    n428
  );


  nor
  g1468
  (
    n1587,
    n265,
    n425,
    n217,
    n178
  );


  xnor
  g1469
  (
    n1179,
    n357,
    n224,
    n510,
    n663
  );


  xor
  g1470
  (
    n817,
    n643,
    n299,
    n338,
    n651
  );


  nor
  g1471
  (
    n752,
    n495,
    n236,
    n575,
    n604
  );


  xnor
  g1472
  (
    n762,
    n297,
    n499,
    n573,
    n543
  );


  nand
  g1473
  (
    n1572,
    n630,
    n352,
    n386,
    n629
  );


  xor
  g1474
  (
    n768,
    n466,
    n514,
    n600,
    n222
  );


  and
  g1475
  (
    n1503,
    n427,
    n661,
    n478,
    n396
  );


  and
  g1476
  (
    n888,
    n643,
    n436,
    n469,
    n369
  );


  xor
  g1477
  (
    n893,
    n511,
    n240,
    n446,
    n617
  );


  nor
  g1478
  (
    n1319,
    n521,
    n258,
    n634,
    n295
  );


  or
  g1479
  (
    n841,
    n285,
    n290,
    n563,
    n488
  );


  xnor
  g1480
  (
    n1539,
    n415,
    n372,
    n457,
    n211
  );


  nor
  g1481
  (
    n748,
    n662,
    n557,
    n519,
    n415
  );


  nor
  g1482
  (
    n1658,
    n385,
    n378,
    n562,
    n558
  );


  nor
  g1483
  (
    n1086,
    n656,
    n454,
    n424,
    n516
  );


  nand
  g1484
  (
    n1107,
    n358,
    n319,
    n324,
    n306
  );


  nand
  g1485
  (
    n822,
    n274,
    n595,
    n518,
    n555
  );


  nor
  g1486
  (
    n1731,
    n454,
    n237,
    n192,
    n180
  );


  or
  g1487
  (
    n1162,
    n351,
    n355,
    n468,
    n416
  );


  xnor
  g1488
  (
    n1556,
    n374,
    n422,
    n410,
    n501
  );


  xor
  g1489
  (
    n755,
    n628,
    n646,
    n487,
    n442
  );


  xor
  g1490
  (
    n1647,
    n427,
    n611,
    n384,
    n245
  );


  or
  g1491
  (
    n716,
    n661,
    n443,
    n609,
    n170
  );


  xor
  g1492
  (
    n1605,
    n181,
    n451,
    n185,
    n541
  );


  or
  g1493
  (
    n1393,
    n338,
    n668,
    n323,
    n538
  );


  nor
  g1494
  (
    n1067,
    n364,
    n254,
    n647,
    n403
  );


  or
  g1495
  (
    n925,
    n606,
    n575,
    n312,
    n554
  );


  nand
  g1496
  (
    n1161,
    n179,
    n183,
    n227,
    n296
  );


  and
  g1497
  (
    n1436,
    n501,
    n366,
    n175,
    n191
  );


  nand
  g1498
  (
    n1217,
    n481,
    n547,
    n490,
    n310
  );


  xor
  g1499
  (
    n997,
    n381,
    n458,
    n528,
    n248
  );


  xnor
  g1500
  (
    n1575,
    n653,
    n401,
    n466,
    n179
  );


  xnor
  g1501
  (
    n1682,
    n245,
    n407,
    n185,
    n592
  );


  xnor
  g1502
  (
    n811,
    n227,
    n266,
    n633,
    n348
  );


  xor
  g1503
  (
    n897,
    n291,
    n421,
    n554,
    n528
  );


  or
  g1504
  (
    n1223,
    n282,
    n278,
    n300,
    n580
  );


  nand
  g1505
  (
    n1281,
    n168,
    n649,
    n626,
    n445
  );


  nand
  g1506
  (
    n1333,
    n312,
    n288,
    n311,
    n645
  );


  or
  g1507
  (
    n1442,
    n314,
    n237,
    n276,
    n509
  );


  and
  g1508
  (
    n674,
    n234,
    n545,
    n459,
    n575
  );


  or
  g1509
  (
    n1721,
    n527,
    n182,
    n380,
    n443
  );


  and
  g1510
  (
    n1409,
    n608,
    n402,
    n642,
    n556
  );


  xnor
  g1511
  (
    n1628,
    n277,
    n569,
    n231,
    n544
  );


  or
  g1512
  (
    KeyWire_0_2,
    n329,
    n273,
    n299,
    n424
  );


  or
  g1513
  (
    n919,
    n395,
    n265,
    n628,
    n287
  );


  nand
  g1514
  (
    n1437,
    n612,
    n219,
    n404,
    n252
  );


  xor
  g1515
  (
    n753,
    n340,
    n657,
    n327,
    n230
  );


  xnor
  g1516
  (
    n710,
    n446,
    n476,
    n522,
    n670
  );


  nor
  g1517
  (
    n1629,
    n591,
    n599,
    n537,
    n425
  );


  nor
  g1518
  (
    n1458,
    n233,
    n444,
    n203,
    n576
  );


  nand
  g1519
  (
    n1367,
    n257,
    n240,
    n623,
    n442
  );


  nand
  g1520
  (
    n1087,
    n170,
    n496,
    n382,
    n186
  );


  or
  g1521
  (
    n1713,
    n173,
    n492,
    n605,
    n630
  );


  xor
  g1522
  (
    n1401,
    n209,
    n404,
    n437,
    n653
  );


  and
  g1523
  (
    n923,
    n259,
    n277,
    n399,
    n316
  );


  nand
  g1524
  (
    n1429,
    n447,
    n170,
    n541,
    n642
  );


  and
  g1525
  (
    n980,
    n527,
    n614,
    n384,
    n578
  );


  nor
  g1526
  (
    n1100,
    n531,
    n580,
    n519,
    n295
  );


  xnor
  g1527
  (
    n1299,
    n662,
    n371,
    n651,
    n343
  );


  xnor
  g1528
  (
    n1595,
    n320,
    n187,
    n459,
    n309
  );


  xor
  g1529
  (
    n792,
    n546,
    n195,
    n291,
    n161
  );


  nor
  g1530
  (
    n1745,
    n494,
    n501,
    n303,
    n560
  );


  nor
  g1531
  (
    n776,
    n584,
    n432,
    n444,
    n477
  );


  nor
  g1532
  (
    n1660,
    n554,
    n170,
    n581,
    n490
  );


  or
  g1533
  (
    n1596,
    n450,
    n336,
    n229,
    n186
  );


  and
  g1534
  (
    n794,
    n399,
    n498,
    n484,
    n616
  );


  nor
  g1535
  (
    n906,
    n536,
    n192,
    n278,
    n586
  );


  nand
  g1536
  (
    n1057,
    n593,
    n368,
    n231,
    n362
  );


  nand
  g1537
  (
    n1050,
    n163,
    n566,
    n474,
    n239
  );


  nand
  g1538
  (
    n810,
    n351,
    n167,
    n526,
    n308
  );


  xor
  g1539
  (
    n859,
    n486,
    n619,
    n171,
    n333
  );


  nor
  g1540
  (
    n1338,
    n633,
    n419,
    n651,
    n359
  );


  or
  g1541
  (
    n1247,
    n553,
    n378,
    n384,
    n645
  );


  xor
  g1542
  (
    n874,
    n640,
    n485,
    n297,
    n571
  );


  nor
  g1543
  (
    n1732,
    n345,
    n217,
    n335,
    n260
  );


  or
  g1544
  (
    n1062,
    n337,
    n578,
    n623,
    n536
  );


  xnor
  g1545
  (
    n924,
    n492,
    n474,
    n190,
    n640
  );


  and
  g1546
  (
    n1537,
    n550,
    n319,
    n272,
    n322
  );


  and
  g1547
  (
    n858,
    n364,
    n222,
    n206,
    n665
  );


  xnor
  g1548
  (
    n1706,
    n449,
    n347,
    n596,
    n311
  );


  or
  g1549
  (
    n1030,
    n400,
    n614,
    n385,
    n357
  );


  xnor
  g1550
  (
    n1700,
    n411,
    n645,
    n467,
    n611
  );


  nor
  g1551
  (
    n1078,
    n388,
    n462,
    n640,
    n657
  );


  and
  g1552
  (
    n1526,
    n428,
    n548,
    n465,
    n517
  );


  xnor
  g1553
  (
    n907,
    n230,
    n532,
    n508,
    n422
  );


  xnor
  g1554
  (
    n931,
    n617,
    n406,
    n409,
    n313
  );


  nand
  g1555
  (
    n1743,
    n216,
    n549,
    n315,
    n229
  );


  nand
  g1556
  (
    n1350,
    n506,
    n562,
    n304,
    n644
  );


  xor
  g1557
  (
    n1320,
    n299,
    n459,
    n444,
    n616
  );


  or
  g1558
  (
    n838,
    n496,
    n535,
    n590,
    n563
  );


  xnor
  g1559
  (
    n1640,
    n240,
    n394,
    n408,
    n403
  );


  or
  g1560
  (
    n791,
    n531,
    n292,
    n247,
    n440
  );


  or
  g1561
  (
    n883,
    n382,
    n309,
    n353,
    n552
  );


  or
  g1562
  (
    n1694,
    n499,
    n671,
    n375,
    n600
  );


  xnor
  g1563
  (
    n1504,
    n298,
    n432,
    n591,
    n587
  );


  and
  g1564
  (
    n1275,
    n546,
    n168,
    n542,
    n427
  );


  and
  g1565
  (
    n1024,
    n604,
    n447,
    n659,
    n505
  );


  and
  g1566
  (
    n1742,
    n393,
    n232,
    n458,
    n664
  );


  xor
  g1567
  (
    n704,
    n563,
    n623,
    n548,
    n411
  );


  and
  g1568
  (
    n774,
    n644,
    n584,
    n574,
    n162
  );


  nand
  g1569
  (
    n1005,
    n215,
    n501,
    n229,
    n560
  );


  xnor
  g1570
  (
    n1313,
    n302,
    n161,
    n221,
    n181
  );


  xor
  g1571
  (
    n1228,
    n477,
    n433,
    n377,
    n669
  );


  xor
  g1572
  (
    n871,
    n539,
    n572,
    n485,
    n329
  );


  xor
  g1573
  (
    n1645,
    n313,
    n623,
    n248,
    n354
  );


  or
  g1574
  (
    n1325,
    n530,
    n314,
    n219,
    n250
  );


  xnor
  g1575
  (
    n1055,
    n521,
    n603,
    n356,
    n201
  );


  nor
  g1576
  (
    n929,
    n529,
    n241,
    n178,
    n472
  );


  xnor
  g1577
  (
    n1479,
    n638,
    n365,
    n269,
    n388
  );


  nand
  g1578
  (
    n901,
    n331,
    n208,
    n468,
    n433
  );


  xor
  g1579
  (
    n865,
    n236,
    n510,
    n584,
    n547
  );


  or
  g1580
  (
    n767,
    n454,
    n293,
    n256,
    n394
  );


  nand
  g1581
  (
    n1208,
    n249,
    n232,
    n294,
    n175
  );


  nand
  g1582
  (
    n1184,
    n354,
    n474,
    n335,
    n366
  );


  xnor
  g1583
  (
    n1091,
    n232,
    n349,
    n173,
    n553
  );


  or
  g1584
  (
    n1196,
    n358,
    n256,
    n177,
    n189
  );


  xnor
  g1585
  (
    n1638,
    n262,
    n622,
    n604,
    n276
  );


  nand
  g1586
  (
    n1124,
    n546,
    n323,
    n650,
    n660
  );


  xor
  g1587
  (
    n1502,
    n165,
    n409,
    n221,
    n202
  );


  nand
  g1588
  (
    n1634,
    n181,
    n626,
    n659,
    n182
  );


  nand
  g1589
  (
    n1446,
    n297,
    n471,
    n455,
    n510
  );


  and
  g1590
  (
    n1019,
    n257,
    n589,
    n576,
    n163
  );


  xor
  g1591
  (
    n1532,
    n494,
    n346,
    n632,
    n652
  );


  xnor
  g1592
  (
    n1174,
    n403,
    n258,
    n221,
    n285
  );


  nor
  g1593
  (
    n1505,
    n368,
    n246,
    n549,
    n298
  );


  or
  g1594
  (
    n1341,
    n192,
    n668,
    n278,
    n255
  );


  or
  g1595
  (
    n847,
    n286,
    n607,
    n650,
    n539
  );


  xnor
  g1596
  (
    n1725,
    n247,
    n598,
    n401,
    n616
  );


  nor
  g1597
  (
    n1300,
    n221,
    n520,
    n577,
    n165
  );


  nor
  g1598
  (
    n993,
    n196,
    n351,
    n269,
    n208
  );


  nand
  g1599
  (
    n713,
    n420,
    n595,
    n606,
    n435
  );


  nor
  g1600
  (
    n1058,
    n218,
    n233,
    n626,
    n429
  );


  nor
  g1601
  (
    KeyWire_0_9,
    n180,
    n302,
    n303,
    n570
  );


  nor
  g1602
  (
    n1106,
    n308,
    n315,
    n178,
    n644
  );


  nand
  g1603
  (
    n1749,
    n172,
    n441,
    n638,
    n356
  );


  xor
  g1604
  (
    n1321,
    n553,
    n378,
    n194,
    n263
  );


  nand
  g1605
  (
    n1075,
    n669,
    n169,
    n183,
    n316
  );


  nor
  g1606
  (
    n898,
    n412,
    n281,
    n512
  );


  and
  g1607
  (
    n1239,
    n375,
    n569,
    n334,
    n611
  );


  xor
  g1608
  (
    n1492,
    n472,
    n456,
    n398,
    n437
  );


  nor
  g1609
  (
    n715,
    n513,
    n406,
    n451,
    n320
  );


  nor
  g1610
  (
    n740,
    n583,
    n371,
    n621,
    n313
  );


  nand
  g1611
  (
    n1428,
    n478,
    n175,
    n597,
    n670
  );


  nor
  g1612
  (
    n1608,
    n506,
    n562,
    n177,
    n563
  );


  xnor
  g1613
  (
    n1261,
    n668,
    n524,
    n448,
    n578
  );


  xor
  g1614
  (
    n1041,
    n302,
    n318,
    n284,
    n261
  );


  xnor
  g1615
  (
    n1040,
    n374,
    n336,
    n261,
    n205
  );


  xor
  g1616
  (
    n736,
    n379,
    n242,
    n266,
    n172
  );


  nor
  g1617
  (
    n1744,
    n464,
    n490,
    n303,
    n270
  );


  xor
  g1618
  (
    n1061,
    n215,
    n573,
    n243,
    n196
  );


  nand
  g1619
  (
    n1471,
    n390,
    n171,
    n566,
    n548
  );


  nand
  g1620
  (
    n1188,
    n344,
    n198,
    n588,
    n387
  );


  xnor
  g1621
  (
    n912,
    n641,
    n173,
    n349,
    n507
  );


  xor
  g1622
  (
    n1380,
    n207,
    n648,
    n191,
    n636
  );


  xnor
  g1623
  (
    n722,
    n305,
    n663,
    n277,
    n163
  );


  nand
  g1624
  (
    n1463,
    n225,
    n330,
    n634,
    n360
  );


  and
  g1625
  (
    n840,
    n333,
    n570,
    n379,
    n294
  );


  xor
  g1626
  (
    n1619,
    n294,
    n637,
    n586,
    n224
  );


  xor
  g1627
  (
    n1093,
    n461,
    n500,
    n355,
    n570
  );


  or
  g1628
  (
    n1108,
    n536,
    n288,
    n617,
    n373
  );


  xor
  g1629
  (
    n916,
    n590,
    n657,
    n200,
    n365
  );


  or
  g1630
  (
    n1506,
    n350,
    n184,
    n557,
    n559
  );


  and
  g1631
  (
    n1027,
    n533,
    n525,
    n264,
    n206
  );


  nand
  g1632
  (
    n1114,
    n275,
    n176,
    n655,
    n249
  );


  or
  g1633
  (
    n1530,
    n633,
    n164,
    n559,
    n392
  );


  or
  g1634
  (
    n1615,
    n567,
    n643,
    n379,
    n408
  );


  xnor
  g1635
  (
    n1491,
    n359,
    n192,
    n430,
    n576
  );


  xnor
  g1636
  (
    n1051,
    n656,
    n630,
    n417,
    n423
  );


  nand
  g1637
  (
    n899,
    n235,
    n436,
    n632,
    n430
  );


  xnor
  g1638
  (
    n783,
    n603,
    n273,
    n197,
    n407
  );


  and
  g1639
  (
    n697,
    n541,
    n555,
    n249,
    n414
  );


  xor
  g1640
  (
    n1398,
    n438,
    n190,
    n337,
    n577
  );


  and
  g1641
  (
    n905,
    n539,
    n250,
    n405,
    n286
  );


  nand
  g1642
  (
    n756,
    n376,
    n475,
    n453,
    n269
  );


  and
  g1643
  (
    n982,
    n551,
    n488,
    n532,
    n383
  );


  xnor
  g1644
  (
    n1295,
    n229,
    n579,
    n242,
    n393
  );


  nor
  g1645
  (
    n1381,
    n256,
    n537,
    n518,
    n185
  );


  nand
  g1646
  (
    n1585,
    n663,
    n587,
    n586,
    n361
  );


  and
  g1647
  (
    n1002,
    n533,
    n495,
    n441,
    n646
  );


  and
  g1648
  (
    n1135,
    n455,
    n169,
    n632,
    n388
  );


  xnor
  g1649
  (
    n1042,
    n507,
    n473,
    n381,
    n397
  );


  nand
  g1650
  (
    n1177,
    n303,
    n487,
    n479,
    n394
  );


  xnor
  g1651
  (
    n1440,
    n325,
    n661,
    n299,
    n639
  );


  and
  g1652
  (
    n1221,
    n305,
    n618,
    n321,
    n178
  );


  and
  g1653
  (
    n968,
    n391,
    n335,
    n454,
    n420
  );


  or
  g1654
  (
    n959,
    n649,
    n251,
    n254,
    n298
  );


  and
  g1655
  (
    n1249,
    n328,
    n177,
    n182,
    n522
  );


  xor
  g1656
  (
    n1105,
    n325,
    n591,
    n386,
    n253
  );


  or
  g1657
  (
    n679,
    n410,
    n334,
    n296,
    n494
  );


  xor
  g1658
  (
    n1185,
    n583,
    n271,
    n622,
    n418
  );


  and
  g1659
  (
    n1738,
    n436,
    n509,
    n552,
    n244
  );


  nand
  g1660
  (
    n1150,
    n504,
    n336,
    n573,
    n217
  );


  and
  g1661
  (
    n1115,
    n506,
    n564,
    n189,
    n575
  );


  and
  g1662
  (
    n940,
    n489,
    n500,
    n166,
    n376
  );


  or
  g1663
  (
    n1623,
    n658,
    n515,
    n523,
    n243
  );


  nor
  g1664
  (
    n851,
    n528,
    n253,
    n637,
    n511
  );


  and
  g1665
  (
    n1597,
    n508,
    n376,
    n308,
    n395
  );


  nand
  g1666
  (
    n1007,
    n569,
    n663,
    n380,
    n213
  );


  xor
  g1667
  (
    n1618,
    n493,
    n642,
    n434,
    n666
  );


  xor
  g1668
  (
    n1191,
    n493,
    n193,
    n462,
    n253
  );


  and
  g1669
  (
    n1034,
    n307,
    n292,
    n259,
    n465
  );


  or
  g1670
  (
    n989,
    n574,
    n254,
    n207,
    n348
  );


  xnor
  g1671
  (
    n803,
    n228,
    n500,
    n615,
    n486
  );


  xnor
  g1672
  (
    n698,
    n279,
    n208,
    n606,
    n300
  );


  xnor
  g1673
  (
    n1023,
    n165,
    n216,
    n235,
    n310
  );


  nand
  g1674
  (
    n998,
    n473,
    n416,
    n369,
    n460
  );


  or
  g1675
  (
    n1159,
    n316,
    n226,
    n631,
    n468
  );


  nor
  g1676
  (
    n1383,
    n458,
    n566,
    n241,
    n607
  );


  nand
  g1677
  (
    n1719,
    n531,
    n620,
    n441,
    n398
  );


  xnor
  g1678
  (
    n1413,
    n609,
    n419,
    n211,
    n204
  );


  xor
  g1679
  (
    n780,
    n289,
    n369,
    n288,
    n293
  );


  xnor
  g1680
  (
    n934,
    n242,
    n626,
    n210,
    n468
  );


  and
  g1681
  (
    n812,
    n669,
    n500,
    n289,
    n491
  );


  xor
  g1682
  (
    n1464,
    n223,
    n250,
    n619,
    n520
  );


  nand
  g1683
  (
    n687,
    n344,
    n312,
    n263,
    n203
  );


  nand
  g1684
  (
    n1548,
    n645,
    n246,
    n611,
    n595
  );


  xor
  g1685
  (
    n813,
    n648,
    n598,
    n261,
    n176
  );


  or
  g1686
  (
    n836,
    n629,
    n646,
    n607,
    n635
  );


  xor
  g1687
  (
    n860,
    n458,
    n486,
    n271,
    n390
  );


  and
  g1688
  (
    n991,
    n419,
    n352,
    n375,
    n594
  );


  xnor
  g1689
  (
    n785,
    n650,
    n660,
    n476,
    n550
  );


  xor
  g1690
  (
    n1054,
    n266,
    n164,
    n293,
    n499
  );


  and
  g1691
  (
    n1222,
    n200,
    n520,
    n225,
    n605
  );


  xnor
  g1692
  (
    n1039,
    n584,
    n394,
    n306,
    n642
  );


  nand
  g1693
  (
    n938,
    n597,
    n176,
    n413,
    n402
  );


  or
  g1694
  (
    n922,
    n667,
    n588,
    n434,
    n227
  );


  and
  g1695
  (
    n1452,
    n578,
    n481,
    n360,
    n379
  );


  nor
  g1696
  (
    n1147,
    n268,
    n489,
    n398,
    n309
  );


  nand
  g1697
  (
    n1136,
    n415,
    n648,
    n493,
    n561
  );


  xnor
  g1698
  (
    n1336,
    n649,
    n295,
    n625,
    n397
  );


  nor
  g1699
  (
    n725,
    n449,
    n609,
    n599,
    n323
  );


  xor
  g1700
  (
    n1287,
    n272,
    n328,
    n317,
    n571
  );


  or
  g1701
  (
    n709,
    n187,
    n187,
    n347,
    n579
  );


  or
  g1702
  (
    n743,
    n224,
    n480,
    n286,
    n430
  );


  xnor
  g1703
  (
    n920,
    n291,
    n559,
    n422,
    n225
  );


  or
  g1704
  (
    n1366,
    n572,
    n620,
    n487,
    n639
  );


  or
  g1705
  (
    n1375,
    n333,
    n372,
    n607,
    n240
  );


  or
  g1706
  (
    n693,
    n199,
    n644,
    n386,
    n461
  );


  xnor
  g1707
  (
    n1020,
    n503,
    n202,
    n301,
    n249
  );


  nor
  g1708
  (
    n950,
    n448,
    n321,
    n521,
    n334
  );


  xnor
  g1709
  (
    n1119,
    n446,
    n273,
    n545,
    n268
  );


  xor
  g1710
  (
    n1552,
    n543,
    n354,
    n203,
    n200
  );


  or
  g1711
  (
    n1565,
    n179,
    n366,
    n193,
    n364
  );


  xor
  g1712
  (
    n765,
    n443,
    n513,
    n339,
    n317
  );


  nor
  g1713
  (
    n868,
    n641,
    n275,
    n647,
    n492
  );


  or
  g1714
  (
    n797,
    n377,
    n319,
    n196,
    n535
  );


  xnor
  g1715
  (
    n1404,
    n534,
    n352,
    n257,
    n568
  );


  xor
  g1716
  (
    n1447,
    n230,
    n161,
    n504,
    n532
  );


  or
  g1717
  (
    n1625,
    n509,
    n524,
    n202,
    n271
  );


  or
  g1718
  (
    n1349,
    n580,
    n641,
    n559,
    n664
  );


  nor
  g1719
  (
    n1753,
    n239,
    n483,
    n333,
    n425
  );


  or
  g1720
  (
    n1111,
    n457,
    n522,
    n342,
    n412
  );


  nand
  g1721
  (
    n1566,
    n396,
    n311,
    n588,
    n414
  );


  xnor
  g1722
  (
    n1430,
    n377,
    n527,
    n195,
    n547
  );


  or
  g1723
  (
    n1828,
    n1411,
    n1125,
    n699,
    n1005
  );


  nor
  g1724
  (
    n1803,
    n1466,
    n1457,
    n1095,
    n1322
  );


  and
  g1725
  (
    n1875,
    n1107,
    n701,
    n1078,
    n764
  );


  nor
  g1726
  (
    n1937,
    n1543,
    n876,
    n1002,
    n1140
  );


  xnor
  g1727
  (
    n1974,
    n697,
    n681,
    n822,
    n1009
  );


  and
  g1728
  (
    n1938,
    n736,
    n1519,
    n944,
    n1077
  );


  or
  g1729
  (
    n1944,
    n1309,
    n1415,
    n1000,
    n1385
  );


  nor
  g1730
  (
    n1895,
    n965,
    n1418,
    n938,
    n1151
  );


  xnor
  g1731
  (
    n1869,
    n1004,
    n783,
    n1093,
    n812
  );


  nor
  g1732
  (
    n1786,
    n1282,
    n1266,
    n759,
    n890
  );


  xor
  g1733
  (
    n1827,
    n1513,
    n1556,
    n1369,
    n927
  );


  or
  g1734
  (
    n1772,
    n904,
    n1485,
    n1269,
    n1067
  );


  xor
  g1735
  (
    n1776,
    n884,
    n1034,
    n1316,
    n709
  );


  nor
  g1736
  (
    n1864,
    n1392,
    n831,
    n1241,
    n1353
  );


  xnor
  g1737
  (
    n1906,
    n939,
    n1390,
    n1131,
    n794
  );


  nand
  g1738
  (
    n1964,
    n1482,
    n1440,
    n870,
    n685
  );


  xnor
  g1739
  (
    n1812,
    n1535,
    n719,
    n1044,
    n982
  );


  xnor
  g1740
  (
    n1867,
    n1033,
    n882,
    n1031,
    n676
  );


  nor
  g1741
  (
    n1760,
    n1202,
    n898,
    n715,
    n718
  );


  nand
  g1742
  (
    n1943,
    n1303,
    n752,
    n1285,
    n1435
  );


  xnor
  g1743
  (
    n1777,
    n1141,
    n855,
    n1356,
    n1366
  );


  xor
  g1744
  (
    n1785,
    n1348,
    n1341,
    n1329,
    n1335
  );


  or
  g1745
  (
    n1890,
    n1120,
    n829,
    n1003,
    n1352
  );


  and
  g1746
  (
    n1947,
    n991,
    n1299,
    n1134,
    n1511
  );


  nor
  g1747
  (
    n1765,
    n802,
    n960,
    n1532,
    n843
  );


  nand
  g1748
  (
    n1914,
    n1110,
    n1247,
    n1340,
    n826
  );


  xnor
  g1749
  (
    n1955,
    n1239,
    n1453,
    n1219,
    n1001
  );


  or
  g1750
  (
    n1782,
    n1458,
    n1441,
    n1200,
    n1289
  );


  nor
  g1751
  (
    n1833,
    n1342,
    n1126,
    n837,
    n1186
  );


  xor
  g1752
  (
    n1800,
    n1379,
    n1150,
    n1307,
    n1063
  );


  nor
  g1753
  (
    n1952,
    n1223,
    n707,
    n1419,
    n780
  );


  nor
  g1754
  (
    n1807,
    n1267,
    n1087,
    n912,
    n952
  );


  xnor
  g1755
  (
    n1797,
    n1483,
    n962,
    n797,
    n1445
  );


  nand
  g1756
  (
    n1961,
    n1117,
    n1400,
    n1235,
    n911
  );


  xnor
  g1757
  (
    n1894,
    n1069,
    n1544,
    n1298,
    n951
  );


  nor
  g1758
  (
    KeyWire_0_7,
    n1011,
    n1060,
    n1128,
    n955
  );


  nor
  g1759
  (
    n1926,
    n1148,
    n909,
    n1270,
    n777
  );


  xnor
  g1760
  (
    n1790,
    n842,
    n1550,
    n770,
    n969
  );


  xor
  g1761
  (
    n1884,
    n1048,
    n1103,
    n1156,
    n1553
  );


  nand
  g1762
  (
    n1927,
    n1066,
    n804,
    n918,
    n1130
  );


  nor
  g1763
  (
    n1769,
    n1030,
    n1104,
    n924,
    n1451
  );


  xor
  g1764
  (
    n1929,
    n1275,
    n1305,
    n992,
    n1055
  );


  nor
  g1765
  (
    n1791,
    n1091,
    n793,
    n728,
    n756
  );


  xnor
  g1766
  (
    n1945,
    n1177,
    n1053,
    n1010,
    n983
  );


  nor
  g1767
  (
    n1792,
    n782,
    n1507,
    n1334,
    n1191
  );


  and
  g1768
  (
    n1868,
    n1430,
    n753,
    n865,
    n1448
  );


  nand
  g1769
  (
    KeyWire_0_15,
    n838,
    n1398,
    n762,
    n1008
  );


  xor
  g1770
  (
    n1789,
    n1509,
    n1173,
    n946,
    n1315
  );


  or
  g1771
  (
    n1768,
    n928,
    n920,
    n1076,
    n1047
  );


  nand
  g1772
  (
    n1842,
    n1070,
    n791,
    n1234,
    n1492
  );


  nor
  g1773
  (
    n1932,
    n925,
    n1163,
    n990,
    n1264
  );


  or
  g1774
  (
    n1784,
    n716,
    n700,
    n808,
    n1115
  );


  nor
  g1775
  (
    n1925,
    n1064,
    n726,
    n1288,
    n806
  );


  nand
  g1776
  (
    n1872,
    n1368,
    n1490,
    n1185,
    n887
  );


  nor
  g1777
  (
    n1761,
    n844,
    n1487,
    n1074,
    n1142
  );


  nor
  g1778
  (
    n1969,
    n1268,
    n795,
    n1508,
    n1488
  );


  nor
  g1779
  (
    n1781,
    n1319,
    n981,
    n1536,
    n828
  );


  and
  g1780
  (
    n1954,
    n908,
    n1549,
    n673,
    n1176
  );


  and
  g1781
  (
    n1770,
    n1438,
    n1478,
    n1479,
    n1024
  );


  xor
  g1782
  (
    n1885,
    n799,
    n760,
    n1221,
    n1263
  );


  xor
  g1783
  (
    n1951,
    n910,
    n926,
    n739,
    n931
  );


  and
  g1784
  (
    n1933,
    n1215,
    n734,
    n1372,
    n1327
  );


  or
  g1785
  (
    n1787,
    n1217,
    n1539,
    n714,
    n1481
  );


  nor
  g1786
  (
    n1907,
    n1073,
    n1542,
    n919,
    n967
  );


  or
  g1787
  (
    n1801,
    n1442,
    n1362,
    n1165,
    n1343
  );


  nor
  g1788
  (
    n1919,
    n901,
    n833,
    n1286,
    n1218
  );


  nand
  g1789
  (
    n1901,
    n1155,
    n1465,
    n1548,
    n906
  );


  xor
  g1790
  (
    n1936,
    n1374,
    n712,
    n773,
    n1265
  );


  xnor
  g1791
  (
    n1826,
    n1522,
    n775,
    n1251,
    n1039
  );


  nor
  g1792
  (
    n1891,
    n1434,
    n1297,
    n1258,
    n1321
  );


  xnor
  g1793
  (
    n1880,
    n1083,
    n1099,
    n1431,
    n819
  );


  or
  g1794
  (
    n1840,
    n1198,
    n824,
    n1059,
    n1138
  );


  nor
  g1795
  (
    n1923,
    n1109,
    n948,
    n805,
    n1377
  );


  nand
  g1796
  (
    n1910,
    n809,
    n1486,
    n1171,
    n866
  );


  xnor
  g1797
  (
    n1930,
    n1456,
    n689,
    n1312,
    n1405
  );


  nand
  g1798
  (
    n1878,
    n1058,
    n1496,
    n1037,
    n933
  );


  nand
  g1799
  (
    n1900,
    n1162,
    n1231,
    n1450,
    n1455
  );


  or
  g1800
  (
    n1892,
    n1132,
    n1273,
    n914,
    n861
  );


  xor
  g1801
  (
    n1928,
    n774,
    n1175,
    n1359,
    n747
  );


  nand
  g1802
  (
    n1897,
    n1524,
    n954,
    n1293,
    n1021
  );


  nor
  g1803
  (
    n1820,
    n1170,
    n1228,
    n684,
    n1245
  );


  or
  g1804
  (
    n1799,
    n690,
    n742,
    n1330,
    n1133
  );


  or
  g1805
  (
    n1845,
    n973,
    n696,
    n1537,
    n1401
  );


  and
  g1806
  (
    n1810,
    n1279,
    n1262,
    n1014,
    n1197
  );


  xnor
  g1807
  (
    n1796,
    n1408,
    n1178,
    n1046,
    n680
  );


  nor
  g1808
  (
    n1822,
    n1404,
    n1506,
    n1236,
    n1546
  );


  nor
  g1809
  (
    n1870,
    n860,
    n953,
    n1308,
    n1261
  );


  xor
  g1810
  (
    n1759,
    n1394,
    n1157,
    n1462,
    n1504
  );


  nand
  g1811
  (
    n1911,
    n1444,
    n1409,
    n897,
    n1291
  );


  xnor
  g1812
  (
    n1905,
    n811,
    n1499,
    n1493,
    n737
  );


  nor
  g1813
  (
    n1946,
    n1439,
    n1244,
    n1213,
    n993
  );


  nand
  g1814
  (
    n1811,
    n1347,
    n1238,
    n871,
    n750
  );


  and
  g1815
  (
    n1798,
    n1233,
    n1025,
    n1056,
    n1407
  );


  nor
  g1816
  (
    n1950,
    n1272,
    n856,
    n1169,
    n1475
  );


  or
  g1817
  (
    n1832,
    n1022,
    n1470,
    n916,
    n1338
  );


  nand
  g1818
  (
    n1831,
    n741,
    n743,
    n731,
    n1295
  );


  nand
  g1819
  (
    n1824,
    n698,
    n823,
    n1274,
    n1443
  );


  xnor
  g1820
  (
    n1848,
    n976,
    n1357,
    n1183,
    n694
  );


  nor
  g1821
  (
    n1939,
    n724,
    n1193,
    n1210,
    n1413
  );


  and
  g1822
  (
    n1918,
    n1437,
    n1154,
    n1512,
    n1380
  );


  nand
  g1823
  (
    n1970,
    n1160,
    n1038,
    n1029,
    n1127
  );


  or
  g1824
  (
    n1802,
    n949,
    n1300,
    n1139,
    n1242
  );


  and
  g1825
  (
    n1876,
    n1480,
    n1187,
    n692,
    n1311
  );


  or
  g1826
  (
    n1865,
    n1360,
    n1510,
    n1211,
    n1015
  );


  nand
  g1827
  (
    n1942,
    n1433,
    n1007,
    n979,
    n853
  );


  xor
  g1828
  (
    n1956,
    n847,
    n1081,
    n917,
    n711
  );


  or
  g1829
  (
    n1843,
    n1079,
    n1153,
    n836,
    n961
  );


  nand
  g1830
  (
    n1757,
    n723,
    n1019,
    n970,
    n1534
  );


  xnor
  g1831
  (
    n1778,
    n1518,
    n1469,
    n825,
    n935
  );


  xnor
  g1832
  (
    n1941,
    n1246,
    n1084,
    n1209,
    n1112
  );


  xor
  g1833
  (
    n1958,
    n1189,
    n1129,
    n929,
    n1318
  );


  or
  g1834
  (
    n1758,
    n846,
    n705,
    n921,
    n980
  );


  xor
  g1835
  (
    n1780,
    n1052,
    n942,
    n1375,
    n1459
  );


  and
  g1836
  (
    n1899,
    n787,
    n1194,
    n851,
    n1461
  );


  xor
  g1837
  (
    n1836,
    n1495,
    n1026,
    n803,
    n796
  );


  xor
  g1838
  (
    n1963,
    n1477,
    n1425,
    n987,
    n1012
  );


  and
  g1839
  (
    n1816,
    n1363,
    n1473,
    n1382,
    n1152
  );


  xnor
  g1840
  (
    n1775,
    n883,
    n1061,
    n1422,
    n978
  );


  xor
  g1841
  (
    n1793,
    n895,
    n1088,
    n1023,
    n757
  );


  xnor
  g1842
  (
    n1808,
    n781,
    n708,
    n720,
    n821
  );


  or
  g1843
  (
    n1771,
    n1500,
    n998,
    n1147,
    n859
  );


  xnor
  g1844
  (
    n1877,
    n1471,
    n784,
    n1224,
    n820
  );


  and
  g1845
  (
    n1904,
    n1158,
    n879,
    n1424,
    n758
  );


  nand
  g1846
  (
    n1830,
    n868,
    n755,
    n999,
    n1119
  );


  nor
  g1847
  (
    n1966,
    n1420,
    n869,
    n679,
    n1460
  );


  and
  g1848
  (
    n1839,
    n1167,
    n971,
    n1136,
    n880
  );


  or
  g1849
  (
    n1852,
    n1421,
    n1230,
    n874,
    n1092
  );


  nor
  g1850
  (
    n1861,
    n1497,
    n1237,
    n1124,
    n1324
  );


  or
  g1851
  (
    n1959,
    n674,
    n761,
    n872,
    n858
  );


  xnor
  g1852
  (
    n1846,
    n1116,
    n801,
    n875,
    n768
  );


  or
  g1853
  (
    n1887,
    n1277,
    n997,
    n767,
    n1317
  );


  nand
  g1854
  (
    n1896,
    n1551,
    n1020,
    n1314,
    n857
  );


  and
  g1855
  (
    n1815,
    n1476,
    n848,
    n922,
    n957
  );


  and
  g1856
  (
    n1774,
    n816,
    n1123,
    n1503,
    n963
  );


  and
  g1857
  (
    n1949,
    n1402,
    n1412,
    n1086,
    n810
  );


  xor
  g1858
  (
    n1809,
    n943,
    n1339,
    n1351,
    n852
  );


  nor
  g1859
  (
    n1849,
    n1166,
    n1057,
    n746,
    n827
  );


  or
  g1860
  (
    n1819,
    n867,
    n1344,
    n1036,
    n1096
  );


  nor
  g1861
  (
    n1940,
    n1468,
    n900,
    n899,
    n1252
  );


  or
  g1862
  (
    n1886,
    n677,
    n1051,
    n958,
    n1065
  );


  nor
  g1863
  (
    n1934,
    n1484,
    n772,
    n1216,
    n989
  );


  and
  g1864
  (
    n1920,
    n1523,
    n1525,
    n779,
    n1035
  );


  nor
  g1865
  (
    n1883,
    n1547,
    n903,
    n1489,
    n1367
  );


  xnor
  g1866
  (
    n1814,
    n721,
    n1208,
    n995,
    n1414
  );


  nor
  g1867
  (
    n1871,
    n1017,
    n873,
    n1101,
    n792
  );


  xor
  g1868
  (
    n1968,
    n1370,
    n1041,
    n1391,
    n854
  );


  or
  g1869
  (
    n1857,
    n1206,
    n940,
    n902,
    n678
  );


  xnor
  g1870
  (
    n1841,
    n1280,
    n1332,
    n1336,
    n710
  );


  xnor
  g1871
  (
    n1863,
    n1199,
    n702,
    n1089,
    n915
  );


  nor
  g1872
  (
    n1851,
    n1174,
    n748,
    n1529,
    n1098
  );


  xnor
  g1873
  (
    n1859,
    n1082,
    n1355,
    n814,
    n1260
  );


  and
  g1874
  (
    n1823,
    n934,
    n1201,
    n786,
    n1517
  );


  xor
  g1875
  (
    n1881,
    n1122,
    n1205,
    n1429,
    n1361
  );


  or
  g1876
  (
    n1957,
    n735,
    n1491,
    n1204,
    n704
  );


  nand
  g1877
  (
    n1804,
    n1278,
    n850,
    n1250,
    n1325
  );


  or
  g1878
  (
    n1975,
    n1384,
    n1555,
    n1304,
    n1257
  );


  nand
  g1879
  (
    n1756,
    n830,
    n1530,
    n1259,
    n945
  );


  and
  g1880
  (
    n1818,
    n751,
    n1521,
    n687,
    n974
  );


  and
  g1881
  (
    n1967,
    n1190,
    n1159,
    n1399,
    n800
  );


  or
  g1882
  (
    n1829,
    n695,
    n894,
    n1214,
    n877
  );


  or
  g1883
  (
    n1971,
    n1393,
    n725,
    n1323,
    n1406
  );


  and
  g1884
  (
    n1873,
    n1331,
    n1386,
    n688,
    n984
  );


  xor
  g1885
  (
    n1893,
    n1149,
    n1527,
    n1387,
    n1164
  );


  nor
  g1886
  (
    n1921,
    n1533,
    n950,
    n947,
    n932
  );


  and
  g1887
  (
    n1912,
    n744,
    n839,
    n1062,
    n675
  );


  nand
  g1888
  (
    n1856,
    n1068,
    n1281,
    n749,
    n683
  );


  xnor
  g1889
  (
    n1835,
    n1220,
    n732,
    n1222,
    n1097
  );


  xnor
  g1890
  (
    n1909,
    n1436,
    n1464,
    n1310,
    n1108
  );


  xnor
  g1891
  (
    n1953,
    n1102,
    n1232,
    n807,
    n1472
  );


  or
  g1892
  (
    n1766,
    n849,
    n1196,
    n1410,
    n1515
  );


  and
  g1893
  (
    n1972,
    n1049,
    n745,
    n729,
    n1114
  );


  nand
  g1894
  (
    n1844,
    n785,
    n1075,
    n1182,
    n1179
  );


  and
  g1895
  (
    n1855,
    n936,
    n1446,
    n1313,
    n727
  );


  nor
  g1896
  (
    n1825,
    n1395,
    n1137,
    n964,
    n864
  );


  xnor
  g1897
  (
    n1834,
    n896,
    n818,
    n923,
    n1294
  );


  nor
  g1898
  (
    n1817,
    n1195,
    n1498,
    n1416,
    n1447
  );


  or
  g1899
  (
    n1853,
    n1243,
    n905,
    n813,
    n754
  );


  and
  g1900
  (
    n1889,
    n1188,
    n790,
    n1463,
    n1301
  );


  and
  g1901
  (
    n1866,
    n1271,
    n988,
    n703,
    n996
  );


  xor
  g1902
  (
    n1858,
    n1143,
    n1094,
    n1432,
    n1105
  );


  xor
  g1903
  (
    n1762,
    n885,
    n1423,
    n1145,
    n1383
  );


  xor
  g1904
  (
    n1850,
    n862,
    n959,
    n1373,
    n771
  );


  xnor
  g1905
  (
    n1962,
    n1276,
    n1388,
    n878,
    n788
  );


  or
  g1906
  (
    n1960,
    n1287,
    n1528,
    n1545,
    n1050
  );


  and
  g1907
  (
    n1794,
    n1505,
    n1520,
    n1516,
    n1474
  );


  and
  g1908
  (
    n1763,
    n713,
    n1080,
    n891,
    n893
  );


  xor
  g1909
  (
    n1805,
    n1292,
    n1172,
    n930,
    n1121
  );


  nand
  g1910
  (
    n1915,
    n1376,
    n1042,
    n722,
    n778
  );


  nand
  g1911
  (
    n1838,
    n1333,
    n1192,
    n776,
    n1502
  );


  or
  g1912
  (
    n1854,
    n1346,
    n1354,
    n845,
    n1349
  );


  nor
  g1913
  (
    n1813,
    n733,
    n1426,
    n789,
    n717
  );


  and
  g1914
  (
    n1795,
    n1161,
    n1350,
    n1146,
    n1552
  );


  nand
  g1915
  (
    n1862,
    n738,
    n1358,
    n1144,
    n1255
  );


  nand
  g1916
  (
    n1888,
    n706,
    n1427,
    n913,
    n886
  );


  xor
  g1917
  (
    n1764,
    n1328,
    n863,
    n1180,
    n1326
  );


  nand
  g1918
  (
    n1773,
    n1027,
    n1296,
    n1302,
    n1203
  );


  nor
  g1919
  (
    n1913,
    n691,
    n1106,
    n1090,
    n730
  );


  nand
  g1920
  (
    n1965,
    n817,
    n682,
    n1514,
    n1054
  );


  or
  g1921
  (
    n1924,
    n986,
    n1118,
    n1541,
    n835
  );


  xnor
  g1922
  (
    n1882,
    n977,
    n1454,
    n1085,
    n1337
  );


  xnor
  g1923
  (
    n1879,
    n1378,
    n889,
    n693,
    n994
  );


  or
  g1924
  (
    n1902,
    n798,
    n1113,
    n1253,
    n1100
  );


  xnor
  g1925
  (
    n1860,
    n1212,
    n1028,
    n1389,
    n1494
  );


  or
  g1926
  (
    n1917,
    n1538,
    n1006,
    n1135,
    n1254
  );


  nand
  g1927
  (
    n1821,
    n763,
    n968,
    n1168,
    n1403
  );


  or
  g1928
  (
    n1788,
    n941,
    n1345,
    n1381,
    n1111
  );


  xnor
  g1929
  (
    n1908,
    n686,
    n888,
    n1043,
    n1467
  );


  xor
  g1930
  (
    n1806,
    n1248,
    n1227,
    n1240,
    n1032
  );


  xnor
  g1931
  (
    n1916,
    n1045,
    n1181,
    n765,
    n1501
  );


  or
  g1932
  (
    n1903,
    n966,
    n1207,
    n1526,
    n740
  );


  nand
  g1933
  (
    n1898,
    n840,
    n815,
    n975,
    n1554
  );


  xor
  g1934
  (
    n1847,
    n1225,
    n841,
    n1531,
    n907
  );


  nand
  g1935
  (
    n1935,
    n956,
    n1417,
    n1016,
    n1452
  );


  nand
  g1936
  (
    n1922,
    n937,
    n1229,
    n1184,
    n1449
  );


  xnor
  g1937
  (
    n1783,
    n769,
    n1397,
    n1072,
    n1365
  );


  nor
  g1938
  (
    n1767,
    n892,
    n1396,
    n1283,
    n766
  );


  and
  g1939
  (
    n1837,
    n1306,
    n1364,
    n834,
    n832
  );


  nand
  g1940
  (
    n1931,
    n1040,
    n1256,
    n1018,
    n1071
  );


  and
  g1941
  (
    n1976,
    n1290,
    n1540,
    n1371,
    n985
  );


  xor
  g1942
  (
    n1874,
    n972,
    n1320,
    n1013,
    n881
  );


  or
  g1943
  (
    n1973,
    n1428,
    n1226,
    n1249,
    n1284
  );


  nand
  g1944
  (
    n1993,
    n1768,
    n1824,
    n1809,
    n1783
  );


  and
  g1945
  (
    n1977,
    n1823,
    n1775,
    n1781,
    n1807
  );


  or
  g1946
  (
    n1978,
    n1808,
    n1759,
    n1761,
    n1773
  );


  nor
  g1947
  (
    n1982,
    n1756,
    n1825,
    n1805,
    n1803
  );


  xor
  g1948
  (
    n1979,
    n1802,
    n1758,
    n1763,
    n1795
  );


  xnor
  g1949
  (
    n1992,
    n1777,
    n1814,
    n1779,
    n1800
  );


  or
  g1950
  (
    n1981,
    n1812,
    n1766,
    n1796,
    n1790
  );


  xnor
  g1951
  (
    n1980,
    n1770,
    n1827,
    n1810,
    n1769
  );


  or
  g1952
  (
    n1985,
    n1806,
    n1811,
    n1797,
    n1801
  );


  or
  g1953
  (
    n1986,
    n1782,
    n1774,
    n1780,
    n1804
  );


  xor
  g1954
  (
    n1983,
    n1776,
    n1784,
    n1760,
    n1787
  );


  nor
  g1955
  (
    n1988,
    n1817,
    n1771,
    n1798,
    n1764
  );


  nand
  g1956
  (
    n1987,
    n1799,
    n1818,
    n1791,
    n1813
  );


  xnor
  g1957
  (
    n1984,
    n1785,
    n1821,
    n1757,
    n1819
  );


  and
  g1958
  (
    n1990,
    n1793,
    n1816,
    n1815,
    n1820
  );


  xnor
  g1959
  (
    n1991,
    n1765,
    n1772,
    n1822,
    n1826
  );


  nand
  g1960
  (
    n1994,
    n1778,
    n1789,
    n1788,
    n1786
  );


  xor
  g1961
  (
    n1989,
    n1762,
    n1792,
    n1767,
    n1794
  );


  nand
  g1962
  (
    n2010,
    n1829,
    n1879,
    n1837,
    n1868
  );


  or
  g1963
  (
    n2005,
    n1876,
    n1866,
    n1832,
    n1869
  );


  or
  g1964
  (
    n2002,
    n1853,
    n1982,
    n1855,
    n1991
  );


  nand
  g1965
  (
    n2001,
    n1988,
    n1987,
    n1849,
    n1872
  );


  and
  g1966
  (
    n2008,
    n1850,
    n1834,
    n1877,
    n1862
  );


  xor
  g1967
  (
    n1995,
    n1860,
    n1992,
    n1993,
    n1843
  );


  and
  g1968
  (
    n2003,
    n1844,
    n1839,
    n1847,
    n1983
  );


  nor
  g1969
  (
    n1997,
    n1864,
    n1833,
    n1977,
    n1989
  );


  nand
  g1970
  (
    n1999,
    n1854,
    n1985,
    n1870,
    n1859
  );


  or
  g1971
  (
    n2011,
    n1842,
    n1828,
    n1835,
    n1986
  );


  xor
  g1972
  (
    n2012,
    n1857,
    n1867,
    n1984,
    n1851
  );


  nor
  g1973
  (
    n2007,
    n1856,
    n1990,
    n1845,
    n1861
  );


  nand
  g1974
  (
    n1998,
    n1846,
    n1880,
    n1831,
    n1978
  );


  xor
  g1975
  (
    n1996,
    n1840,
    n1848,
    n1830,
    n1881
  );


  and
  g1976
  (
    n2004,
    n1873,
    n1980,
    n1865,
    n1994
  );


  nand
  g1977
  (
    n2006,
    n1878,
    n1852,
    n1836,
    n1838
  );


  xnor
  g1978
  (
    n2009,
    n1841,
    n1863,
    n1874,
    n1979
  );


  xnor
  g1979
  (
    n2000,
    n1858,
    n1871,
    n1981,
    n1875
  );


  buf
  g1980
  (
    n2013,
    n1566
  );


  buf
  g1981
  (
    n2019,
    n1558
  );


  not
  g1982
  (
    n2020,
    n1557
  );


  buf
  g1983
  (
    n2018,
    n1996
  );


  not
  g1984
  (
    n2021,
    n1560
  );


  nor
  g1985
  (
    n2014,
    n1997,
    n1559,
    n1996
  );


  nand
  g1986
  (
    n2017,
    n1995,
    n1996,
    n1563
  );


  nand
  g1987
  (
    n2022,
    n1564,
    n1995,
    n1562
  );


  xor
  g1988
  (
    n2015,
    n1995,
    n1561,
    n1997
  );


  and
  g1989
  (
    n2016,
    n1996,
    n1565,
    n1995
  );


  buf
  g1990
  (
    n2029,
    n2021
  );


  buf
  g1991
  (
    n2023,
    n2013
  );


  not
  g1992
  (
    n2028,
    n1885
  );


  not
  g1993
  (
    n2025,
    n1569
  );


  buf
  g1994
  (
    n2026,
    n2019
  );


  not
  g1995
  (
    n2027,
    n2014
  );


  or
  g1996
  (
    n2024,
    n1567,
    n2017,
    n2015,
    n1883
  );


  xnor
  g1997
  (
    n2031,
    n2020,
    n1568,
    n1884,
    n1571
  );


  nor
  g1998
  (
    n2030,
    n2018,
    n1882,
    n2016,
    n1570
  );


  buf
  g1999
  (
    n2034,
    n1573
  );


  buf
  g2000
  (
    n2033,
    n2023
  );


  nand
  g2001
  (
    n2032,
    n1574,
    n1572,
    n2025,
    n2024
  );


  xnor
  g2002
  (
    n2036,
    n1576,
    n2033
  );


  nand
  g2003
  (
    n2035,
    n1575,
    n2032
  );


  nor
  g2004
  (
    n2037,
    n1888,
    n1886,
    n2035,
    n1887
  );


  buf
  g2005
  (
    n2039,
    n2037
  );


  buf
  g2006
  (
    n2038,
    n2037
  );


  buf
  g2007
  (
    n2042,
    n2039
  );


  not
  g2008
  (
    n2041,
    n2038
  );


  not
  g2009
  (
    n2044,
    n2038
  );


  not
  g2010
  (
    n2046,
    n2038
  );


  not
  g2011
  (
    n2043,
    n2039
  );


  not
  g2012
  (
    n2047,
    n2039
  );


  buf
  g2013
  (
    n2040,
    n2038
  );


  not
  g2014
  (
    n2045,
    n2039
  );


  xnor
  g2015
  (
    n2054,
    n1890,
    n2026,
    n2046
  );


  xnor
  g2016
  (
    n2048,
    n2047,
    n2029,
    n2041
  );


  xnor
  g2017
  (
    n2049,
    n1891,
    n2027,
    n2030,
    n2046
  );


  nand
  g2018
  (
    n2050,
    n1889,
    n2029,
    n2047,
    n2031
  );


  nand
  g2019
  (
    n2053,
    n2043,
    n2042,
    n2045,
    n2030
  );


  and
  g2020
  (
    n2051,
    n2046,
    n2030,
    n2044
  );


  xor
  g2021
  (
    n2052,
    n2040,
    n2029,
    n2031,
    n2028
  );


  not
  g2022
  (
    n2056,
    n2052
  );


  xor
  g2023
  (
    n2055,
    n2051,
    n2053,
    n1577
  );


  or
  g2024
  (
    n2057,
    n2050,
    n2054,
    n2031,
    n1578
  );


  and
  g2025
  (
    n2058,
    n1898,
    n1892
  );


  xor
  g2026
  (
    n2059,
    n2055,
    n1895,
    n1899,
    n2057
  );


  and
  g2027
  (
    n2060,
    n1896,
    n2057,
    n2034
  );


  xnor
  g2028
  (
    n2061,
    n1893,
    n1894,
    n2056,
    n1897
  );


  not
  g2029
  (
    n2066,
    n1582
  );


  or
  g2030
  (
    n2064,
    n2047,
    n2061
  );


  xnor
  g2031
  (
    n2063,
    n2059,
    n1579,
    n672,
    n2047
  );


  and
  g2032
  (
    n2062,
    n2036,
    n2058,
    n1581,
    n2060
  );


  nor
  g2033
  (
    n2065,
    n1580,
    n672
  );


  xor
  g2034
  (
    n2067,
    n1591,
    n1586,
    n2065,
    n1593
  );


  nand
  g2035
  (
    n2070,
    n2064,
    n1587,
    n2063,
    n1583
  );


  and
  g2036
  (
    n2069,
    n1589,
    n1584,
    n2066,
    n1590
  );


  xor
  g2037
  (
    n2068,
    n1588,
    n1585,
    n1594,
    n1592
  );


  and
  g2038
  (
    n2071,
    n2070,
    n1907,
    n1910,
    n1901
  );


  and
  g2039
  (
    n2072,
    n1914,
    n1921,
    n1922,
    n2067
  );


  nor
  g2040
  (
    n2078,
    n1911,
    n1917,
    n1920,
    n1900
  );


  xor
  g2041
  (
    n2076,
    n1913,
    n1902,
    n2069,
    n1903
  );


  nor
  g2042
  (
    n2073,
    n1918,
    n2069,
    n1915,
    n1906
  );


  nor
  g2043
  (
    n2075,
    n1916,
    n2068,
    n1909,
    n1904
  );


  nor
  g2044
  (
    n2074,
    n1908,
    n2070,
    n1905
  );


  and
  g2045
  (
    n2077,
    n1912,
    n1923,
    n2069,
    n1919
  );


  xnor
  g2046
  (
    n2081,
    n2076,
    n2077,
    n2075,
    n1597
  );


  or
  g2047
  (
    n2082,
    n1596,
    n1603,
    n1606,
    n1595
  );


  nand
  g2048
  (
    n2079,
    n1599,
    n1604,
    n1601,
    n1600
  );


  nor
  g2049
  (
    n2080,
    n1602,
    n1605,
    n1598,
    n2074
  );


  nand
  g2050
  (
    n2084,
    n1607,
    n1612,
    n1610,
    n1609
  );


  and
  g2051
  (
    n2083,
    n1611,
    n1608,
    n2081,
    n2082
  );


  buf
  g2052
  (
    n2085,
    n2084
  );


  not
  g2053
  (
    n2087,
    n2084
  );


  buf
  g2054
  (
    n2092,
    n2083
  );


  buf
  g2055
  (
    n2091,
    n2083
  );


  not
  g2056
  (
    n2089,
    n2084
  );


  buf
  g2057
  (
    n2088,
    n2083
  );


  nor
  g2058
  (
    n2086,
    n1925,
    n1927
  );


  or
  g2059
  (
    n2090,
    n1926,
    n2083,
    n1924,
    n2084
  );


  nor
  g2060
  (
    n2120,
    n2092,
    n2086
  );


  nor
  g2061
  (
    n2112,
    n2092,
    n1931
  );


  nor
  g2062
  (
    n2094,
    n1941,
    n1950
  );


  xor
  g2063
  (
    n2119,
    n2085,
    n1949
  );


  nand
  g2064
  (
    n2101,
    n1613,
    n1620
  );


  xnor
  g2065
  (
    n2113,
    n2091,
    n2092
  );


  xor
  g2066
  (
    n2107,
    n1952,
    n2091
  );


  and
  g2067
  (
    n2122,
    n1933,
    n1936
  );


  xnor
  g2068
  (
    n2109,
    n2090,
    n1614
  );


  xnor
  g2069
  (
    n2104,
    n1954,
    n1943
  );


  nand
  g2070
  (
    n2118,
    n1618,
    n1942
  );


  xor
  g2071
  (
    n2097,
    n1615,
    n2087
  );


  xor
  g2072
  (
    n2110,
    n1951,
    n1938
  );


  or
  g2073
  (
    n2116,
    n1955,
    n2091
  );


  nand
  g2074
  (
    n2099,
    n1940,
    n1947
  );


  nor
  g2075
  (
    n2108,
    n2085,
    n1934
  );


  nor
  g2076
  (
    n2111,
    n1944,
    n2085
  );


  nand
  g2077
  (
    n2093,
    n2088,
    n2087
  );


  or
  g2078
  (
    n2098,
    n2091,
    n1946
  );


  or
  g2079
  (
    n2106,
    n1619,
    n1957
  );


  xnor
  g2080
  (
    n2123,
    n2090,
    n2088
  );


  nor
  g2081
  (
    n2124,
    n2088,
    n2086
  );


  xor
  g2082
  (
    n2096,
    n1959,
    n2090
  );


  and
  g2083
  (
    n2117,
    n1929,
    n1958
  );


  nand
  g2084
  (
    n2114,
    n2092,
    n1953
  );


  xor
  g2085
  (
    n2121,
    n2089,
    n1935
  );


  nor
  g2086
  (
    n2103,
    n1617,
    n1616
  );


  or
  g2087
  (
    n2105,
    n2086,
    n1956
  );


  xnor
  g2088
  (
    n2100,
    n1930,
    n2087,
    n1948,
    n2086
  );


  and
  g2089
  (
    n2102,
    n1932,
    n2089,
    n1939,
    n2085
  );


  nor
  g2090
  (
    n2095,
    n1937,
    n2090,
    n2088,
    n2089
  );


  and
  g2091
  (
    n2115,
    n1945,
    n1928,
    n2087,
    n2089
  );


  buf
  g2092
  (
    n2147,
    n2008
  );


  not
  g2093
  (
    n2168,
    n2003
  );


  not
  g2094
  (
    n2153,
    n2121
  );


  not
  g2095
  (
    n2251,
    n2098
  );


  not
  g2096
  (
    n2148,
    n2003
  );


  buf
  g2097
  (
    n2134,
    n2123
  );


  not
  g2098
  (
    n2180,
    n2095
  );


  buf
  g2099
  (
    n2149,
    n2006
  );


  not
  g2100
  (
    n2170,
    n2006
  );


  not
  g2101
  (
    n2189,
    n2121
  );


  buf
  g2102
  (
    n2141,
    n2102
  );


  buf
  g2103
  (
    n2204,
    n1625
  );


  not
  g2104
  (
    n2211,
    n2001
  );


  buf
  g2105
  (
    n2240,
    n2106
  );


  buf
  g2106
  (
    n2249,
    n2094
  );


  buf
  g2107
  (
    n2209,
    n2119
  );


  not
  g2108
  (
    n2194,
    n2000
  );


  not
  g2109
  (
    n2139,
    n1632
  );


  buf
  g2110
  (
    n2238,
    n2117
  );


  not
  g2111
  (
    n2222,
    n2107
  );


  buf
  g2112
  (
    n2233,
    n2001
  );


  not
  g2113
  (
    n2129,
    n2093
  );


  not
  g2114
  (
    n2126,
    n2120
  );


  buf
  g2115
  (
    n2236,
    n2106
  );


  buf
  g2116
  (
    n2181,
    n2109
  );


  buf
  g2117
  (
    n2224,
    n2004
  );


  buf
  g2118
  (
    n2192,
    n2007
  );


  buf
  g2119
  (
    n2205,
    n2114
  );


  buf
  g2120
  (
    n2128,
    n2006
  );


  not
  g2121
  (
    n2230,
    n2006
  );


  buf
  g2122
  (
    n2164,
    n1630
  );


  not
  g2123
  (
    n2174,
    n2107
  );


  buf
  g2124
  (
    n2203,
    n2007
  );


  buf
  g2125
  (
    n2228,
    n2111
  );


  not
  g2126
  (
    n2132,
    n2119
  );


  not
  g2127
  (
    n2213,
    n2113
  );


  not
  g2128
  (
    n2138,
    n2009
  );


  not
  g2129
  (
    n2140,
    n2110
  );


  not
  g2130
  (
    n2166,
    n2112
  );


  not
  g2131
  (
    n2183,
    n2104
  );


  buf
  g2132
  (
    n2159,
    n2004
  );


  buf
  g2133
  (
    n2198,
    n2124
  );


  not
  g2134
  (
    n2235,
    n2115
  );


  not
  g2135
  (
    n2136,
    n2099
  );


  not
  g2136
  (
    n2229,
    n2100
  );


  buf
  g2137
  (
    n2185,
    n2104
  );


  not
  g2138
  (
    n2163,
    n2124
  );


  buf
  g2139
  (
    n2145,
    n2116
  );


  not
  g2140
  (
    n2169,
    n2118
  );


  not
  g2141
  (
    n2161,
    n2097
  );


  buf
  g2142
  (
    n2176,
    n2119
  );


  not
  g2143
  (
    n2154,
    n2093
  );


  buf
  g2144
  (
    n2207,
    n2118
  );


  not
  g2145
  (
    n2220,
    n2100
  );


  buf
  g2146
  (
    n2237,
    n2095
  );


  buf
  g2147
  (
    n2171,
    n2122
  );


  not
  g2148
  (
    n2208,
    n2094
  );


  not
  g2149
  (
    n2227,
    n2098
  );


  buf
  g2150
  (
    n2216,
    n1628
  );


  buf
  g2151
  (
    n2210,
    n2094
  );


  not
  g2152
  (
    n2156,
    n2112
  );


  buf
  g2153
  (
    n2223,
    n2005
  );


  not
  g2154
  (
    n2167,
    n2106
  );


  buf
  g2155
  (
    n2142,
    n2107
  );


  not
  g2156
  (
    n2218,
    n2120
  );


  buf
  g2157
  (
    n2195,
    n2110
  );


  buf
  g2158
  (
    n2152,
    n2001
  );


  buf
  g2159
  (
    n2125,
    n2113
  );


  buf
  g2160
  (
    n2162,
    n2000
  );


  not
  g2161
  (
    n2244,
    n1624
  );


  buf
  g2162
  (
    n2186,
    n2104
  );


  not
  g2163
  (
    n2242,
    n2005
  );


  not
  g2164
  (
    n2243,
    n2100
  );


  buf
  g2165
  (
    n2187,
    n2009
  );


  not
  g2166
  (
    n2248,
    n2119
  );


  buf
  g2167
  (
    n2202,
    n2002
  );


  not
  g2168
  (
    n2172,
    n2112
  );


  buf
  g2169
  (
    n2196,
    n2102
  );


  not
  g2170
  (
    n2137,
    n2011
  );


  not
  g2171
  (
    n2155,
    n2010
  );


  not
  g2172
  (
    n2247,
    n2123
  );


  not
  g2173
  (
    n2250,
    n1998
  );


  not
  g2174
  (
    n2157,
    n2096
  );


  not
  g2175
  (
    n2217,
    n2111
  );


  buf
  g2176
  (
    KeyWire_0_1,
    n2103
  );


  buf
  g2177
  (
    n2241,
    n2108
  );


  not
  g2178
  (
    n2131,
    n2104
  );


  not
  g2179
  (
    n2199,
    n2115
  );


  buf
  g2180
  (
    n2177,
    n2101
  );


  buf
  g2181
  (
    n2143,
    n1997
  );


  not
  g2182
  (
    n2221,
    n2123
  );


  not
  g2183
  (
    n2184,
    n2002
  );


  buf
  g2184
  (
    n2130,
    n2005
  );


  not
  g2185
  (
    n2127,
    n2096
  );


  buf
  g2186
  (
    n2146,
    n1997
  );


  not
  g2187
  (
    n2252,
    n2103
  );


  not
  g2188
  (
    n2193,
    n2108
  );


  buf
  g2189
  (
    n2151,
    n2121
  );


  not
  g2190
  (
    n2219,
    n1999
  );


  buf
  g2191
  (
    n2182,
    n2102
  );


  not
  g2192
  (
    n2239,
    n2101
  );


  not
  g2193
  (
    n2160,
    n2010
  );


  not
  g2194
  (
    n2165,
    n2000
  );


  or
  g2195
  (
    n2191,
    n1627,
    n2008,
    n2114,
    n2101
  );


  or
  g2196
  (
    n2150,
    n2122,
    n2108,
    n2095,
    n2113
  );


  xnor
  g2197
  (
    n2144,
    n2100,
    n2111,
    n2105,
    n2004
  );


  nor
  g2198
  (
    n2135,
    n2096,
    n2011,
    n2124,
    n2107
  );


  xnor
  g2199
  (
    n2188,
    n2097,
    n2109,
    n1621,
    n2105
  );


  nand
  g2200
  (
    n2173,
    n2097,
    n2110,
    n2011,
    n2003
  );


  xnor
  g2201
  (
    n2201,
    n1998,
    n1999,
    n2115
  );


  nor
  g2202
  (
    n2234,
    n2093,
    n2116,
    n2122,
    n2002
  );


  xor
  g2203
  (
    n2231,
    n2120,
    n2099,
    n2109,
    n2003
  );


  nand
  g2204
  (
    n2175,
    n2103,
    n2008,
    n1999,
    n2106
  );


  and
  g2205
  (
    n2215,
    n2009,
    n2114,
    n2007,
    n2093
  );


  nor
  g2206
  (
    n2245,
    n2012,
    n2122,
    n2103,
    n2098
  );


  nand
  g2207
  (
    n2226,
    n2116,
    n2110,
    n2102,
    n2008
  );


  and
  g2208
  (
    n2225,
    n1629,
    n1633,
    n1622,
    n2000
  );


  xnor
  g2209
  (
    n2232,
    n2012,
    n1631,
    n2095,
    n1998
  );


  nand
  g2210
  (
    n2179,
    n2094,
    n2010,
    n2009,
    n2012
  );


  xnor
  g2211
  (
    n2246,
    n2109,
    n1623,
    n2113,
    n2001
  );


  or
  g2212
  (
    n2133,
    n2117,
    n2120,
    n2105,
    n2124
  );


  nor
  g2213
  (
    n2190,
    n2121,
    n2004,
    n2114,
    n2002
  );


  or
  g2214
  (
    n2214,
    n2096,
    n2099,
    n2097,
    n1998
  );


  xor
  g2215
  (
    n2178,
    n2099,
    n1634,
    n2098,
    n2118
  );


  nand
  g2216
  (
    n2158,
    n1626,
    n2011,
    n2101,
    n2117
  );


  nor
  g2217
  (
    n2212,
    n2005,
    n2111,
    n2108,
    n2116
  );


  nor
  g2218
  (
    n2200,
    n1999,
    n2118,
    n2010,
    n2123
  );


  and
  g2219
  (
    n2206,
    n2117,
    n2007,
    n2105,
    n2112
  );


  buf
  g2220
  (
    n2293,
    n2252
  );


  buf
  g2221
  (
    n2609,
    n2211
  );


  buf
  g2222
  (
    n2585,
    n1640
  );


  buf
  g2223
  (
    n2467,
    n2235
  );


  buf
  g2224
  (
    n2262,
    n2135
  );


  not
  g2225
  (
    n2740,
    n2231
  );


  buf
  g2226
  (
    n2438,
    n2171
  );


  not
  g2227
  (
    n2679,
    n2222
  );


  buf
  g2228
  (
    n2541,
    n2172
  );


  not
  g2229
  (
    n2457,
    n2157
  );


  not
  g2230
  (
    n2633,
    n2228
  );


  buf
  g2231
  (
    n2329,
    n2169
  );


  not
  g2232
  (
    n2295,
    n2142
  );


  not
  g2233
  (
    n2628,
    n2215
  );


  not
  g2234
  (
    n2462,
    n2199
  );


  not
  g2235
  (
    n2713,
    n2125
  );


  not
  g2236
  (
    n2602,
    n2239
  );


  buf
  g2237
  (
    n2537,
    n2180
  );


  buf
  g2238
  (
    n2607,
    n2242
  );


  not
  g2239
  (
    n2440,
    n2131
  );


  buf
  g2240
  (
    n2398,
    n2252
  );


  buf
  g2241
  (
    n2664,
    n2221
  );


  not
  g2242
  (
    n2512,
    n2190
  );


  buf
  g2243
  (
    n2568,
    n2239
  );


  buf
  g2244
  (
    n2556,
    n1649
  );


  buf
  g2245
  (
    n2708,
    n2174
  );


  buf
  g2246
  (
    n2463,
    n2238
  );


  not
  g2247
  (
    n2487,
    n2198
  );


  not
  g2248
  (
    n2582,
    n2189
  );


  buf
  g2249
  (
    n2753,
    n2159
  );


  not
  g2250
  (
    n2322,
    n2216
  );


  not
  g2251
  (
    n2751,
    n2224
  );


  buf
  g2252
  (
    n2533,
    n2238
  );


  buf
  g2253
  (
    n2428,
    n2153
  );


  not
  g2254
  (
    n2334,
    n2147
  );


  buf
  g2255
  (
    n2673,
    n2150
  );


  not
  g2256
  (
    n2763,
    n2148
  );


  not
  g2257
  (
    n2565,
    n2171
  );


  buf
  g2258
  (
    n2307,
    n2151
  );


  buf
  g2259
  (
    n2729,
    n1647
  );


  buf
  g2260
  (
    n2693,
    n2152
  );


  buf
  g2261
  (
    n2577,
    n2214
  );


  buf
  g2262
  (
    n2518,
    n1635
  );


  buf
  g2263
  (
    n2504,
    n2161
  );


  buf
  g2264
  (
    n2759,
    n2132
  );


  not
  g2265
  (
    n2430,
    n2127
  );


  buf
  g2266
  (
    n2553,
    n1644
  );


  buf
  g2267
  (
    n2682,
    n2235
  );


  buf
  g2268
  (
    n2285,
    n2185
  );


  not
  g2269
  (
    n2323,
    n2128
  );


  buf
  g2270
  (
    n2555,
    n2178
  );


  not
  g2271
  (
    n2516,
    n2219
  );


  buf
  g2272
  (
    n2371,
    n2145
  );


  buf
  g2273
  (
    n2671,
    n2183
  );


  buf
  g2274
  (
    n2324,
    n2204
  );


  not
  g2275
  (
    n2275,
    n2212
  );


  buf
  g2276
  (
    n2596,
    n2195
  );


  buf
  g2277
  (
    n2492,
    n2220
  );


  buf
  g2278
  (
    n2279,
    n2201
  );


  buf
  g2279
  (
    n2717,
    n2190
  );


  buf
  g2280
  (
    n2645,
    n2154
  );


  not
  g2281
  (
    n2380,
    n2167
  );


  buf
  g2282
  (
    n2444,
    n2154
  );


  not
  g2283
  (
    n2394,
    n2182
  );


  buf
  g2284
  (
    n2372,
    n2251
  );


  buf
  g2285
  (
    n2375,
    n2177
  );


  not
  g2286
  (
    n2571,
    n2247
  );


  not
  g2287
  (
    n2574,
    n2190
  );


  buf
  g2288
  (
    n2485,
    n2168
  );


  buf
  g2289
  (
    n2406,
    n2186
  );


  buf
  g2290
  (
    n2362,
    n2211
  );


  buf
  g2291
  (
    n2344,
    n2242
  );


  not
  g2292
  (
    n2413,
    n2206
  );


  not
  g2293
  (
    n2545,
    n2178
  );


  not
  g2294
  (
    n2655,
    n2219
  );


  buf
  g2295
  (
    n2578,
    n2155
  );


  buf
  g2296
  (
    n2643,
    n2169
  );


  buf
  g2297
  (
    n2525,
    n2181
  );


  buf
  g2298
  (
    n2477,
    n2225
  );


  not
  g2299
  (
    n2583,
    n2217
  );


  not
  g2300
  (
    n2675,
    n2208
  );


  buf
  g2301
  (
    n2297,
    n2138
  );


  not
  g2302
  (
    n2374,
    n2208
  );


  not
  g2303
  (
    n2738,
    n2184
  );


  buf
  g2304
  (
    n2662,
    n2182
  );


  buf
  g2305
  (
    n2426,
    n2125
  );


  buf
  g2306
  (
    n2456,
    n1638
  );


  not
  g2307
  (
    n2657,
    n2225
  );


  not
  g2308
  (
    n2700,
    n2195
  );


  not
  g2309
  (
    n2598,
    n2144
  );


  buf
  g2310
  (
    n2678,
    n2219
  );


  buf
  g2311
  (
    n2706,
    n2163
  );


  not
  g2312
  (
    n2734,
    n2241
  );


  buf
  g2313
  (
    n2475,
    n2131
  );


  buf
  g2314
  (
    n2563,
    n2187
  );


  buf
  g2315
  (
    n2658,
    n1639
  );


  not
  g2316
  (
    n2442,
    n2126
  );


  not
  g2317
  (
    n2466,
    n2247
  );


  not
  g2318
  (
    n2646,
    n2202
  );


  buf
  g2319
  (
    n2317,
    n2237
  );


  not
  g2320
  (
    n2315,
    n2245
  );


  not
  g2321
  (
    n2336,
    n2158
  );


  buf
  g2322
  (
    n2617,
    n2248
  );


  buf
  g2323
  (
    n2507,
    n2200
  );


  not
  g2324
  (
    n2411,
    n2156
  );


  not
  g2325
  (
    n2669,
    n2186
  );


  not
  g2326
  (
    n2592,
    n2164
  );


  not
  g2327
  (
    n2291,
    n2196
  );


  not
  g2328
  (
    n2625,
    n2137
  );


  not
  g2329
  (
    n2342,
    n2230
  );


  not
  g2330
  (
    n2381,
    n2153
  );


  buf
  g2331
  (
    n2539,
    n2252
  );


  buf
  g2332
  (
    n2757,
    n2207
  );


  not
  g2333
  (
    n2668,
    n2209
  );


  not
  g2334
  (
    n2520,
    n2132
  );


  buf
  g2335
  (
    n2735,
    n2134
  );


  buf
  g2336
  (
    n2292,
    n2181
  );


  buf
  g2337
  (
    n2366,
    n2160
  );


  not
  g2338
  (
    n2500,
    n2185
  );


  not
  g2339
  (
    n2273,
    n2133
  );


  buf
  g2340
  (
    n2640,
    n2173
  );


  buf
  g2341
  (
    n2459,
    n2203
  );


  buf
  g2342
  (
    n2441,
    n2144
  );


  not
  g2343
  (
    n2272,
    n2219
  );


  buf
  g2344
  (
    n2259,
    n2188
  );


  not
  g2345
  (
    n2427,
    n2187
  );


  buf
  g2346
  (
    n2491,
    n2207
  );


  buf
  g2347
  (
    n2328,
    n2204
  );


  not
  g2348
  (
    n2732,
    n2136
  );


  not
  g2349
  (
    n2690,
    n2239
  );


  not
  g2350
  (
    n2761,
    n2136
  );


  buf
  g2351
  (
    n2730,
    n2161
  );


  not
  g2352
  (
    n2672,
    n2227
  );


  buf
  g2353
  (
    n2719,
    n2175
  );


  buf
  g2354
  (
    n2281,
    n2217
  );


  buf
  g2355
  (
    n2451,
    n2226
  );


  not
  g2356
  (
    n2268,
    n2146
  );


  not
  g2357
  (
    n2499,
    n2167
  );


  not
  g2358
  (
    n2649,
    n2197
  );


  buf
  g2359
  (
    n2721,
    n2179
  );


  buf
  g2360
  (
    n2595,
    n2240
  );


  not
  g2361
  (
    n2439,
    n2200
  );


  buf
  g2362
  (
    n2599,
    n2196
  );


  not
  g2363
  (
    n2663,
    n2138
  );


  not
  g2364
  (
    n2471,
    n2176
  );


  buf
  g2365
  (
    n2405,
    n2192
  );


  not
  g2366
  (
    n2755,
    n2168
  );


  not
  g2367
  (
    n2589,
    n2142
  );


  buf
  g2368
  (
    n2635,
    n2145
  );


  not
  g2369
  (
    n2529,
    n2226
  );


  not
  g2370
  (
    n2603,
    n2140
  );


  not
  g2371
  (
    n2530,
    n2141
  );


  buf
  g2372
  (
    n2497,
    n2172
  );


  buf
  g2373
  (
    n2739,
    n2222
  );


  not
  g2374
  (
    n2483,
    n2143
  );


  buf
  g2375
  (
    n2549,
    n2178
  );


  not
  g2376
  (
    n2579,
    n2134
  );


  buf
  g2377
  (
    n2376,
    n2244
  );


  buf
  g2378
  (
    n2552,
    n2251
  );


  not
  g2379
  (
    n2289,
    n2243
  );


  not
  g2380
  (
    n2567,
    n2176
  );


  buf
  g2381
  (
    n2685,
    n2188
  );


  buf
  g2382
  (
    n2660,
    n2213
  );


  buf
  g2383
  (
    n2514,
    n2236
  );


  not
  g2384
  (
    n2384,
    n2231
  );


  not
  g2385
  (
    n2355,
    n2130
  );


  buf
  g2386
  (
    n2697,
    n2177
  );


  buf
  g2387
  (
    n2652,
    n2158
  );


  buf
  g2388
  (
    n2495,
    n2135
  );


  not
  g2389
  (
    n2415,
    n2249
  );


  not
  g2390
  (
    n2310,
    n2175
  );


  buf
  g2391
  (
    n2526,
    n2169
  );


  buf
  g2392
  (
    n2330,
    n2229
  );


  buf
  g2393
  (
    n2647,
    n2164
  );


  not
  g2394
  (
    n2350,
    n2149
  );


  not
  g2395
  (
    n2496,
    n2133
  );


  not
  g2396
  (
    n2443,
    n2214
  );


  not
  g2397
  (
    n2365,
    n2198
  );


  buf
  g2398
  (
    n2546,
    n2207
  );


  buf
  g2399
  (
    n2624,
    n1960
  );


  buf
  g2400
  (
    n2290,
    n1961
  );


  not
  g2401
  (
    n2667,
    n2248
  );


  buf
  g2402
  (
    n2488,
    n2199
  );


  buf
  g2403
  (
    n2432,
    n2129
  );


  buf
  g2404
  (
    n2725,
    n2131
  );


  not
  g2405
  (
    n2403,
    n2238
  );


  buf
  g2406
  (
    n2691,
    n2230
  );


  buf
  g2407
  (
    n2360,
    n2183
  );


  not
  g2408
  (
    n2666,
    n2242
  );


  buf
  g2409
  (
    n2511,
    n2160
  );


  buf
  g2410
  (
    n2524,
    n2154
  );


  buf
  g2411
  (
    n2267,
    n2167
  );


  buf
  g2412
  (
    n2299,
    n2146
  );


  not
  g2413
  (
    n2611,
    n2163
  );


  buf
  g2414
  (
    n2348,
    n1653
  );


  buf
  g2415
  (
    n2745,
    n2150
  );


  not
  g2416
  (
    n2543,
    n2173
  );


  buf
  g2417
  (
    n2561,
    n2232
  );


  buf
  g2418
  (
    n2733,
    n1652
  );


  not
  g2419
  (
    n2622,
    n2233
  );


  buf
  g2420
  (
    n2493,
    n2216
  );


  not
  g2421
  (
    n2593,
    n2223
  );


  not
  g2422
  (
    n2631,
    n2127
  );


  buf
  g2423
  (
    n2349,
    n2203
  );


  not
  g2424
  (
    n2490,
    n2201
  );


  buf
  g2425
  (
    n2363,
    n2146
  );


  not
  g2426
  (
    n2659,
    n2193
  );


  buf
  g2427
  (
    n2620,
    n2209
  );


  not
  g2428
  (
    n2276,
    n2222
  );


  buf
  g2429
  (
    n2287,
    n2208
  );


  not
  g2430
  (
    n2606,
    n2162
  );


  buf
  g2431
  (
    n2385,
    n2179
  );


  not
  g2432
  (
    n2446,
    n2174
  );


  buf
  g2433
  (
    n2338,
    n2232
  );


  not
  g2434
  (
    n2562,
    n2195
  );


  not
  g2435
  (
    n2709,
    n2194
  );


  buf
  g2436
  (
    n2308,
    n1650
  );


  not
  g2437
  (
    n2551,
    n2223
  );


  buf
  g2438
  (
    n2354,
    n2225
  );


  buf
  g2439
  (
    n2627,
    n2139
  );


  not
  g2440
  (
    n2752,
    n2179
  );


  not
  g2441
  (
    n2754,
    n2210
  );


  not
  g2442
  (
    n2277,
    n2227
  );


  not
  g2443
  (
    n2351,
    n2212
  );


  buf
  g2444
  (
    n2470,
    n2200
  );


  buf
  g2445
  (
    n2610,
    n1637
  );


  buf
  g2446
  (
    n2736,
    n2246
  );


  not
  g2447
  (
    n2332,
    n2237
  );


  buf
  g2448
  (
    n2472,
    n2204
  );


  not
  g2449
  (
    n2455,
    n2126
  );


  not
  g2450
  (
    n2409,
    n2216
  );


  not
  g2451
  (
    n2465,
    n1648
  );


  not
  g2452
  (
    n2296,
    n2135
  );


  not
  g2453
  (
    n2361,
    n2224
  );


  buf
  g2454
  (
    n2270,
    n2173
  );


  not
  g2455
  (
    n2648,
    n2147
  );


  not
  g2456
  (
    n2588,
    n2231
  );


  not
  g2457
  (
    n2261,
    n2132
  );


  not
  g2458
  (
    n2639,
    n2206
  );


  not
  g2459
  (
    n2377,
    n2137
  );


  buf
  g2460
  (
    n2764,
    n2248
  );


  not
  g2461
  (
    n2305,
    n2180
  );


  buf
  g2462
  (
    n2744,
    n2144
  );


  not
  g2463
  (
    n2353,
    n2190
  );


  buf
  g2464
  (
    n2557,
    n2180
  );


  not
  g2465
  (
    n2653,
    n2199
  );


  not
  g2466
  (
    n2309,
    n1642
  );


  buf
  g2467
  (
    n2417,
    n2247
  );


  not
  g2468
  (
    n2570,
    n2222
  );


  buf
  g2469
  (
    n2656,
    n2193
  );


  not
  g2470
  (
    n2550,
    n2192
  );


  buf
  g2471
  (
    n2630,
    n2125
  );


  buf
  g2472
  (
    n2325,
    n2168
  );


  not
  g2473
  (
    n2758,
    n2170
  );


  buf
  g2474
  (
    n2703,
    n2211
  );


  buf
  g2475
  (
    n2489,
    n2142
  );


  not
  g2476
  (
    n2688,
    n2249
  );


  buf
  g2477
  (
    n2498,
    n2235
  );


  not
  g2478
  (
    n2601,
    n2225
  );


  not
  g2479
  (
    n2367,
    n2217
  );


  not
  g2480
  (
    n2704,
    n2139
  );


  not
  g2481
  (
    n2674,
    n2193
  );


  buf
  g2482
  (
    n2312,
    n1636
  );


  not
  g2483
  (
    n2683,
    n2128
  );


  not
  g2484
  (
    n2760,
    n2237
  );


  buf
  g2485
  (
    n2743,
    n2078
  );


  not
  g2486
  (
    n2711,
    n2167
  );


  not
  g2487
  (
    n2425,
    n2230
  );


  not
  g2488
  (
    n2343,
    n2160
  );


  not
  g2489
  (
    n2536,
    n2198
  );


  not
  g2490
  (
    n2254,
    n2201
  );


  buf
  g2491
  (
    n2587,
    n2205
  );


  not
  g2492
  (
    n2386,
    n2245
  );


  not
  g2493
  (
    n2522,
    n2174
  );


  not
  g2494
  (
    n2638,
    n2234
  );


  not
  g2495
  (
    n2686,
    n2218
  );


  buf
  g2496
  (
    n2508,
    n2166
  );


  not
  g2497
  (
    n2301,
    n2159
  );


  not
  g2498
  (
    n2597,
    n2184
  );


  buf
  g2499
  (
    n2347,
    n2130
  );


  not
  g2500
  (
    n2604,
    n2180
  );


  buf
  g2501
  (
    n2715,
    n2165
  );


  not
  g2502
  (
    n2723,
    n2221
  );


  not
  g2503
  (
    n2445,
    n2183
  );


  buf
  g2504
  (
    n2707,
    n2191
  );


  buf
  g2505
  (
    n2594,
    n2209
  );


  buf
  g2506
  (
    n2756,
    n2191
  );


  buf
  g2507
  (
    n2559,
    n2155
  );


  buf
  g2508
  (
    n2554,
    n2242
  );


  buf
  g2509
  (
    n2728,
    n2031
  );


  not
  g2510
  (
    n2605,
    n2187
  );


  not
  g2511
  (
    n2357,
    n2228
  );


  buf
  g2512
  (
    n2534,
    n2162
  );


  not
  g2513
  (
    n2373,
    n2184
  );


  not
  g2514
  (
    n2505,
    n2178
  );


  not
  g2515
  (
    n2564,
    n2156
  );


  buf
  g2516
  (
    n2590,
    n2129
  );


  buf
  g2517
  (
    n2431,
    n2215
  );


  buf
  g2518
  (
    n2651,
    n2128
  );


  not
  g2519
  (
    n2341,
    n2189
  );


  not
  g2520
  (
    n2661,
    n2226
  );


  buf
  g2521
  (
    n2421,
    n2187
  );


  buf
  g2522
  (
    n2391,
    n2169
  );


  not
  g2523
  (
    n2288,
    n2192
  );


  buf
  g2524
  (
    n2412,
    n2159
  );


  not
  g2525
  (
    n2448,
    n2133
  );


  not
  g2526
  (
    n2701,
    n2246
  );


  not
  g2527
  (
    n2320,
    n2194
  );


  buf
  g2528
  (
    n2665,
    n2127
  );


  buf
  g2529
  (
    n2687,
    n2241
  );


  not
  g2530
  (
    n2473,
    n2241
  );


  not
  g2531
  (
    n2644,
    n2170
  );


  buf
  g2532
  (
    n2558,
    n2250
  );


  buf
  g2533
  (
    n2454,
    n2217
  );


  buf
  g2534
  (
    n2684,
    n2234
  );


  buf
  g2535
  (
    n2304,
    n2230
  );


  not
  g2536
  (
    n2702,
    n2185
  );


  not
  g2537
  (
    n2540,
    n2143
  );


  buf
  g2538
  (
    n2548,
    n2162
  );


  buf
  g2539
  (
    n2333,
    n2149
  );


  not
  g2540
  (
    n2718,
    n2172
  );


  buf
  g2541
  (
    n2510,
    n2153
  );


  buf
  g2542
  (
    n2544,
    n2149
  );


  buf
  g2543
  (
    n2314,
    n2240
  );


  not
  g2544
  (
    n2460,
    n2129
  );


  buf
  g2545
  (
    n2437,
    n2125
  );


  buf
  g2546
  (
    n2689,
    n2188
  );


  buf
  g2547
  (
    n2313,
    n2228
  );


  not
  g2548
  (
    n2318,
    n2145
  );


  buf
  g2549
  (
    n2694,
    n2158
  );


  buf
  g2550
  (
    n2748,
    n2227
  );


  not
  g2551
  (
    n2284,
    n2143
  );


  not
  g2552
  (
    n2634,
    n2182
  );


  buf
  g2553
  (
    n2591,
    n2149
  );


  buf
  g2554
  (
    n2345,
    n2189
  );


  not
  g2555
  (
    n2632,
    n2143
  );


  not
  g2556
  (
    n2629,
    n2241
  );


  not
  g2557
  (
    n2265,
    n2232
  );


  not
  g2558
  (
    n2538,
    n2224
  );


  not
  g2559
  (
    n2294,
    n2236
  );


  buf
  g2560
  (
    n2464,
    n2144
  );


  not
  g2561
  (
    n2714,
    n2234
  );


  not
  g2562
  (
    n2419,
    n2155
  );


  buf
  g2563
  (
    n2390,
    n2132
  );


  buf
  g2564
  (
    n2468,
    n2231
  );


  buf
  g2565
  (
    n2263,
    n2135
  );


  not
  g2566
  (
    n2346,
    n2165
  );


  not
  g2567
  (
    n2452,
    n2151
  );


  buf
  g2568
  (
    n2614,
    n2218
  );


  not
  g2569
  (
    n2527,
    n2137
  );


  buf
  g2570
  (
    n2306,
    n2240
  );


  buf
  g2571
  (
    n2741,
    n2168
  );


  buf
  g2572
  (
    n2260,
    n2155
  );


  not
  g2573
  (
    n2316,
    n2204
  );


  buf
  g2574
  (
    KeyWire_0_10,
    n2197
  );


  buf
  g2575
  (
    n2303,
    n2234
  );


  not
  g2576
  (
    n2337,
    n2229
  );


  not
  g2577
  (
    n2257,
    n2154
  );


  buf
  g2578
  (
    n2712,
    n2166
  );


  not
  g2579
  (
    n2716,
    n2161
  );


  not
  g2580
  (
    n2408,
    n2246
  );


  not
  g2581
  (
    n2650,
    n2147
  );


  not
  g2582
  (
    n2681,
    n2131
  );


  not
  g2583
  (
    n2387,
    n2179
  );


  not
  g2584
  (
    n2358,
    n2211
  );


  buf
  g2585
  (
    n2388,
    n2233
  );


  buf
  g2586
  (
    n2392,
    n2248
  );


  buf
  g2587
  (
    n2531,
    n2141
  );


  not
  g2588
  (
    n2258,
    n2213
  );


  not
  g2589
  (
    n2420,
    n2150
  );


  not
  g2590
  (
    n2331,
    n2186
  );


  not
  g2591
  (
    n2429,
    n2243
  );


  buf
  g2592
  (
    n2560,
    n2129
  );


  buf
  g2593
  (
    n2502,
    n2140
  );


  not
  g2594
  (
    n2433,
    n2136
  );


  not
  g2595
  (
    n2699,
    n2185
  );


  buf
  g2596
  (
    n2282,
    n2148
  );


  not
  g2597
  (
    n2519,
    n2166
  );


  not
  g2598
  (
    n2696,
    n2176
  );


  buf
  g2599
  (
    n2423,
    n2184
  );


  not
  g2600
  (
    n2547,
    n2186
  );


  not
  g2601
  (
    n2750,
    n2152
  );


  buf
  g2602
  (
    n2621,
    n2250
  );


  buf
  g2603
  (
    n2422,
    n2205
  );


  not
  g2604
  (
    n2608,
    n2215
  );


  buf
  g2605
  (
    n2370,
    n2245
  );


  buf
  g2606
  (
    n2396,
    n2191
  );


  not
  g2607
  (
    n2399,
    n2172
  );


  buf
  g2608
  (
    n2737,
    n2151
  );


  not
  g2609
  (
    n2509,
    n2220
  );


  buf
  g2610
  (
    n2517,
    n2249
  );


  not
  g2611
  (
    n2436,
    n2165
  );


  not
  g2612
  (
    n2747,
    n2141
  );


  not
  g2613
  (
    n2654,
    n2173
  );


  not
  g2614
  (
    n2298,
    n2175
  );


  buf
  g2615
  (
    n2528,
    n2171
  );


  buf
  g2616
  (
    n2494,
    n2220
  );


  not
  g2617
  (
    n2383,
    n2212
  );


  not
  g2618
  (
    n2569,
    n2139
  );


  not
  g2619
  (
    n2615,
    n2193
  );


  buf
  g2620
  (
    n2724,
    n2197
  );


  not
  g2621
  (
    n2352,
    n2251
  );


  buf
  g2622
  (
    n2486,
    n2147
  );


  buf
  g2623
  (
    n2480,
    n2236
  );


  buf
  g2624
  (
    n2379,
    n2175
  );


  buf
  g2625
  (
    n2523,
    n2223
  );


  buf
  g2626
  (
    n2680,
    n2194
  );


  buf
  g2627
  (
    n2576,
    n2236
  );


  not
  g2628
  (
    n2584,
    n2249
  );


  not
  g2629
  (
    n2311,
    n2244
  );


  not
  g2630
  (
    n2676,
    n2181
  );


  buf
  g2631
  (
    n2636,
    n2215
  );


  not
  g2632
  (
    n2449,
    n2229
  );


  buf
  g2633
  (
    n2300,
    n2157
  );


  buf
  g2634
  (
    n2501,
    n2134
  );


  buf
  g2635
  (
    n2705,
    n2244
  );


  not
  g2636
  (
    n2255,
    n2164
  );


  not
  g2637
  (
    n2407,
    n2199
  );


  buf
  g2638
  (
    n2612,
    n2157
  );


  buf
  g2639
  (
    n2280,
    n2196
  );


  buf
  g2640
  (
    n2450,
    n2233
  );


  buf
  g2641
  (
    n2731,
    n2223
  );


  not
  g2642
  (
    n2484,
    n2201
  );


  buf
  g2643
  (
    n2359,
    n1651
  );


  buf
  g2644
  (
    n2469,
    n2163
  );


  not
  g2645
  (
    n2503,
    n2162
  );


  buf
  g2646
  (
    n2424,
    n2233
  );


  not
  g2647
  (
    n2478,
    n2128
  );


  not
  g2648
  (
    n2368,
    n2213
  );


  not
  g2649
  (
    n2397,
    n2192
  );


  buf
  g2650
  (
    n2695,
    n2239
  );


  buf
  g2651
  (
    n2521,
    n2127
  );


  not
  g2652
  (
    n2616,
    n2235
  );


  buf
  g2653
  (
    n2326,
    n2158
  );


  buf
  g2654
  (
    n2474,
    n2214
  );


  buf
  g2655
  (
    n2575,
    n2152
  );


  not
  g2656
  (
    n2572,
    n2198
  );


  buf
  g2657
  (
    n2573,
    n2134
  );


  buf
  g2658
  (
    n2410,
    n2237
  );


  not
  g2659
  (
    n2340,
    n2145
  );


  buf
  g2660
  (
    n2746,
    n2165
  );


  not
  g2661
  (
    n2482,
    n2140
  );


  not
  g2662
  (
    n2600,
    n2137
  );


  not
  g2663
  (
    n2580,
    n2170
  );


  buf
  g2664
  (
    n2586,
    n2191
  );


  not
  g2665
  (
    n2749,
    n2210
  );


  not
  g2666
  (
    n2461,
    n2157
  );


  buf
  g2667
  (
    n2335,
    n2142
  );


  buf
  g2668
  (
    n2641,
    n2163
  );


  buf
  g2669
  (
    n2269,
    n2166
  );


  buf
  g2670
  (
    n2286,
    n2243
  );


  buf
  g2671
  (
    n2619,
    n2221
  );


  buf
  g2672
  (
    n2476,
    n2139
  );


  buf
  g2673
  (
    n2513,
    n2251
  );


  not
  g2674
  (
    n2710,
    n2156
  );


  buf
  g2675
  (
    n2264,
    n2140
  );


  buf
  g2676
  (
    n2266,
    n2153
  );


  not
  g2677
  (
    n2481,
    n2194
  );


  not
  g2678
  (
    n2566,
    n2203
  );


  not
  g2679
  (
    n2637,
    n2210
  );


  not
  g2680
  (
    n2256,
    n2164
  );


  buf
  g2681
  (
    n2274,
    n2126
  );


  buf
  g2682
  (
    n2742,
    n2200
  );


  not
  g2683
  (
    n2623,
    n2203
  );


  not
  g2684
  (
    n2626,
    n2216
  );


  buf
  g2685
  (
    n2698,
    n2247
  );


  buf
  g2686
  (
    n2418,
    n2229
  );


  buf
  g2687
  (
    n2302,
    n2224
  );


  not
  g2688
  (
    n2479,
    n2250
  );


  not
  g2689
  (
    n2642,
    n2148
  );


  not
  g2690
  (
    n2720,
    n2156
  );


  not
  g2691
  (
    n2542,
    n1643
  );


  not
  g2692
  (
    n2762,
    n2141
  );


  buf
  g2693
  (
    n2692,
    n2171
  );


  not
  g2694
  (
    n2416,
    n2250
  );


  buf
  g2695
  (
    n2378,
    n2202
  );


  buf
  g2696
  (
    n2395,
    n2183
  );


  buf
  g2697
  (
    n2364,
    n2218
  );


  not
  g2698
  (
    n2581,
    n2148
  );


  buf
  g2699
  (
    n2453,
    n2195
  );


  buf
  g2700
  (
    n2458,
    n2160
  );


  not
  g2701
  (
    n2722,
    n2244
  );


  buf
  g2702
  (
    n2532,
    n2170
  );


  buf
  g2703
  (
    n2726,
    n2214
  );


  buf
  g2704
  (
    n2278,
    n2138
  );


  buf
  g2705
  (
    n2271,
    n1646
  );


  not
  g2706
  (
    n2434,
    n2151
  );


  not
  g2707
  (
    n2677,
    n2130
  );


  not
  g2708
  (
    n2339,
    n2138
  );


  not
  g2709
  (
    n2515,
    n2252
  );


  not
  g2710
  (
    n2414,
    n2182
  );


  not
  g2711
  (
    n2401,
    n2202
  );


  not
  g2712
  (
    n2400,
    n2221
  );


  buf
  g2713
  (
    n2613,
    n1645
  );


  not
  g2714
  (
    n2327,
    n2181
  );


  not
  g2715
  (
    n2535,
    n2243
  );


  buf
  g2716
  (
    n2321,
    n2177
  );


  not
  g2717
  (
    n2382,
    n2227
  );


  not
  g2718
  (
    n2404,
    n2159
  );


  not
  g2719
  (
    n2402,
    n2197
  );


  not
  g2720
  (
    n2253,
    n2189
  );


  not
  g2721
  (
    n2319,
    n2218
  );


  buf
  g2722
  (
    n2435,
    n2205
  );


  buf
  g2723
  (
    n2447,
    n1654
  );


  or
  g2724
  (
    n2356,
    n2209,
    n2161,
    n2176,
    n2212
  );


  and
  g2725
  (
    n2283,
    n2245,
    n2210,
    n2205,
    n2150
  );


  nor
  g2726
  (
    n2389,
    n2220,
    n2146,
    n2174,
    n2202
  );


  nand
  g2727
  (
    n2369,
    n2208,
    n2206,
    n2177,
    n2130
  );


  and
  g2728
  (
    n2393,
    n2240,
    n2226,
    n2246,
    n2213
  );


  xnor
  g2729
  (
    n2506,
    n2126,
    n2136,
    n2228,
    n2188
  );


  nor
  g2730
  (
    n2670,
    n2196,
    n1641,
    n2133,
    n2206
  );


  or
  g2731
  (
    n2618,
    n2152,
    n2232,
    n2207,
    n2238
  );


  nor
  g2732
  (
    n2859,
    n2582,
    n2546,
    n2627,
    n2559
  );


  and
  g2733
  (
    n2811,
    n2493,
    n2623,
    n2421,
    n2576
  );


  nor
  g2734
  (
    n2784,
    n2615,
    n2481,
    n2459,
    n2655
  );


  and
  g2735
  (
    n2840,
    n2379,
    n2403,
    n2463,
    n2609
  );


  or
  g2736
  (
    n2787,
    n2458,
    n2264,
    n2362,
    n2344
  );


  nand
  g2737
  (
    n2837,
    n2543,
    n2305,
    n2423,
    n2420
  );


  nor
  g2738
  (
    n2769,
    n2378,
    n2658,
    n2397,
    n2622
  );


  and
  g2739
  (
    n2819,
    n2331,
    n2439,
    n2614,
    n2485
  );


  or
  g2740
  (
    n2779,
    n2292,
    n2516,
    n2451,
    n2585
  );


  nor
  g2741
  (
    n2798,
    n2406,
    n2646,
    n2638,
    n2389
  );


  nor
  g2742
  (
    n2846,
    n2293,
    n2474,
    n2309,
    n2257
  );


  nor
  g2743
  (
    n2785,
    n2360,
    n2259,
    n2492,
    n2637
  );


  xnor
  g2744
  (
    n2813,
    n2284,
    n2444,
    n2280,
    n2351
  );


  nand
  g2745
  (
    n2847,
    n2395,
    n1656,
    n2364,
    n2412
  );


  and
  g2746
  (
    n2795,
    n2579,
    n2393,
    n2301,
    n2556
  );


  and
  g2747
  (
    n2807,
    n2290,
    n2618,
    n2594,
    n2617
  );


  xnor
  g2748
  (
    n2781,
    n2296,
    n2324,
    n2508,
    n2599
  );


  or
  g2749
  (
    n2841,
    n2447,
    n2565,
    n2587,
    n2619
  );


  xor
  g2750
  (
    n2780,
    n2430,
    n2448,
    n2503,
    n2457
  );


  nand
  g2751
  (
    n2831,
    n2521,
    n2610,
    n2352,
    n2367
  );


  nand
  g2752
  (
    n2860,
    n1655,
    n2538,
    n2537,
    n2648
  );


  xnor
  g2753
  (
    n2797,
    n2564,
    n2612,
    n2639,
    n2480
  );


  nor
  g2754
  (
    n2852,
    n2468,
    n2471,
    n2476,
    n2555
  );


  nor
  g2755
  (
    n2839,
    n2385,
    n2449,
    n2401,
    n2548
  );


  nor
  g2756
  (
    n2792,
    n2445,
    n2414,
    n2542,
    n2526
  );


  and
  g2757
  (
    n2803,
    n2495,
    n2308,
    n2349,
    n2632
  );


  or
  g2758
  (
    n2842,
    n2452,
    n2507,
    n2377,
    n2398
  );


  nand
  g2759
  (
    n2865,
    n2381,
    n2600,
    n2390,
    n2645
  );


  nor
  g2760
  (
    n2849,
    n2396,
    n2580,
    n2533,
    n2402
  );


  nor
  g2761
  (
    n2802,
    n2336,
    n2373,
    n2383,
    n2274
  );


  xnor
  g2762
  (
    n2825,
    n2473,
    n2583,
    n2434,
    n2314
  );


  nor
  g2763
  (
    n2818,
    n2568,
    n2653,
    n2591,
    n2654
  );


  nand
  g2764
  (
    n2790,
    n2604,
    n2354,
    n2269,
    n2392
  );


  nand
  g2765
  (
    n2799,
    n2484,
    n2522,
    n2291,
    n2608
  );


  xnor
  g2766
  (
    n2844,
    n2295,
    n2404,
    n2416,
    n2371
  );


  and
  g2767
  (
    n2776,
    n2338,
    n2577,
    n2483,
    n2299
  );


  xnor
  g2768
  (
    n2773,
    n2302,
    n2359,
    n2270,
    n2271
  );


  xor
  g2769
  (
    n2793,
    n2550,
    n2426,
    n2524,
    n2642
  );


  xor
  g2770
  (
    n2835,
    n2418,
    n2334,
    n2549,
    n2281
  );


  xor
  g2771
  (
    n2765,
    n2551,
    n2429,
    n2509,
    n2286
  );


  xnor
  g2772
  (
    n2854,
    n2656,
    n2268,
    n2438,
    n2643
  );


  nand
  g2773
  (
    n2855,
    n2333,
    n2254,
    n2282,
    n2456
  );


  xnor
  g2774
  (
    n2834,
    n2624,
    n2307,
    n2394,
    n2558
  );


  nor
  g2775
  (
    n2832,
    n2278,
    n2477,
    n2313,
    n2424
  );


  and
  g2776
  (
    n2794,
    n2479,
    n2365,
    n2650,
    n2342
  );


  or
  g2777
  (
    n2808,
    n2419,
    n2328,
    n2285,
    n2529
  );


  xor
  g2778
  (
    n2774,
    n2561,
    n2625,
    n2486,
    n2279
  );


  or
  g2779
  (
    n2827,
    n2415,
    n2356,
    n2567,
    n2320
  );


  nor
  g2780
  (
    n2806,
    n2540,
    n2647,
    n2649,
    n2417
  );


  xnor
  g2781
  (
    n2824,
    n2571,
    n2287,
    n2462,
    n2534
  );


  nor
  g2782
  (
    n2775,
    n2541,
    n2512,
    n2312,
    n2488
  );


  or
  g2783
  (
    n2848,
    n2425,
    n2482,
    n2363,
    n2531
  );


  nand
  g2784
  (
    n2843,
    n2528,
    n2496,
    n2464,
    n2358
  );


  xor
  g2785
  (
    n2815,
    n2437,
    n2337,
    n2640,
    n2586
  );


  xor
  g2786
  (
    n2856,
    n2311,
    n2554,
    n2317,
    n2478
  );


  or
  g2787
  (
    n2820,
    n2511,
    n2409,
    n2602,
    n2345
  );


  xor
  g2788
  (
    n2853,
    n2323,
    n2316,
    n2440,
    n2380
  );


  and
  g2789
  (
    n2845,
    n2273,
    n2500,
    n2575,
    n2369
  );


  nand
  g2790
  (
    n2783,
    n2494,
    n2466,
    n2453,
    n2319
  );


  nor
  g2791
  (
    n2777,
    n2501,
    n2350,
    n2498,
    n2408
  );


  xnor
  g2792
  (
    n2823,
    n2450,
    n2298,
    n2353,
    n2589
  );


  nand
  g2793
  (
    n2801,
    n2515,
    n2569,
    n2326,
    n2261
  );


  and
  g2794
  (
    n2778,
    n2297,
    n2304,
    n2256,
    n2562
  );


  or
  g2795
  (
    n2858,
    n2346,
    n2399,
    n2283,
    n2634
  );


  xnor
  g2796
  (
    n2830,
    n2597,
    n2518,
    n2581,
    n2321
  );


  xor
  g2797
  (
    n2833,
    n2441,
    n2276,
    n2631,
    n2388
  );


  and
  g2798
  (
    n2791,
    n2446,
    n2536,
    n2387,
    n2327
  );


  nand
  g2799
  (
    n2862,
    n2407,
    n2595,
    n2405,
    n2596
  );


  and
  g2800
  (
    n2817,
    n2348,
    n2303,
    n2384,
    n2400
  );


  nor
  g2801
  (
    n2826,
    n2544,
    n2578,
    n2598,
    n2435
  );


  and
  g2802
  (
    n2767,
    n2374,
    n2588,
    n2294,
    n2530
  );


  and
  g2803
  (
    n2800,
    n2563,
    n2330,
    n2566,
    n2487
  );


  and
  g2804
  (
    n2828,
    n2436,
    n2545,
    n2465,
    n2603
  );


  and
  g2805
  (
    n2809,
    n2490,
    n2620,
    n2635,
    n2611
  );


  and
  g2806
  (
    n2782,
    n2343,
    n2584,
    n2266,
    n2499
  );


  nand
  g2807
  (
    n2770,
    n2657,
    n2329,
    n2652,
    n2527
  );


  nor
  g2808
  (
    n2796,
    n2422,
    n2376,
    n2318,
    n2306
  );


  nor
  g2809
  (
    n2857,
    n2491,
    n2552,
    n2590,
    n2535
  );


  xnor
  g2810
  (
    KeyWire_0_13,
    n2570,
    n2489,
    n2633,
    n2300
  );


  nand
  g2811
  (
    n2864,
    n2475,
    n2253,
    n2255,
    n2454
  );


  or
  g2812
  (
    n2822,
    n2593,
    n2411,
    n2413,
    n2267
  );


  xor
  g2813
  (
    n2821,
    n2428,
    n2340,
    n2601,
    n2628
  );


  xnor
  g2814
  (
    n2861,
    n2382,
    n2460,
    n2510,
    n2505
  );


  and
  g2815
  (
    n2788,
    n2520,
    n2467,
    n2347,
    n2514
  );


  nand
  g2816
  (
    n2829,
    n2277,
    n2557,
    n2572,
    n2525
  );


  xor
  g2817
  (
    n2814,
    n2262,
    n2339,
    n2539,
    n2472
  );


  nand
  g2818
  (
    n2851,
    n2432,
    n2470,
    n2497,
    n2626
  );


  and
  g2819
  (
    n2786,
    n2433,
    n2272,
    n2651,
    n2532
  );


  nand
  g2820
  (
    n2850,
    n2605,
    n2370,
    n2455,
    n2355
  );


  xnor
  g2821
  (
    n2816,
    n2506,
    n2613,
    n2513,
    n2386
  );


  nand
  g2822
  (
    n2866,
    n2265,
    n2519,
    n2621,
    n2517
  );


  nand
  g2823
  (
    n2771,
    n2372,
    n2641,
    n2275,
    n2547
  );


  nor
  g2824
  (
    n2789,
    n2431,
    n2616,
    n2325,
    n2361
  );


  or
  g2825
  (
    n2838,
    n2553,
    n2410,
    n2442,
    n2502
  );


  xnor
  g2826
  (
    n2772,
    n2560,
    n2258,
    n2289,
    n2375
  );


  nand
  g2827
  (
    n2768,
    n2263,
    n2629,
    n2574,
    n2644
  );


  and
  g2828
  (
    n2804,
    n2592,
    n2573,
    n2391,
    n2504
  );


  and
  g2829
  (
    n2812,
    n2443,
    n2461,
    n2523,
    n2335
  );


  and
  g2830
  (
    n2810,
    n2332,
    n2630,
    n2636,
    n2288
  );


  nor
  g2831
  (
    n2863,
    n2322,
    n2366,
    n2427,
    n2368
  );


  or
  g2832
  (
    n2836,
    n2607,
    n2315,
    n2357,
    n2469
  );


  nor
  g2833
  (
    n2766,
    n2341,
    n2310,
    n2606,
    n2260
  );


  buf
  g2834
  (
    n2867,
    n2768
  );


  buf
  g2835
  (
    n2870,
    n2765
  );


  buf
  g2836
  (
    n2869,
    n2767
  );


  not
  g2837
  (
    n2868,
    n2766
  );


  and
  g2838
  (
    n2872,
    n2867,
    n2772,
    n2771,
    n2868
  );


  nand
  g2839
  (
    n2871,
    n2773,
    n2774,
    n2770,
    n2769
  );


  xor
  g2840
  (
    n2875,
    n1969,
    n1964,
    n1970,
    n1967
  );


  xor
  g2841
  (
    n2873,
    n2872,
    n2872,
    n1971,
    n1966
  );


  xnor
  g2842
  (
    n2874,
    n1973,
    n1965,
    n1968,
    n2871
  );


  and
  g2843
  (
    n2876,
    n1972,
    n1962,
    n1963,
    n2872
  );


  or
  g2844
  (
    n2878,
    n2777,
    n2780,
    n2778,
    n2775
  );


  nor
  g2845
  (
    n2877,
    n2779,
    n2874,
    n2776,
    n2873
  );


  buf
  g2846
  (
    n2882,
    n2878
  );


  buf
  g2847
  (
    n2883,
    n2878
  );


  not
  g2848
  (
    n2879,
    n2877
  );


  not
  g2849
  (
    n2880,
    n2878
  );


  not
  g2850
  (
    n2881,
    n2878
  );


  and
  g2851
  (
    n2884,
    n2783,
    n2879,
    n2781,
    n2784
  );


  and
  g2852
  (
    n2885,
    n2782,
    n2880,
    n2879
  );


  buf
  g2853
  (
    n2887,
    n2884
  );


  buf
  g2854
  (
    n2890,
    n2885
  );


  buf
  g2855
  (
    n2886,
    n2885
  );


  not
  g2856
  (
    n2889,
    n2885
  );


  buf
  g2857
  (
    n2888,
    n2885
  );


  xnor
  g2858
  (
    n2893,
    n1974,
    n2876,
    n2880
  );


  xor
  g2859
  (
    n2894,
    n2789,
    n2876,
    n2889,
    n2870
  );


  nor
  g2860
  (
    n2892,
    n2790,
    n2887,
    n2875,
    n2876
  );


  and
  g2861
  (
    n2891,
    n2890,
    n2787,
    n2788,
    n2875
  );


  or
  g2862
  (
    n2896,
    n2791,
    n2890,
    n2886,
    n2875
  );


  xnor
  g2863
  (
    n2897,
    n2785,
    n2786,
    n1657,
    n2888
  );


  or
  g2864
  (
    n2895,
    n1975,
    n2022,
    n2869,
    n2890
  );


  buf
  g2865
  (
    n2899,
    n2897
  );


  buf
  g2866
  (
    n2900,
    n2895
  );


  not
  g2867
  (
    n2898,
    n2896
  );


  nand
  g2868
  (
    n2901,
    n2898,
    n2881
  );


  xor
  g2869
  (
    n2902,
    n2898,
    n2881
  );


  not
  g2870
  (
    n2903,
    n2882
  );


  nor
  g2871
  (
    n2905,
    n2901,
    n2902
  );


  xor
  g2872
  (
    n2904,
    n2902,
    n2882
  );


  xor
  g2873
  (
    n2906,
    n2882,
    n2883,
    n2903
  );


  nor
  g2874
  (
    n2908,
    n1976,
    n2012,
    n2906,
    n2904
  );


  xnor
  g2875
  (
    n2907,
    n2792,
    n2794,
    n2906,
    n2793
  );


  buf
  g2876
  (
    n2910,
    n2907
  );


  not
  g2877
  (
    n2912,
    n2908
  );


  buf
  g2878
  (
    n2914,
    n2908
  );


  not
  g2879
  (
    n2913,
    n2907
  );


  buf
  g2880
  (
    n2911,
    n2908
  );


  buf
  g2881
  (
    n2909,
    n2907
  );


  and
  g2882
  (
    n2921,
    n2851,
    n2821,
    n2799,
    n2863
  );


  nand
  g2883
  (
    n2938,
    n2801,
    n2910,
    n2912,
    n2914
  );


  nand
  g2884
  (
    n2920,
    n2803,
    n2808,
    n2822,
    n2814
  );


  xor
  g2885
  (
    n2934,
    n2910,
    n2857,
    n2842,
    n2862
  );


  or
  g2886
  (
    n2930,
    n2834,
    n2861,
    n2815,
    n2913
  );


  or
  g2887
  (
    n2927,
    n2795,
    n2859,
    n2911,
    n2852
  );


  nor
  g2888
  (
    n2928,
    n2860,
    n2865,
    n2817,
    n2810
  );


  and
  g2889
  (
    n2922,
    n2853,
    n2829,
    n2839,
    n2844
  );


  xor
  g2890
  (
    n2929,
    n2830,
    n2824,
    n2912,
    n2827
  );


  nor
  g2891
  (
    n2926,
    n2909,
    n2909,
    n2864,
    n2914
  );


  xor
  g2892
  (
    n2936,
    n2838,
    n2910,
    n2911,
    n2800
  );


  nor
  g2893
  (
    n2937,
    n2804,
    n2812,
    n2825,
    n2858
  );


  or
  g2894
  (
    n2923,
    n2832,
    n2866,
    n2913,
    n2914
  );


  and
  g2895
  (
    n2918,
    n2835,
    n2909,
    n2912,
    n2850
  );


  nor
  g2896
  (
    n2925,
    n2798,
    n2854,
    n2813,
    n2855
  );


  xor
  g2897
  (
    n2915,
    n2805,
    n2909,
    n2912,
    n2797
  );


  xor
  g2898
  (
    n2917,
    n2833,
    n2837,
    n2826,
    n2845
  );


  and
  g2899
  (
    n2932,
    n2843,
    n2913,
    n2914,
    n2911
  );


  nand
  g2900
  (
    n2931,
    n2809,
    n2823,
    n2811,
    n2818
  );


  nand
  g2901
  (
    n2933,
    n2807,
    n2841,
    n2848,
    n2816
  );


  xor
  g2902
  (
    n2919,
    n2911,
    n2840,
    n2849,
    n2836
  );


  nor
  g2903
  (
    n2924,
    n2846,
    n2831,
    n2828,
    n2796
  );


  xnor
  g2904
  (
    n2916,
    n2802,
    n2913,
    n2820,
    n2856
  );


  or
  g2905
  (
    n2935,
    n2819,
    n2806,
    n2847,
    n2910
  );


  nor
  g2906
  (
    n2952,
    n1755,
    n2713,
    n2930,
    n2933
  );


  or
  g2907
  (
    n3005,
    n1733,
    n2934,
    n2746,
    n1705
  );


  nor
  g2908
  (
    n2998,
    n2900,
    n2701,
    n2932,
    n2754
  );


  xnor
  g2909
  (
    n2975,
    n2937,
    n2900,
    n2740,
    n1692
  );


  xnor
  g2910
  (
    n2988,
    n1669,
    n1710,
    n1753,
    n1673
  );


  nor
  g2911
  (
    n2953,
    n2937,
    n1702,
    n2757,
    n2930
  );


  xor
  g2912
  (
    n2966,
    n2691,
    n2937,
    n2899,
    n2927
  );


  or
  g2913
  (
    n2963,
    n1667,
    n2662,
    n1675,
    n2935
  );


  xor
  g2914
  (
    n2976,
    n2734,
    n2900,
    n2715,
    n1742
  );


  xor
  g2915
  (
    n2965,
    n2932,
    n1699,
    n1751,
    n1743
  );


  nor
  g2916
  (
    n2949,
    n1661,
    n1668,
    n1720,
    n2931
  );


  xnor
  g2917
  (
    n3006,
    n1717,
    n1731,
    n2929,
    n1721
  );


  or
  g2918
  (
    n3000,
    n2686,
    n2689,
    n2933,
    n2720
  );


  xor
  g2919
  (
    n2979,
    n2922,
    n1674,
    n1672,
    n1671
  );


  nand
  g2920
  (
    n3011,
    n2924,
    n1747,
    n1679,
    n2925
  );


  xor
  g2921
  (
    n2989,
    n2687,
    n2932,
    n1727,
    n2899
  );


  xnor
  g2922
  (
    n2992,
    n2927,
    n1722,
    n1663,
    n2756
  );


  xnor
  g2923
  (
    n2969,
    n2899,
    n2898,
    n2707,
    n2755
  );


  xor
  g2924
  (
    n3010,
    n2709,
    n2936,
    n2926,
    n1670
  );


  xnor
  g2925
  (
    n2973,
    n1741,
    n2921,
    n1748,
    n2917
  );


  xnor
  g2926
  (
    n2981,
    n2708,
    n2738,
    n2726,
    n2728
  );


  xor
  g2927
  (
    n2990,
    n2744,
    n1689,
    n2718,
    n2710
  );


  xor
  g2928
  (
    n2939,
    n2922,
    n1740,
    n2883,
    n2927
  );


  nor
  g2929
  (
    n2982,
    n2743,
    n2883,
    n2938,
    n2698
  );


  or
  g2930
  (
    n2980,
    n2902,
    n2763,
    n1676,
    n2664
  );


  xor
  g2931
  (
    n3001,
    n2681,
    n1660,
    n2699,
    n2930
  );


  or
  g2932
  (
    n3007,
    n2672,
    n2723,
    n2764,
    n2762
  );


  and
  g2933
  (
    n2946,
    n1704,
    n1723,
    n1662,
    n2930
  );


  nand
  g2934
  (
    n2983,
    n2925,
    n2706,
    n2712,
    n2731
  );


  and
  g2935
  (
    n3013,
    n2717,
    n2683,
    n2763
  );


  xnor
  g2936
  (
    n3004,
    n2935,
    n2670,
    n2938,
    n2936
  );


  and
  g2937
  (
    n2964,
    n2928,
    n2673,
    n2661,
    n2666
  );


  nand
  g2938
  (
    n2987,
    n1735,
    n1746,
    n2695,
    n1697
  );


  xnor
  g2939
  (
    n2972,
    n2703,
    n2925,
    n1700,
    n2926
  );


  nor
  g2940
  (
    n2956,
    n2722,
    n2747,
    n2915,
    n2763
  );


  nand
  g2941
  (
    n2950,
    n2936,
    n2929,
    n1745,
    n2753
  );


  nand
  g2942
  (
    n2957,
    n2759,
    n2719,
    n2923,
    n2922
  );


  and
  g2943
  (
    n2997,
    n2764,
    n1683,
    n2933,
    n2694
  );


  and
  g2944
  (
    n2968,
    n2685,
    n1734,
    n2711,
    n2674
  );


  nor
  g2945
  (
    n3012,
    n2925,
    n2928,
    n1696,
    n2902
  );


  xor
  g2946
  (
    n2999,
    n1694,
    n2725,
    n2936,
    n2737
  );


  and
  g2947
  (
    n2960,
    n1682,
    n2663,
    n2916,
    n2671
  );


  or
  g2948
  (
    n2958,
    n1724,
    n2923,
    n1680,
    n1678
  );


  nand
  g2949
  (
    n2993,
    n2667,
    n2675,
    n2752,
    n1666
  );


  xnor
  g2950
  (
    n2955,
    n2660,
    n2923,
    n2678,
    n2730
  );


  nand
  g2951
  (
    n3008,
    n1711,
    n1687,
    n2668,
    n2690
  );


  nand
  g2952
  (
    n2961,
    n1664,
    n2932,
    n1738,
    n2700
  );


  nand
  g2953
  (
    n2986,
    n2679,
    n1752,
    n2692,
    n1725
  );


  and
  g2954
  (
    n3009,
    n1690,
    n1739,
    n1728,
    n2905
  );


  or
  g2955
  (
    n2985,
    n2677,
    n2739,
    n2688,
    n2898
  );


  or
  g2956
  (
    n2991,
    n2684,
    n1665,
    n1719,
    n2727
  );


  and
  g2957
  (
    n3003,
    n1750,
    n2732,
    n2931,
    n1749
  );


  xor
  g2958
  (
    n2974,
    n2716,
    n2704,
    n2721,
    n2669
  );


  nor
  g2959
  (
    n2954,
    n2938,
    n1732,
    n2937,
    n2924
  );


  nor
  g2960
  (
    n2944,
    n2696,
    n2931,
    n1714,
    n2926
  );


  and
  g2961
  (
    n2995,
    n1729,
    n2933,
    n1686,
    n2924
  );


  and
  g2962
  (
    n2947,
    n2714,
    n1703,
    n1695,
    n2758
  );


  nor
  g2963
  (
    n2967,
    n2741,
    n2934,
    n2931,
    n2920
  );


  and
  g2964
  (
    n2941,
    n2735,
    n2924,
    n1712,
    n1698
  );


  xnor
  g2965
  (
    n2962,
    n1658,
    n2751,
    n1744,
    n2927
  );


  nand
  g2966
  (
    n2977,
    n2748,
    n1685,
    n1691,
    n2724
  );


  nand
  g2967
  (
    n2970,
    n2919,
    n2745,
    n1726,
    n2899
  );


  nor
  g2968
  (
    n2971,
    n2935,
    n2702,
    n2760,
    n2736
  );


  xor
  g2969
  (
    n2942,
    n2934,
    n2929,
    n2926,
    n1718
  );


  nand
  g2970
  (
    n2994,
    n2729,
    n1715,
    n2764,
    n1706
  );


  xor
  g2971
  (
    n3002,
    n2659,
    n1693,
    n1688,
    n1684
  );


  nand
  g2972
  (
    n2959,
    n1708,
    n2749,
    n2697,
    n2929
  );


  nor
  g2973
  (
    n2940,
    n1701,
    n1736,
    n1659,
    n2680
  );


  nand
  g2974
  (
    n2945,
    n2742,
    n2682,
    n2693,
    n2928
  );


  or
  g2975
  (
    n2978,
    n1730,
    n2764,
    n2934,
    n1713
  );


  nand
  g2976
  (
    n2948,
    n2733,
    n2928,
    n2705,
    n2935
  );


  or
  g2977
  (
    n2996,
    n2761,
    n2938,
    n1716,
    n2923
  );


  nand
  g2978
  (
    n2943,
    n1707,
    n1754,
    n2918,
    n2922
  );


  xnor
  g2979
  (
    n2984,
    n1681,
    n2750,
    n1677,
    n2665
  );


  xor
  g2980
  (
    n2951,
    n1737,
    n2900,
    n1709,
    n2676
  );


  xor
  g2981
  (
    n3017,
    n2976,
    n3000,
    n2986,
    n3013
  );


  and
  g2982
  (
    n3031,
    n2950,
    n2956,
    n2948,
    n2965
  );


  and
  g2983
  (
    n3019,
    n2963,
    n2996,
    n2968,
    n2951
  );


  xnor
  g2984
  (
    n3030,
    n2981,
    n3013,
    n2993,
    n2958
  );


  xnor
  g2985
  (
    n3015,
    n2957,
    n3003,
    n2972,
    n3005
  );


  nor
  g2986
  (
    n3014,
    n3010,
    n2946,
    n3002,
    n2990
  );


  xor
  g2987
  (
    n3025,
    n2995,
    n2977,
    n2945,
    n2979
  );


  nand
  g2988
  (
    n3023,
    n2953,
    n2984,
    n2949,
    n2997
  );


  nand
  g2989
  (
    n3029,
    n3001,
    n3008,
    n2973,
    n3013
  );


  nor
  g2990
  (
    n3028,
    n2985,
    n2992,
    n2982,
    n2940
  );


  and
  g2991
  (
    n3026,
    n2961,
    n2952,
    n2970,
    n2971
  );


  xnor
  g2992
  (
    n3032,
    n2959,
    n2974,
    n3006,
    n2991
  );


  xor
  g2993
  (
    n3020,
    n2960,
    n2975,
    n2969,
    n2943
  );


  xor
  g2994
  (
    n3022,
    n2983,
    n2994,
    n2967,
    n2941
  );


  nand
  g2995
  (
    n3024,
    n3012,
    n2998,
    n2988,
    n2944
  );


  nor
  g2996
  (
    n3016,
    n2942,
    n3007,
    n2964,
    n3011
  );


  xor
  g2997
  (
    n3021,
    n3004,
    n2966,
    n2978,
    n2999
  );


  xnor
  g2998
  (
    n3027,
    n2955,
    n2954,
    n2962,
    n2989
  );


  and
  g2999
  (
    n3018,
    n3009,
    n2980,
    n2947,
    n2987
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1693,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n2197,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n846,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1182,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1652,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n1653,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n750,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1779,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n729,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n1568,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n2727,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n88,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n192,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n2805,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1244,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1948,
    KeyNOTWire_0_15
  );


endmodule

