// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_387_1118 written by SynthGen on 2021/05/24 19:47:35
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_387_1118 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n175, n170, n167, n159, n166, n151, n174, n160,
 n157, n152, n173, n182, n162, n169, n406, n408,
 n407, n409, n411, n410);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24;

output n175, n170, n167, n159, n166, n151, n174, n160,
 n157, n152, n173, n182, n162, n169, n406, n408,
 n407, n409, n411, n410;

wire n25, n26, n27, n28, n29, n30, n31, n32,
 n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n153, n154,
 n155, n156, n158, n161, n163, n164, n165, n168,
 n171, n172, n176, n177, n178, n179, n180, n181,
 n183, n184, n185, n186, n187, n188, n189, n190,
 n191, n192, n193, n194, n195, n196, n197, n198,
 n199, n200, n201, n202, n203, n204, n205, n206,
 n207, n208, n209, n210, n211, n212, n213, n214,
 n215, n216, n217, n218, n219, n220, n221, n222,
 n223, n224, n225, n226, n227, n228, n229, n230,
 n231, n232, n233, n234, n235, n236, n237, n238,
 n239, n240, n241, n242, n243, n244, n245, n246,
 n247, n248, n249, n250, n251, n252, n253, n254,
 n255, n256, n257, n258, n259, n260, n261, n262,
 n263, n264, n265, n266, n267, n268, n269, n270,
 n271, n272, n273, n274, n275, n276, n277, n278,
 n279, n280, n281, n282, n283, n284, n285, n286,
 n287, n288, n289, n290, n291, n292, n293, n294,
 n295, n296, n297, n298, n299, n300, n301, n302,
 n303, n304, n305, n306, n307, n308, n309, n310,
 n311, n312, n313, n314, n315, n316, n317, n318,
 n319, n320, n321, n322, n323, n324, n325, n326,
 n327, n328, n329, n330, n331, n332, n333, n334,
 n335, n336, n337, n338, n339, n340, n341, n342,
 n343, n344, n345, n346, n347, n348, n349, n350,
 n351, n352, n353, n354, n355, n356, n357, n358,
 n359, n360, n361, n362, n363, n364, n365, n366,
 n367, n368, n369, n370, n371, n372, n373, n374,
 n375, n376, n377, n378, n379, n380, n381, n382,
 n383, n384, n385, n386, n387, n388, n389, n390,
 n391, n392, n393, n394, n395, n396, n397, n398,
 n399, n400, n401, n402, n403, n404, n405;

not  g0 (n66, n9);
buf  g1 (n41, n11);
not  g2 (n43, n16);
not  g3 (n45, n20);
not  g4 (n62, n14);
buf  g5 (n35, n15);
not  g6 (n61, n4);
not  g7 (n69, n4);
not  g8 (n58, n17);
not  g9 (n96, n11);
buf  g10 (n80, n22);
buf  g11 (n57, n6);
buf  g12 (n91, n18);
buf  g13 (n30, n5);
not  g14 (n67, n10);
buf  g15 (n38, n16);
not  g16 (n25, n8);
not  g17 (n60, n17);
buf  g18 (n74, n19);
buf  g19 (n100, n13);
not  g20 (n83, n14);
not  g21 (n98, n23);
not  g22 (n32, n20);
not  g23 (n99, n6);
not  g24 (n85, n15);
not  g25 (n54, n7);
buf  g26 (n75, n8);
not  g27 (n48, n10);
not  g28 (n49, n23);
buf  g29 (n97, n10);
not  g30 (n87, n6);
not  g31 (n81, n20);
buf  g32 (n70, n13);
not  g33 (n28, n18);
buf  g34 (n36, n5);
buf  g35 (n42, n12);
not  g36 (n92, n9);
not  g37 (n89, n8);
buf  g38 (n47, n23);
buf  g39 (n40, n9);
not  g40 (n84, n20);
not  g41 (n55, n15);
not  g42 (n26, n19);
buf  g43 (n72, n21);
not  g44 (n63, n11);
not  g45 (n39, n21);
not  g46 (n46, n16);
not  g47 (n102, n19);
not  g48 (n37, n13);
not  g49 (n65, n18);
not  g50 (n44, n17);
not  g51 (n82, n22);
not  g52 (n27, n1);
buf  g53 (n90, n14);
buf  g54 (n68, n2);
buf  g55 (n86, n19);
buf  g56 (n95, n18);
not  g57 (n56, n11);
not  g58 (n73, n7);
buf  g59 (n31, n7);
buf  g60 (n64, n22);
buf  g61 (n29, n7);
not  g62 (n78, n21);
buf  g63 (n76, n14);
buf  g64 (n79, n3);
not  g65 (n101, n12);
not  g66 (n88, n9);
buf  g67 (n34, n13);
not  g68 (n50, n12);
not  g69 (n53, n10);
buf  g70 (n52, n21);
not  g71 (n71, n12);
not  g72 (n77, n15);
not  g73 (n51, n6);
not  g74 (n33, n16);
not  g75 (n59, n8);
not  g76 (n94, n17);
not  g77 (n93, n22);
buf  g78 (n143, n28);
not  g79 (n147, n61);
not  g80 (n113, n67);
buf  g81 (n132, n44);
not  g82 (n107, n32);
buf  g83 (n140, n27);
buf  g84 (n130, n43);
not  g85 (n137, n56);
not  g86 (n135, n70);
not  g87 (n114, n58);
buf  g88 (n127, n64);
not  g89 (n112, n39);
not  g90 (n104, n55);
buf  g91 (n105, n59);
not  g92 (n111, n36);
buf  g93 (n148, n71);
buf  g94 (n146, n42);
buf  g95 (n118, n30);
buf  g96 (n123, n34);
not  g97 (n124, n50);
buf  g98 (n109, n48);
not  g99 (n106, n54);
buf  g100 (n149, n33);
not  g101 (n122, n60);
buf  g102 (n131, n35);
not  g103 (n117, n49);
buf  g104 (n134, n46);
not  g105 (n121, n69);
buf  g106 (n136, n37);
not  g107 (n128, n38);
buf  g108 (n115, n29);
buf  g109 (n150, n51);
buf  g110 (n120, n63);
buf  g111 (n103, n68);
buf  g112 (n116, n40);
not  g113 (n144, n31);
buf  g114 (n142, n62);
not  g115 (n119, n52);
not  g116 (n138, n72);
not  g117 (n139, n41);
not  g118 (n108, n26);
buf  g119 (n141, n53);
not  g120 (n125, n65);
buf  g121 (n133, n57);
not  g122 (n145, n25);
not  g123 (n110, n47);
not  g124 (n129, n66);
buf  g125 (n126, n45);
not  g126 (n153, n116);
buf  g127 (n155, n146);
not  g128 (n172, n135);
not  g129 (n163, n124);
not  g130 (n177, n138);
buf  g131 (n168, n137);
buf  g132 (n179, n121);
not  g133 (n161, n148);
not  g134 (n167, n145);
not  g135 (n176, n141);
not  g136 (n175, n143);
not  g137 (n152, n108);
not  g138 (n165, n139);
not  g139 (n166, n149);
buf  g140 (n178, n127);
buf  g141 (n151, n128);
not  g142 (n169, n150);
buf  g143 (n170, n133);
not  g144 (n173, n118);
not  g145 (n159, n103);
buf  g146 (n180, n136);
buf  g147 (n181, n140);
buf  g148 (n156, n114);
buf  g149 (n154, n110);
not  g150 (n164, n104);
buf  g151 (n162, n130);
and  g152 (n160, n117, n105);
xnor g153 (n158, n142, n144, n113, n106);
xnor g154 (n174, n131, n123, n129, n115);
or   g155 (n171, n119, n107, n125, n111);
and  g156 (n157, n126, n132, n120, n147);
and  g157 (n182, n134, n109, n112, n122);
not  g158 (n197, n81);
not  g159 (n189, n175);
buf  g160 (n192, n165);
not  g161 (n198, n172);
not  g162 (n186, n77);
buf  g163 (n184, n75);
buf  g164 (n195, n170);
buf  g165 (n200, n173);
buf  g166 (n199, n171);
buf  g167 (n193, n169);
not  g168 (n191, n174);
not  g169 (n190, n179);
buf  g170 (n183, n176);
buf  g171 (n187, n167);
nand g172 (n196, n80, n168);
or   g173 (n188, n177, n74, n79, n178);
xnor g174 (n185, n78, n180, n76, n73);
xor  g175 (n194, n182, n166, n181, n150);
buf  g176 (n202, n188);
buf  g177 (n210, n186);
not  g178 (n209, n189);
buf  g179 (n203, n193);
not  g180 (n211, n192);
buf  g181 (n205, n183);
buf  g182 (n201, n187);
buf  g183 (n204, n185);
buf  g184 (n208, n191);
not  g185 (n206, n190);
buf  g186 (n207, n184);
buf  g187 (n222, n205);
not  g188 (n246, n201);
buf  g189 (n252, n202);
not  g190 (n234, n209);
buf  g191 (n244, n207);
buf  g192 (n245, n202);
buf  g193 (n214, n202);
not  g194 (n248, n211);
not  g195 (n243, n207);
buf  g196 (n215, n209);
not  g197 (n216, n194);
not  g198 (n213, n205);
not  g199 (n219, n206);
buf  g200 (n229, n206);
not  g201 (n237, n203);
buf  g202 (n227, n205);
buf  g203 (n225, n207);
not  g204 (n233, n205);
not  g205 (n242, n204);
not  g206 (n241, n206);
not  g207 (n228, n204);
not  g208 (n236, n204);
buf  g209 (n232, n203);
not  g210 (n253, n209);
buf  g211 (n255, n210);
not  g212 (n247, n207);
not  g213 (n238, n209);
not  g214 (n239, n203);
buf  g215 (n226, n203);
buf  g216 (n224, n206);
not  g217 (n249, n201);
not  g218 (n212, n210);
not  g219 (n217, n208);
buf  g220 (n230, n202);
buf  g221 (n231, n211);
buf  g222 (n221, n208);
not  g223 (n250, n194);
not  g224 (n218, n208);
not  g225 (n251, n201);
not  g226 (n220, n204);
not  g227 (n235, n210);
buf  g228 (n223, n210);
buf  g229 (n240, n201);
nor  g230 (n254, n208, n211);
buf  g231 (n260, n231);
buf  g232 (n264, n215);
buf  g233 (n268, n224);
not  g234 (n256, n212);
not  g235 (n266, n226);
buf  g236 (n262, n228);
buf  g237 (n270, n218);
not  g238 (n257, n230);
buf  g239 (n273, n229);
not  g240 (n272, n223);
not  g241 (n265, n222);
buf  g242 (n267, n225);
not  g243 (n269, n217);
not  g244 (n271, n213);
buf  g245 (n259, n216);
buf  g246 (n275, n221);
buf  g247 (n261, n227);
not  g248 (n258, n219);
not  g249 (n263, n214);
buf  g250 (n274, n220);
not  g251 (n314, n263);
buf  g252 (n288, n247);
buf  g253 (n309, n264);
not  g254 (n319, n266);
not  g255 (n330, n253);
buf  g256 (n303, n238);
buf  g257 (n287, n97);
buf  g258 (n285, n264);
not  g259 (n276, n195);
buf  g260 (n304, n83);
buf  g261 (n298, n241);
not  g262 (n320, n260);
not  g263 (n315, n244);
buf  g264 (n317, n263);
not  g265 (n310, n254);
buf  g266 (n333, n195);
not  g267 (n295, n246);
buf  g268 (n318, n236);
buf  g269 (n292, n92);
buf  g270 (n301, n265);
buf  g271 (n323, n82);
not  g272 (n300, n196);
buf  g273 (n279, n268);
not  g274 (n296, n263);
not  g275 (n302, n253);
buf  g276 (n313, n253);
not  g277 (n328, n270);
buf  g278 (n307, n259);
buf  g279 (n311, n251);
not  g280 (n334, n271);
buf  g281 (n327, n271);
not  g282 (n299, n245);
not  g283 (n297, n256);
not  g284 (n290, n249);
nor  g285 (n277, n240, n250, n272);
xnor g286 (n329, n266, n270, n275, n249);
nor  g287 (n332, n89, n274, n242, n233);
and  g288 (n293, n272, n267, n268);
xnor g289 (n286, n269, n252, n262, n99);
and  g290 (n322, n273, n101, n196, n237);
xnor g291 (n321, n98, n272, n95, n250);
xor  g292 (n324, n266, n264, n250, n195);
xnor g293 (n278, n96, n274, n253);
or   g294 (n284, n197, n243, n102, n195);
xnor g295 (n335, n271, n232, n248, n252);
nand g296 (n289, n254, n251, n258, n273);
nor  g297 (n325, n251, n100, n235, n271);
and  g298 (n316, n197, n275, n250, n270);
and  g299 (n281, n265, n197, n252, n251);
nand g300 (n312, n86, n268, n267, n94);
nor  g301 (n306, n198, n196, n254, n267);
nor  g302 (n283, n257, n249, n93);
xor  g303 (n305, n269, n263, n90, n275);
xor  g304 (n331, n88, n265, n274, n239);
or   g305 (n282, n262, n84, n85, n273);
and  g306 (n326, n194, n261, n197, n264);
nor  g307 (n294, n254, n196, n267, n265);
xnor g308 (n291, n275, n273, n252, n87);
and  g309 (n280, n91, n266, n198, n270);
nor  g310 (n308, n234, n194, n269);
nor  g311 (n368, n330, n306, n326, n329);
nor  g312 (n362, n295, n317, n298, n324);
and  g313 (n364, n276, n286, n298, n310);
nor  g314 (n386, n333, n288, n311, n322);
xor  g315 (n338, n303, n286, n294);
xnor g316 (n348, n312, n329, n299, n327);
nand g317 (n346, n323, n291, n320, n328);
xnor g318 (n347, n279, n296, n331, n310);
and  g319 (n383, n321, n302, n255, n287);
nor  g320 (n337, n305, n291, n328, n325);
xor  g321 (n387, n327, n287, n295, n302);
and  g322 (n378, n295, n332, n322, n282);
nor  g323 (n342, n312, n285, n280, n325);
xnor g324 (n372, n323, n320, n307, n335);
xor  g325 (n370, n324, n319, n301, n289);
or   g326 (n391, n314, n299, n305, n278);
nor  g327 (n363, n286, n317, n303, n324);
nand g328 (n361, n306, n290, n281);
and  g329 (n341, n284, n325, n301, n320);
xnor g330 (n376, n311, n314, n302, n307);
nand g331 (n379, n304, n329, n293, n294);
xnor g332 (n351, n321, n292, n313, n332);
xnor g333 (n373, n335, n308, n333, n316);
xnor g334 (n381, n324, n289, n316, n293);
nand g335 (n336, n327, n305, n283, n322);
xor  g336 (n390, n307, n299, n301, n288);
xor  g337 (n354, n334, n255, n294, n331);
and  g338 (n340, n298, n300, n332, n296);
nand g339 (n343, n335, n331, n297, n289);
nand g340 (n350, n317, n24, n286, n314);
nor  g341 (n366, n284, n313, n307, n323);
nand g342 (n382, n317, n326, n303, n318);
xnor g343 (n344, n297, n296, n283, n295);
xor  g344 (n380, n292, n309, n308, n24);
xor  g345 (n357, n288, n291, n293, n304);
nor  g346 (n359, n312, n318, n292, n255);
xnor g347 (n360, n311, n316, n321);
xnor g348 (n375, n285, n315, n319, n331);
nand g349 (n339, n304, n313, n287, n308);
xor  g350 (n367, n326, n292, n330, n300);
xor  g351 (n358, n332, n309, n306, n334);
nor  g352 (n374, n319, n300, n310, n277);
nand g353 (n352, n334, n297, n301, n325);
and  g354 (n389, n24, n318, n315, n291);
or   g355 (n384, n308, n288, n289, n328);
xnor g356 (n353, n297, n330, n309, n290);
nand g357 (n355, n296, n305, n309, n313);
and  g358 (n369, n328, n300, n24, n326);
and  g359 (n388, n303, n285, n333, n293);
and  g360 (n371, n323, n23, n298, n304);
xor  g361 (n356, n299, n334, n318, n330);
and  g362 (n377, n320, n333, n287, n329);
nand g363 (n385, n335, n255, n312, n315);
and  g364 (n349, n322, n314, n310, n315);
xor  g365 (n365, n302, n290, n327, n306);
xor  g366 (n345, n319, n311, n316, n285);
or   g367 (n399, n345, n364, n360, n377);
or   g368 (n392, n337, n378, n340, n344);
nand g369 (n401, n356, n341, n389, n384);
xnor g370 (n405, n370, n348, n358, n373);
nor  g371 (n403, n379, n359, n390, n363);
xnor g372 (n398, n346, n380, n342, n367);
nand g373 (n397, n355, n374, n383, n369);
nor  g374 (n393, n339, n354, n361, n382);
nand g375 (n404, n388, n347, n357, n336);
and  g376 (n394, n385, n343, n349, n387);
nand g377 (n402, n368, n352, n350, n386);
nand g378 (n396, n372, n375, n366, n353);
or   g379 (n400, n338, n362, n351, n365);
xnor g380 (n395, n371, n376, n381, n391);
and  g381 (n409, n394, n402, n200, n395);
or   g382 (n408, n401, n200, n199, n403);
and  g383 (n411, n397, n393, n392, n198);
nor  g384 (n407, n200, n396, n199, n404);
and  g385 (n410, n198, n199, n200, n398);
nor  g386 (n406, n199, n399, n405, n400);
endmodule
