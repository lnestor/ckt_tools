

module Stat_1789_21_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n732,
  n813,
  n1808,
  n1797,
  n1792,
  n1798,
  n1810,
  n1796,
  n1811,
  n1804,
  n1787,
  n1807,
  n1814,
  n1786,
  n1794,
  n1812,
  n1789,
  n1790,
  n1791,
  n1799,
  n1795,
  n1805,
  n1800,
  n1801,
  n1788,
  n1803,
  n1806,
  n1793,
  n1813,
  n1802,
  n1809,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n732;
  output n813;
  output n1808;
  output n1797;
  output n1792;
  output n1798;
  output n1810;
  output n1796;
  output n1811;
  output n1804;
  output n1787;
  output n1807;
  output n1814;
  output n1786;
  output n1794;
  output n1812;
  output n1789;
  output n1790;
  output n1791;
  output n1799;
  output n1795;
  output n1805;
  output n1800;
  output n1801;
  output n1788;
  output n1803;
  output n1806;
  output n1793;
  output n1813;
  output n1802;
  output n1809;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  not
  g0
  (
    n98,
    n4
  );


  not
  g1
  (
    n26,
    n3
  );


  buf
  g2
  (
    n48,
    n20
  );


  not
  g3
  (
    n32,
    n13
  );


  not
  g4
  (
    n71,
    n19
  );


  buf
  g5
  (
    n64,
    n5
  );


  buf
  g6
  (
    n43,
    n14
  );


  not
  g7
  (
    n100,
    n1
  );


  buf
  g8
  (
    n89,
    n5
  );


  not
  g9
  (
    n44,
    n10
  );


  not
  g10
  (
    n55,
    n19
  );


  not
  g11
  (
    n35,
    n8
  );


  buf
  g12
  (
    n91,
    n12
  );


  not
  g13
  (
    n52,
    n6
  );


  not
  g14
  (
    n95,
    n15
  );


  not
  g15
  (
    n46,
    n21
  );


  not
  g16
  (
    n103,
    n18
  );


  buf
  g17
  (
    n36,
    n18
  );


  not
  g18
  (
    n60,
    n3
  );


  not
  g19
  (
    n56,
    n8
  );


  buf
  g20
  (
    n94,
    n19
  );


  buf
  g21
  (
    n31,
    n17
  );


  not
  g22
  (
    n61,
    n15
  );


  buf
  g23
  (
    n58,
    n11
  );


  not
  g24
  (
    n77,
    n16
  );


  buf
  g25
  (
    n39,
    n14
  );


  buf
  g26
  (
    n66,
    n18
  );


  buf
  g27
  (
    n87,
    n2
  );


  not
  g28
  (
    n99,
    n20
  );


  not
  g29
  (
    n93,
    n4
  );


  buf
  g30
  (
    n65,
    n11
  );


  buf
  g31
  (
    n84,
    n10
  );


  buf
  g32
  (
    n57,
    n15
  );


  buf
  g33
  (
    n73,
    n3
  );


  buf
  g34
  (
    n74,
    n17
  );


  buf
  g35
  (
    n50,
    n5
  );


  buf
  g36
  (
    n78,
    n9
  );


  not
  g37
  (
    n67,
    n16
  );


  buf
  g38
  (
    KeyWire_0_19,
    n7
  );


  buf
  g39
  (
    n51,
    n14
  );


  not
  g40
  (
    n34,
    n10
  );


  buf
  g41
  (
    n28,
    n1
  );


  not
  g42
  (
    n62,
    n7
  );


  buf
  g43
  (
    n47,
    n11
  );


  not
  g44
  (
    n41,
    n5
  );


  not
  g45
  (
    n85,
    n18
  );


  buf
  g46
  (
    n30,
    n7
  );


  buf
  g47
  (
    n80,
    n2
  );


  buf
  g48
  (
    n81,
    n4
  );


  buf
  g49
  (
    n101,
    n16
  );


  not
  g50
  (
    n53,
    n13
  );


  not
  g51
  (
    n42,
    n6
  );


  not
  g52
  (
    n45,
    n10
  );


  not
  g53
  (
    n33,
    n4
  );


  buf
  g54
  (
    n27,
    n3
  );


  not
  g55
  (
    n38,
    n11
  );


  not
  g56
  (
    n83,
    n8
  );


  not
  g57
  (
    n102,
    n15
  );


  not
  g58
  (
    n49,
    n8
  );


  buf
  g59
  (
    n90,
    n9
  );


  not
  g60
  (
    n63,
    n20
  );


  buf
  g61
  (
    n106,
    n17
  );


  buf
  g62
  (
    n96,
    n14
  );


  not
  g63
  (
    n86,
    n17
  );


  buf
  g64
  (
    n37,
    n12
  );


  buf
  g65
  (
    n75,
    n9
  );


  buf
  g66
  (
    n40,
    n2
  );


  buf
  g67
  (
    n82,
    n13
  );


  not
  g68
  (
    n88,
    n6
  );


  not
  g69
  (
    n54,
    n1
  );


  buf
  g70
  (
    n69,
    n20
  );


  buf
  g71
  (
    KeyWire_0_5,
    n7
  );


  buf
  g72
  (
    n97,
    n6
  );


  buf
  g73
  (
    n68,
    n19
  );


  buf
  g74
  (
    n76,
    n12
  );


  not
  g75
  (
    n70,
    n9
  );


  buf
  g76
  (
    n105,
    n12
  );


  buf
  g77
  (
    n59,
    n13
  );


  buf
  g78
  (
    KeyWire_0_27,
    n2
  );


  not
  g79
  (
    n79,
    n16
  );


  not
  g80
  (
    n72,
    n1
  );


  not
  g81
  (
    n214,
    n73
  );


  buf
  g82
  (
    n159,
    n42
  );


  not
  g83
  (
    n186,
    n79
  );


  not
  g84
  (
    n373,
    n102
  );


  not
  g85
  (
    n344,
    n76
  );


  buf
  g86
  (
    n405,
    n63
  );


  not
  g87
  (
    n364,
    n74
  );


  not
  g88
  (
    n394,
    n37
  );


  not
  g89
  (
    n162,
    n39
  );


  buf
  g90
  (
    n340,
    n92
  );


  not
  g91
  (
    n294,
    n68
  );


  buf
  g92
  (
    n234,
    n57
  );


  not
  g93
  (
    n332,
    n27
  );


  buf
  g94
  (
    n257,
    n47
  );


  not
  g95
  (
    n318,
    n72
  );


  not
  g96
  (
    n163,
    n49
  );


  buf
  g97
  (
    n360,
    n67
  );


  not
  g98
  (
    n131,
    n71
  );


  not
  g99
  (
    n237,
    n76
  );


  not
  g100
  (
    n115,
    n31
  );


  not
  g101
  (
    n156,
    n57
  );


  not
  g102
  (
    n208,
    n77
  );


  not
  g103
  (
    n111,
    n95
  );


  not
  g104
  (
    n225,
    n74
  );


  buf
  g105
  (
    n406,
    n61
  );


  not
  g106
  (
    n414,
    n50
  );


  not
  g107
  (
    n302,
    n67
  );


  buf
  g108
  (
    n253,
    n101
  );


  buf
  g109
  (
    n236,
    n54
  );


  not
  g110
  (
    n321,
    n60
  );


  not
  g111
  (
    n217,
    n75
  );


  buf
  g112
  (
    n140,
    n55
  );


  not
  g113
  (
    n410,
    n99
  );


  buf
  g114
  (
    n325,
    n81
  );


  buf
  g115
  (
    n351,
    n73
  );


  not
  g116
  (
    n285,
    n42
  );


  buf
  g117
  (
    n215,
    n30
  );


  not
  g118
  (
    n232,
    n90
  );


  not
  g119
  (
    n395,
    n45
  );


  buf
  g120
  (
    n280,
    n85
  );


  not
  g121
  (
    n187,
    n81
  );


  buf
  g122
  (
    n164,
    n49
  );


  buf
  g123
  (
    n135,
    n93
  );


  not
  g124
  (
    n370,
    n68
  );


  buf
  g125
  (
    n390,
    n48
  );


  not
  g126
  (
    n388,
    n42
  );


  buf
  g127
  (
    n313,
    n36
  );


  not
  g128
  (
    n362,
    n61
  );


  buf
  g129
  (
    n261,
    n55
  );


  not
  g130
  (
    n396,
    n83
  );


  buf
  g131
  (
    n377,
    n28
  );


  not
  g132
  (
    n165,
    n92
  );


  buf
  g133
  (
    n178,
    n31
  );


  buf
  g134
  (
    KeyWire_0_15,
    n59
  );


  buf
  g135
  (
    n315,
    n53
  );


  not
  g136
  (
    n407,
    n95
  );


  buf
  g137
  (
    n317,
    n26
  );


  not
  g138
  (
    n250,
    n27
  );


  buf
  g139
  (
    n244,
    n77
  );


  not
  g140
  (
    n322,
    n85
  );


  buf
  g141
  (
    n326,
    n54
  );


  buf
  g142
  (
    n352,
    n102
  );


  buf
  g143
  (
    n306,
    n70
  );


  buf
  g144
  (
    n116,
    n43
  );


  not
  g145
  (
    n350,
    n77
  );


  not
  g146
  (
    n266,
    n75
  );


  buf
  g147
  (
    n147,
    n54
  );


  buf
  g148
  (
    n144,
    n88
  );


  not
  g149
  (
    n305,
    n65
  );


  buf
  g150
  (
    n193,
    n82
  );


  buf
  g151
  (
    n122,
    n32
  );


  not
  g152
  (
    n158,
    n59
  );


  buf
  g153
  (
    n132,
    n88
  );


  buf
  g154
  (
    n386,
    n78
  );


  not
  g155
  (
    n320,
    n28
  );


  buf
  g156
  (
    n278,
    n97
  );


  buf
  g157
  (
    n153,
    n89
  );


  buf
  g158
  (
    n287,
    n26
  );


  buf
  g159
  (
    n281,
    n95
  );


  buf
  g160
  (
    n372,
    n91
  );


  not
  g161
  (
    n363,
    n70
  );


  buf
  g162
  (
    n251,
    n57
  );


  buf
  g163
  (
    n355,
    n35
  );


  not
  g164
  (
    n114,
    n63
  );


  buf
  g165
  (
    n110,
    n47
  );


  buf
  g166
  (
    n272,
    n90
  );


  not
  g167
  (
    n269,
    n51
  );


  not
  g168
  (
    n284,
    n80
  );


  not
  g169
  (
    n310,
    n39
  );


  not
  g170
  (
    n231,
    n64
  );


  not
  g171
  (
    n233,
    n78
  );


  buf
  g172
  (
    n229,
    n67
  );


  buf
  g173
  (
    n401,
    n58
  );


  buf
  g174
  (
    n262,
    n81
  );


  buf
  g175
  (
    n338,
    n59
  );


  buf
  g176
  (
    n190,
    n84
  );


  not
  g177
  (
    n341,
    n37
  );


  buf
  g178
  (
    n346,
    n74
  );


  buf
  g179
  (
    n380,
    n53
  );


  buf
  g180
  (
    n169,
    n39
  );


  not
  g181
  (
    n299,
    n93
  );


  buf
  g182
  (
    n197,
    n80
  );


  buf
  g183
  (
    n282,
    n44
  );


  buf
  g184
  (
    n289,
    n48
  );


  not
  g185
  (
    n277,
    n33
  );


  not
  g186
  (
    n118,
    n97
  );


  buf
  g187
  (
    n182,
    n45
  );


  not
  g188
  (
    n271,
    n48
  );


  not
  g189
  (
    n398,
    n70
  );


  buf
  g190
  (
    n167,
    n96
  );


  buf
  g191
  (
    n195,
    n33
  );


  buf
  g192
  (
    n378,
    n97
  );


  not
  g193
  (
    n241,
    n46
  );


  buf
  g194
  (
    n374,
    n50
  );


  not
  g195
  (
    n113,
    n34
  );


  not
  g196
  (
    n335,
    n41
  );


  not
  g197
  (
    n146,
    n29
  );


  not
  g198
  (
    n411,
    n86
  );


  not
  g199
  (
    n336,
    n29
  );


  buf
  g200
  (
    n154,
    n56
  );


  buf
  g201
  (
    n356,
    n78
  );


  buf
  g202
  (
    n379,
    n99
  );


  buf
  g203
  (
    n218,
    n79
  );


  buf
  g204
  (
    n412,
    n60
  );


  not
  g205
  (
    n267,
    n98
  );


  not
  g206
  (
    n143,
    n44
  );


  not
  g207
  (
    n201,
    n42
  );


  not
  g208
  (
    n188,
    n34
  );


  buf
  g209
  (
    n183,
    n89
  );


  not
  g210
  (
    n124,
    n84
  );


  not
  g211
  (
    n137,
    n63
  );


  buf
  g212
  (
    n358,
    n48
  );


  buf
  g213
  (
    n357,
    n62
  );


  buf
  g214
  (
    n328,
    n56
  );


  buf
  g215
  (
    n181,
    n38
  );


  not
  g216
  (
    n226,
    n47
  );


  buf
  g217
  (
    n168,
    n51
  );


  not
  g218
  (
    n296,
    n91
  );


  buf
  g219
  (
    n397,
    n29
  );


  not
  g220
  (
    n354,
    n90
  );


  not
  g221
  (
    n275,
    n69
  );


  buf
  g222
  (
    n141,
    n75
  );


  not
  g223
  (
    n298,
    n85
  );


  buf
  g224
  (
    n133,
    n38
  );


  not
  g225
  (
    KeyWire_0_18,
    n30
  );


  buf
  g226
  (
    n273,
    n81
  );


  buf
  g227
  (
    n265,
    n96
  );


  buf
  g228
  (
    n136,
    n36
  );


  buf
  g229
  (
    n368,
    n66
  );


  buf
  g230
  (
    n112,
    n100
  );


  not
  g231
  (
    n120,
    n96
  );


  not
  g232
  (
    n199,
    n63
  );


  buf
  g233
  (
    n129,
    n84
  );


  buf
  g234
  (
    n301,
    n88
  );


  buf
  g235
  (
    n107,
    n40
  );


  not
  g236
  (
    n319,
    n34
  );


  buf
  g237
  (
    n185,
    n52
  );


  buf
  g238
  (
    n160,
    n43
  );


  not
  g239
  (
    n216,
    n92
  );


  not
  g240
  (
    n139,
    n27
  );


  buf
  g241
  (
    n327,
    n37
  );


  not
  g242
  (
    n400,
    n101
  );


  not
  g243
  (
    n258,
    n73
  );


  buf
  g244
  (
    n180,
    n53
  );


  buf
  g245
  (
    n399,
    n28
  );


  not
  g246
  (
    n393,
    n98
  );


  not
  g247
  (
    n324,
    n32
  );


  not
  g248
  (
    n375,
    n82
  );


  buf
  g249
  (
    n347,
    n72
  );


  not
  g250
  (
    n308,
    n58
  );


  buf
  g251
  (
    n295,
    n80
  );


  buf
  g252
  (
    n176,
    n31
  );


  buf
  g253
  (
    n245,
    n86
  );


  buf
  g254
  (
    n246,
    n30
  );


  not
  g255
  (
    n259,
    n95
  );


  buf
  g256
  (
    n290,
    n89
  );


  buf
  g257
  (
    n145,
    n73
  );


  not
  g258
  (
    n337,
    n58
  );


  buf
  g259
  (
    n151,
    n26
  );


  buf
  g260
  (
    n148,
    n54
  );


  not
  g261
  (
    n307,
    n87
  );


  buf
  g262
  (
    n309,
    n46
  );


  not
  g263
  (
    n369,
    n84
  );


  buf
  g264
  (
    n198,
    n52
  );


  buf
  g265
  (
    n171,
    n76
  );


  buf
  g266
  (
    n409,
    n27
  );


  buf
  g267
  (
    n387,
    n80
  );


  not
  g268
  (
    n256,
    n53
  );


  not
  g269
  (
    n239,
    n33
  );


  buf
  g270
  (
    n196,
    n65
  );


  buf
  g271
  (
    n300,
    n55
  );


  buf
  g272
  (
    n219,
    n61
  );


  buf
  g273
  (
    n138,
    n26
  );


  buf
  g274
  (
    n184,
    n98
  );


  buf
  g275
  (
    n345,
    n77
  );


  not
  g276
  (
    n384,
    n68
  );


  buf
  g277
  (
    n402,
    n99
  );


  not
  g278
  (
    n211,
    n93
  );


  not
  g279
  (
    n210,
    n62
  );


  not
  g280
  (
    n312,
    n102
  );


  not
  g281
  (
    n274,
    n94
  );


  not
  g282
  (
    n297,
    n91
  );


  buf
  g283
  (
    n123,
    n76
  );


  buf
  g284
  (
    n150,
    n46
  );


  buf
  g285
  (
    n126,
    n64
  );


  not
  g286
  (
    n125,
    n41
  );


  not
  g287
  (
    n252,
    n87
  );


  not
  g288
  (
    n365,
    n44
  );


  buf
  g289
  (
    n209,
    n79
  );


  buf
  g290
  (
    n170,
    n44
  );


  buf
  g291
  (
    n108,
    n101
  );


  buf
  g292
  (
    n238,
    n56
  );


  buf
  g293
  (
    n109,
    n41
  );


  not
  g294
  (
    n329,
    n86
  );


  not
  g295
  (
    n349,
    n94
  );


  not
  g296
  (
    n127,
    n99
  );


  buf
  g297
  (
    n367,
    n50
  );


  not
  g298
  (
    n204,
    n43
  );


  buf
  g299
  (
    n194,
    n101
  );


  not
  g300
  (
    n221,
    n64
  );


  buf
  g301
  (
    n268,
    n71
  );


  buf
  g302
  (
    n334,
    n33
  );


  not
  g303
  (
    n189,
    n43
  );


  buf
  g304
  (
    n291,
    n96
  );


  not
  g305
  (
    n292,
    n45
  );


  buf
  g306
  (
    n413,
    n85
  );


  buf
  g307
  (
    n383,
    n91
  );


  buf
  g308
  (
    n227,
    n71
  );


  not
  g309
  (
    n128,
    n75
  );


  buf
  g310
  (
    n228,
    n83
  );


  not
  g311
  (
    n382,
    n66
  );


  not
  g312
  (
    n175,
    n86
  );


  not
  g313
  (
    n260,
    n97
  );


  buf
  g314
  (
    n119,
    n92
  );


  not
  g315
  (
    n279,
    n49
  );


  not
  g316
  (
    n179,
    n56
  );


  buf
  g317
  (
    n359,
    n59
  );


  buf
  g318
  (
    n166,
    n62
  );


  buf
  g319
  (
    n371,
    n30
  );


  buf
  g320
  (
    n304,
    n66
  );


  buf
  g321
  (
    n323,
    n60
  );


  not
  g322
  (
    n348,
    n47
  );


  not
  g323
  (
    n263,
    n64
  );


  not
  g324
  (
    n255,
    n71
  );


  not
  g325
  (
    n288,
    n67
  );


  buf
  g326
  (
    n283,
    n46
  );


  buf
  g327
  (
    n264,
    n57
  );


  not
  g328
  (
    n331,
    n65
  );


  not
  g329
  (
    n254,
    n88
  );


  buf
  g330
  (
    n121,
    n98
  );


  not
  g331
  (
    n391,
    n38
  );


  buf
  g332
  (
    n408,
    n35
  );


  not
  g333
  (
    n361,
    n50
  );


  not
  g334
  (
    n314,
    n52
  );


  not
  g335
  (
    n155,
    n83
  );


  not
  g336
  (
    n200,
    n49
  );


  not
  g337
  (
    n213,
    n32
  );


  not
  g338
  (
    n316,
    n82
  );


  not
  g339
  (
    n230,
    n94
  );


  not
  g340
  (
    n249,
    n29
  );


  not
  g341
  (
    KeyWire_0_24,
    n51
  );


  not
  g342
  (
    n333,
    n36
  );


  buf
  g343
  (
    KeyWire_0_6,
    n78
  );


  buf
  g344
  (
    n243,
    n69
  );


  buf
  g345
  (
    n343,
    n83
  );


  buf
  g346
  (
    n224,
    n36
  );


  buf
  g347
  (
    n276,
    n52
  );


  buf
  g348
  (
    n235,
    n39
  );


  buf
  g349
  (
    n311,
    n55
  );


  not
  g350
  (
    n286,
    n41
  );


  buf
  g351
  (
    n242,
    n35
  );


  buf
  g352
  (
    n223,
    n69
  );


  not
  g353
  (
    n389,
    n37
  );


  not
  g354
  (
    n149,
    n58
  );


  buf
  g355
  (
    n330,
    n74
  );


  buf
  g356
  (
    n202,
    n102
  );


  buf
  g357
  (
    n117,
    n100
  );


  buf
  g358
  (
    n339,
    n28
  );


  not
  g359
  (
    n203,
    n60
  );


  not
  g360
  (
    n248,
    n38
  );


  not
  g361
  (
    n220,
    n100
  );


  not
  g362
  (
    n222,
    n72
  );


  buf
  g363
  (
    n134,
    n87
  );


  not
  g364
  (
    n385,
    n31
  );


  buf
  g365
  (
    n270,
    n90
  );


  not
  g366
  (
    n173,
    n61
  );


  buf
  g367
  (
    n392,
    n79
  );


  buf
  g368
  (
    n142,
    n51
  );


  not
  g369
  (
    n381,
    n72
  );


  buf
  g370
  (
    n212,
    n32
  );


  not
  g371
  (
    n152,
    n94
  );


  buf
  g372
  (
    n161,
    n35
  );


  buf
  g373
  (
    n172,
    n62
  );


  buf
  g374
  (
    n192,
    n69
  );


  buf
  g375
  (
    n366,
    n40
  );


  buf
  g376
  (
    n207,
    n66
  );


  buf
  g377
  (
    n247,
    n100
  );


  not
  g378
  (
    n174,
    n34
  );


  not
  g379
  (
    n130,
    n70
  );


  buf
  g380
  (
    n376,
    n40
  );


  buf
  g381
  (
    n240,
    n45
  );


  not
  g382
  (
    n205,
    n65
  );


  buf
  g383
  (
    n191,
    n40
  );


  not
  g384
  (
    n353,
    n89
  );


  not
  g385
  (
    n303,
    n87
  );


  not
  g386
  (
    n206,
    n93
  );


  not
  g387
  (
    n157,
    n82
  );


  buf
  g388
  (
    n177,
    n68
  );


  buf
  g389
  (
    n423,
    n340
  );


  not
  g390
  (
    n680,
    n21
  );


  not
  g391
  (
    n431,
    n167
  );


  buf
  g392
  (
    n512,
    n364
  );


  not
  g393
  (
    n445,
    n226
  );


  buf
  g394
  (
    n440,
    n367
  );


  not
  g395
  (
    n521,
    n322
  );


  not
  g396
  (
    n520,
    n203
  );


  buf
  g397
  (
    n470,
    n201
  );


  not
  g398
  (
    n502,
    n154
  );


  buf
  g399
  (
    n637,
    n183
  );


  buf
  g400
  (
    n618,
    n363
  );


  not
  g401
  (
    n464,
    n357
  );


  not
  g402
  (
    n657,
    n376
  );


  not
  g403
  (
    n534,
    n384
  );


  not
  g404
  (
    n463,
    n339
  );


  buf
  g405
  (
    n623,
    n321
  );


  not
  g406
  (
    n640,
    n373
  );


  buf
  g407
  (
    n533,
    n130
  );


  buf
  g408
  (
    n660,
    n133
  );


  not
  g409
  (
    n418,
    n314
  );


  not
  g410
  (
    n519,
    n282
  );


  not
  g411
  (
    n621,
    n334
  );


  buf
  g412
  (
    n528,
    n349
  );


  not
  g413
  (
    n585,
    n268
  );


  not
  g414
  (
    n659,
    n241
  );


  not
  g415
  (
    n508,
    n343
  );


  not
  g416
  (
    n617,
    n375
  );


  not
  g417
  (
    n551,
    n209
  );


  buf
  g418
  (
    n525,
    n338
  );


  not
  g419
  (
    n554,
    n219
  );


  not
  g420
  (
    n557,
    n362
  );


  not
  g421
  (
    n609,
    n366
  );


  buf
  g422
  (
    n648,
    n340
  );


  not
  g423
  (
    n583,
    n290
  );


  not
  g424
  (
    n449,
    n378
  );


  not
  g425
  (
    n604,
    n347
  );


  buf
  g426
  (
    n523,
    n166
  );


  buf
  g427
  (
    n596,
    n143
  );


  not
  g428
  (
    n529,
    n199
  );


  buf
  g429
  (
    n608,
    n341
  );


  not
  g430
  (
    n480,
    n309
  );


  not
  g431
  (
    n441,
    n207
  );


  buf
  g432
  (
    n575,
    n22
  );


  buf
  g433
  (
    n550,
    n312
  );


  buf
  g434
  (
    n587,
    n381
  );


  buf
  g435
  (
    n457,
    n177
  );


  not
  g436
  (
    n496,
    n267
  );


  buf
  g437
  (
    n438,
    n289
  );


  not
  g438
  (
    n573,
    n238
  );


  buf
  g439
  (
    n670,
    n296
  );


  not
  g440
  (
    n421,
    n379
  );


  buf
  g441
  (
    n600,
    n369
  );


  not
  g442
  (
    n510,
    n202
  );


  not
  g443
  (
    n630,
    n370
  );


  not
  g444
  (
    n579,
    n375
  );


  buf
  g445
  (
    n539,
    n169
  );


  buf
  g446
  (
    n627,
    n351
  );


  buf
  g447
  (
    n432,
    n360
  );


  not
  g448
  (
    n668,
    n382
  );


  not
  g449
  (
    n461,
    n377
  );


  not
  g450
  (
    n607,
    n264
  );


  not
  g451
  (
    n576,
    n379
  );


  not
  g452
  (
    n645,
    n337
  );


  buf
  g453
  (
    n499,
    n320
  );


  not
  g454
  (
    n527,
    n266
  );


  not
  g455
  (
    n631,
    n23
  );


  not
  g456
  (
    n515,
    n338
  );


  buf
  g457
  (
    n633,
    n336
  );


  buf
  g458
  (
    n484,
    n131
  );


  buf
  g459
  (
    n435,
    n375
  );


  not
  g460
  (
    n543,
    n189
  );


  buf
  g461
  (
    n634,
    n237
  );


  buf
  g462
  (
    n590,
    n280
  );


  not
  g463
  (
    n507,
    n347
  );


  not
  g464
  (
    n462,
    n344
  );


  buf
  g465
  (
    n558,
    n160
  );


  xnor
  g466
  (
    n584,
    n346,
    n385
  );


  or
  g467
  (
    n531,
    n134,
    n210
  );


  nor
  g468
  (
    n615,
    n381,
    n255
  );


  nor
  g469
  (
    n620,
    n185,
    n145
  );


  and
  g470
  (
    n514,
    n370,
    n384
  );


  or
  g471
  (
    n493,
    n363,
    n369
  );


  not
  g472
  (
    n629,
    n386
  );


  and
  g473
  (
    n429,
    n284,
    n277
  );


  nand
  g474
  (
    KeyWire_0_2,
    n142,
    n120
  );


  nor
  g475
  (
    n536,
    n371,
    n125
  );


  nor
  g476
  (
    n610,
    n136,
    n366
  );


  xor
  g477
  (
    n419,
    n353,
    n317
  );


  nand
  g478
  (
    n522,
    n345,
    n371
  );


  nor
  g479
  (
    n549,
    n372,
    n362
  );


  or
  g480
  (
    n665,
    n360,
    n150
  );


  nand
  g481
  (
    n427,
    n339,
    n368
  );


  xor
  g482
  (
    n597,
    n355,
    n371
  );


  or
  g483
  (
    n572,
    n383,
    n301
  );


  or
  g484
  (
    n489,
    n386,
    n369
  );


  xnor
  g485
  (
    n478,
    n387,
    n257
  );


  and
  g486
  (
    n471,
    n374,
    n376
  );


  or
  g487
  (
    n428,
    n365,
    n311
  );


  nand
  g488
  (
    n458,
    n192,
    n223
  );


  nor
  g489
  (
    n562,
    n157,
    n351
  );


  xnor
  g490
  (
    n453,
    n112,
    n308
  );


  and
  g491
  (
    n425,
    n113,
    n378
  );


  or
  g492
  (
    n564,
    n366,
    n336
  );


  and
  g493
  (
    n555,
    n332,
    n211
  );


  nand
  g494
  (
    n658,
    n186,
    n107
  );


  xnor
  g495
  (
    n437,
    n364,
    n251
  );


  nor
  g496
  (
    n448,
    n170,
    n368
  );


  and
  g497
  (
    n469,
    n354,
    n151
  );


  xor
  g498
  (
    n628,
    n368,
    n22
  );


  nand
  g499
  (
    n612,
    n147,
    n262
  );


  or
  g500
  (
    n433,
    n109,
    n357
  );


  xor
  g501
  (
    n663,
    n294,
    n263
  );


  or
  g502
  (
    n532,
    n325,
    n214
  );


  nor
  g503
  (
    n439,
    n122,
    n349
  );


  and
  g504
  (
    n481,
    n353,
    n234
  );


  xnor
  g505
  (
    n662,
    n132,
    n377
  );


  nor
  g506
  (
    n467,
    n356,
    n24
  );


  nand
  g507
  (
    n599,
    n138,
    n345
  );


  xnor
  g508
  (
    n544,
    n127,
    n247
  );


  nor
  g509
  (
    n446,
    n337,
    n359
  );


  and
  g510
  (
    n614,
    n358,
    n378
  );


  nand
  g511
  (
    n415,
    n231,
    n243
  );


  xor
  g512
  (
    n676,
    n286,
    n25
  );


  and
  g513
  (
    n625,
    n353,
    n114
  );


  xor
  g514
  (
    n538,
    n213,
    n345
  );


  and
  g515
  (
    n483,
    n323,
    n362
  );


  xor
  g516
  (
    n568,
    n222,
    n337
  );


  or
  g517
  (
    n547,
    n346,
    n135
  );


  or
  g518
  (
    n566,
    n22,
    n341
  );


  or
  g519
  (
    n571,
    n291,
    n144
  );


  xnor
  g520
  (
    n513,
    n342,
    n364
  );


  xnor
  g521
  (
    n451,
    n358,
    n272
  );


  and
  g522
  (
    n635,
    n252,
    n117
  );


  xor
  g523
  (
    n516,
    n292,
    n298
  );


  nor
  g524
  (
    n485,
    n191,
    n274
  );


  xnor
  g525
  (
    n651,
    n240,
    n229
  );


  xor
  g526
  (
    n491,
    n355,
    n340
  );


  xnor
  g527
  (
    n580,
    n141,
    n174
  );


  and
  g528
  (
    n541,
    n236,
    n385
  );


  nor
  g529
  (
    n501,
    n279,
    n352
  );


  and
  g530
  (
    n653,
    n355,
    n357
  );


  and
  g531
  (
    n490,
    n380,
    n363
  );


  nor
  g532
  (
    n626,
    n198,
    n359
  );


  nand
  g533
  (
    n518,
    n357,
    n381
  );


  and
  g534
  (
    n540,
    n377,
    n360
  );


  nor
  g535
  (
    n506,
    n348,
    n146
  );


  xor
  g536
  (
    n473,
    n352,
    n230
  );


  xnor
  g537
  (
    n588,
    n361,
    n197
  );


  and
  g538
  (
    n595,
    n140,
    n23
  );


  xor
  g539
  (
    n416,
    n233,
    n128
  );


  and
  g540
  (
    n561,
    n350,
    n347
  );


  xor
  g541
  (
    n477,
    n370,
    n386
  );


  and
  g542
  (
    n619,
    n361,
    n270
  );


  or
  g543
  (
    n553,
    n341,
    n24
  );


  nor
  g544
  (
    n589,
    n365,
    n361
  );


  xnor
  g545
  (
    n505,
    n108,
    n288
  );


  nor
  g546
  (
    n678,
    n121,
    n355
  );


  xnor
  g547
  (
    n509,
    n180,
    n24
  );


  nand
  g548
  (
    n581,
    n342,
    n22
  );


  or
  g549
  (
    n592,
    n354,
    n158
  );


  xor
  g550
  (
    n430,
    n129,
    n367
  );


  or
  g551
  (
    n422,
    n245,
    n336
  );


  xnor
  g552
  (
    n652,
    n356,
    n338
  );


  or
  g553
  (
    KeyWire_0_3,
    n220,
    n382
  );


  nand
  g554
  (
    n643,
    n353,
    n149
  );


  nand
  g555
  (
    n524,
    n153,
    n281
  );


  and
  g556
  (
    n601,
    n344,
    n253
  );


  and
  g557
  (
    n603,
    n232,
    n350
  );


  xnor
  g558
  (
    KeyWire_0_12,
    n261,
    n249
  );


  nand
  g559
  (
    n563,
    n319,
    n387
  );


  or
  g560
  (
    n622,
    n139,
    n228
  );


  nand
  g561
  (
    n569,
    n224,
    n354
  );


  or
  g562
  (
    n556,
    n380,
    n259
  );


  xor
  g563
  (
    n475,
    n118,
    n218
  );


  nor
  g564
  (
    n460,
    n111,
    n343
  );


  nor
  g565
  (
    n466,
    n244,
    n376
  );


  nand
  g566
  (
    n632,
    n119,
    n116
  );


  xor
  g567
  (
    n482,
    n307,
    n379
  );


  and
  g568
  (
    n577,
    n356,
    n235
  );


  nor
  g569
  (
    n639,
    n315,
    n273
  );


  or
  g570
  (
    n679,
    n351,
    n363
  );


  xnor
  g571
  (
    KeyWire_0_0,
    n217,
    n227
  );


  xnor
  g572
  (
    n655,
    n373,
    n164
  );


  or
  g573
  (
    n638,
    n179,
    n328
  );


  or
  g574
  (
    n530,
    n316,
    n349
  );


  xnor
  g575
  (
    n594,
    n348,
    n193
  );


  and
  g576
  (
    n605,
    n374,
    n278
  );


  and
  g577
  (
    n677,
    n380,
    n171
  );


  xor
  g578
  (
    n616,
    n350,
    n342
  );


  nand
  g579
  (
    n548,
    n384,
    n126
  );


  nand
  g580
  (
    n472,
    n225,
    n297
  );


  nand
  g581
  (
    n517,
    n124,
    n313
  );


  xor
  g582
  (
    n426,
    n381,
    n123
  );


  nand
  g583
  (
    n545,
    n250,
    n383
  );


  and
  g584
  (
    n444,
    n354,
    n172
  );


  or
  g585
  (
    n646,
    n299,
    n156
  );


  nand
  g586
  (
    n447,
    n359,
    n165
  );


  nand
  g587
  (
    n669,
    n276,
    n364
  );


  or
  g588
  (
    n420,
    n385,
    n348
  );


  and
  g589
  (
    n450,
    n194,
    n181
  );


  nand
  g590
  (
    n500,
    n336,
    n372
  );


  xnor
  g591
  (
    n611,
    n326,
    n205
  );


  xnor
  g592
  (
    n574,
    n248,
    n347
  );


  nand
  g593
  (
    n537,
    n344,
    n374
  );


  nor
  g594
  (
    n492,
    n366,
    n331
  );


  nand
  g595
  (
    n497,
    n358,
    n303
  );


  or
  g596
  (
    n495,
    n372,
    n379
  );


  xor
  g597
  (
    n641,
    n190,
    n293
  );


  nand
  g598
  (
    n624,
    n348,
    n175
  );


  nand
  g599
  (
    n442,
    n341,
    n352
  );


  or
  g600
  (
    n649,
    n283,
    n23
  );


  and
  g601
  (
    n644,
    n162,
    n21
  );


  nor
  g602
  (
    n417,
    n342,
    n346
  );


  or
  g603
  (
    n613,
    n387,
    n375
  );


  and
  g604
  (
    n465,
    n373,
    n365
  );


  xor
  g605
  (
    n666,
    n152,
    n358
  );


  xor
  g606
  (
    n675,
    n110,
    n327
  );


  nor
  g607
  (
    n476,
    n195,
    n337
  );


  nand
  g608
  (
    n456,
    n335,
    n200
  );


  xor
  g609
  (
    n560,
    n285,
    n168
  );


  nand
  g610
  (
    n494,
    n318,
    n159
  );


  xor
  g611
  (
    n591,
    n305,
    n265
  );


  xnor
  g612
  (
    n602,
    n176,
    n148
  );


  or
  g613
  (
    n526,
    n365,
    n345
  );


  nand
  g614
  (
    n503,
    n25,
    n275
  );


  and
  g615
  (
    n504,
    n188,
    n304
  );


  nor
  g616
  (
    n459,
    n383,
    n260
  );


  xor
  g617
  (
    n443,
    n161,
    n324
  );


  nor
  g618
  (
    n455,
    n378,
    n196
  );


  xor
  g619
  (
    n661,
    n339,
    n383
  );


  nor
  g620
  (
    n667,
    n374,
    n350
  );


  and
  g621
  (
    n606,
    n258,
    n212
  );


  xnor
  g622
  (
    n567,
    n340,
    n343
  );


  xnor
  g623
  (
    n674,
    n182,
    n362
  );


  or
  g624
  (
    n570,
    n300,
    n215
  );


  and
  g625
  (
    n656,
    n385,
    n206
  );


  xnor
  g626
  (
    n479,
    n271,
    n346
  );


  xor
  g627
  (
    n474,
    n370,
    n344
  );


  xor
  g628
  (
    n582,
    n382,
    n367
  );


  and
  g629
  (
    n636,
    n356,
    n163
  );


  nand
  g630
  (
    n511,
    n269,
    n216
  );


  xor
  g631
  (
    n654,
    n352,
    n306
  );


  nand
  g632
  (
    n488,
    n254,
    n367
  );


  nor
  g633
  (
    n542,
    n369,
    n295
  );


  nand
  g634
  (
    n487,
    n373,
    n349
  );


  xnor
  g635
  (
    n424,
    n239,
    n25
  );


  xor
  g636
  (
    n486,
    n377,
    n204
  );


  and
  g637
  (
    n672,
    n178,
    n184
  );


  and
  g638
  (
    n664,
    n351,
    n359
  );


  and
  g639
  (
    n535,
    n246,
    n256
  );


  xnor
  g640
  (
    n468,
    n187,
    n115
  );


  nand
  g641
  (
    n498,
    n242,
    n23
  );


  and
  g642
  (
    n559,
    n376,
    n339
  );


  xnor
  g643
  (
    n452,
    n333,
    n360
  );


  nand
  g644
  (
    n578,
    n380,
    n310
  );


  nor
  g645
  (
    KeyWire_0_25,
    n21,
    n173
  );


  xnor
  g646
  (
    n598,
    n384,
    n24
  );


  xor
  g647
  (
    n671,
    n372,
    n208
  );


  nor
  g648
  (
    n552,
    n302,
    n368
  );


  xnor
  g649
  (
    n673,
    n221,
    n387
  );


  nor
  g650
  (
    n565,
    n343,
    n137
  );


  or
  g651
  (
    n642,
    n329,
    n155
  );


  or
  g652
  (
    n436,
    n330,
    n361
  );


  xnor
  g653
  (
    n454,
    n382,
    n287
  );


  xnor
  g654
  (
    n650,
    n338,
    n371
  );


  buf
  g655
  (
    n686,
    n422
  );


  not
  g656
  (
    n687,
    n106
  );


  buf
  g657
  (
    n690,
    n105
  );


  not
  g658
  (
    n694,
    n103
  );


  buf
  g659
  (
    n695,
    n420
  );


  buf
  g660
  (
    n691,
    n417
  );


  buf
  g661
  (
    n696,
    n103
  );


  buf
  g662
  (
    n692,
    n104
  );


  buf
  g663
  (
    n681,
    n421
  );


  not
  g664
  (
    n693,
    n106
  );


  and
  g665
  (
    n684,
    n430,
    n426
  );


  xor
  g666
  (
    n688,
    n415,
    n104,
    n106,
    n428
  );


  xor
  g667
  (
    n683,
    n105,
    n424,
    n418,
    n416
  );


  xnor
  g668
  (
    n682,
    n427,
    n423,
    n103
  );


  xnor
  g669
  (
    n689,
    n425,
    n429,
    n419,
    n106
  );


  nand
  g670
  (
    n685,
    n104,
    n105
  );


  xor
  g671
  (
    n699,
    n388,
    n388,
    n391,
    n687
  );


  or
  g672
  (
    n698,
    n682,
    n394,
    n689
  );


  nand
  g673
  (
    n705,
    n390,
    n395,
    n393,
    n681
  );


  nor
  g674
  (
    n697,
    n392,
    n396
  );


  or
  g675
  (
    n708,
    n390,
    n392,
    n394,
    n685
  );


  or
  g676
  (
    n704,
    n389,
    n388,
    n683,
    n686
  );


  or
  g677
  (
    n707,
    n393,
    n395,
    n389,
    n391
  );


  or
  g678
  (
    KeyWire_0_26,
    n395,
    n692,
    n390
  );


  xor
  g679
  (
    n701,
    n394,
    n389,
    n690,
    n691
  );


  or
  g680
  (
    n703,
    n396,
    n391,
    n389,
    n392
  );


  xor
  g681
  (
    n706,
    n688,
    n393,
    n388,
    n391
  );


  or
  g682
  (
    n700,
    n684,
    n392,
    n395,
    n393
  );


  not
  g683
  (
    n716,
    n703
  );


  buf
  g684
  (
    n712,
    n700
  );


  buf
  g685
  (
    n719,
    n432
  );


  buf
  g686
  (
    n713,
    n437
  );


  not
  g687
  (
    n715,
    n704
  );


  buf
  g688
  (
    n714,
    n434
  );


  not
  g689
  (
    n710,
    n702
  );


  buf
  g690
  (
    n718,
    n703
  );


  nor
  g691
  (
    n709,
    n703,
    n436
  );


  nand
  g692
  (
    n717,
    n698,
    n431,
    n433,
    n703
  );


  and
  g693
  (
    n711,
    n701,
    n697,
    n435,
    n699
  );


  nand
  g694
  (
    n721,
    n717,
    n718,
    n715,
    n439
  );


  or
  g695
  (
    n722,
    n397,
    n467,
    n715,
    n480
  );


  nand
  g696
  (
    n728,
    n469,
    n455,
    n463,
    n495
  );


  nor
  g697
  (
    n727,
    n494,
    n714,
    n474,
    n695
  );


  and
  g698
  (
    n741,
    n718,
    n696,
    n484,
    n496
  );


  or
  g699
  (
    n731,
    n486,
    n397,
    n693,
    n466
  );


  nand
  g700
  (
    n744,
    n460,
    n461,
    n452,
    n696
  );


  nand
  g701
  (
    n742,
    n473,
    n447,
    n481,
    n454
  );


  xor
  g702
  (
    n736,
    n451,
    n438,
    n695,
    n499
  );


  nand
  g703
  (
    n735,
    n710,
    n483,
    n711,
    n493
  );


  xor
  g704
  (
    n723,
    n712,
    n716,
    n445,
    n492
  );


  xnor
  g705
  (
    n726,
    n716,
    n446,
    n397,
    n695
  );


  nand
  g706
  (
    n746,
    n458,
    n465,
    n471,
    n468
  );


  or
  g707
  (
    n743,
    n714,
    n478,
    n476,
    n497
  );


  xnor
  g708
  (
    n720,
    n449,
    n489,
    n444,
    n490
  );


  nand
  g709
  (
    n734,
    n470,
    n715,
    n718
  );


  and
  g710
  (
    n739,
    n503,
    n717,
    n464,
    n716
  );


  xnor
  g711
  (
    n729,
    n448,
    n443,
    n716,
    n479
  );


  nand
  g712
  (
    n732,
    n456,
    n482,
    n718,
    n453
  );


  xor
  g713
  (
    n733,
    n488,
    n397,
    n472,
    n440
  );


  nor
  g714
  (
    n725,
    n477,
    n450,
    n717,
    n696
  );


  nand
  g715
  (
    n738,
    n502,
    n462,
    n709,
    n719
  );


  xnor
  g716
  (
    n745,
    n694,
    n719,
    n504,
    n713
  );


  xor
  g717
  (
    n740,
    n459,
    n717,
    n719,
    n457
  );


  and
  g718
  (
    n730,
    n696,
    n441,
    n475,
    n719
  );


  xor
  g719
  (
    n737,
    n487,
    n695,
    n500,
    n498
  );


  xor
  g720
  (
    n724,
    n501,
    n485,
    n442,
    n491
  );


  not
  g721
  (
    n749,
    n726
  );


  buf
  g722
  (
    n755,
    n729
  );


  buf
  g723
  (
    n753,
    n736
  );


  buf
  g724
  (
    n763,
    n731
  );


  buf
  g725
  (
    n751,
    n733
  );


  not
  g726
  (
    n762,
    n721
  );


  buf
  g727
  (
    n758,
    n723
  );


  not
  g728
  (
    n747,
    n725
  );


  not
  g729
  (
    n764,
    n734
  );


  buf
  g730
  (
    n750,
    n738
  );


  not
  g731
  (
    n757,
    n727
  );


  buf
  g732
  (
    n761,
    n735
  );


  buf
  g733
  (
    n760,
    n728
  );


  buf
  g734
  (
    n754,
    n732
  );


  not
  g735
  (
    n756,
    n737
  );


  buf
  g736
  (
    n748,
    n722
  );


  not
  g737
  (
    KeyWire_0_30,
    n724
  );


  buf
  g738
  (
    n752,
    n730
  );


  not
  g739
  (
    n784,
    n761
  );


  buf
  g740
  (
    n801,
    n761
  );


  buf
  g741
  (
    n777,
    n401
  );


  not
  g742
  (
    n770,
    n757
  );


  buf
  g743
  (
    n783,
    n763
  );


  not
  g744
  (
    n790,
    n760
  );


  not
  g745
  (
    n788,
    n758
  );


  buf
  g746
  (
    n798,
    n753
  );


  not
  g747
  (
    n778,
    n402
  );


  buf
  g748
  (
    n772,
    n749
  );


  not
  g749
  (
    n773,
    n757
  );


  buf
  g750
  (
    n774,
    n747
  );


  not
  g751
  (
    n791,
    n401
  );


  buf
  g752
  (
    n765,
    n400
  );


  buf
  g753
  (
    n793,
    n398
  );


  xnor
  g754
  (
    n781,
    n756,
    n751,
    n760
  );


  nor
  g755
  (
    n787,
    n752,
    n752,
    n401,
    n750
  );


  nand
  g756
  (
    n794,
    n753,
    n741,
    n399,
    n760
  );


  xor
  g757
  (
    n767,
    n759,
    n763,
    n758,
    n750
  );


  or
  g758
  (
    n768,
    n749,
    n754,
    n758,
    n750
  );


  or
  g759
  (
    n776,
    n762,
    n506,
    n513,
    n756
  );


  or
  g760
  (
    n775,
    n747,
    n756,
    n402,
    n752
  );


  and
  g761
  (
    n771,
    n747,
    n753,
    n754,
    n761
  );


  nor
  g762
  (
    n797,
    n758,
    n514,
    n743,
    n753
  );


  xnor
  g763
  (
    n766,
    n742,
    n401,
    n755,
    n507
  );


  or
  g764
  (
    n789,
    n762,
    n759,
    n739
  );


  nand
  g765
  (
    n802,
    n748,
    n763,
    n751,
    n402
  );


  or
  g766
  (
    n799,
    n755,
    n398,
    n403,
    n509
  );


  and
  g767
  (
    n769,
    n761,
    n755,
    n754
  );


  nand
  g768
  (
    n792,
    n752,
    n750,
    n400,
    n762
  );


  xnor
  g769
  (
    n782,
    n511,
    n400,
    n749,
    n505
  );


  xor
  g770
  (
    n779,
    n740,
    n508,
    n398,
    n402
  );


  or
  g771
  (
    n786,
    n751,
    n399,
    n756,
    n763
  );


  nor
  g772
  (
    n785,
    n510,
    n512,
    n398,
    n747
  );


  nand
  g773
  (
    n795,
    n754,
    n760,
    n748,
    n762
  );


  xnor
  g774
  (
    n800,
    n403,
    n399,
    n759
  );


  or
  g775
  (
    n780,
    n748,
    n757,
    n403,
    n751
  );


  xnor
  g776
  (
    n796,
    n400,
    n748,
    n749,
    n757
  );


  buf
  g777
  (
    n803,
    n766
  );


  and
  g778
  (
    n804,
    n744,
    n746,
    n765,
    n745
  );


  or
  g779
  (
    n805,
    n803,
    n764
  );


  not
  g780
  (
    n807,
    n805
  );


  not
  g781
  (
    n806,
    n805
  );


  buf
  g782
  (
    n810,
    n516
  );


  not
  g783
  (
    n812,
    n804
  );


  not
  g784
  (
    n811,
    n518
  );


  xnor
  g785
  (
    n809,
    n515,
    n807
  );


  nand
  g786
  (
    n808,
    n806,
    n807,
    n517
  );


  buf
  g787
  (
    n819,
    n810
  );


  buf
  g788
  (
    n816,
    n809
  );


  not
  g789
  (
    n815,
    n809
  );


  buf
  g790
  (
    n818,
    n808
  );


  buf
  g791
  (
    n814,
    n808
  );


  buf
  g792
  (
    n820,
    n810
  );


  not
  g793
  (
    n817,
    n808
  );


  not
  g794
  (
    n821,
    n809
  );


  buf
  g795
  (
    n822,
    n808
  );


  buf
  g796
  (
    n813,
    n809
  );


  xnor
  g797
  (
    n828,
    n818,
    n523,
    n815,
    n821
  );


  nor
  g798
  (
    n824,
    n536,
    n545,
    n534,
    n544
  );


  xor
  g799
  (
    n825,
    n535,
    n532,
    n531,
    n541
  );


  or
  g800
  (
    n829,
    n526,
    n537,
    n521,
    n529
  );


  nand
  g801
  (
    n826,
    n816,
    n530,
    n817,
    n539
  );


  and
  g802
  (
    n831,
    n520,
    n819,
    n528,
    n814
  );


  xnor
  g803
  (
    n830,
    n527,
    n540,
    n522,
    n820
  );


  nand
  g804
  (
    n827,
    n525,
    n524,
    n822,
    n542
  );


  or
  g805
  (
    n823,
    n519,
    n533,
    n543,
    n538
  );


  not
  g806
  (
    n837,
    n831
  );


  not
  g807
  (
    n866,
    n823
  );


  not
  g808
  (
    n863,
    n825
  );


  not
  g809
  (
    n834,
    n553
  );


  buf
  g810
  (
    n845,
    n775
  );


  buf
  g811
  (
    n852,
    n826
  );


  buf
  g812
  (
    n846,
    n812
  );


  buf
  g813
  (
    n840,
    n550
  );


  not
  g814
  (
    n857,
    n829
  );


  not
  g815
  (
    n851,
    n830
  );


  buf
  g816
  (
    n865,
    n552
  );


  not
  g817
  (
    n833,
    n811
  );


  buf
  g818
  (
    n858,
    n824
  );


  buf
  g819
  (
    n838,
    n825
  );


  not
  g820
  (
    n835,
    n551
  );


  not
  g821
  (
    n848,
    n811
  );


  not
  g822
  (
    n855,
    n824
  );


  buf
  g823
  (
    n849,
    n810
  );


  not
  g824
  (
    n844,
    n823
  );


  buf
  g825
  (
    n843,
    n829
  );


  buf
  g826
  (
    n847,
    n812
  );


  not
  g827
  (
    n867,
    n767
  );


  not
  g828
  (
    n856,
    n549
  );


  buf
  g829
  (
    n854,
    n811
  );


  buf
  g830
  (
    n861,
    n810
  );


  not
  g831
  (
    n864,
    n827
  );


  xnor
  g832
  (
    n862,
    n823,
    n831
  );


  xnor
  g833
  (
    n850,
    n548,
    n824,
    n768,
    n547
  );


  xnor
  g834
  (
    n841,
    n826,
    n830,
    n827,
    n825
  );


  and
  g835
  (
    n860,
    n811,
    n824,
    n826,
    n825
  );


  nor
  g836
  (
    n853,
    n831,
    n772,
    n546,
    n829
  );


  xor
  g837
  (
    n832,
    n831,
    n828,
    n812,
    n830
  );


  nor
  g838
  (
    n842,
    n704,
    n830,
    n829,
    n827
  );


  nand
  g839
  (
    n839,
    n769,
    n774,
    n773,
    n812
  );


  or
  g840
  (
    n836,
    n826,
    n828,
    n770
  );


  nor
  g841
  (
    n859,
    n771,
    n823,
    n827,
    n828
  );


  buf
  g842
  (
    n879,
    n777
  );


  buf
  g843
  (
    KeyWire_0_11,
    n848
  );


  not
  g844
  (
    n926,
    n867
  );


  not
  g845
  (
    n909,
    n864
  );


  buf
  g846
  (
    n976,
    n834
  );


  not
  g847
  (
    n987,
    n847
  );


  buf
  g848
  (
    n941,
    n866
  );


  buf
  g849
  (
    n882,
    n849
  );


  not
  g850
  (
    n903,
    n861
  );


  not
  g851
  (
    n982,
    n708
  );


  buf
  g852
  (
    n991,
    n832
  );


  not
  g853
  (
    n955,
    n841
  );


  not
  g854
  (
    n930,
    n705
  );


  not
  g855
  (
    n887,
    n863
  );


  buf
  g856
  (
    n888,
    n572
  );


  not
  g857
  (
    n949,
    n839
  );


  not
  g858
  (
    n884,
    n565
  );


  not
  g859
  (
    n914,
    n866
  );


  not
  g860
  (
    n973,
    n705
  );


  buf
  g861
  (
    n996,
    n708
  );


  buf
  g862
  (
    n872,
    n858
  );


  buf
  g863
  (
    n871,
    n836
  );


  not
  g864
  (
    n934,
    n834
  );


  buf
  g865
  (
    n947,
    n845
  );


  buf
  g866
  (
    n883,
    n856
  );


  buf
  g867
  (
    n945,
    n859
  );


  buf
  g868
  (
    n998,
    n861
  );


  not
  g869
  (
    n951,
    n854
  );


  buf
  g870
  (
    n877,
    n846
  );


  buf
  g871
  (
    n969,
    n834
  );


  buf
  g872
  (
    n894,
    n559
  );


  not
  g873
  (
    n1002,
    n852
  );


  not
  g874
  (
    n965,
    n837
  );


  not
  g875
  (
    n876,
    n866
  );


  buf
  g876
  (
    n978,
    n863
  );


  buf
  g877
  (
    n992,
    n849
  );


  buf
  g878
  (
    n921,
    n706
  );


  buf
  g879
  (
    n964,
    n850
  );


  buf
  g880
  (
    n920,
    n574
  );


  buf
  g881
  (
    n1003,
    n706
  );


  not
  g882
  (
    n923,
    n782
  );


  buf
  g883
  (
    n886,
    n857
  );


  not
  g884
  (
    n984,
    n569
  );


  not
  g885
  (
    n891,
    n837
  );


  not
  g886
  (
    n977,
    n844
  );


  buf
  g887
  (
    n1009,
    n832
  );


  buf
  g888
  (
    n927,
    n568
  );


  buf
  g889
  (
    n988,
    n849
  );


  not
  g890
  (
    n972,
    n860
  );


  buf
  g891
  (
    n939,
    n851
  );


  not
  g892
  (
    KeyWire_0_9,
    n851
  );


  buf
  g893
  (
    n1000,
    n854
  );


  not
  g894
  (
    n997,
    n848
  );


  buf
  g895
  (
    n1004,
    n859
  );


  buf
  g896
  (
    n981,
    n862
  );


  not
  g897
  (
    n980,
    n707
  );


  buf
  g898
  (
    n986,
    n840
  );


  buf
  g899
  (
    n954,
    n858
  );


  not
  g900
  (
    n875,
    n833
  );


  not
  g901
  (
    n916,
    n832
  );


  buf
  g902
  (
    n904,
    n845
  );


  not
  g903
  (
    n924,
    n554
  );


  buf
  g904
  (
    n898,
    n566
  );


  not
  g905
  (
    n943,
    n853
  );


  not
  g906
  (
    n975,
    n865
  );


  buf
  g907
  (
    n878,
    n570
  );


  buf
  g908
  (
    n967,
    n707
  );


  not
  g909
  (
    n1011,
    n865
  );


  buf
  g910
  (
    n942,
    n861
  );


  buf
  g911
  (
    n966,
    n837
  );


  buf
  g912
  (
    n918,
    n864
  );


  not
  g913
  (
    n881,
    n846
  );


  not
  g914
  (
    n953,
    n776
  );


  not
  g915
  (
    n938,
    n833
  );


  buf
  g916
  (
    n912,
    n846
  );


  not
  g917
  (
    n985,
    n555
  );


  buf
  g918
  (
    n913,
    n844
  );


  buf
  g919
  (
    n994,
    n834
  );


  buf
  g920
  (
    n910,
    n708
  );


  not
  g921
  (
    n963,
    n833
  );


  not
  g922
  (
    n962,
    n707
  );


  buf
  g923
  (
    n873,
    n849
  );


  buf
  g924
  (
    n897,
    n842
  );


  buf
  g925
  (
    n911,
    n844
  );


  not
  g926
  (
    n957,
    n857
  );


  buf
  g927
  (
    n959,
    n840
  );


  buf
  g928
  (
    n915,
    n856
  );


  buf
  g929
  (
    n922,
    n856
  );


  not
  g930
  (
    n907,
    n838
  );


  buf
  g931
  (
    n1006,
    n859
  );


  buf
  g932
  (
    n905,
    n843
  );


  not
  g933
  (
    n940,
    n850
  );


  buf
  g934
  (
    n919,
    n706
  );


  not
  g935
  (
    n956,
    n706
  );


  not
  g936
  (
    n958,
    n705
  );


  buf
  g937
  (
    n892,
    n867
  );


  buf
  g938
  (
    n979,
    n838
  );


  buf
  g939
  (
    n890,
    n863
  );


  buf
  g940
  (
    n1007,
    n558
  );


  not
  g941
  (
    n989,
    n864
  );


  buf
  g942
  (
    n932,
    n845
  );


  buf
  g943
  (
    n995,
    n840
  );


  buf
  g944
  (
    n928,
    n842
  );


  buf
  g945
  (
    n908,
    n561
  );


  not
  g946
  (
    n974,
    n847
  );


  buf
  g947
  (
    n906,
    n835
  );


  not
  g948
  (
    n889,
    n858
  );


  buf
  g949
  (
    n899,
    n864
  );


  not
  g950
  (
    n870,
    n846
  );


  buf
  g951
  (
    n993,
    n780
  );


  buf
  g952
  (
    n895,
    n854
  );


  not
  g953
  (
    n874,
    n865
  );


  not
  g954
  (
    n1010,
    n841
  );


  buf
  g955
  (
    n885,
    n839
  );


  not
  g956
  (
    n983,
    n852
  );


  not
  g957
  (
    n970,
    n844
  );


  buf
  g958
  (
    n902,
    n836
  );


  buf
  g959
  (
    n961,
    n860
  );


  buf
  g960
  (
    n971,
    n832
  );


  not
  g961
  (
    n968,
    n865
  );


  buf
  g962
  (
    n893,
    n835
  );


  nor
  g963
  (
    n1005,
    n867,
    n839,
    n843
  );


  nor
  g964
  (
    n880,
    n851,
    n855,
    n845
  );


  nand
  g965
  (
    n960,
    n857,
    n567,
    n847
  );


  nor
  g966
  (
    n1008,
    n848,
    n853,
    n862
  );


  or
  g967
  (
    n952,
    n858,
    n835,
    n850
  );


  nand
  g968
  (
    n1001,
    n838,
    n843,
    n781
  );


  nor
  g969
  (
    n990,
    n563,
    n855,
    n835
  );


  nor
  g970
  (
    n999,
    n851,
    n708,
    n850
  );


  xor
  g971
  (
    n936,
    n564,
    n778,
    n852
  );


  xnor
  g972
  (
    n931,
    n571,
    n840,
    n556
  );


  xor
  g973
  (
    n896,
    n860,
    n862,
    n843
  );


  nor
  g974
  (
    n917,
    n837,
    n842,
    n855
  );


  xnor
  g975
  (
    n901,
    n847,
    n573,
    n836
  );


  xor
  g976
  (
    n933,
    n861,
    n562,
    n707
  );


  nand
  g977
  (
    n937,
    n705,
    n867,
    n855
  );


  and
  g978
  (
    n869,
    n704,
    n856,
    n842
  );


  xor
  g979
  (
    n948,
    n857,
    n848,
    n853
  );


  or
  g980
  (
    n929,
    n862,
    n779,
    n841
  );


  xnor
  g981
  (
    n946,
    n704,
    n838,
    n852
  );


  nor
  g982
  (
    n900,
    n854,
    n859,
    n836
  );


  nor
  g983
  (
    n950,
    n860,
    n839,
    n560
  );


  xor
  g984
  (
    n944,
    n557,
    n863,
    n866
  );


  nand
  g985
  (
    n925,
    n841,
    n833,
    n853
  );


  not
  g986
  (
    n1405,
    n895
  );


  not
  g987
  (
    n1053,
    n880
  );


  not
  g988
  (
    n1439,
    n917
  );


  buf
  g989
  (
    n1332,
    n900
  );


  not
  g990
  (
    n1071,
    n976
  );


  not
  g991
  (
    n1432,
    n873
  );


  not
  g992
  (
    n1016,
    n913
  );


  not
  g993
  (
    n1233,
    n969
  );


  not
  g994
  (
    n1401,
    n884
  );


  not
  g995
  (
    n1171,
    n931
  );


  buf
  g996
  (
    n1040,
    n872
  );


  not
  g997
  (
    n1074,
    n929
  );


  buf
  g998
  (
    n1279,
    n922
  );


  not
  g999
  (
    n1065,
    n786
  );


  buf
  g1000
  (
    n1215,
    n930
  );


  not
  g1001
  (
    n1093,
    n966
  );


  buf
  g1002
  (
    n1387,
    n901
  );


  not
  g1003
  (
    n1273,
    n891
  );


  buf
  g1004
  (
    n1277,
    n896
  );


  buf
  g1005
  (
    n1120,
    n890
  );


  buf
  g1006
  (
    KeyWire_0_14,
    n976
  );


  buf
  g1007
  (
    n1445,
    n955
  );


  not
  g1008
  (
    n1404,
    n887
  );


  buf
  g1009
  (
    n1292,
    n784
  );


  not
  g1010
  (
    n1343,
    n918
  );


  not
  g1011
  (
    n1235,
    n975
  );


  buf
  g1012
  (
    n1122,
    n947
  );


  buf
  g1013
  (
    n1386,
    n870
  );


  buf
  g1014
  (
    n1348,
    n974
  );


  buf
  g1015
  (
    n1360,
    n906
  );


  buf
  g1016
  (
    n1399,
    n890
  );


  not
  g1017
  (
    n1059,
    n941
  );


  not
  g1018
  (
    n1443,
    n885
  );


  not
  g1019
  (
    n1154,
    n916
  );


  buf
  g1020
  (
    n1186,
    n963
  );


  not
  g1021
  (
    n1448,
    n919
  );


  buf
  g1022
  (
    n1114,
    n905
  );


  not
  g1023
  (
    n1018,
    n914
  );


  not
  g1024
  (
    n1052,
    n954
  );


  buf
  g1025
  (
    n1376,
    n960
  );


  not
  g1026
  (
    n1125,
    n890
  );


  buf
  g1027
  (
    n1103,
    n919
  );


  not
  g1028
  (
    n1287,
    n921
  );


  not
  g1029
  (
    n1095,
    n927
  );


  not
  g1030
  (
    n1340,
    n912
  );


  not
  g1031
  (
    n1198,
    n951
  );


  not
  g1032
  (
    n1226,
    n930
  );


  buf
  g1033
  (
    n1364,
    n916
  );


  buf
  g1034
  (
    n1222,
    n930
  );


  buf
  g1035
  (
    n1159,
    n957
  );


  not
  g1036
  (
    n1436,
    n891
  );


  buf
  g1037
  (
    n1110,
    n879
  );


  not
  g1038
  (
    n1419,
    n955
  );


  buf
  g1039
  (
    n1179,
    n889
  );


  buf
  g1040
  (
    n1423,
    n948
  );


  buf
  g1041
  (
    n1308,
    n881
  );


  buf
  g1042
  (
    n1409,
    n949
  );


  not
  g1043
  (
    n1070,
    n880
  );


  buf
  g1044
  (
    n1144,
    n892
  );


  buf
  g1045
  (
    n1037,
    n936
  );


  buf
  g1046
  (
    n1310,
    n959
  );


  buf
  g1047
  (
    n1377,
    n969
  );


  not
  g1048
  (
    n1145,
    n791
  );


  buf
  g1049
  (
    n1341,
    n901
  );


  not
  g1050
  (
    n1265,
    n968
  );


  buf
  g1051
  (
    n1302,
    n909
  );


  buf
  g1052
  (
    n1101,
    n937
  );


  buf
  g1053
  (
    n1225,
    n899
  );


  not
  g1054
  (
    n1098,
    n911
  );


  buf
  g1055
  (
    n1282,
    n912
  );


  not
  g1056
  (
    n1418,
    n935
  );


  buf
  g1057
  (
    n1355,
    n925
  );


  buf
  g1058
  (
    n1437,
    n953
  );


  not
  g1059
  (
    n1421,
    n876
  );


  buf
  g1060
  (
    n1441,
    n941
  );


  not
  g1061
  (
    n1150,
    n931
  );


  buf
  g1062
  (
    n1396,
    n889
  );


  buf
  g1063
  (
    n1232,
    n908
  );


  buf
  g1064
  (
    n1061,
    n790
  );


  not
  g1065
  (
    n1172,
    n896
  );


  buf
  g1066
  (
    n1251,
    n949
  );


  not
  g1067
  (
    n1047,
    n796
  );


  not
  g1068
  (
    n1076,
    n877
  );


  not
  g1069
  (
    n1033,
    n907
  );


  buf
  g1070
  (
    n1391,
    n897
  );


  not
  g1071
  (
    n1178,
    n971
  );


  buf
  g1072
  (
    n1353,
    n964
  );


  buf
  g1073
  (
    n1211,
    n917
  );


  buf
  g1074
  (
    n1240,
    n934
  );


  not
  g1075
  (
    n1081,
    n872
  );


  not
  g1076
  (
    n1109,
    n974
  );


  buf
  g1077
  (
    n1088,
    n975
  );


  not
  g1078
  (
    n1392,
    n905
  );


  not
  g1079
  (
    n1147,
    n944
  );


  not
  g1080
  (
    n1393,
    n918
  );


  buf
  g1081
  (
    n1077,
    n945
  );


  buf
  g1082
  (
    n1176,
    n891
  );


  buf
  g1083
  (
    n1424,
    n962
  );


  not
  g1084
  (
    n1256,
    n875
  );


  buf
  g1085
  (
    n1291,
    n952
  );


  not
  g1086
  (
    n1119,
    n922
  );


  buf
  g1087
  (
    n1136,
    n976
  );


  not
  g1088
  (
    n1371,
    n871
  );


  not
  g1089
  (
    n1411,
    n970
  );


  not
  g1090
  (
    n1168,
    n940
  );


  buf
  g1091
  (
    n1135,
    n920
  );


  buf
  g1092
  (
    n1347,
    n951
  );


  buf
  g1093
  (
    n1227,
    n924
  );


  not
  g1094
  (
    n1152,
    n879
  );


  not
  g1095
  (
    n1231,
    n868
  );


  not
  g1096
  (
    n1362,
    n883
  );


  not
  g1097
  (
    n1415,
    n937
  );


  not
  g1098
  (
    n1045,
    n964
  );


  not
  g1099
  (
    n1300,
    n908
  );


  buf
  g1100
  (
    n1202,
    n893
  );


  buf
  g1101
  (
    n1158,
    n938
  );


  buf
  g1102
  (
    n1034,
    n885
  );


  buf
  g1103
  (
    n1189,
    n932
  );


  buf
  g1104
  (
    n1163,
    n920
  );


  buf
  g1105
  (
    n1299,
    n944
  );


  not
  g1106
  (
    n1195,
    n967
  );


  buf
  g1107
  (
    n1280,
    n874
  );


  not
  g1108
  (
    n1124,
    n933
  );


  buf
  g1109
  (
    n1048,
    n950
  );


  not
  g1110
  (
    n1126,
    n946
  );


  buf
  g1111
  (
    n1138,
    n920
  );


  buf
  g1112
  (
    n1284,
    n912
  );


  not
  g1113
  (
    n1293,
    n897
  );


  not
  g1114
  (
    n1151,
    n954
  );


  buf
  g1115
  (
    n1434,
    n868
  );


  not
  g1116
  (
    n1329,
    n943
  );


  not
  g1117
  (
    n1191,
    n802
  );


  buf
  g1118
  (
    n1378,
    n945
  );


  not
  g1119
  (
    n1260,
    n928
  );


  buf
  g1120
  (
    n1236,
    n961
  );


  buf
  g1121
  (
    n1400,
    n868
  );


  buf
  g1122
  (
    n1449,
    n898
  );


  not
  g1123
  (
    n1199,
    n882
  );


  buf
  g1124
  (
    n1438,
    n943
  );


  buf
  g1125
  (
    n1013,
    n886
  );


  not
  g1126
  (
    n1352,
    n909
  );


  not
  g1127
  (
    n1116,
    n950
  );


  not
  g1128
  (
    n1139,
    n913
  );


  buf
  g1129
  (
    n1219,
    n879
  );


  not
  g1130
  (
    n1181,
    n876
  );


  buf
  g1131
  (
    n1369,
    n925
  );


  not
  g1132
  (
    n1406,
    n959
  );


  not
  g1133
  (
    n1326,
    n932
  );


  not
  g1134
  (
    n1257,
    n869
  );


  buf
  g1135
  (
    n1224,
    n914
  );


  not
  g1136
  (
    n1366,
    n937
  );


  not
  g1137
  (
    n1204,
    n799
  );


  buf
  g1138
  (
    n1363,
    n893
  );


  not
  g1139
  (
    n1241,
    n918
  );


  buf
  g1140
  (
    n1270,
    n939
  );


  not
  g1141
  (
    n1111,
    n962
  );


  buf
  g1142
  (
    n1177,
    n966
  );


  buf
  g1143
  (
    n1313,
    n902
  );


  not
  g1144
  (
    n1056,
    n875
  );


  not
  g1145
  (
    n1019,
    n972
  );


  buf
  g1146
  (
    n1155,
    n883
  );


  not
  g1147
  (
    n1373,
    n938
  );


  buf
  g1148
  (
    n1078,
    n942
  );


  not
  g1149
  (
    n1267,
    n958
  );


  not
  g1150
  (
    KeyWire_0_4,
    n919
  );


  buf
  g1151
  (
    n1022,
    n910
  );


  not
  g1152
  (
    n1190,
    n957
  );


  not
  g1153
  (
    n1440,
    n881
  );


  not
  g1154
  (
    n1390,
    n902
  );


  buf
  g1155
  (
    n1239,
    n873
  );


  not
  g1156
  (
    n1200,
    n928
  );


  not
  g1157
  (
    n1068,
    n902
  );


  not
  g1158
  (
    n1220,
    n878
  );


  not
  g1159
  (
    n1294,
    n911
  );


  buf
  g1160
  (
    n1201,
    n975
  );


  buf
  g1161
  (
    n1115,
    n946
  );


  buf
  g1162
  (
    n1254,
    n900
  );


  not
  g1163
  (
    n1160,
    n888
  );


  buf
  g1164
  (
    KeyWire_0_16,
    n788
  );


  buf
  g1165
  (
    n1237,
    n932
  );


  not
  g1166
  (
    n1245,
    n957
  );


  not
  g1167
  (
    n1407,
    n960
  );


  not
  g1168
  (
    n1342,
    n940
  );


  not
  g1169
  (
    n1130,
    n943
  );


  buf
  g1170
  (
    n1197,
    n800
  );


  not
  g1171
  (
    n1137,
    n949
  );


  buf
  g1172
  (
    n1031,
    n962
  );


  not
  g1173
  (
    n1205,
    n881
  );


  buf
  g1174
  (
    n1039,
    n942
  );


  not
  g1175
  (
    n1085,
    n873
  );


  buf
  g1176
  (
    n1242,
    n926
  );


  not
  g1177
  (
    n1305,
    n930
  );


  buf
  g1178
  (
    n1314,
    n894
  );


  not
  g1179
  (
    n1338,
    n960
  );


  buf
  g1180
  (
    n1425,
    n924
  );


  not
  g1181
  (
    n1261,
    n895
  );


  not
  g1182
  (
    n1249,
    n927
  );


  not
  g1183
  (
    n1266,
    n883
  );


  buf
  g1184
  (
    n1075,
    n880
  );


  buf
  g1185
  (
    KeyWire_0_22,
    n941
  );


  not
  g1186
  (
    n1167,
    n963
  );


  not
  g1187
  (
    n1134,
    n798
  );


  not
  g1188
  (
    n1107,
    n973
  );


  buf
  g1189
  (
    n1194,
    n964
  );


  buf
  g1190
  (
    n1214,
    n923
  );


  not
  g1191
  (
    n1187,
    n933
  );


  not
  g1192
  (
    n1322,
    n905
  );


  not
  g1193
  (
    n1183,
    n875
  );


  buf
  g1194
  (
    n1025,
    n887
  );


  buf
  g1195
  (
    n1028,
    n928
  );


  buf
  g1196
  (
    n1316,
    n888
  );


  buf
  g1197
  (
    n1024,
    n797
  );


  buf
  g1198
  (
    n1382,
    n899
  );


  not
  g1199
  (
    n1248,
    n909
  );


  buf
  g1200
  (
    n1062,
    n883
  );


  buf
  g1201
  (
    n1264,
    n909
  );


  not
  g1202
  (
    n1097,
    n933
  );


  not
  g1203
  (
    n1099,
    n963
  );


  buf
  g1204
  (
    n1096,
    n884
  );


  not
  g1205
  (
    KeyWire_0_13,
    n947
  );


  buf
  g1206
  (
    n1243,
    n977
  );


  buf
  g1207
  (
    n1083,
    n783
  );


  buf
  g1208
  (
    n1394,
    n926
  );


  not
  g1209
  (
    n1427,
    n892
  );


  not
  g1210
  (
    n1203,
    n917
  );


  not
  g1211
  (
    n1296,
    n878
  );


  buf
  g1212
  (
    n1223,
    n928
  );


  not
  g1213
  (
    n1327,
    n972
  );


  buf
  g1214
  (
    n1315,
    n933
  );


  not
  g1215
  (
    n1412,
    n964
  );


  buf
  g1216
  (
    n1209,
    n879
  );


  not
  g1217
  (
    n1370,
    n939
  );


  buf
  g1218
  (
    n1361,
    n896
  );


  buf
  g1219
  (
    n1351,
    n880
  );


  buf
  g1220
  (
    n1234,
    n960
  );


  buf
  g1221
  (
    n1082,
    n962
  );


  buf
  g1222
  (
    n1298,
    n907
  );


  buf
  g1223
  (
    n1323,
    n870
  );


  not
  g1224
  (
    n1311,
    n894
  );


  not
  g1225
  (
    n1238,
    n959
  );


  not
  g1226
  (
    n1131,
    n912
  );


  buf
  g1227
  (
    n1210,
    n926
  );


  buf
  g1228
  (
    n1337,
    n898
  );


  buf
  g1229
  (
    n1247,
    n886
  );


  buf
  g1230
  (
    n1417,
    n897
  );


  not
  g1231
  (
    n1356,
    n971
  );


  buf
  g1232
  (
    n1208,
    n876
  );


  buf
  g1233
  (
    n1143,
    n918
  );


  buf
  g1234
  (
    n1334,
    n904
  );


  not
  g1235
  (
    n1346,
    n888
  );


  buf
  g1236
  (
    n1108,
    n869
  );


  buf
  g1237
  (
    n1379,
    n947
  );


  buf
  g1238
  (
    n1029,
    n973
  );


  buf
  g1239
  (
    KeyWire_0_23,
    n936
  );


  buf
  g1240
  (
    n1429,
    n935
  );


  buf
  g1241
  (
    n1023,
    n900
  );


  not
  g1242
  (
    n1169,
    n936
  );


  not
  g1243
  (
    n1184,
    n954
  );


  buf
  g1244
  (
    n1193,
    n967
  );


  buf
  g1245
  (
    n1035,
    n900
  );


  not
  g1246
  (
    n1185,
    n949
  );


  buf
  g1247
  (
    n1170,
    n963
  );


  buf
  g1248
  (
    n1212,
    n952
  );


  not
  g1249
  (
    n1206,
    n938
  );


  buf
  g1250
  (
    n1258,
    n948
  );


  buf
  g1251
  (
    n1051,
    n898
  );


  buf
  g1252
  (
    n1066,
    n874
  );


  buf
  g1253
  (
    n1063,
    n914
  );


  buf
  g1254
  (
    n1207,
    n871
  );


  not
  g1255
  (
    n1057,
    n942
  );


  buf
  g1256
  (
    n1050,
    n884
  );


  not
  g1257
  (
    n1192,
    n887
  );


  not
  g1258
  (
    n1303,
    n886
  );


  buf
  g1259
  (
    n1398,
    n956
  );


  buf
  g1260
  (
    n1272,
    n878
  );


  buf
  g1261
  (
    n1344,
    n929
  );


  not
  g1262
  (
    n1149,
    n876
  );


  buf
  g1263
  (
    n1426,
    n893
  );


  not
  g1264
  (
    n1345,
    n789
  );


  buf
  g1265
  (
    n1049,
    n968
  );


  buf
  g1266
  (
    n1320,
    n870
  );


  not
  g1267
  (
    n1140,
    n921
  );


  buf
  g1268
  (
    n1244,
    n892
  );


  not
  g1269
  (
    n1067,
    n925
  );


  buf
  g1270
  (
    n1161,
    n961
  );


  buf
  g1271
  (
    n1165,
    n958
  );


  not
  g1272
  (
    n1064,
    n925
  );


  not
  g1273
  (
    n1414,
    n882
  );


  not
  g1274
  (
    n1321,
    n965
  );


  not
  g1275
  (
    n1397,
    n906
  );


  not
  g1276
  (
    n1444,
    n872
  );


  buf
  g1277
  (
    KeyWire_0_1,
    n889
  );


  buf
  g1278
  (
    n1105,
    n972
  );


  not
  g1279
  (
    n1286,
    n793
  );


  not
  g1280
  (
    n1036,
    n870
  );


  not
  g1281
  (
    n1175,
    n923
  );


  buf
  g1282
  (
    n1042,
    n946
  );


  not
  g1283
  (
    n1295,
    n955
  );


  buf
  g1284
  (
    n1044,
    n958
  );


  buf
  g1285
  (
    n1148,
    n903
  );


  not
  g1286
  (
    n1112,
    n894
  );


  not
  g1287
  (
    n1038,
    n954
  );


  buf
  g1288
  (
    n1127,
    n801
  );


  buf
  g1289
  (
    n1312,
    n795
  );


  not
  g1290
  (
    n1094,
    n881
  );


  buf
  g1291
  (
    n1281,
    n961
  );


  buf
  g1292
  (
    n1317,
    n972
  );


  not
  g1293
  (
    n1372,
    n923
  );


  not
  g1294
  (
    n1269,
    n945
  );


  not
  g1295
  (
    n1402,
    n919
  );


  not
  g1296
  (
    n1055,
    n885
  );


  buf
  g1297
  (
    n1188,
    n887
  );


  not
  g1298
  (
    n1446,
    n929
  );


  not
  g1299
  (
    n1246,
    n951
  );


  not
  g1300
  (
    n1365,
    n927
  );


  buf
  g1301
  (
    n1413,
    n902
  );


  buf
  g1302
  (
    n1278,
    n907
  );


  not
  g1303
  (
    n1420,
    n904
  );


  not
  g1304
  (
    n1174,
    n875
  );


  buf
  g1305
  (
    n1180,
    n940
  );


  buf
  g1306
  (
    n1276,
    n939
  );


  buf
  g1307
  (
    n1408,
    n965
  );


  not
  g1308
  (
    n1084,
    n913
  );


  not
  g1309
  (
    n1091,
    n889
  );


  not
  g1310
  (
    n1079,
    n976
  );


  buf
  g1311
  (
    n1389,
    n952
  );


  buf
  g1312
  (
    n1026,
    n969
  );


  not
  g1313
  (
    n1325,
    n973
  );


  not
  g1314
  (
    n1309,
    n934
  );


  buf
  g1315
  (
    n1217,
    n885
  );


  buf
  g1316
  (
    n1306,
    n974
  );


  buf
  g1317
  (
    n1021,
    n950
  );


  not
  g1318
  (
    n1173,
    n787
  );


  buf
  g1319
  (
    n1032,
    n901
  );


  not
  g1320
  (
    n1395,
    n944
  );


  buf
  g1321
  (
    n1153,
    n936
  );


  buf
  g1322
  (
    n1041,
    n794
  );


  not
  g1323
  (
    n1142,
    n898
  );


  buf
  g1324
  (
    n1403,
    n899
  );


  buf
  g1325
  (
    n1357,
    n970
  );


  not
  g1326
  (
    n1339,
    n914
  );


  not
  g1327
  (
    n1213,
    n944
  );


  not
  g1328
  (
    n1080,
    n884
  );


  buf
  g1329
  (
    n1014,
    n904
  );


  buf
  g1330
  (
    n1350,
    n882
  );


  buf
  g1331
  (
    n1388,
    n895
  );


  buf
  g1332
  (
    n1253,
    n910
  );


  buf
  g1333
  (
    n1228,
    n946
  );


  buf
  g1334
  (
    n1335,
    n961
  );


  not
  g1335
  (
    n1162,
    n897
  );


  buf
  g1336
  (
    n1072,
    n956
  );


  not
  g1337
  (
    n1087,
    n935
  );


  buf
  g1338
  (
    n1442,
    n917
  );


  not
  g1339
  (
    n1146,
    n916
  );


  buf
  g1340
  (
    KeyWire_0_21,
    n890
  );


  not
  g1341
  (
    n1090,
    n908
  );


  buf
  g1342
  (
    n1123,
    n973
  );


  not
  g1343
  (
    n1290,
    n903
  );


  buf
  g1344
  (
    n1196,
    n905
  );


  buf
  g1345
  (
    n1216,
    n957
  );


  buf
  g1346
  (
    n1289,
    n891
  );


  buf
  g1347
  (
    n1086,
    n906
  );


  not
  g1348
  (
    n1331,
    n915
  );


  not
  g1349
  (
    n1383,
    n894
  );


  buf
  g1350
  (
    n1100,
    n950
  );


  not
  g1351
  (
    n1118,
    n951
  );


  not
  g1352
  (
    n1128,
    n948
  );


  not
  g1353
  (
    n1319,
    n903
  );


  buf
  g1354
  (
    n1318,
    n974
  );


  buf
  g1355
  (
    n1030,
    n935
  );


  not
  g1356
  (
    n1447,
    n911
  );


  not
  g1357
  (
    n1330,
    n886
  );


  buf
  g1358
  (
    n1375,
    n911
  );


  not
  g1359
  (
    n1324,
    n895
  );


  not
  g1360
  (
    n1046,
    n901
  );


  buf
  g1361
  (
    n1141,
    n913
  );


  not
  g1362
  (
    n1328,
    n916
  );


  buf
  g1363
  (
    n1133,
    n921
  );


  not
  g1364
  (
    n1121,
    n948
  );


  buf
  g1365
  (
    n1435,
    n969
  );


  buf
  g1366
  (
    n1164,
    n970
  );


  not
  g1367
  (
    n1359,
    n908
  );


  buf
  g1368
  (
    n1255,
    n943
  );


  not
  g1369
  (
    n1304,
    n931
  );


  not
  g1370
  (
    n1092,
    n882
  );


  buf
  g1371
  (
    n1104,
    n924
  );


  not
  g1372
  (
    n1422,
    n924
  );


  buf
  g1373
  (
    n1182,
    n896
  );


  buf
  g1374
  (
    n1374,
    n922
  );


  buf
  g1375
  (
    n1252,
    n869
  );


  not
  g1376
  (
    n1230,
    n977
  );


  buf
  g1377
  (
    n1349,
    n910
  );


  not
  g1378
  (
    n1166,
    n968
  );


  buf
  g1379
  (
    n1054,
    n932
  );


  buf
  g1380
  (
    n1271,
    n934
  );


  not
  g1381
  (
    n1218,
    n967
  );


  buf
  g1382
  (
    n1333,
    n785
  );


  buf
  g1383
  (
    n1336,
    n868
  );


  not
  g1384
  (
    n1129,
    n575
  );


  buf
  g1385
  (
    n1431,
    n971
  );


  not
  g1386
  (
    n1381,
    n892
  );


  buf
  g1387
  (
    n1073,
    n956
  );


  not
  g1388
  (
    n1416,
    n970
  );


  buf
  g1389
  (
    n1221,
    n922
  );


  buf
  g1390
  (
    n1275,
    n966
  );


  buf
  g1391
  (
    n1060,
    n926
  );


  not
  g1392
  (
    n1027,
    n952
  );


  not
  g1393
  (
    n1043,
    n927
  );


  buf
  g1394
  (
    n1132,
    n975
  );


  buf
  g1395
  (
    n1058,
    n953
  );


  buf
  g1396
  (
    n1301,
    n956
  );


  buf
  g1397
  (
    n1307,
    n921
  );


  buf
  g1398
  (
    n1367,
    n920
  );


  buf
  g1399
  (
    n1106,
    n878
  );


  not
  g1400
  (
    n1250,
    n965
  );


  not
  g1401
  (
    n1384,
    n966
  );


  buf
  g1402
  (
    n1157,
    n792
  );


  buf
  g1403
  (
    n1288,
    n965
  );


  not
  g1404
  (
    n1102,
    n953
  );


  buf
  g1405
  (
    n1069,
    n945
  );


  not
  g1406
  (
    n1020,
    n910
  );


  not
  g1407
  (
    n1354,
    n904
  );


  buf
  g1408
  (
    n1113,
    n937
  );


  buf
  g1409
  (
    n1017,
    n934
  );


  buf
  g1410
  (
    n1368,
    n942
  );


  not
  g1411
  (
    n1262,
    n953
  );


  not
  g1412
  (
    n1156,
    n959
  );


  buf
  g1413
  (
    n1229,
    n941
  );


  not
  g1414
  (
    n1012,
    n871
  );


  not
  g1415
  (
    n1433,
    n888
  );


  not
  g1416
  (
    n1297,
    n877
  );


  xor
  g1417
  (
    n1268,
    n915,
    n877,
    n967,
    n903
  );


  nor
  g1418
  (
    n1259,
    n907,
    n923,
    n872,
    n968
  );


  or
  g1419
  (
    n1263,
    n958,
    n871,
    n874,
    n938
  );


  xor
  g1420
  (
    n1385,
    n874,
    n873,
    n971,
    n929
  );


  nor
  g1421
  (
    n1274,
    n940,
    n915,
    n955,
    n877
  );


  or
  g1422
  (
    n1117,
    n931,
    n893,
    n869,
    n906
  );


  xor
  g1423
  (
    n1285,
    n939,
    n915,
    n899,
    n947
  );


  or
  g1424
  (
    n1608,
    n1379,
    n1407,
    n1329,
    n1445
  );


  nand
  g1425
  (
    n1540,
    n1294,
    n1354,
    n1337,
    n405
  );


  xnor
  g1426
  (
    n1606,
    n1381,
    n408,
    n1331,
    n1226
  );


  xor
  g1427
  (
    n1662,
    n1361,
    n1392,
    n1048,
    n1346
  );


  nand
  g1428
  (
    n1456,
    n1326,
    n1350,
    n1399,
    n1166
  );


  nor
  g1429
  (
    n1622,
    n1041,
    n1237,
    n1374,
    n1443
  );


  nand
  g1430
  (
    n1464,
    n1445,
    n1035,
    n1136,
    n1377
  );


  or
  g1431
  (
    n1586,
    n1373,
    n1353,
    n1243,
    n1059
  );


  or
  g1432
  (
    n1504,
    n1362,
    n1398,
    n1078
  );


  nor
  g1433
  (
    n1522,
    n1424,
    n1175,
    n1303,
    n1173
  );


  nand
  g1434
  (
    n1570,
    n1393,
    n1403,
    n404
  );


  xor
  g1435
  (
    n1519,
    n1380,
    n1055,
    n1188,
    n1049
  );


  or
  g1436
  (
    n1530,
    n1060,
    n1415,
    n1342,
    n1109
  );


  nor
  g1437
  (
    n1491,
    n1367,
    n1413,
    n1326,
    n1369
  );


  nand
  g1438
  (
    n1602,
    n1427,
    n1079,
    n1318,
    n1252
  );


  or
  g1439
  (
    n1494,
    n1424,
    n1351,
    n1401,
    n1371
  );


  xnor
  g1440
  (
    n1474,
    n1388,
    n1402,
    n1253,
    n1082
  );


  xnor
  g1441
  (
    n1511,
    n1215,
    n1414,
    n1108,
    n1428
  );


  or
  g1442
  (
    n1481,
    n1220,
    n1099,
    n1287,
    n1116
  );


  nor
  g1443
  (
    n1476,
    n1132,
    n406,
    n1158,
    n1364
  );


  nand
  g1444
  (
    n1607,
    n1344,
    n1389,
    n764,
    n1168
  );


  nand
  g1445
  (
    n1613,
    n1229,
    n1402,
    n1437,
    n1413
  );


  and
  g1446
  (
    n1551,
    n1160,
    n1337,
    n1053,
    n1409
  );


  xnor
  g1447
  (
    n1643,
    n407,
    n1310,
    n1193,
    n1300
  );


  xor
  g1448
  (
    n1584,
    n1352,
    n1305,
    n1395,
    n1430
  );


  or
  g1449
  (
    n1610,
    n1114,
    n1354,
    n1030,
    n1024
  );


  xnor
  g1450
  (
    n1512,
    n1447,
    n412,
    n1297,
    n1421
  );


  nor
  g1451
  (
    n1495,
    n1027,
    n1380,
    n1343,
    n1368
  );


  nand
  g1452
  (
    n1486,
    n1375,
    n1313,
    n1380,
    n1401
  );


  xor
  g1453
  (
    n1660,
    n408,
    n1042,
    n1301,
    n1090
  );


  xor
  g1454
  (
    n1574,
    n1236,
    n1444,
    n1437,
    n1095
  );


  and
  g1455
  (
    n1462,
    n1306,
    n1203,
    n1213,
    n1348
  );


  xor
  g1456
  (
    n1638,
    n409,
    n1323,
    n1398,
    n1334
  );


  xor
  g1457
  (
    n1509,
    n1410,
    n1349,
    n1164,
    n1043
  );


  or
  g1458
  (
    n1536,
    n1376,
    n1420,
    n1432,
    n411
  );


  nor
  g1459
  (
    n1668,
    n1401,
    n1322,
    n1415,
    n1386
  );


  xor
  g1460
  (
    n1630,
    n1316,
    n1385,
    n1374,
    n1433
  );


  xnor
  g1461
  (
    n1533,
    n1382,
    n1299,
    n1034,
    n1391
  );


  or
  g1462
  (
    n1580,
    n1330,
    n1426,
    n1428,
    n1269
  );


  nor
  g1463
  (
    n1455,
    n1293,
    n1142,
    n1087,
    n1396
  );


  nor
  g1464
  (
    n1598,
    n1438,
    n1126,
    n1389,
    n1442
  );


  or
  g1465
  (
    n1488,
    n1267,
    n1091,
    n1376,
    n1355
  );


  nand
  g1466
  (
    n1605,
    n1391,
    n1112,
    n405,
    n1397
  );


  nor
  g1467
  (
    n1581,
    n1412,
    n1438,
    n1342,
    n1373
  );


  and
  g1468
  (
    n1567,
    n1419,
    n410,
    n1250,
    n1223
  );


  or
  g1469
  (
    n1590,
    n1406,
    n1408,
    n1425,
    n1421
  );


  xor
  g1470
  (
    n1634,
    n1178,
    n1444,
    n1192,
    n1172
  );


  xnor
  g1471
  (
    n1480,
    n412,
    n1424,
    n1359,
    n1037
  );


  nor
  g1472
  (
    n1585,
    n1384,
    n1380,
    n1446,
    n1352
  );


  or
  g1473
  (
    n1669,
    n1084,
    n1359,
    n1354,
    n1272
  );


  xor
  g1474
  (
    n1629,
    n1350,
    n1131,
    n1033,
    n1384
  );


  nor
  g1475
  (
    n1554,
    n1357,
    n1032,
    n404,
    n407
  );


  and
  g1476
  (
    n1492,
    n1254,
    n1230,
    n1329,
    n1232
  );


  or
  g1477
  (
    n1604,
    n1423,
    n1122,
    n1441,
    n1054
  );


  or
  g1478
  (
    n1478,
    n1357,
    n1362,
    n1249,
    n1377
  );


  xnor
  g1479
  (
    n1487,
    n1156,
    n1150,
    n1094,
    n1337
  );


  nand
  g1480
  (
    KeyWire_0_20,
    n1210,
    n1361,
    n1231,
    n1341
  );


  or
  g1481
  (
    n1620,
    n1443,
    n1330,
    n1426,
    n1355
  );


  nor
  g1482
  (
    n1468,
    n1330,
    n1277,
    n1296,
    n1308
  );


  xnor
  g1483
  (
    n1661,
    n1420,
    n1358,
    n1382,
    n1335
  );


  nand
  g1484
  (
    n1452,
    n1264,
    n1266,
    n1363,
    n1336
  );


  or
  g1485
  (
    n1517,
    n1187,
    n1341,
    n1319,
    n1322
  );


  and
  g1486
  (
    n1609,
    n1437,
    n1425,
    n1422,
    n1361
  );


  or
  g1487
  (
    n1624,
    n1446,
    n1397,
    n1370,
    n403
  );


  or
  g1488
  (
    n1472,
    n1386,
    n1433,
    n1211,
    n1340
  );


  xnor
  g1489
  (
    n1612,
    n1260,
    n1387,
    n1372,
    n1329
  );


  xnor
  g1490
  (
    n1556,
    n1410,
    n1434,
    n1022,
    n1040
  );


  nand
  g1491
  (
    n1475,
    n1367,
    n1416,
    n1390,
    n1436
  );


  nor
  g1492
  (
    n1550,
    n1413,
    n1089,
    n1343,
    n1367
  );


  nand
  g1493
  (
    n1600,
    n1434,
    n1270,
    n1093,
    n1333
  );


  nand
  g1494
  (
    n1461,
    n409,
    n1410,
    n1352,
    n1438
  );


  and
  g1495
  (
    n1628,
    n1015,
    n1246,
    n1278,
    n1367
  );


  and
  g1496
  (
    n1647,
    n413,
    n1137,
    n1419,
    n1359
  );


  xor
  g1497
  (
    n1641,
    n1292,
    n1373,
    n1085,
    n1344
  );


  or
  g1498
  (
    n1565,
    n1239,
    n1346,
    n1233,
    n1338
  );


  and
  g1499
  (
    n1483,
    n1191,
    n1419,
    n1351,
    n1199
  );


  xor
  g1500
  (
    n1657,
    n1348,
    n1407,
    n1409,
    n1014
  );


  nand
  g1501
  (
    n1619,
    n1381,
    n1097,
    n1449,
    n411
  );


  xor
  g1502
  (
    n1557,
    n1445,
    n1256,
    n1325
  );


  nor
  g1503
  (
    n1592,
    n1346,
    n1110,
    n1436,
    n1363
  );


  and
  g1504
  (
    n1646,
    n1274,
    n1334,
    n1381,
    n1415
  );


  and
  g1505
  (
    n1460,
    n1422,
    n1412,
    n1314,
    n1426
  );


  or
  g1506
  (
    n1531,
    n1386,
    n1373,
    n1433,
    n1123
  );


  and
  g1507
  (
    n1513,
    n1135,
    n1208,
    n1088,
    n1159
  );


  and
  g1508
  (
    n1591,
    n1376,
    n1328,
    n1395,
    n1275
  );


  nor
  g1509
  (
    n1489,
    n1324,
    n1155,
    n411,
    n1398
  );


  xnor
  g1510
  (
    n1572,
    n1242,
    n1216,
    n1081,
    n1405
  );


  nand
  g1511
  (
    n1649,
    n1382,
    n414,
    n1261,
    n1435
  );


  xnor
  g1512
  (
    n1599,
    n1438,
    n1430,
    n1441,
    n1360
  );


  xor
  g1513
  (
    n1485,
    n1363,
    n1371,
    n1430,
    n1255
  );


  xor
  g1514
  (
    n1508,
    n1432,
    n410,
    n1379,
    n406
  );


  xnor
  g1515
  (
    n1469,
    n1333,
    n1434,
    n1375,
    n1038
  );


  nor
  g1516
  (
    n1593,
    n1393,
    n1385,
    n1422,
    n1449
  );


  or
  g1517
  (
    n1479,
    n1416,
    n1446,
    n1432,
    n1241
  );


  nor
  g1518
  (
    n1666,
    n1334,
    n1394,
    n1421,
    n409
  );


  xor
  g1519
  (
    n1526,
    n1086,
    n1138,
    n1284,
    n1348
  );


  nor
  g1520
  (
    n1579,
    n1448,
    n404,
    n1411,
    n1282
  );


  xnor
  g1521
  (
    n1532,
    n414,
    n1377,
    n1396,
    n1298
  );


  xor
  g1522
  (
    n1515,
    n1387,
    n1434,
    n1194,
    n1202
  );


  xor
  g1523
  (
    n1516,
    n1317,
    n1416,
    n1435,
    n1447
  );


  nor
  g1524
  (
    n1603,
    n1356,
    n1184,
    n1257,
    n1349
  );


  xor
  g1525
  (
    n1514,
    n1141,
    n1336,
    n1064,
    n1347
  );


  and
  g1526
  (
    n1503,
    n1397,
    n1174,
    n1104,
    n1074
  );


  xor
  g1527
  (
    n1625,
    n1335,
    n1338,
    n1117,
    n1427
  );


  xor
  g1528
  (
    KeyWire_0_17,
    n1418,
    n1347,
    n1406,
    n1383
  );


  nand
  g1529
  (
    n1496,
    n1324,
    n1448,
    n1383,
    n1344
  );


  nand
  g1530
  (
    n1663,
    n1197,
    n1190,
    n1056,
    n1440
  );


  nor
  g1531
  (
    n1537,
    n406,
    n1345,
    n1385,
    n1339
  );


  and
  g1532
  (
    n1467,
    n1368,
    n1355,
    n1050,
    n1402
  );


  nor
  g1533
  (
    n1538,
    n1395,
    n1370,
    n1442,
    n411
  );


  or
  g1534
  (
    n1547,
    n1385,
    n1047,
    n1262,
    n407
  );


  or
  g1535
  (
    n1654,
    n1394,
    n1212,
    n409,
    n1279
  );


  nor
  g1536
  (
    n1539,
    n1365,
    n1428,
    n1360,
    n1280
  );


  nand
  g1537
  (
    n1470,
    n1346,
    n1423,
    n1425,
    n1371
  );


  or
  g1538
  (
    n1573,
    n1340,
    n1436,
    n1318,
    n1240
  );


  nor
  g1539
  (
    n1623,
    n1115,
    n1439,
    n1320,
    n1409
  );


  xnor
  g1540
  (
    n1458,
    n1389,
    n1157,
    n1339,
    n1393
  );


  nor
  g1541
  (
    n1527,
    n1376,
    n1390,
    n414,
    n1331
  );


  xnor
  g1542
  (
    n1571,
    n1039,
    n1384,
    n1066,
    n1165
  );


  xnor
  g1543
  (
    n1520,
    n1320,
    n1447,
    n1444,
    n1375
  );


  and
  g1544
  (
    n1626,
    n1238,
    n1205,
    n1403,
    n1320
  );


  nand
  g1545
  (
    n1543,
    n1391,
    n1189,
    n404,
    n1312
  );


  and
  g1546
  (
    n1597,
    n1439,
    n1403,
    n1442,
    n1198
  );


  xnor
  g1547
  (
    n1450,
    n1392,
    n1263,
    n1448,
    n1133
  );


  nor
  g1548
  (
    n1528,
    n1358,
    n1143,
    n1057,
    n1347
  );


  nand
  g1549
  (
    n1658,
    n1227,
    n1375,
    n1268,
    n1445
  );


  xor
  g1550
  (
    n1463,
    n1319,
    n1302,
    n1356,
    n1387
  );


  nor
  g1551
  (
    n1640,
    n1072,
    n1345,
    n1291,
    n1031
  );


  xor
  g1552
  (
    n1558,
    n1012,
    n405,
    n1358,
    n1326
  );


  xor
  g1553
  (
    n1655,
    n1444,
    n405,
    n1338,
    n1068
  );


  nor
  g1554
  (
    n1529,
    n1423,
    n1364,
    n1404,
    n1222
  );


  and
  g1555
  (
    n1525,
    n413,
    n1368,
    n1389,
    n1374
  );


  and
  g1556
  (
    n1562,
    n1083,
    n1321,
    n1361
  );


  and
  g1557
  (
    n1555,
    n1111,
    n1219,
    n1167,
    n1106
  );


  xnor
  g1558
  (
    n1542,
    n1364,
    n1076,
    n1319,
    n1378
  );


  nor
  g1559
  (
    n1477,
    n1431,
    n1429,
    n1182,
    n1286
  );


  nor
  g1560
  (
    n1521,
    n1186,
    n1207,
    n1371,
    n1171
  );


  or
  g1561
  (
    n1583,
    n1345,
    n1147,
    n1431,
    n1446
  );


  xor
  g1562
  (
    n1621,
    n1407,
    n1388,
    n1443,
    n1353
  );


  xor
  g1563
  (
    n1577,
    n1204,
    n1315,
    n1342,
    n1323
  );


  xor
  g1564
  (
    n1553,
    n1335,
    n1420,
    n1181,
    n1439
  );


  nand
  g1565
  (
    n1664,
    n1146,
    n1394,
    n1423,
    n1323
  );


  nand
  g1566
  (
    KeyWire_0_29,
    n1214,
    n1139,
    n1070,
    n1400
  );


  xnor
  g1567
  (
    n1465,
    n1311,
    n1046,
    n1392,
    n1063
  );


  xor
  g1568
  (
    n1650,
    n1351,
    n1320,
    n1429,
    n1378
  );


  or
  g1569
  (
    n1588,
    n1356,
    n1449,
    n1101,
    n1045
  );


  xnor
  g1570
  (
    n1594,
    n1307,
    n1162,
    n1319,
    n1366
  );


  xnor
  g1571
  (
    n1482,
    n412,
    n1369,
    n1358,
    n1365
  );


  or
  g1572
  (
    n1611,
    n1405,
    n1325,
    n1327,
    n1151
  );


  or
  g1573
  (
    n1559,
    n1285,
    n1416,
    n1410,
    n1412
  );


  xnor
  g1574
  (
    n1665,
    n1288,
    n1447,
    n1357,
    n1185
  );


  nor
  g1575
  (
    n1500,
    n1183,
    n1390,
    n1383,
    n1071
  );


  xor
  g1576
  (
    n1471,
    n1096,
    n1321,
    n1360,
    n410
  );


  xnor
  g1577
  (
    n1639,
    n1224,
    n1417,
    n1382,
    n1077
  );


  nand
  g1578
  (
    n1451,
    n1379,
    n1247,
    n1443,
    n1427
  );


  or
  g1579
  (
    n1457,
    n1356,
    n1121,
    n1366,
    n1435
  );


  and
  g1580
  (
    n1617,
    n1339,
    n1340,
    n1118,
    n1195
  );


  xor
  g1581
  (
    n1645,
    n1366,
    n1152,
    n1422,
    n1245
  );


  or
  g1582
  (
    n1576,
    n1304,
    n1399,
    n1332,
    n1413
  );


  nor
  g1583
  (
    n1548,
    n1153,
    n413,
    n1370,
    n1345
  );


  and
  g1584
  (
    n1631,
    n1418,
    n1441,
    n1359,
    n1429
  );


  xnor
  g1585
  (
    n1642,
    n1391,
    n1028,
    n1092,
    n1324
  );


  nand
  g1586
  (
    n1578,
    n1384,
    n1362,
    n1349,
    n1154
  );


  xnor
  g1587
  (
    n1505,
    n1388,
    n1248,
    n1283,
    n1414
  );


  nor
  g1588
  (
    n1644,
    n1439,
    n1330,
    n1145,
    n1333
  );


  xor
  g1589
  (
    n1566,
    n1429,
    n1036,
    n1200,
    n1365
  );


  xnor
  g1590
  (
    n1546,
    n1328,
    n1228,
    n1427,
    n1324
  );


  xnor
  g1591
  (
    n1490,
    n1180,
    n1400,
    n1281,
    n1052
  );


  nand
  g1592
  (
    n1552,
    n1103,
    n408,
    n1370,
    n1425
  );


  xor
  g1593
  (
    n1659,
    n1404,
    n1318,
    n1343,
    n1405
  );


  and
  g1594
  (
    n1564,
    n1401,
    n1020,
    n1128,
    n1323
  );


  nor
  g1595
  (
    n1596,
    n1259,
    n1426,
    n1328,
    n1349
  );


  xor
  g1596
  (
    n1618,
    n1105,
    n1411,
    n1067,
    n1433
  );


  nor
  g1597
  (
    n1563,
    n1290,
    n1430,
    n1399,
    n1125
  );


  xnor
  g1598
  (
    n1632,
    n1432,
    n1402,
    n1169,
    n1424
  );


  nand
  g1599
  (
    n1523,
    n1061,
    n1016,
    n1351,
    n1322
  );


  nor
  g1600
  (
    n1541,
    n1418,
    n1129,
    n1069,
    n1353
  );


  nand
  g1601
  (
    n1575,
    n1415,
    n1018,
    n1414,
    n1396
  );


  nor
  g1602
  (
    n1535,
    n1406,
    n1179,
    n1289,
    n1340
  );


  xor
  g1603
  (
    n1454,
    n1336,
    n1341,
    n1436,
    n1431
  );


  nand
  g1604
  (
    n1466,
    n1419,
    n1388,
    n1163,
    n1177
  );


  xnor
  g1605
  (
    n1615,
    n1244,
    n1209,
    n410,
    n1417
  );


  or
  g1606
  (
    n1493,
    n1341,
    n1044,
    n1107,
    n1393
  );


  and
  g1607
  (
    KeyWire_0_8,
    n1383,
    n1372,
    n1417,
    n1448
  );


  xnor
  g1608
  (
    n1497,
    n1295,
    n1404,
    n408,
    n1357
  );


  and
  g1609
  (
    n1506,
    n1337,
    n1196,
    n1075,
    n1201
  );


  nand
  g1610
  (
    n1616,
    n1221,
    n1134,
    n1409,
    n1343
  );


  nand
  g1611
  (
    n1636,
    n1338,
    n1322,
    n1234,
    n1386
  );


  xor
  g1612
  (
    n1453,
    n1206,
    n1344,
    n1051,
    n1149
  );


  xnor
  g1613
  (
    n1510,
    n1414,
    n1342,
    n1364,
    n1362
  );


  xnor
  g1614
  (
    n1633,
    n1327,
    n1251,
    n1437,
    n1332
  );


  and
  g1615
  (
    n1459,
    n1119,
    n1347,
    n1021,
    n1408
  );


  xnor
  g1616
  (
    n1589,
    n1258,
    n1372,
    n1235,
    n1273
  );


  xor
  g1617
  (
    n1484,
    n1399,
    n1335,
    n1411,
    n1417
  );


  nor
  g1618
  (
    n1507,
    n1326,
    n1161,
    n1442,
    n1392
  );


  or
  g1619
  (
    n1667,
    n1013,
    n413,
    n1026,
    n1406
  );


  and
  g1620
  (
    n1656,
    n1363,
    n412,
    n406,
    n1377
  );


  xnor
  g1621
  (
    n1652,
    n1408,
    n1265,
    n1225,
    n1058
  );


  xor
  g1622
  (
    n1534,
    n1348,
    n1332,
    n1120,
    n1440
  );


  or
  g1623
  (
    n1498,
    n1062,
    n407,
    n1327,
    n1127
  );


  xnor
  g1624
  (
    n1582,
    n1449,
    n1400,
    n1144,
    n1331
  );


  nor
  g1625
  (
    n1501,
    n1435,
    n1366,
    n1073,
    n1394
  );


  xor
  g1626
  (
    n1524,
    n1113,
    n1333,
    n1327,
    n1336
  );


  xnor
  g1627
  (
    n1637,
    n1404,
    n1418,
    n1440,
    n414
  );


  or
  g1628
  (
    n1549,
    n1102,
    n1130,
    n1140,
    n1381
  );


  nand
  g1629
  (
    n1518,
    n1328,
    n1353,
    n1431,
    n1350
  );


  xnor
  g1630
  (
    n1560,
    n1350,
    n1100,
    n1321,
    n1098
  );


  xor
  g1631
  (
    n1544,
    n1355,
    n1412,
    n1331,
    n1407
  );


  xor
  g1632
  (
    n1499,
    n1405,
    n1329,
    n1390,
    n1148
  );


  xnor
  g1633
  (
    n1648,
    n1080,
    n1325,
    n1440,
    n1176
  );


  xnor
  g1634
  (
    n1502,
    n1395,
    n1411,
    n1276,
    n1309
  );


  xnor
  g1635
  (
    n1635,
    n1372,
    n1365,
    n1408,
    n1396
  );


  and
  g1636
  (
    n1569,
    n1354,
    n1360,
    n1420,
    n1170
  );


  nand
  g1637
  (
    n1587,
    n1017,
    n1379,
    n1421,
    n1397
  );


  xor
  g1638
  (
    n1595,
    n1400,
    n1124,
    n1217,
    n1023
  );


  xnor
  g1639
  (
    n1614,
    n1374,
    n1029,
    n1339,
    n1369
  );


  xnor
  g1640
  (
    n1545,
    n1369,
    n1378,
    n1352,
    n1387
  );


  xnor
  g1641
  (
    n1473,
    n1428,
    n1019,
    n1065,
    n1368
  );


  and
  g1642
  (
    n1601,
    n1441,
    n1218,
    n1378,
    n1332
  );


  xor
  g1643
  (
    n1651,
    n1025,
    n1334,
    n1271,
    n1318
  );


  nand
  g1644
  (
    n1711,
    n988,
    n1468,
    n586,
    n1599
  );


  nand
  g1645
  (
    n1785,
    n1513,
    n1549,
    n658,
    n984
  );


  xnor
  g1646
  (
    n1755,
    n1553,
    n991,
    n1467,
    n662
  );


  nand
  g1647
  (
    n1708,
    n1582,
    n986,
    n1011,
    n1584
  );


  or
  g1648
  (
    n1758,
    n1494,
    n1519,
    n993,
    n1545
  );


  or
  g1649
  (
    n1727,
    n643,
    n618,
    n1565,
    n1509
  );


  nand
  g1650
  (
    n1783,
    n1613,
    n640,
    n1664,
    n1542
  );


  xnor
  g1651
  (
    n1709,
    n1548,
    n1635,
    n676,
    n978
  );


  or
  g1652
  (
    n1706,
    n1003,
    n641,
    n1008,
    n603
  );


  nor
  g1653
  (
    n1683,
    n1591,
    n1500,
    n1653,
    n611
  );


  or
  g1654
  (
    n1705,
    n985,
    n626,
    n1463,
    n1562
  );


  xnor
  g1655
  (
    n1738,
    n1596,
    n1489,
    n624,
    n588
  );


  and
  g1656
  (
    n1740,
    n989,
    n1010,
    n988,
    n1640
  );


  nand
  g1657
  (
    n1739,
    n1006,
    n1004,
    n1649,
    n1540
  );


  xnor
  g1658
  (
    n1774,
    n1641,
    n1496,
    n655,
    n997
  );


  and
  g1659
  (
    n1750,
    n1660,
    n1531,
    n25,
    n1469
  );


  or
  g1660
  (
    n1722,
    n1002,
    n1650,
    n1538,
    n1566
  );


  nand
  g1661
  (
    n1742,
    n1657,
    n606,
    n986,
    n1667
  );


  or
  g1662
  (
    n1672,
    n667,
    n1007,
    n1011,
    n981
  );


  xnor
  g1663
  (
    n1745,
    n578,
    n1004,
    n1662,
    n1005
  );


  xnor
  g1664
  (
    n1733,
    n990,
    n597,
    n1010,
    n581
  );


  and
  g1665
  (
    n1763,
    n595,
    n1619,
    n1011,
    n633
  );


  nand
  g1666
  (
    n1737,
    n1585,
    n1006,
    n1505,
    n1465
  );


  and
  g1667
  (
    n1715,
    n1511,
    n625,
    n620,
    n1456
  );


  nor
  g1668
  (
    n1781,
    n1637,
    n1668,
    n617,
    n998
  );


  xor
  g1669
  (
    n1710,
    n982,
    n1654,
    n607,
    n1452
  );


  and
  g1670
  (
    n1707,
    n644,
    n1479,
    n1478,
    n637
  );


  nand
  g1671
  (
    n1718,
    n1554,
    n1002,
    n1007,
    n991
  );


  and
  g1672
  (
    n1768,
    n1524,
    n1559,
    n1503,
    n656
  );


  nand
  g1673
  (
    n1712,
    n977,
    n1665,
    n1539,
    n991
  );


  nand
  g1674
  (
    n1761,
    n608,
    n982,
    n996,
    n989
  );


  xnor
  g1675
  (
    n1700,
    n1610,
    n1517,
    n987
  );


  and
  g1676
  (
    n1744,
    n1570,
    n1564,
    n989,
    n1647
  );


  nand
  g1677
  (
    n1779,
    n1615,
    n993,
    n990,
    n1481
  );


  nand
  g1678
  (
    n1696,
    n1627,
    n1508,
    n1666,
    n621
  );


  xnor
  g1679
  (
    n1720,
    n1008,
    n1636,
    n1626,
    n1609
  );


  xnor
  g1680
  (
    n1757,
    n1464,
    n674,
    n987,
    n1560
  );


  xor
  g1681
  (
    KeyWire_0_28,
    n1003,
    n1583,
    n1638,
    n1620
  );


  xor
  g1682
  (
    n1725,
    n600,
    n649,
    n661,
    n989
  );


  xor
  g1683
  (
    n1671,
    n1472,
    n1006,
    n665,
    n1614
  );


  nor
  g1684
  (
    n1759,
    n1482,
    n592,
    n1527,
    n1491
  );


  or
  g1685
  (
    n1762,
    n1574,
    n985,
    n1008,
    n636
  );


  nand
  g1686
  (
    n1678,
    n987,
    n1611,
    n1612,
    n1617
  );


  xnor
  g1687
  (
    n1699,
    n657,
    n1561,
    n634,
    n1470
  );


  or
  g1688
  (
    n1682,
    n1498,
    n978,
    n673,
    n1529
  );


  and
  g1689
  (
    n1775,
    n1628,
    n994,
    n986,
    n981
  );


  nand
  g1690
  (
    n1728,
    n1644,
    n1450,
    n1483,
    n619
  );


  nand
  g1691
  (
    n1769,
    n576,
    n998,
    n997,
    n1504
  );


  nand
  g1692
  (
    n1770,
    n996,
    n591,
    n1485,
    n638
  );


  xnor
  g1693
  (
    n1680,
    n1466,
    n1629,
    n1000,
    n1579
  );


  or
  g1694
  (
    n1734,
    n994,
    n1008,
    n601,
    n1009
  );


  or
  g1695
  (
    n1723,
    n1005,
    n594,
    n623,
    n1010
  );


  xnor
  g1696
  (
    n1674,
    n1551,
    n629,
    n998,
    n1490
  );


  nor
  g1697
  (
    n1686,
    n639,
    n1663,
    n1004,
    n1618
  );


  and
  g1698
  (
    n1765,
    n1001,
    n1606,
    n1646,
    n1525
  );


  xnor
  g1699
  (
    n1704,
    n1546,
    n983,
    n1578,
    n614
  );


  nor
  g1700
  (
    n1756,
    n1534,
    n1571,
    n1616,
    n1652
  );


  xnor
  g1701
  (
    n1675,
    n664,
    n622,
    n1645,
    n1556
  );


  or
  g1702
  (
    n1749,
    n980,
    n1597,
    n984,
    n598
  );


  xor
  g1703
  (
    n1726,
    n1002,
    n1604,
    n1651,
    n582
  );


  nand
  g1704
  (
    n1784,
    n993,
    n1528,
    n613,
    n663
  );


  xor
  g1705
  (
    n1746,
    n584,
    n1594,
    n1009,
    n1526
  );


  nand
  g1706
  (
    n1670,
    n1510,
    n651,
    n983,
    n1633
  );


  and
  g1707
  (
    n1717,
    n1555,
    n1639,
    n993,
    n670
  );


  xor
  g1708
  (
    n1676,
    n1622,
    n615,
    n1580,
    n1669
  );


  xnor
  g1709
  (
    n1684,
    n646,
    n1514,
    n1497,
    n1567
  );


  xor
  g1710
  (
    n1764,
    n1004,
    n1006,
    n981,
    n1592
  );


  nor
  g1711
  (
    n1782,
    n1575,
    n983,
    n986,
    n1486
  );


  xnor
  g1712
  (
    n1689,
    n1544,
    n587,
    n988,
    n1461
  );


  nand
  g1713
  (
    n1777,
    n585,
    n1516,
    n1598,
    n602
  );


  xor
  g1714
  (
    n1703,
    n995,
    n1521,
    n981,
    n612
  );


  xor
  g1715
  (
    n1719,
    n1501,
    n1007,
    n679,
    n642
  );


  and
  g1716
  (
    n1694,
    n1520,
    n979,
    n1523,
    n593
  );


  and
  g1717
  (
    n1731,
    n1588,
    n1001,
    n1605,
    n660
  );


  xnor
  g1718
  (
    n1741,
    n1648,
    n997,
    n1000,
    n982
  );


  nand
  g1719
  (
    n1751,
    n979,
    n680,
    n990,
    n1547
  );


  nand
  g1720
  (
    n1673,
    n1507,
    n1625,
    n1522,
    n1631
  );


  xnor
  g1721
  (
    n1729,
    n1624,
    n999,
    n1576,
    n1002
  );


  nor
  g1722
  (
    n1776,
    n995,
    n1495,
    n671,
    n985
  );


  nand
  g1723
  (
    n1685,
    n627,
    n1518,
    n979,
    n677
  );


  nand
  g1724
  (
    n1773,
    n1535,
    n1642,
    n653,
    n1460
  );


  or
  g1725
  (
    n1736,
    n1593,
    n992,
    n1480
  );


  and
  g1726
  (
    n1679,
    n984,
    n994,
    n583,
    n1623
  );


  nand
  g1727
  (
    n1691,
    n635,
    n1543,
    n605,
    n1603
  );


  nand
  g1728
  (
    n1772,
    n599,
    n1608,
    n997,
    n1005
  );


  xnor
  g1729
  (
    n1701,
    n666,
    n1451,
    n1632,
    n994
  );


  nor
  g1730
  (
    n1698,
    n998,
    n1661,
    n1009,
    n628
  );


  or
  g1731
  (
    n1681,
    n1573,
    n1488,
    n1586,
    n1552
  );


  nor
  g1732
  (
    n1732,
    n1010,
    n1656,
    n1634,
    n1590
  );


  or
  g1733
  (
    n1778,
    n580,
    n1457,
    n999,
    n590
  );


  or
  g1734
  (
    n1713,
    n985,
    n1499,
    n1474,
    n579
  );


  nor
  g1735
  (
    n1695,
    n1487,
    n1587,
    n632,
    n1550
  );


  nor
  g1736
  (
    n1714,
    n980,
    n648,
    n1000,
    n630
  );


  or
  g1737
  (
    n1743,
    n647,
    n596,
    n982,
    n1536
  );


  or
  g1738
  (
    n1752,
    n1600,
    n678,
    n672,
    n650
  );


  nand
  g1739
  (
    n1688,
    n1484,
    n1493,
    n995,
    n1532
  );


  or
  g1740
  (
    n1766,
    n604,
    n645,
    n1009,
    n652
  );


  xnor
  g1741
  (
    n1697,
    n1471,
    n1643,
    n996,
    n1515
  );


  nor
  g1742
  (
    n1760,
    n1005,
    n654,
    n978,
    n1602
  );


  nor
  g1743
  (
    n1780,
    n609,
    n992,
    n1655,
    n999
  );


  or
  g1744
  (
    n1716,
    n1581,
    n669,
    n1512,
    n577
  );


  nor
  g1745
  (
    n1748,
    n1572,
    n610,
    n1000,
    n1530
  );


  nand
  g1746
  (
    n1771,
    n977,
    n1455,
    n1621,
    n631
  );


  xor
  g1747
  (
    n1692,
    n1454,
    n1475,
    n1011,
    n1558
  );


  and
  g1748
  (
    n1754,
    n1476,
    n616,
    n1659,
    n1569
  );


  or
  g1749
  (
    n1724,
    n1453,
    n1003,
    n1630,
    n589
  );


  nor
  g1750
  (
    n1747,
    n1533,
    n1537,
    n1459,
    n1601
  );


  nand
  g1751
  (
    n1690,
    n999,
    n659,
    n984,
    n1492
  );


  nand
  g1752
  (
    n1721,
    n1506,
    n1477,
    n983,
    n988
  );


  nand
  g1753
  (
    n1767,
    n1595,
    n995,
    n990,
    n1001
  );


  or
  g1754
  (
    n1753,
    n996,
    n675,
    n1563,
    n1568
  );


  and
  g1755
  (
    n1730,
    n1589,
    n1001,
    n1557,
    n1502
  );


  or
  g1756
  (
    n1693,
    n1577,
    n991,
    n980,
    n1462
  );


  xnor
  g1757
  (
    n1702,
    n668,
    n1607,
    n1473,
    n980
  );


  xnor
  g1758
  (
    KeyWire_0_31,
    n978,
    n1003,
    n1658,
    n1007
  );


  xnor
  g1759
  (
    n1735,
    n979,
    n1458,
    n992,
    n1541
  );


  nor
  g1760
  (
    n1814,
    n1723,
    n1694,
    n1707,
    n1705
  );


  xor
  g1761
  (
    n1812,
    n1675,
    n1722,
    n1746,
    n1716
  );


  nor
  g1762
  (
    n1795,
    n1703,
    n1682,
    n1720,
    n1709
  );


  nand
  g1763
  (
    n1805,
    n1696,
    n1727,
    n1752,
    n1699
  );


  nor
  g1764
  (
    n1798,
    n1728,
    n1686,
    n1739,
    n1767
  );


  xor
  g1765
  (
    n1810,
    n1743,
    n1678,
    n1714,
    n1744
  );


  nand
  g1766
  (
    n1794,
    n1681,
    n1742,
    n1734,
    n1670
  );


  nand
  g1767
  (
    n1806,
    n1779,
    n1735,
    n1680,
    n1730
  );


  nand
  g1768
  (
    n1804,
    n1689,
    n1704,
    n1695,
    n1749
  );


  xnor
  g1769
  (
    n1786,
    n1731,
    n1691,
    n1778,
    n1777
  );


  xnor
  g1770
  (
    n1796,
    n1761,
    n1685,
    n1721,
    n1718
  );


  xor
  g1771
  (
    n1789,
    n1679,
    n1780,
    n1762,
    n1759
  );


  xnor
  g1772
  (
    KeyWire_0_10,
    n1671,
    n1683,
    n1755,
    n1783
  );


  nor
  g1773
  (
    n1808,
    n1764,
    n1753,
    n1748,
    n1784
  );


  xnor
  g1774
  (
    n1813,
    n1733,
    n1757,
    n1729,
    n1732
  );


  xnor
  g1775
  (
    KeyWire_0_7,
    n1747,
    n1756,
    n1774,
    n1677
  );


  and
  g1776
  (
    n1790,
    n1684,
    n1754,
    n1700,
    n1697
  );


  or
  g1777
  (
    n1787,
    n1773,
    n1710,
    n1775,
    n1688
  );


  nand
  g1778
  (
    n1801,
    n1706,
    n1769,
    n1750,
    n1776
  );


  or
  g1779
  (
    n1792,
    n1672,
    n1726,
    n1738,
    n1768
  );


  xnor
  g1780
  (
    n1809,
    n1771,
    n1673,
    n1674,
    n1693
  );


  xor
  g1781
  (
    n1788,
    n1717,
    n1702,
    n1741,
    n1760
  );


  and
  g1782
  (
    n1791,
    n1711,
    n1782,
    n1698,
    n1690
  );


  xnor
  g1783
  (
    n1793,
    n1719,
    n1736,
    n1765,
    n1758
  );


  or
  g1784
  (
    n1797,
    n1737,
    n1751,
    n1772,
    n1725
  );


  and
  g1785
  (
    n1799,
    n1713,
    n1770,
    n1740,
    n1676
  );


  nor
  g1786
  (
    n1811,
    n1785,
    n1766,
    n1715,
    n1763
  );


  and
  g1787
  (
    n1803,
    n1692,
    n1712,
    n1781,
    n1701
  );


  nand
  g1788
  (
    n1800,
    n1724,
    n1687,
    n1708,
    n1745
  );


  xor
  KeyGate_0_0
  (
    n593,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n1430,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n434,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n586,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1283,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n92,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n404,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1802,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n1627,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n935,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n1807,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n868,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n546,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1380,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n1015,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n342,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1089,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1561,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n293,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n104,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1653,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1358,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n1410,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n1428,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n403,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n647,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n702,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n29,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1687,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n1568,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n759,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n1677,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

