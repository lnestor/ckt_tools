// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_177_411 written by SynthGen on 2021/05/24 19:47:13
module Stat_177_411( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18,
 nCHANGED, n192, n187, n186, n177, n194, n189, n190,
 n195, n180, n184, n185, n179, n188, n178, n176,
 n193, n191, n181, n183, n182);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18;

output nCHANGED, n192, n187, n186, n177, n194, n189, n190,
 n195, n180, n184, n185, n179, n188, n178, n176,
 n193, n191, n181, n183, n182;

wire n19, n20, n21, n22, n23, n24, n25, n26,
 n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175;

not  g0 (n35, n12);
buf  g1 (n29, n9);
not  g2 (n34, n7);
not  g3 (n25, n6);
not  g4 (n33, n5);
not  g5 (n27, n17);
not  g6 (n26, n16);
buf  g7 (n28, n2);
buf  g8 (n30, n8);
not  g9 (n22, n3);
buf  g10 (n23, n18);
buf  g11 (n19, n14);
not  g12 (n32, n13);
buf  g13 (n21, n15);
buf  g14 (n31, n4);
buf  g15 (n24, n10);
buf  g16 (n20, n11);
buf  g17 (n90, n20);
buf  g18 (n96, n34);
buf  g19 (n46, n25);
buf  g20 (n99, n19);
not  g21 (n77, n35);
buf  g22 (n68, n27);
not  g23 (n64, n23);
not  g24 (n40, n31);
not  g25 (n66, n34);
buf  g26 (n70, n28);
buf  g27 (n63, n26);
buf  g28 (n50, n24);
not  g29 (n81, n25);
not  g30 (n86, n25);
buf  g31 (n41, n24);
not  g32 (n53, n32);
not  g33 (n73, n35);
not  g34 (n55, n19);
buf  g35 (n57, n21);
buf  g36 (n78, n29);
buf  g37 (n79, n30);
buf  g38 (n44, n33);
not  g39 (n60, n20);
buf  g40 (n59, n33);
not  g41 (n65, n21);
buf  g42 (n103, n22);
not  g43 (n97, n26);
buf  g44 (n47, n26);
buf  g45 (n88, n33);
not  g46 (n89, n25);
buf  g47 (n56, n34);
not  g48 (n51, n19);
not  g49 (n93, n30);
buf  g50 (n91, n27);
not  g51 (n95, n24);
buf  g52 (n100, n32);
buf  g53 (n98, n30);
buf  g54 (n58, n22);
not  g55 (n101, n23);
buf  g56 (n74, n32);
buf  g57 (n80, n35);
not  g58 (n76, n27);
not  g59 (n83, n20);
not  g60 (n67, n23);
buf  g61 (n42, n23);
buf  g62 (n36, n22);
buf  g63 (n75, n29);
buf  g64 (n61, n28);
not  g65 (n54, n34);
not  g66 (n49, n21);
buf  g67 (n85, n30);
buf  g68 (n84, n31);
buf  g69 (n62, n31);
not  g70 (n102, n20);
buf  g71 (n43, n29);
buf  g72 (n92, n35);
buf  g73 (n52, n24);
buf  g74 (n39, n29);
not  g75 (n45, n28);
not  g76 (n94, n27);
buf  g77 (n69, n31);
buf  g78 (n82, n28);
buf  g79 (n71, n33);
buf  g80 (n38, n19);
buf  g81 (n48, n21);
buf  g82 (n37, n26);
not  g83 (n87, n32);
not  g84 (n72, n22);
nor  g85 (n115, n52, n102, n64);
nand g86 (n153, n94, n56, n79);
xor  g87 (n116, n41, n96, n43);
or   g88 (n112, n82, n57, n96);
xnor g89 (n161, n64, n82, n93);
or   g90 (n120, n62, n94, n70);
or   g91 (n149, n44, n38, n60);
nor  g92 (n171, n58, n93, n51);
nor  g93 (n129, n95, n103, n56);
or   g94 (n165, n78, n86, n70);
or   g95 (n108, n101, n37, n52);
and  g96 (n172, n91, n92, n67);
xnor g97 (n169, n100, n45, n59);
nand g98 (n131, n93, n80, n102);
xnor g99 (n134, n91, n50, n76);
xnor g100 (n166, n80, n55, n52);
nand g101 (n158, n62, n97, n54, n66);
xor  g102 (n156, n61, n90, n36, n82);
and  g103 (n152, n92, n45, n36, n54);
or   g104 (n163, n102, n73, n44, n74);
xnor g105 (n136, n43, n77, n76, n99);
and  g106 (n170, n100, n95, n69, n70);
xnor g107 (n144, n54, n42, n81, n98);
xor  g108 (n130, n40, n82, n51, n85);
and  g109 (n140, n77, n48, n78, n96);
nand g110 (n141, n42, n72, n47, n78);
or   g111 (n133, n66, n89, n100, n39);
nor  g112 (n164, n48, n72, n38, n49);
and  g113 (n162, n103, n84, n53, n58);
or   g114 (n122, n72, n92, n81, n43);
xor  g115 (n142, n48, n68, n56, n42);
xor  g116 (n132, n50, n72, n41, n98);
nand g117 (n135, n68, n54, n69, n88);
and  g118 (n148, n51, n55, n63);
nand g119 (n126, n61, n68, n64, n74);
nor  g120 (n137, n37, n83, n89, n97);
xor  g121 (n118, n36, n71, n95, n44);
xor  g122 (n168, n101, n39, n94, n96);
or   g123 (n109, n87, n50, n69, n37);
nand g124 (n104, n76, n66, n93, n85);
nand g125 (n110, n40, n99, n76, n67);
nand g126 (n160, n90, n46, n65, n47);
or   g127 (n117, n65, n83, n50, n89);
xor  g128 (n123, n88, n71, n97, n83);
and  g129 (n143, n75, n62, n85, n38);
nand g130 (n147, n85, n59, n65, n46);
or   g131 (n119, n57, n40, n69, n91);
nor  g132 (n154, n99, n53, n73, n59);
xnor g133 (n125, n95, n97, n77, n63);
xor  g134 (n167, n83, n80, n86, n87);
nor  g135 (n127, n55, n58, n60, n61);
nor  g136 (n173, n41, n57, n71, n36);
xnor g137 (n146, n66, n101, n74, n78);
xor  g138 (n157, n39, n51, n84, n49);
nor  g139 (n151, n46, n88, n65, n40);
or   g140 (n124, n86, n58, n101, n87);
and  g141 (n139, n60, n94, n73, n81);
and  g142 (n113, n48, n87, n90, n47);
xnor g143 (n128, n91, n68, n102, n37);
nor  g144 (n155, n49, n79, n90, n52);
or   g145 (n106, n88, n63, n73, n60);
nor  g146 (n175, n98, n45, n53, n74);
or   g147 (n145, n61, n70, n75);
nand g148 (n107, n64, n59, n79, n43);
nand g149 (n105, n45, n92, n41, n84);
nor  g150 (n150, n71, n100, n49, n57);
or   g151 (n174, n98, n84, n67, n46);
nand g152 (n114, n56, n81, n89, n53);
xor  g153 (n111, n42, n103, n86);
xor  g154 (n159, n38, n99, n44, n75);
or   g155 (n138, n77, n79, n63, n62);
nand g156 (n121, n67, n47, n39, n80);
not  g157 (n183, n119);
not  g158 (n188, n122);
and  g159 (n194, n162, n126);
nand g160 (n195, n104, n164, n151, n123);
and  g161 (n189, n173, n141, n161, n145);
or   g162 (n186, n148, n131, n128, n139);
nor  g163 (n184, n112, n165, n153, n149);
nor  g164 (n177, n171, n174, n113, n160);
xnor g165 (n187, n155, n134, n117, n137);
nor  g166 (n181, n105, n142, n138, n132);
nor  g167 (n176, n154, n146, n166, n135);
or   g168 (n193, n129, n152, n156, n116);
or   g169 (n179, n130, n169, n127, n114);
xnor g170 (n178, n168, n118, n144, n163);
or   g171 (n190, n109, n111, n110, n108);
or   g172 (n180, n115, n157, n133, n124);
and  g173 (n182, n140, n121, n150, n159);
or   g174 (n192, n120, n167, n147, n136);
nor  g175 (n191, n125, n107, n175, n170);
and  g176 (n185, n106, n172, n158, n143);
buf g177 (nCHANGED, n13);
endmodule
