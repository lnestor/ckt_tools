

module Stat_100_58
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n108,
  n113,
  n110,
  n105,
  n128,
  n129,
  n131,
  n107,
  n122,
  n118,
  n115,
  n127,
  n130,
  n121,
  n102,
  n103,
  n106,
  n132,
  n124,
  n104,
  n125,
  n119,
  n123,
  n116,
  n117,
  n120,
  n109,
  n126,
  n101,
  n114,
  n111,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  output n112;
  output n108;
  output n113;
  output n110;
  output n105;
  output n128;
  output n129;
  output n131;
  output n107;
  output n122;
  output n118;
  output n115;
  output n127;
  output n130;
  output n121;
  output n102;
  output n103;
  output n106;
  output n132;
  output n124;
  output n104;
  output n125;
  output n119;
  output n123;
  output n116;
  output n117;
  output n120;
  output n109;
  output n126;
  output n101;
  output n114;
  output n111;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;

  buf
  g0
  (
    KeyWire_0_27,
    n17
  );


  not
  g1
  (
    n53,
    n16
  );


  buf
  g2
  (
    KeyWire_0_4,
    n13
  );


  not
  g3
  (
    n45,
    n13
  );


  buf
  g4
  (
    n66,
    n10
  );


  not
  g5
  (
    n49,
    n12
  );


  not
  g6
  (
    n67,
    n16
  );


  buf
  g7
  (
    n58,
    n9
  );


  not
  g8
  (
    KeyWire_0_25,
    n15
  );


  buf
  g9
  (
    KeyWire_0_22,
    n17
  );


  buf
  g10
  (
    n61,
    n14
  );


  buf
  g11
  (
    n50,
    n18
  );


  buf
  g12
  (
    KeyWire_0_10,
    n1
  );


  not
  g13
  (
    n40,
    n14
  );


  buf
  g14
  (
    KeyWire_0_18,
    n18
  );


  not
  g15
  (
    n43,
    n5
  );


  buf
  g16
  (
    n55,
    n19
  );


  not
  g17
  (
    n48,
    n17
  );


  not
  g18
  (
    n52,
    n11
  );


  not
  g19
  (
    n65,
    n16
  );


  buf
  g20
  (
    n47,
    n9
  );


  not
  g21
  (
    n62,
    n11
  );


  not
  g22
  (
    KeyWire_0_7,
    n8
  );


  not
  g23
  (
    KeyWire_0_6,
    n11
  );


  buf
  g24
  (
    KeyWire_0_17,
    n4
  );


  buf
  g25
  (
    KeyWire_0_11,
    n12
  );


  not
  g26
  (
    KeyWire_0_28,
    n3
  );


  not
  g27
  (
    n36,
    n12
  );


  buf
  g28
  (
    n34,
    n19
  );


  buf
  g29
  (
    KeyWire_0_24,
    n6
  );


  buf
  g30
  (
    n68,
    n9
  );


  not
  g31
  (
    n37,
    n13
  );


  buf
  g32
  (
    n69,
    n18
  );


  buf
  g33
  (
    KeyWire_0_23,
    n2
  );


  buf
  g34
  (
    n33,
    n7
  );


  not
  g35
  (
    KeyWire_0_26,
    n15
  );


  buf
  g36
  (
    n59,
    n15
  );


  not
  g37
  (
    n51,
    n10
  );


  buf
  g38
  (
    n54,
    n14
  );


  buf
  g39
  (
    n60,
    n10
  );


  buf
  g40
  (
    n77,
    n37
  );


  buf
  g41
  (
    n76,
    n40
  );


  buf
  g42
  (
    n80,
    n38
  );


  buf
  g43
  (
    KeyWire_0_2,
    n34
  );


  not
  g44
  (
    KeyWire_0_20,
    n36
  );


  buf
  g45
  (
    KeyWire_0_19,
    n40
  );


  not
  g46
  (
    n79,
    n35
  );


  nor
  g47
  (
    n73,
    n33,
    n39,
    n40
  );


  buf
  g48
  (
    n82,
    n73
  );


  not
  g49
  (
    n84,
    n75
  );


  not
  g50
  (
    KeyWire_0_30,
    n74
  );


  not
  g51
  (
    n85,
    n77
  );


  not
  g52
  (
    n81,
    n76
  );


  nand
  g53
  (
    n96,
    n22,
    n80,
    n81,
    n27
  );


  and
  g54
  (
    n98,
    n32,
    n21,
    n84
  );


  xnor
  g55
  (
    n91,
    n24,
    n78,
    n27,
    n20
  );


  xnor
  g56
  (
    KeyWire_0_31,
    n30,
    n85,
    n32
  );


  nand
  g57
  (
    n88,
    n19,
    n25,
    n84,
    n24
  );


  nor
  g58
  (
    n97,
    n22,
    n84,
    n32,
    n21
  );


  xnor
  g59
  (
    n100,
    n85,
    n29,
    n23,
    n82
  );


  xor
  g60
  (
    n93,
    n80,
    n83,
    n31,
    n81
  );


  xor
  g61
  (
    n94,
    n82,
    n31,
    n27
  );


  xor
  g62
  (
    n86,
    n22,
    n25,
    n83,
    n26
  );


  nand
  g63
  (
    n87,
    n30,
    n30,
    n25,
    n20
  );


  and
  g64
  (
    n89,
    n23,
    n26,
    n83,
    n82
  );


  and
  g65
  (
    KeyWire_0_0,
    n20,
    n79,
    n28,
    n29
  );


  nor
  g66
  (
    n95,
    n23,
    n26,
    n29,
    n24
  );


  or
  g67
  (
    KeyWire_0_1,
    n81,
    n28,
    n80
  );


  nor
  g68
  (
    n121,
    n44,
    n65,
    n56,
    n63
  );


  and
  g69
  (
    n108,
    n59,
    n52,
    n45,
    n72
  );


  xor
  g70
  (
    n126,
    n67,
    n62,
    n86,
    n98
  );


  and
  g71
  (
    KeyWire_0_12,
    n49,
    n59,
    n65,
    n55
  );


  or
  g72
  (
    n109,
    n93,
    n69,
    n96
  );


  nand
  g73
  (
    n132,
    n54,
    n70,
    n92,
    n58
  );


  xor
  g74
  (
    KeyWire_0_3,
    n69,
    n43,
    n94,
    n62
  );


  and
  g75
  (
    n125,
    n95,
    n61,
    n93,
    n42
  );


  xor
  g76
  (
    n129,
    n53,
    n59,
    n60,
    n54
  );


  or
  g77
  (
    n130,
    n94,
    n51,
    n64,
    n66
  );


  nand
  g78
  (
    KeyWire_0_21,
    n46,
    n57,
    n92,
    n47
  );


  xnor
  g79
  (
    KeyWire_0_8,
    n93,
    n72,
    n98,
    n71
  );


  or
  g80
  (
    n107,
    n56,
    n97,
    n50,
    n64
  );


  nor
  g81
  (
    n122,
    n42,
    n55,
    n53,
    n63
  );


  and
  g82
  (
    KeyWire_0_14,
    n52,
    n100,
    n97,
    n91
  );


  nor
  g83
  (
    n114,
    n99,
    n94,
    n100,
    n57
  );


  nor
  g84
  (
    n110,
    n98,
    n45,
    n69,
    n61
  );


  or
  g85
  (
    KeyWire_0_15,
    n95,
    n70,
    n87,
    n68
  );


  xor
  g86
  (
    KeyWire_0_5,
    n50,
    n49,
    n43,
    n71
  );


  and
  g87
  (
    n104,
    n48,
    n56,
    n67,
    n51
  );


  or
  g88
  (
    n131,
    n61,
    n41,
    n90,
    n70
  );


  xnor
  g89
  (
    n118,
    n48,
    n62,
    n64,
    n57
  );


  and
  g90
  (
    n113,
    n50,
    n51,
    n44,
    n41
  );


  xor
  g91
  (
    n120,
    n45,
    n66,
    n49,
    n99
  );


  nand
  g92
  (
    KeyWire_0_9,
    n60,
    n52,
    n42,
    n97
  );


  nand
  g93
  (
    n115,
    n96,
    n68,
    n65,
    n63
  );


  and
  g94
  (
    KeyWire_0_13,
    n71,
    n67,
    n89,
    n53
  );


  nor
  g95
  (
    n128,
    n66,
    n72,
    n55,
    n100
  );


  or
  g96
  (
    n117,
    n46,
    n68,
    n43,
    n47
  );


  or
  g97
  (
    n101,
    n58,
    n41,
    n95,
    n54
  );


  nand
  g98
  (
    KeyWire_0_16,
    n44,
    n88,
    n58,
    n60
  );


  nor
  g99
  (
    KeyWire_0_29,
    n48,
    n99,
    n47,
    n46
  );


  xnor
  KeyGate_0_0
  (
    n90,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n92,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n78,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n106,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n70,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n111,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n56,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n41,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n119,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n105,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n71,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n35,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n123,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n112,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n116,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n102,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n127,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n39,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n72,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n74,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n75,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n124,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n42,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n44,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n57,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n46,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n64,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n63,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n38,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n103,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n83,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n99,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

