// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_225 written by SynthGen on 2021/04/05 11:23:26
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_225 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1718, n1775, n1764, n1758, n1765, n1755, n1773, n1750,
 n1768, n1757, n1769, n1771, n1748, n1759, n1751, n1749,
 n1770, n1754, n1762, n1804, n1797, n1802, n1791, n1806,
 n1789, n1801, n2030, n2031, n2029, n2027, n2028, n2032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1718, n1775, n1764, n1758, n1765, n1755, n1773, n1750,
 n1768, n1757, n1769, n1771, n1748, n1759, n1751, n1749,
 n1770, n1754, n1762, n1804, n1797, n1802, n1791, n1806,
 n1789, n1801, n2030, n2031, n2029, n2027, n2028, n2032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
 n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
 n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
 n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
 n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
 n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
 n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
 n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
 n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
 n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
 n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
 n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
 n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
 n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
 n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
 n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
 n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
 n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
 n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
 n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
 n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
 n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
 n1713, n1714, n1715, n1716, n1717, n1719, n1720, n1721,
 n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
 n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
 n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
 n1746, n1747, n1752, n1753, n1756, n1760, n1761, n1763,
 n1766, n1767, n1772, n1774, n1776, n1777, n1778, n1779,
 n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
 n1788, n1790, n1792, n1793, n1794, n1795, n1796, n1798,
 n1799, n1800, n1803, n1805, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
 n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986,
 n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
 n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
 n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
 n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
 n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026;

buf  g0 (n79, n13);
buf  g1 (n57, n12);
not  g2 (n104, n11);
buf  g3 (n77, n24);
buf  g4 (n50, n30);
not  g5 (n93, n12);
not  g6 (n111, n30);
buf  g7 (n124, n26);
not  g8 (n116, n5);
buf  g9 (n53, n22);
buf  g10 (n56, n26);
buf  g11 (n101, n20);
buf  g12 (n86, n18);
not  g13 (n113, n9);
not  g14 (n45, n31);
not  g15 (n78, n17);
buf  g16 (n81, n32);
not  g17 (n135, n17);
not  g18 (n76, n5);
buf  g19 (n89, n18);
not  g20 (n142, n3);
buf  g21 (n147, n14);
not  g22 (n34, n1);
buf  g23 (n133, n28);
not  g24 (n84, n25);
not  g25 (n95, n17);
not  g26 (n117, n15);
buf  g27 (n106, n16);
buf  g28 (n62, n13);
buf  g29 (n150, n8);
buf  g30 (n107, n29);
not  g31 (n52, n26);
buf  g32 (n127, n6);
buf  g33 (n80, n16);
not  g34 (n156, n31);
not  g35 (n83, n6);
not  g36 (n87, n31);
buf  g37 (n47, n7);
not  g38 (n75, n25);
not  g39 (n139, n20);
not  g40 (n136, n11);
not  g41 (n69, n21);
not  g42 (n61, n19);
buf  g43 (n132, n2);
buf  g44 (n126, n16);
not  g45 (n43, n12);
buf  g46 (n120, n11);
buf  g47 (n99, n27);
not  g48 (n42, n7);
buf  g49 (n130, n28);
not  g50 (n158, n24);
buf  g51 (n144, n27);
not  g52 (n148, n25);
not  g53 (n145, n29);
buf  g54 (n102, n21);
not  g55 (n129, n1);
not  g56 (n154, n5);
buf  g57 (n74, n21);
not  g58 (n36, n15);
buf  g59 (n63, n4);
buf  g60 (n151, n13);
not  g61 (n88, n30);
buf  g62 (n155, n18);
buf  g63 (n68, n4);
buf  g64 (n123, n3);
not  g65 (n149, n14);
buf  g66 (n67, n10);
buf  g67 (n122, n24);
buf  g68 (n118, n1);
not  g69 (n90, n19);
not  g70 (n109, n29);
not  g71 (n114, n31);
not  g72 (n58, n32);
not  g73 (n51, n10);
buf  g74 (n35, n17);
not  g75 (n140, n24);
buf  g76 (n105, n29);
not  g77 (n100, n14);
buf  g78 (n41, n12);
buf  g79 (n54, n23);
not  g80 (n131, n21);
buf  g81 (n152, n4);
buf  g82 (n115, n6);
buf  g83 (n40, n19);
not  g84 (n143, n25);
buf  g85 (n72, n28);
not  g86 (n39, n7);
buf  g87 (n153, n3);
buf  g88 (n73, n32);
not  g89 (n46, n9);
not  g90 (n94, n22);
not  g91 (n48, n20);
not  g92 (n38, n13);
buf  g93 (n138, n18);
not  g94 (n71, n8);
not  g95 (n110, n14);
buf  g96 (n119, n3);
not  g97 (n49, n22);
buf  g98 (n108, n15);
buf  g99 (n98, n27);
buf  g100 (n128, n10);
not  g101 (n160, n9);
not  g102 (n97, n4);
buf  g103 (n65, n11);
not  g104 (n112, n15);
not  g105 (n159, n16);
not  g106 (n85, n9);
not  g107 (n91, n22);
not  g108 (n134, n28);
buf  g109 (n44, n8);
buf  g110 (n125, n7);
buf  g111 (n66, n2);
not  g112 (n82, n6);
buf  g113 (n103, n1);
buf  g114 (n70, n2);
buf  g115 (n137, n23);
not  g116 (n37, n32);
buf  g117 (n96, n26);
not  g118 (n60, n10);
buf  g119 (n33, n23);
buf  g120 (n141, n8);
buf  g121 (n146, n23);
buf  g122 (n121, n2);
not  g123 (n55, n27);
not  g124 (n157, n5);
not  g125 (n92, n20);
not  g126 (n64, n19);
not  g127 (n59, n30);
buf  g128 (n630, n119);
buf  g129 (n490, n149);
not  g130 (n650, n81);
not  g131 (n453, n41);
not  g132 (n208, n50);
not  g133 (n593, n40);
not  g134 (n309, n105);
not  g135 (n380, n147);
not  g136 (n649, n126);
buf  g137 (n358, n101);
not  g138 (n646, n145);
buf  g139 (n245, n43);
not  g140 (n241, n46);
not  g141 (n297, n99);
not  g142 (n510, n80);
not  g143 (n509, n152);
buf  g144 (n577, n83);
not  g145 (n240, n91);
not  g146 (n169, n33);
not  g147 (n399, n134);
buf  g148 (n261, n147);
not  g149 (n415, n54);
not  g150 (n653, n66);
not  g151 (n525, n119);
buf  g152 (n352, n54);
not  g153 (n536, n130);
buf  g154 (n391, n154);
buf  g155 (n591, n155);
not  g156 (n171, n120);
not  g157 (n366, n79);
buf  g158 (n269, n66);
buf  g159 (n183, n152);
not  g160 (n596, n67);
buf  g161 (n424, n49);
not  g162 (n557, n68);
buf  g163 (n329, n91);
buf  g164 (n361, n139);
not  g165 (n512, n113);
buf  g166 (n317, n107);
buf  g167 (n461, n46);
not  g168 (n579, n120);
buf  g169 (n634, n50);
buf  g170 (n396, n79);
not  g171 (n242, n64);
not  g172 (n548, n68);
buf  g173 (n544, n73);
buf  g174 (n587, n104);
buf  g175 (n389, n77);
buf  g176 (n530, n108);
not  g177 (n243, n41);
buf  g178 (n501, n97);
not  g179 (n231, n54);
buf  g180 (n522, n127);
not  g181 (n449, n92);
not  g182 (n246, n112);
buf  g183 (n372, n143);
not  g184 (n661, n40);
not  g185 (n534, n142);
not  g186 (n635, n38);
buf  g187 (n494, n38);
not  g188 (n194, n43);
buf  g189 (n450, n159);
not  g190 (n344, n42);
not  g191 (n437, n71);
buf  g192 (n333, n130);
buf  g193 (n316, n150);
buf  g194 (n489, n108);
buf  g195 (n373, n148);
buf  g196 (n527, n42);
buf  g197 (n405, n38);
not  g198 (n216, n40);
not  g199 (n561, n55);
not  g200 (n293, n100);
buf  g201 (n495, n158);
buf  g202 (n448, n63);
buf  g203 (n488, n135);
buf  g204 (n300, n124);
buf  g205 (n563, n120);
not  g206 (n395, n69);
buf  g207 (n416, n33);
not  g208 (n457, n142);
buf  g209 (n638, n64);
buf  g210 (n601, n95);
not  g211 (n475, n158);
buf  g212 (n647, n126);
buf  g213 (n408, n140);
not  g214 (n386, n120);
not  g215 (n622, n75);
not  g216 (n428, n106);
not  g217 (n545, n105);
not  g218 (n432, n139);
buf  g219 (n324, n76);
buf  g220 (n521, n135);
not  g221 (n303, n89);
not  g222 (n190, n82);
not  g223 (n403, n54);
buf  g224 (n631, n140);
not  g225 (n398, n61);
buf  g226 (n346, n61);
not  g227 (n652, n34);
not  g228 (n304, n90);
buf  g229 (n247, n68);
not  g230 (n538, n86);
not  g231 (n263, n132);
not  g232 (n255, n57);
not  g233 (n497, n68);
buf  g234 (n307, n128);
not  g235 (n272, n98);
buf  g236 (n185, n95);
not  g237 (n586, n124);
buf  g238 (n262, n39);
buf  g239 (n340, n158);
not  g240 (n610, n44);
not  g241 (n665, n79);
buf  g242 (n574, n137);
buf  g243 (n221, n135);
buf  g244 (n573, n70);
not  g245 (n655, n36);
not  g246 (n259, n158);
not  g247 (n543, n129);
buf  g248 (n524, n114);
buf  g249 (n420, n38);
not  g250 (n302, n89);
not  g251 (n628, n131);
not  g252 (n659, n103);
buf  g253 (n287, n41);
buf  g254 (n315, n155);
not  g255 (n611, n114);
buf  g256 (n220, n64);
not  g257 (n321, n99);
not  g258 (n257, n47);
buf  g259 (n618, n83);
buf  g260 (n180, n50);
not  g261 (n376, n130);
buf  g262 (n199, n123);
buf  g263 (n514, n94);
buf  g264 (n248, n150);
buf  g265 (n452, n48);
not  g266 (n583, n146);
not  g267 (n170, n75);
buf  g268 (n230, n93);
buf  g269 (n417, n88);
not  g270 (n513, n83);
buf  g271 (n589, n57);
not  g272 (n662, n86);
not  g273 (n546, n157);
buf  g274 (n533, n78);
not  g275 (n163, n141);
buf  g276 (n474, n138);
not  g277 (n312, n73);
buf  g278 (n350, n85);
not  g279 (n167, n111);
not  g280 (n277, n125);
buf  g281 (n639, n67);
buf  g282 (n336, n88);
buf  g283 (n296, n150);
buf  g284 (n466, n85);
buf  g285 (n294, n139);
not  g286 (n581, n102);
not  g287 (n603, n45);
not  g288 (n164, n82);
buf  g289 (n479, n132);
buf  g290 (n195, n98);
buf  g291 (n175, n37);
buf  g292 (n496, n86);
buf  g293 (n556, n114);
buf  g294 (n595, n84);
buf  g295 (n560, n59);
not  g296 (n658, n116);
not  g297 (n569, n47);
not  g298 (n644, n110);
buf  g299 (n298, n44);
buf  g300 (n590, n110);
not  g301 (n555, n106);
buf  g302 (n584, n74);
buf  g303 (n267, n98);
not  g304 (n279, n35);
not  g305 (n425, n89);
buf  g306 (n431, n92);
not  g307 (n162, n87);
buf  g308 (n455, n71);
not  g309 (n367, n39);
not  g310 (n290, n59);
not  g311 (n381, n140);
buf  g312 (n582, n143);
buf  g313 (n283, n69);
buf  g314 (n327, n126);
buf  g315 (n305, n122);
not  g316 (n365, n57);
buf  g317 (n531, n63);
not  g318 (n423, n141);
not  g319 (n224, n44);
buf  g320 (n244, n97);
buf  g321 (n619, n140);
buf  g322 (n440, n110);
buf  g323 (n223, n39);
buf  g324 (n460, n149);
not  g325 (n471, n109);
buf  g326 (n377, n147);
not  g327 (n478, n154);
buf  g328 (n498, n98);
buf  g329 (n613, n62);
buf  g330 (n552, n111);
buf  g331 (n492, n48);
buf  g332 (n189, n160);
buf  g333 (n566, n35);
not  g334 (n617, n133);
not  g335 (n233, n84);
not  g336 (n249, n122);
not  g337 (n390, n104);
not  g338 (n620, n56);
buf  g339 (n239, n89);
not  g340 (n414, n153);
buf  g341 (n339, n136);
not  g342 (n627, n109);
not  g343 (n483, n130);
buf  g344 (n371, n55);
not  g345 (n282, n56);
buf  g346 (n656, n82);
not  g347 (n385, n78);
not  g348 (n193, n45);
buf  g349 (n480, n40);
not  g350 (n671, n152);
not  g351 (n491, n35);
buf  g352 (n331, n86);
buf  g353 (n217, n125);
buf  g354 (n228, n145);
buf  g355 (n559, n112);
buf  g356 (n549, n155);
not  g357 (n486, n51);
buf  g358 (n337, n116);
buf  g359 (n310, n87);
buf  g360 (n651, n69);
buf  g361 (n429, n100);
not  g362 (n402, n60);
not  g363 (n571, n157);
not  g364 (n181, n139);
buf  g365 (n172, n137);
not  g366 (n565, n74);
not  g367 (n532, n67);
not  g368 (n487, n90);
buf  g369 (n258, n116);
buf  g370 (n251, n81);
buf  g371 (n516, n147);
not  g372 (n477, n118);
buf  g373 (n553, n63);
not  g374 (n614, n118);
buf  g375 (n467, n70);
not  g376 (n214, n150);
not  g377 (n347, n77);
buf  g378 (n187, n45);
buf  g379 (n179, n60);
buf  g380 (n482, n119);
not  g381 (n433, n46);
buf  g382 (n355, n53);
not  g383 (n550, n109);
buf  g384 (n551, n62);
not  g385 (n218, n157);
not  g386 (n541, n144);
buf  g387 (n438, n141);
buf  g388 (n197, n132);
buf  g389 (n353, n93);
not  g390 (n222, n44);
buf  g391 (n446, n112);
not  g392 (n237, n74);
not  g393 (n354, n81);
buf  g394 (n278, n111);
not  g395 (n418, n117);
not  g396 (n273, n119);
buf  g397 (n539, n73);
not  g398 (n174, n156);
not  g399 (n363, n108);
not  g400 (n323, n52);
buf  g401 (n568, n154);
buf  g402 (n667, n71);
not  g403 (n529, n100);
not  g404 (n572, n160);
not  g405 (n654, n72);
not  g406 (n427, n154);
not  g407 (n280, n123);
not  g408 (n642, n105);
buf  g409 (n342, n115);
not  g410 (n328, n151);
buf  g411 (n301, n59);
not  g412 (n286, n108);
buf  g413 (n200, n124);
not  g414 (n463, n36);
buf  g415 (n275, n58);
buf  g416 (n444, n55);
buf  g417 (n469, n91);
not  g418 (n599, n96);
not  g419 (n515, n95);
not  g420 (n306, n48);
buf  g421 (n641, n87);
buf  g422 (n349, n113);
buf  g423 (n413, n133);
buf  g424 (n575, n59);
not  g425 (n669, n141);
not  g426 (n215, n80);
not  g427 (n314, n61);
buf  g428 (n409, n101);
not  g429 (n341, n116);
buf  g430 (n626, n74);
buf  g431 (n188, n72);
buf  g432 (n394, n101);
not  g433 (n345, n88);
buf  g434 (n284, n137);
buf  g435 (n412, n47);
not  g436 (n260, n110);
not  g437 (n558, n123);
not  g438 (n600, n53);
buf  g439 (n351, n100);
not  g440 (n547, n73);
buf  g441 (n210, n71);
not  g442 (n660, n34);
not  g443 (n459, n51);
not  g444 (n447, n34);
not  g445 (n484, n148);
buf  g446 (n338, n55);
buf  g447 (n493, n36);
not  g448 (n192, n156);
buf  g449 (n410, n46);
not  g450 (n481, n131);
not  g451 (n624, n125);
not  g452 (n426, n53);
not  g453 (n211, n134);
buf  g454 (n332, n134);
buf  g455 (n364, n48);
buf  g456 (n313, n127);
not  g457 (n178, n65);
not  g458 (n252, n118);
not  g459 (n203, n136);
buf  g460 (n213, n79);
buf  g461 (n209, n43);
not  g462 (n406, n152);
not  g463 (n504, n50);
buf  g464 (n456, n81);
buf  g465 (n201, n93);
buf  g466 (n308, n109);
not  g467 (n625, n102);
not  g468 (n421, n49);
buf  g469 (n540, n42);
buf  g470 (n401, n66);
not  g471 (n205, n80);
not  g472 (n335, n66);
buf  g473 (n292, n149);
not  g474 (n567, n64);
not  g475 (n508, n63);
not  g476 (n161, n126);
buf  g477 (n322, n62);
not  g478 (n206, n144);
not  g479 (n640, n43);
not  g480 (n570, n65);
not  g481 (n378, n37);
buf  g482 (n562, n127);
not  g483 (n604, n80);
not  g484 (n334, n115);
buf  g485 (n535, n41);
buf  g486 (n472, n107);
not  g487 (n368, n115);
buf  g488 (n256, n112);
buf  g489 (n254, n60);
not  g490 (n615, n121);
not  g491 (n598, n56);
buf  g492 (n528, n131);
buf  g493 (n219, n84);
buf  g494 (n623, n121);
not  g495 (n443, n117);
buf  g496 (n451, n149);
not  g497 (n436, n131);
not  g498 (n576, n58);
not  g499 (n374, n117);
not  g500 (n379, n67);
buf  g501 (n476, n36);
not  g502 (n311, n76);
not  g503 (n276, n53);
buf  g504 (n473, n57);
buf  g505 (n404, n90);
buf  g506 (n434, n142);
buf  g507 (n503, n160);
buf  g508 (n176, n136);
buf  g509 (n168, n102);
buf  g510 (n362, n135);
buf  g511 (n411, n106);
not  g512 (n435, n69);
buf  g513 (n166, n138);
buf  g514 (n445, n82);
buf  g515 (n578, n51);
not  g516 (n648, n157);
not  g517 (n225, n148);
not  g518 (n318, n103);
buf  g519 (n606, n144);
not  g520 (n182, n94);
buf  g521 (n645, n99);
not  g522 (n238, n132);
buf  g523 (n173, n65);
not  g524 (n186, n153);
buf  g525 (n668, n96);
not  g526 (n271, n137);
buf  g527 (n207, n146);
buf  g528 (n580, n117);
buf  g529 (n348, n106);
not  g530 (n594, n56);
not  g531 (n454, n124);
not  g532 (n554, n77);
not  g533 (n357, n145);
buf  g534 (n226, n72);
buf  g535 (n266, n58);
buf  g536 (n375, n70);
not  g537 (n330, n123);
buf  g538 (n419, n151);
not  g539 (n523, n84);
buf  g540 (n537, n95);
buf  g541 (n439, n60);
not  g542 (n281, n92);
buf  g543 (n462, n113);
not  g544 (n442, n87);
buf  g545 (n458, n76);
buf  g546 (n383, n156);
not  g547 (n250, n49);
not  g548 (n485, n118);
buf  g549 (n326, n136);
not  g550 (n519, n88);
buf  g551 (n387, n47);
not  g552 (n253, n35);
not  g553 (n621, n62);
not  g554 (n597, n143);
not  g555 (n370, n115);
buf  g556 (n212, n96);
not  g557 (n198, n144);
not  g558 (n191, n101);
not  g559 (n184, n94);
buf  g560 (n236, n151);
buf  g561 (n356, n143);
buf  g562 (n670, n159);
not  g563 (n382, n51);
not  g564 (n607, n102);
buf  g565 (n288, n128);
not  g566 (n204, n45);
buf  g567 (n500, n90);
buf  g568 (n360, n104);
not  g569 (n384, n142);
buf  g570 (n588, n134);
not  g571 (n325, n138);
buf  g572 (n585, n70);
buf  g573 (n369, n128);
not  g574 (n227, n78);
not  g575 (n470, n85);
not  g576 (n608, n52);
not  g577 (n468, n133);
buf  g578 (n320, n65);
not  g579 (n502, n52);
not  g580 (n609, n121);
buf  g581 (n664, n85);
not  g582 (n643, n146);
buf  g583 (n520, n156);
buf  g584 (n518, n133);
buf  g585 (n629, n76);
buf  g586 (n264, n97);
not  g587 (n526, n34);
not  g588 (n232, n145);
buf  g589 (n441, n104);
buf  g590 (n657, n153);
not  g591 (n602, n33);
not  g592 (n636, n121);
not  g593 (n430, n49);
buf  g594 (n592, n159);
not  g595 (n343, n155);
buf  g596 (n616, n113);
not  g597 (n177, n99);
not  g598 (n234, n83);
buf  g599 (n270, n122);
buf  g600 (n393, n94);
not  g601 (n229, n91);
not  g602 (n612, n129);
buf  g603 (n511, n92);
buf  g604 (n295, n151);
not  g605 (n299, n77);
buf  g606 (n165, n58);
not  g607 (n637, n75);
not  g608 (n359, n146);
buf  g609 (n285, n148);
buf  g610 (n388, n52);
not  g611 (n397, n122);
buf  g612 (n392, n107);
not  g613 (n633, n129);
buf  g614 (n465, n37);
buf  g615 (n666, n33);
not  g616 (n542, n129);
not  g617 (n632, n107);
not  g618 (n265, n93);
not  g619 (n319, n103);
buf  g620 (n422, n39);
buf  g621 (n605, n61);
buf  g622 (n274, n72);
buf  g623 (n506, n159);
buf  g624 (n400, n114);
buf  g625 (n196, n128);
not  g626 (n268, n78);
not  g627 (n505, n37);
buf  g628 (n517, n96);
buf  g629 (n235, n153);
not  g630 (n407, n75);
buf  g631 (n507, n103);
buf  g632 (n202, n105);
not  g633 (n499, n160);
buf  g634 (n672, n138);
not  g635 (n663, n42);
buf  g636 (n289, n127);
not  g637 (n464, n125);
buf  g638 (n291, n97);
buf  g639 (n564, n111);
not  g640 (n700, n534);
buf  g641 (n773, n174);
not  g642 (n954, n345);
not  g643 (n1071, n273);
buf  g644 (n1008, n486);
not  g645 (n955, n421);
not  g646 (n763, n185);
not  g647 (n999, n524);
buf  g648 (n968, n375);
buf  g649 (n894, n422);
not  g650 (n809, n403);
buf  g651 (n729, n483);
buf  g652 (n1053, n298);
buf  g653 (n829, n382);
buf  g654 (n1003, n314);
not  g655 (n753, n428);
buf  g656 (n693, n516);
buf  g657 (n915, n536);
not  g658 (n797, n476);
buf  g659 (n767, n354);
not  g660 (n877, n467);
not  g661 (n690, n319);
buf  g662 (n985, n200);
buf  g663 (n959, n442);
not  g664 (n1041, n446);
not  g665 (n851, n285);
buf  g666 (n852, n208);
not  g667 (n1015, n242);
buf  g668 (n794, n368);
buf  g669 (n918, n272);
not  g670 (n715, n514);
buf  g671 (n726, n187);
buf  g672 (n1032, n253);
buf  g673 (n764, n463);
buf  g674 (n783, n209);
buf  g675 (n822, n231);
buf  g676 (n1021, n348);
buf  g677 (n845, n513);
buf  g678 (n774, n262);
not  g679 (n1045, n457);
not  g680 (n1027, n183);
buf  g681 (n953, n184);
not  g682 (n1054, n502);
not  g683 (n923, n531);
buf  g684 (n727, n468);
buf  g685 (n675, n373);
not  g686 (n880, n460);
buf  g687 (n867, n214);
not  g688 (n697, n286);
buf  g689 (n758, n432);
not  g690 (n738, n244);
buf  g691 (n1055, n230);
buf  g692 (n835, n473);
not  g693 (n1058, n414);
not  g694 (n1011, n453);
buf  g695 (n824, n362);
not  g696 (n722, n290);
buf  g697 (n1001, n498);
not  g698 (n814, n533);
not  g699 (n733, n255);
buf  g700 (n864, n393);
buf  g701 (n673, n211);
not  g702 (n1067, n515);
not  g703 (n833, n287);
not  g704 (n868, n392);
not  g705 (n747, n279);
not  g706 (n1046, n485);
not  g707 (n866, n249);
buf  g708 (n831, n376);
not  g709 (n889, n497);
buf  g710 (n930, n283);
buf  g711 (n805, n266);
buf  g712 (n964, n365);
not  g713 (n859, n271);
not  g714 (n1004, n532);
buf  g715 (n960, n327);
not  g716 (n827, n363);
buf  g717 (n744, n216);
buf  g718 (n854, n213);
buf  g719 (n749, n347);
not  g720 (n736, n530);
not  g721 (n810, n454);
not  g722 (n1009, n529);
not  g723 (n993, n406);
not  g724 (n931, n234);
not  g725 (n890, n201);
not  g726 (n1035, n489);
buf  g727 (n912, n461);
buf  g728 (n790, n338);
buf  g729 (n987, n504);
buf  g730 (n755, n371);
buf  g731 (n849, n381);
not  g732 (n881, n436);
not  g733 (n936, n202);
buf  g734 (n883, n512);
buf  g735 (n1013, n344);
not  g736 (n832, n491);
not  g737 (n788, n500);
buf  g738 (n1048, n204);
buf  g739 (n910, n260);
buf  g740 (n806, n387);
not  g741 (n847, n434);
buf  g742 (n1020, n488);
not  g743 (n804, n303);
buf  g744 (n989, n440);
buf  g745 (n1034, n189);
buf  g746 (n841, n477);
buf  g747 (n737, n337);
not  g748 (n780, n278);
not  g749 (n958, n173);
buf  g750 (n679, n317);
not  g751 (n1060, n296);
buf  g752 (n893, n443);
buf  g753 (n1023, n197);
buf  g754 (n978, n530);
buf  g755 (n696, n384);
buf  g756 (n922, n340);
not  g757 (n948, n289);
not  g758 (n848, n163);
buf  g759 (n969, n417);
not  g760 (n1002, n388);
not  g761 (n967, n261);
not  g762 (n1063, n179);
buf  g763 (n1044, n475);
not  g764 (n981, n229);
buf  g765 (n975, n207);
not  g766 (n798, n455);
not  g767 (n909, n535);
not  g768 (n811, n325);
buf  g769 (n911, n495);
buf  g770 (n863, n236);
not  g771 (n1018, n537);
buf  g772 (n1049, n416);
buf  g773 (n1037, n539);
buf  g774 (n896, n427);
buf  g775 (n762, n452);
not  g776 (n1069, n263);
buf  g777 (n674, n525);
buf  g778 (n1025, n302);
buf  g779 (n872, n171);
not  g780 (n971, n245);
not  g781 (n916, n275);
buf  g782 (n775, n259);
buf  g783 (n997, n175);
not  g784 (n897, n445);
not  g785 (n898, n458);
not  g786 (n904, n482);
buf  g787 (n940, n520);
buf  g788 (n836, n356);
buf  g789 (n907, n248);
not  g790 (n875, n450);
buf  g791 (n908, n394);
not  g792 (n839, n324);
not  g793 (n965, n526);
not  g794 (n741, n479);
not  g795 (n692, n227);
not  g796 (n1012, n243);
buf  g797 (n678, n168);
not  g798 (n956, n210);
buf  g799 (n941, n540);
buf  g800 (n751, n519);
buf  g801 (n998, n374);
buf  g802 (n884, n469);
buf  g803 (n947, n385);
buf  g804 (n717, n369);
buf  g805 (n681, n306);
not  g806 (n921, n328);
not  g807 (n823, n320);
not  g808 (n800, n499);
not  g809 (n702, n508);
not  g810 (n807, n444);
buf  g811 (n757, n531);
not  g812 (n1072, n294);
buf  g813 (n996, n330);
not  g814 (n705, n219);
not  g815 (n802, n258);
buf  g816 (n988, n527);
buf  g817 (n906, n507);
not  g818 (n920, n424);
not  g819 (n808, n170);
buf  g820 (n719, n288);
not  g821 (n934, n386);
not  g822 (n878, n191);
buf  g823 (n879, n308);
buf  g824 (n903, n505);
not  g825 (n830, n542);
buf  g826 (n976, n493);
buf  g827 (n787, n291);
buf  g828 (n682, n496);
buf  g829 (n932, n233);
buf  g830 (n984, n355);
buf  g831 (n957, n358);
not  g832 (n815, n465);
not  g833 (n778, n537);
buf  g834 (n687, n437);
not  g835 (n951, n357);
not  g836 (n739, n478);
not  g837 (n943, n380);
buf  g838 (n905, n256);
buf  g839 (n861, n218);
buf  g840 (n791, n538);
buf  g841 (n703, n269);
not  g842 (n695, n309);
buf  g843 (n1014, n438);
not  g844 (n748, n349);
not  g845 (n944, n223);
buf  g846 (n735, n529);
not  g847 (n761, n400);
not  g848 (n677, n359);
not  g849 (n723, n509);
buf  g850 (n980, n284);
not  g851 (n837, n487);
not  g852 (n777, n198);
buf  g853 (n718, n164);
not  g854 (n754, n402);
buf  g855 (n684, n464);
not  g856 (n768, n447);
not  g857 (n694, n451);
not  g858 (n874, n532);
buf  g859 (n942, n226);
buf  g860 (n766, n398);
not  g861 (n1059, n351);
buf  g862 (n732, n448);
buf  g863 (n812, n293);
not  g864 (n742, n503);
not  g865 (n986, n490);
not  g866 (n913, n364);
buf  g867 (n825, n439);
buf  g868 (n745, n339);
buf  g869 (n821, n276);
buf  g870 (n779, n366);
not  g871 (n970, n212);
buf  g872 (n994, n313);
not  g873 (n983, n418);
buf  g874 (n1064, n221);
buf  g875 (n873, n301);
not  g876 (n853, n166);
not  g877 (n979, n350);
not  g878 (n728, n295);
not  g879 (n899, n199);
buf  g880 (n928, n188);
not  g881 (n707, n270);
not  g882 (n721, n176);
buf  g883 (n1061, n312);
buf  g884 (n796, n186);
buf  g885 (n731, n541);
buf  g886 (n973, n472);
buf  g887 (n961, n419);
buf  g888 (n743, n523);
buf  g889 (n933, n220);
buf  g890 (n992, n430);
buf  g891 (n869, n336);
buf  g892 (n816, n280);
buf  g893 (n1016, n449);
buf  g894 (n871, n470);
buf  g895 (n1039, n541);
buf  g896 (n1066, n367);
not  g897 (n756, n435);
buf  g898 (n1030, n372);
not  g899 (n730, n177);
not  g900 (n919, n360);
not  g901 (n803, n192);
buf  g902 (n887, n322);
not  g903 (n1062, n361);
not  g904 (n925, n534);
buf  g905 (n760, n161);
buf  g906 (n1005, n539);
buf  g907 (n713, n235);
not  g908 (n949, n182);
buf  g909 (n819, n307);
not  g910 (n888, n407);
not  g911 (n750, n390);
not  g912 (n876, n169);
buf  g913 (n1000, n533);
buf  g914 (n937, n190);
buf  g915 (n846, n335);
not  g916 (n710, n389);
not  g917 (n1033, n353);
buf  g918 (n686, n540);
not  g919 (n1026, n459);
buf  g920 (n704, n250);
not  g921 (n711, n343);
not  g922 (n850, n492);
not  g923 (n716, n501);
buf  g924 (n1010, n441);
buf  g925 (n862, n535);
buf  g926 (n844, n517);
not  g927 (n901, n254);
not  g928 (n691, n267);
buf  g929 (n1029, n429);
not  g930 (n902, n195);
buf  g931 (n963, n274);
not  g932 (n927, n456);
buf  g933 (n689, n332);
not  g934 (n740, n480);
buf  g935 (n882, n425);
buf  g936 (n900, n412);
buf  g937 (n792, n474);
buf  g938 (n685, n240);
buf  g939 (n725, n224);
not  g940 (n772, n215);
not  g941 (n966, n178);
buf  g942 (n1068, n510);
buf  g943 (n746, n405);
not  g944 (n843, n318);
not  g945 (n1047, n399);
buf  g946 (n891, n206);
not  g947 (n813, n238);
buf  g948 (n683, n423);
not  g949 (n840, n408);
not  g950 (n1022, n391);
not  g951 (n860, n162);
buf  g952 (n781, n401);
buf  g953 (n770, n536);
buf  g954 (n771, n257);
buf  g955 (n1056, n481);
buf  g956 (n1040, n506);
not  g957 (n995, n232);
buf  g958 (n817, n310);
buf  g959 (n769, n377);
buf  g960 (n950, n528);
buf  g961 (n1065, n265);
buf  g962 (n820, n352);
not  g963 (n699, n341);
buf  g964 (n1050, n433);
buf  g965 (n782, n172);
buf  g966 (n789, n378);
buf  g967 (n680, n526);
buf  g968 (n982, n471);
not  g969 (n962, n268);
not  g970 (n924, n282);
not  g971 (n856, n297);
not  g972 (n676, n181);
buf  g973 (n795, n518);
not  g974 (n945, n299);
buf  g975 (n935, n311);
not  g976 (n776, n300);
buf  g977 (n885, n241);
not  g978 (n734, n346);
buf  g979 (n720, n521);
buf  g980 (n991, n194);
not  g981 (n1043, n522);
not  g982 (n708, n304);
buf  g983 (n842, n383);
not  g984 (n865, n409);
buf  g985 (n714, n395);
buf  g986 (n1006, n397);
buf  g987 (n1052, n484);
not  g988 (n1057, n203);
buf  g989 (n1042, n431);
buf  g990 (n818, n370);
buf  g991 (n886, n247);
buf  g992 (n1028, n277);
buf  g993 (n857, n426);
buf  g994 (n946, n411);
buf  g995 (n855, n329);
buf  g996 (n929, n225);
buf  g997 (n1024, n334);
buf  g998 (n938, n281);
buf  g999 (n765, n228);
buf  g1000 (n826, n323);
not  g1001 (n1036, n413);
not  g1002 (n917, n511);
buf  g1003 (n759, n305);
not  g1004 (n926, n239);
buf  g1005 (n914, n415);
buf  g1006 (n801, n462);
not  g1007 (n834, n252);
buf  g1008 (n870, n180);
buf  g1009 (n972, n196);
buf  g1010 (n892, n538);
not  g1011 (n895, n165);
not  g1012 (n784, n326);
buf  g1013 (n990, n342);
buf  g1014 (n752, n410);
buf  g1015 (n709, n331);
not  g1016 (n1007, n525);
not  g1017 (n1019, n217);
buf  g1018 (n1017, n193);
not  g1019 (n838, n527);
not  g1020 (n701, n420);
buf  g1021 (n724, n396);
buf  g1022 (n1031, n292);
buf  g1023 (n977, n466);
not  g1024 (n698, n222);
not  g1025 (n688, n237);
not  g1026 (n1070, n494);
not  g1027 (n799, n528);
not  g1028 (n786, n315);
buf  g1029 (n706, n246);
not  g1030 (n1038, n321);
not  g1031 (n974, n333);
not  g1032 (n952, n524);
buf  g1033 (n828, n167);
buf  g1034 (n712, n379);
buf  g1035 (n793, n264);
not  g1036 (n939, n316);
not  g1037 (n1051, n404);
buf  g1038 (n858, n205);
not  g1039 (n785, n251);
buf  g1040 (n1239, n738);
not  g1041 (n1274, n545);
not  g1042 (n1203, n570);
buf  g1043 (n1317, n1003);
buf  g1044 (n1342, n562);
not  g1045 (n1398, n679);
buf  g1046 (n1314, n838);
buf  g1047 (n1090, n596);
not  g1048 (n1305, n736);
buf  g1049 (n1256, n573);
not  g1050 (n1230, n590);
not  g1051 (n1341, n914);
buf  g1052 (n1293, n761);
not  g1053 (n1108, n564);
not  g1054 (n1073, n723);
not  g1055 (n1202, n1056);
buf  g1056 (n1158, n606);
buf  g1057 (n1119, n629);
not  g1058 (n1287, n623);
buf  g1059 (n1289, n1026);
not  g1060 (n1312, n568);
not  g1061 (n1360, n581);
buf  g1062 (n1179, n690);
not  g1063 (n1213, n543);
not  g1064 (n1078, n605);
not  g1065 (n1214, n1058);
not  g1066 (n1217, n903);
buf  g1067 (n1306, n926);
not  g1068 (n1221, n837);
buf  g1069 (n1376, n759);
buf  g1070 (n1304, n592);
not  g1071 (n1327, n577);
buf  g1072 (n1125, n937);
not  g1073 (n1294, n884);
not  g1074 (n1261, n825);
not  g1075 (n1393, n801);
buf  g1076 (n1083, n985);
not  g1077 (n1345, n606);
not  g1078 (n1207, n994);
not  g1079 (n1133, n607);
not  g1080 (n1338, n809);
buf  g1081 (n1173, n919);
not  g1082 (n1286, n1014);
not  g1083 (n1150, n885);
not  g1084 (n1302, n799);
buf  g1085 (n1372, n869);
buf  g1086 (n1243, n592);
not  g1087 (n1394, n932);
not  g1088 (n1124, n865);
buf  g1089 (n1153, n943);
not  g1090 (n1268, n558);
buf  g1091 (n1363, n864);
buf  g1092 (n1195, n610);
not  g1093 (n1190, n620);
not  g1094 (n1186, n599);
buf  g1095 (n1318, n603);
buf  g1096 (n1323, n621);
not  g1097 (n1188, n565);
buf  g1098 (n1194, n606);
buf  g1099 (n1353, n629);
not  g1100 (n1187, n897);
buf  g1101 (n1298, n879);
buf  g1102 (n1132, n548);
buf  g1103 (n1311, n682);
not  g1104 (n1365, n577);
buf  g1105 (n1369, n609);
buf  g1106 (n1351, n629);
not  g1107 (n1334, n728);
buf  g1108 (n1180, n614);
buf  g1109 (n1301, n575);
not  g1110 (n1216, n1030);
not  g1111 (n1185, n585);
buf  g1112 (n1160, n700);
buf  g1113 (n1210, n706);
buf  g1114 (n1196, n617);
not  g1115 (n1247, n600);
buf  g1116 (n1115, n992);
not  g1117 (n1355, n552);
not  g1118 (n1350, n588);
buf  g1119 (n1399, n621);
not  g1120 (n1255, n603);
not  g1121 (n1152, n750);
buf  g1122 (n1076, n712);
not  g1123 (n1277, n1025);
not  g1124 (n1122, n715);
not  g1125 (n1401, n563);
not  g1126 (n1381, n583);
not  g1127 (n1390, n1018);
not  g1128 (n1326, n610);
buf  g1129 (n1181, n576);
buf  g1130 (n1165, n611);
buf  g1131 (n1085, n588);
buf  g1132 (n1114, n891);
buf  g1133 (n1263, n615);
not  g1134 (n1144, n569);
buf  g1135 (n1379, n751);
not  g1136 (n1198, n900);
not  g1137 (n1176, n616);
buf  g1138 (n1143, n777);
buf  g1139 (n1370, n595);
buf  g1140 (n1319, n842);
not  g1141 (n1266, n560);
not  g1142 (n1206, n708);
not  g1143 (n1248, n957);
not  g1144 (n1358, n716);
not  g1145 (n1264, n574);
buf  g1146 (n1405, n959);
not  g1147 (n1250, n603);
not  g1148 (n1244, n1007);
buf  g1149 (n1192, n836);
buf  g1150 (n1077, n1015);
not  g1151 (n1320, n566);
buf  g1152 (n1356, n599);
not  g1153 (n1303, n752);
buf  g1154 (n1183, n1021);
buf  g1155 (n1099, n590);
buf  g1156 (n1283, n946);
buf  g1157 (n1328, n581);
not  g1158 (n1082, n1048);
buf  g1159 (n1092, n729);
not  g1160 (n1253, n560);
buf  g1161 (n1251, n969);
buf  g1162 (n1271, n857);
not  g1163 (n1138, n907);
not  g1164 (n1290, n810);
buf  g1165 (n1219, n798);
buf  g1166 (n1307, n727);
buf  g1167 (n1313, n621);
not  g1168 (n1162, n1041);
buf  g1169 (n1166, n827);
buf  g1170 (n1134, n570);
not  g1171 (n1352, n899);
buf  g1172 (n1205, n623);
not  g1173 (n1081, n734);
not  g1174 (n1086, n867);
not  g1175 (n1171, n614);
not  g1176 (n1238, n622);
buf  g1177 (n1330, n1053);
buf  g1178 (n1074, n576);
not  g1179 (n1172, n630);
not  g1180 (n1235, n692);
buf  g1181 (n1103, n905);
not  g1182 (n1224, n840);
not  g1183 (n1107, n619);
not  g1184 (n1395, n719);
not  g1185 (n1105, n894);
not  g1186 (n1333, n1010);
buf  g1187 (n1362, n846);
not  g1188 (n1371, n1055);
not  g1189 (n1299, n954);
buf  g1190 (n1391, n859);
buf  g1191 (n1109, n1000);
not  g1192 (n1111, n978);
buf  g1193 (n1354, n596);
buf  g1194 (n1339, n561);
buf  g1195 (n1278, n695);
not  g1196 (n1149, n592);
buf  g1197 (n1265, n902);
not  g1198 (n1335, n966);
not  g1199 (n1329, n841);
not  g1200 (n1367, n601);
buf  g1201 (n1118, n595);
buf  g1202 (n1136, n990);
buf  g1203 (n1240, n627);
not  g1204 (n1154, n549);
buf  g1205 (n1392, n680);
buf  g1206 (n1110, n698);
buf  g1207 (n1249, n862);
buf  g1208 (n1408, n845);
not  g1209 (n1101, n898);
not  g1210 (n1383, n1060);
not  g1211 (n1388, n1032);
buf  g1212 (n1084, n594);
buf  g1213 (n1325, n588);
not  g1214 (n1373, n604);
not  g1215 (n1361, n748);
buf  g1216 (n1273, n764);
not  g1217 (n1331, n811);
buf  g1218 (n1182, n558);
not  g1219 (n1223, n820);
buf  g1220 (n1272, n938);
buf  g1221 (n1100, n830);
buf  g1222 (n1275, n718);
not  g1223 (n1117, n585);
buf  g1224 (n1113, n624);
buf  g1225 (n1232, n623);
not  g1226 (n1102, n711);
buf  g1227 (n1245, n707);
not  g1228 (n1170, n609);
buf  g1229 (n1141, n694);
buf  g1230 (n1157, n852);
not  g1231 (n1279, n565);
not  g1232 (n1226, n608);
not  g1233 (n1262, n772);
buf  g1234 (n1295, n551);
buf  g1235 (n1079, n593);
buf  g1236 (n1116, n832);
not  g1237 (n1292, n574);
not  g1238 (n1280, n602);
not  g1239 (n1155, n601);
buf  g1240 (n1169, n747);
buf  g1241 (n1106, n818);
not  g1242 (n1343, n815);
buf  g1243 (n1258, n873);
buf  g1244 (n1241, n568);
buf  g1245 (n1231, n785);
buf  g1246 (n1296, n930);
not  g1247 (n1112, n1006);
buf  g1248 (n1297, n602);
buf  g1249 (n1178, n1051);
xnor g1250 (n1387, n742, n575);
xor  g1251 (n1167, n618, n596, n550, n620);
or   g1252 (n1212, n574, n923, n880, n1020);
nand g1253 (n1344, n631, n626, n545, n915);
xor  g1254 (n1075, n1027, n563, n721, n586);
nand g1255 (n1322, n553, n807, n566, n568);
xnor g1256 (n1254, n1009, n861, n724, n887);
xor  g1257 (n1346, n886, n678, n1036, n586);
or   g1258 (n1159, n816, n617, n975, n583);
and  g1259 (n1140, n717, n980, n1013, n608);
xor  g1260 (n1337, n570, n1042, n593, n605);
nand g1261 (n1161, n1044, n765, n560, n584);
xor  g1262 (n1189, n851, n600, n940, n740);
and  g1263 (n1229, n949, n597, n604, n850);
or   g1264 (n1128, n780, n703, n572, n1031);
xor  g1265 (n1242, n1046, n619, n624, n582);
nand g1266 (n1097, n1038, n753, n591, n843);
or   g1267 (n1281, n554, n1057, n689, n560);
nand g1268 (n1403, n855, n770, n598, n555);
xnor g1269 (n1168, n769, n577, n589, n854);
or   g1270 (n1347, n677, n573, n626, n584);
and  g1271 (n1409, n589, n918, n627, n792);
xnor g1272 (n1094, n609, n699, n1040, n702);
or   g1273 (n1359, n741, n601, n627, n578);
or   g1274 (n1267, n995, n797, n986, n758);
nor  g1275 (n1123, n916, n1024, n1059, n565);
xor  g1276 (n1121, n555, n629, n691, n547);
nand g1277 (n1375, n587, n1028, n973, n1029);
nand g1278 (n1321, n585, n970, n872, n876);
and  g1279 (n1237, n1005, n953, n630, n598);
nand g1280 (n1259, n543, n599, n906, n612);
xor  g1281 (n1236, n562, n860, n625, n1019);
nor  g1282 (n1201, n624, n768, n877, n583);
nand g1283 (n1300, n609, n910, n762, n613);
xor  g1284 (n1252, n882, n596, n971, n561);
xnor g1285 (n1131, n1050, n989, n697, n582);
xnor g1286 (n1386, n709, n788, n773, n968);
xnor g1287 (n1276, n604, n802, n608, n909);
or   g1288 (n1389, n1039, n890, n796, n547);
or   g1289 (n1324, n839, n813, n590, n591);
xor  g1290 (n1406, n573, n600, n579, n1047);
nor  g1291 (n1126, n996, n1004, n616, n722);
nand g1292 (n1377, n1023, n559, n988, n610);
or   g1293 (n1095, n1016, n912, n853, n917);
xnor g1294 (n1228, n725, n558, n812, n567);
nor  g1295 (n1404, n870, n952, n566, n615);
or   g1296 (n1089, n904, n597, n922, n929);
xor  g1297 (n1349, n763, n618, n571, n972);
xnor g1298 (n1316, n866, n1022, n720, n548);
xnor g1299 (n1220, n605, n630, n1012, n580);
nor  g1300 (n1315, n607, n620, n939, n774);
xnor g1301 (n1098, n550, n951, n594, n626);
or   g1302 (n1285, n616, n806, n829, n684);
nand g1303 (n1257, n618, n618, n622, n587);
or   g1304 (n1209, n673, n546, n579, n961);
nand g1305 (n1348, n793, n569, n881);
nand g1306 (n1407, n606, n625, n602, n598);
nor  g1307 (n1080, n749, n705, n626, n562);
nand g1308 (n1087, n575, n828, n566, n592);
nand g1309 (n1215, n760, n779, n790, n557);
or   g1310 (n1291, n831, n874, n544, n675);
and  g1311 (n1135, n580, n745, n617, n1052);
nand g1312 (n1184, n1054, n572, n931, n735);
xor  g1313 (n1309, n603, n947, n579, n974);
or   g1314 (n1233, n928, n571, n1017, n803);
xor  g1315 (n1127, n567, n743, n948, n580);
nand g1316 (n1175, n579, n936, n889, n800);
xnor g1317 (n1104, n895, n920, n559, n833);
and  g1318 (n1384, n896, n542, n925, n775);
and  g1319 (n1368, n622, n814, n688, n614);
nor  g1320 (n1129, n578, n977, n559, n781);
nor  g1321 (n1284, n569, n693, n732, n597);
nand g1322 (n1396, n623, n616, n962, n630);
xor  g1323 (n1282, n1049, n1033, n611, n587);
nor  g1324 (n1091, n935, n556, n1034, n1001);
nor  g1325 (n1310, n563, n888, n967, n584);
xor  g1326 (n1208, n613, n822, n982, n608);
nor  g1327 (n1191, n856, n588, n627, n1063);
xnor g1328 (n1139, n624, n578, n782, n871);
and  g1329 (n1142, n901, n805, n737, n776);
nor  g1330 (n1308, n614, n546, n963, n1002);
and  g1331 (n1222, n921, n625, n564, n934);
or   g1332 (n1364, n704, n600, n744, n585);
and  g1333 (n1148, n561, n981, n746, n754);
nand g1334 (n1374, n683, n848, n726, n984);
xnor g1335 (n1174, n933, n549, n858, n784);
and  g1336 (n1146, n574, n612, n983, n976);
xnor g1337 (n1193, n710, n586, n826, n787);
or   g1338 (n1332, n942, n821, n835, n687);
nand g1339 (n1385, n583, n615, n571, n572);
xnor g1340 (n1260, n573, n958, n587, n553);
xnor g1341 (n1199, n950, n575, n733, n927);
and  g1342 (n1204, n610, n544, n756, n991);
xor  g1343 (n1156, n619, n1043, n674, n696);
nor  g1344 (n1096, n789, n778, n713, n586);
and  g1345 (n1177, n834, n631, n577, n595);
and  g1346 (n1378, n617, n589, n701, n551);
nand g1347 (n1093, n960, n582, n911, n599);
xor  g1348 (n1234, n611, n844, n1008, n757);
or   g1349 (n1397, n924, n999, n681, n730);
xnor g1350 (n1088, n628, n823, n739, n731);
xor  g1351 (n1120, n572, n987, n621, n558);
and  g1352 (n1382, n590, n613, n941, n593);
nand g1353 (n1340, n993, n628, n998, n783);
nor  g1354 (n1366, n686, n567, n571);
nand g1355 (n1147, n561, n554, n628, n564);
xor  g1356 (n1227, n564, n997, n578, n1035);
or   g1357 (n1200, n611, n582, n594, n868);
nand g1358 (n1211, n965, n1061, n685, n956);
or   g1359 (n1269, n755, n615, n620, n619);
and  g1360 (n1137, n595, n604, n808, n622);
xnor g1361 (n1218, n557, n570, n1011, n607);
or   g1362 (n1246, n847, n591, n979, n568);
xor  g1363 (n1145, n1037, n824, n584, n607);
or   g1364 (n1225, n605, n791, n804, n1045);
and  g1365 (n1357, n767, n795, n676, n594);
or   g1366 (n1130, n612, n883, n559, n892);
and  g1367 (n1400, n576, n849, n955, n581);
xnor g1368 (n1288, n878, n593, n601, n786);
xnor g1369 (n1163, n863, n714, n625, n552);
xnor g1370 (n1164, n598, n964, n913, n563);
nor  g1371 (n1151, n556, n612, n613, n908);
or   g1372 (n1380, n771, n576, n565, n817);
nor  g1373 (n1336, n794, n819, n597, n589);
nand g1374 (n1270, n944, n893, n945, n602);
nor  g1375 (n1402, n581, n591, n875, n562);
or   g1376 (n1197, n1062, n766, n628, n580);
not  g1377 (n1411, n1074);
not  g1378 (n1410, n1073);
not  g1379 (n1418, n1410);
not  g1380 (n1416, n1411);
buf  g1381 (n1417, n1410);
not  g1382 (n1412, n1411);
not  g1383 (n1413, n1411);
not  g1384 (n1415, n1410);
buf  g1385 (n1414, n1410);
not  g1386 (n1419, n1411);
buf  g1387 (n1427, n1419);
buf  g1388 (n1430, n1412);
not  g1389 (n1445, n1415);
not  g1390 (n1446, n1416);
buf  g1391 (n1432, n1412);
not  g1392 (n1424, n1417);
buf  g1393 (n1442, n1418);
buf  g1394 (n1423, n1418);
not  g1395 (n1443, n1419);
buf  g1396 (n1451, n1417);
not  g1397 (n1448, n1413);
buf  g1398 (n1450, n1417);
not  g1399 (n1439, n1416);
not  g1400 (n1429, n1416);
buf  g1401 (n1431, n1419);
not  g1402 (n1437, n1413);
not  g1403 (n1420, n1414);
not  g1404 (n1425, n1413);
buf  g1405 (n1441, n1412);
not  g1406 (n1428, n1412);
buf  g1407 (n1438, n1415);
not  g1408 (n1422, n1415);
buf  g1409 (n1433, n1414);
buf  g1410 (n1434, n1416);
buf  g1411 (n1421, n1419);
buf  g1412 (n1435, n1413);
not  g1413 (n1436, n1414);
buf  g1414 (n1447, n1418);
buf  g1415 (n1440, n1415);
not  g1416 (n1449, n1417);
not  g1417 (n1426, n1414);
not  g1418 (n1444, n1418);
buf  g1419 (n1492, n1434);
not  g1420 (n1488, n1437);
not  g1421 (n1474, n1426);
not  g1422 (n1479, n1426);
not  g1423 (n1531, n1428);
buf  g1424 (n1483, n1422);
not  g1425 (n1491, n1092);
buf  g1426 (n1485, n1439);
buf  g1427 (n1481, n1079);
not  g1428 (n1522, n1432);
not  g1429 (n1528, n1431);
not  g1430 (n1482, n1105);
buf  g1431 (n1517, n1420);
not  g1432 (n1454, n1103);
buf  g1433 (n1525, n1076);
buf  g1434 (n1470, n1436);
buf  g1435 (n1530, n1436);
buf  g1436 (n1521, n1428);
not  g1437 (n1456, n1087);
not  g1438 (n1455, n1421);
not  g1439 (n1499, n1090);
not  g1440 (n1509, n1432);
buf  g1441 (n1480, n1110);
buf  g1442 (n1501, n1433);
not  g1443 (n1452, n1437);
not  g1444 (n1496, n1422);
not  g1445 (n1510, n1425);
not  g1446 (n1465, n1083);
buf  g1447 (n1506, n1437);
buf  g1448 (n1511, n1104);
buf  g1449 (n1489, n1107);
buf  g1450 (n1512, n1423);
buf  g1451 (n1497, n1427);
buf  g1452 (n1498, n1102);
not  g1453 (n1494, n1429);
buf  g1454 (n1500, n1427);
not  g1455 (n1463, n1429);
not  g1456 (n1507, n1100);
not  g1457 (n1487, n1075);
buf  g1458 (n1453, n1428);
buf  g1459 (n1459, n1429);
not  g1460 (n1526, n1112);
not  g1461 (n1493, n1438);
not  g1462 (n1515, n1426);
buf  g1463 (n1516, n1427);
buf  g1464 (n1490, n1425);
not  g1465 (n1462, n1081);
buf  g1466 (n1527, n1094);
buf  g1467 (n1529, n1420);
buf  g1468 (n1457, n1437);
buf  g1469 (n1514, n1420);
buf  g1470 (n1513, n1430);
buf  g1471 (n1471, n1082);
buf  g1472 (n1508, n1430);
not  g1473 (n1473, n1429);
buf  g1474 (n1468, n1424);
not  g1475 (n1518, n1089);
not  g1476 (n1484, n1431);
not  g1477 (n1460, n1435);
not  g1478 (n1464, n1435);
not  g1479 (n1475, n1434);
not  g1480 (n1505, n1439);
buf  g1481 (n1519, n1430);
buf  g1482 (n1476, n1099);
buf  g1483 (n1495, n1433);
not  g1484 (n1469, n1084);
nand g1485 (n1461, n1424, n1421, n1078);
nand g1486 (n1503, n1427, n1428, n1424);
nor  g1487 (n1524, n1106, n1095, n1433, n1085);
nor  g1488 (n1523, n1091, n1431, n1109, n1436);
and  g1489 (n1478, n1432, n1439, n1098, n1088);
xor  g1490 (n1458, n1093, n1101, n1438, n1435);
nor  g1491 (n1486, n1421, n1114, n1433, n1080);
xor  g1492 (n1466, n1430, n1434, n1432);
xor  g1493 (n1477, n1096, n1423, n1420, n1113);
nand g1494 (n1472, n1436, n1086, n1077, n1422);
or   g1495 (n1467, n1423, n1424, n1438, n1426);
xor  g1496 (n1504, n1421, n1422, n1425);
xor  g1497 (n1520, n1435, n1108, n1111, n1423);
xor  g1498 (n1502, n1438, n1439, n1431, n1097);
buf  g1499 (n1603, n1475);
buf  g1500 (n1580, n1458);
not  g1501 (n1600, n1458);
not  g1502 (n1563, n1464);
not  g1503 (n1565, n1468);
not  g1504 (n1572, n1452);
buf  g1505 (n1553, n1461);
not  g1506 (n1560, n1457);
buf  g1507 (n1559, n1469);
not  g1508 (n1557, n1470);
buf  g1509 (n1545, n1455);
buf  g1510 (n1574, n1474);
not  g1511 (n1558, n1461);
buf  g1512 (n1570, n1476);
buf  g1513 (n1575, n1463);
not  g1514 (n1583, n1462);
buf  g1515 (n1599, n1473);
not  g1516 (n1541, n1476);
buf  g1517 (n1589, n1458);
buf  g1518 (n1571, n1461);
buf  g1519 (n1601, n1471);
not  g1520 (n1594, n1453);
buf  g1521 (n1536, n1472);
not  g1522 (n1587, n1115);
buf  g1523 (n1591, n1476);
buf  g1524 (n1547, n1457);
not  g1525 (n1538, n1117);
buf  g1526 (n1554, n1453);
buf  g1527 (n1567, n1468);
buf  g1528 (n1562, n1467);
not  g1529 (n1555, n1474);
not  g1530 (n1576, n1471);
buf  g1531 (n1537, n1468);
buf  g1532 (n1566, n1467);
buf  g1533 (n1581, n1460);
buf  g1534 (n1564, n1463);
not  g1535 (n1535, n1457);
not  g1536 (n1579, n1455);
buf  g1537 (n1533, n1478);
buf  g1538 (n1532, n1452);
not  g1539 (n1577, n1456);
not  g1540 (n1604, n1464);
buf  g1541 (n1550, n1474);
not  g1542 (n1573, n1466);
not  g1543 (n1539, n1477);
not  g1544 (n1543, n1469);
buf  g1545 (n1534, n1463);
not  g1546 (n1596, n1473);
not  g1547 (n1548, n1469);
buf  g1548 (n1542, n1460);
not  g1549 (n1540, n1463);
buf  g1550 (n1546, n1476);
buf  g1551 (n1585, n1472);
buf  g1552 (n1578, n1453);
buf  g1553 (n1569, n1459);
not  g1554 (n1584, n1475);
buf  g1555 (n1593, n1455);
buf  g1556 (n1590, n1454);
not  g1557 (n1598, n1473);
buf  g1558 (n1586, n1465);
not  g1559 (n1556, n1465);
xor  g1560 (n1588, n1116, n1465, n1477);
nand g1561 (n1561, n1470, n1464, n1475);
and  g1562 (n1595, n1457, n1460, n1473, n1455);
xnor g1563 (n1549, n1454, n1462, n1477, n1460);
xor  g1564 (n1552, n1456, n1459, n1467, n1453);
nand g1565 (n1568, n1472, n1466, n1461, n1467);
or   g1566 (n1597, n1462, n1471, n1456, n1468);
and  g1567 (n1551, n1470, n1454, n1477, n1466);
or   g1568 (n1602, n1456, n1454, n1452, n1471);
nor  g1569 (n1592, n1459, n1452, n1469, n1474);
nand g1570 (n1582, n1466, n1462, n1464, n1465);
and  g1571 (n1544, n1470, n1472, n1458, n1459);
not  g1572 (n1679, n1132);
not  g1573 (n1646, n1586);
buf  g1574 (n1658, n1511);
buf  g1575 (n1686, n1492);
not  g1576 (n1607, n1126);
buf  g1577 (n1609, n1517);
buf  g1578 (n1653, n1512);
not  g1579 (n1635, n1494);
not  g1580 (n1696, n1554);
not  g1581 (n1689, n1524);
not  g1582 (n1608, n1580);
not  g1583 (n1637, n1545);
buf  g1584 (n1684, n1491);
buf  g1585 (n1639, n1522);
not  g1586 (n1663, n1566);
buf  g1587 (n1627, n1586);
not  g1588 (n1638, n1507);
buf  g1589 (n1659, n1589);
not  g1590 (n1629, n1511);
not  g1591 (n1662, n1501);
and  g1592 (n1687, n1481, n1524, n1492, n1129);
and  g1593 (n1676, n1509, n1478, n1555, n1523);
nand g1594 (n1693, n1507, n1584, n1581, n1514);
xnor g1595 (n1672, n1519, n1490, n1526, n1478);
nand g1596 (n1669, n1482, n1494, n1512, n1496);
or   g1597 (n1652, n1571, n1485, n1505, n1483);
or   g1598 (n1690, n1505, n1493, n1508, n1492);
or   g1599 (n1614, n1501, n1496, n1514, n1587);
nor  g1600 (n1622, n1520, n1499, n1490, n1567);
xnor g1601 (n1680, n1503, n1122, n1121, n1480);
nand g1602 (n1677, n1479, n1481, n1583, n1534);
and  g1603 (n1628, n1529, n1510, n1487, n1584);
xor  g1604 (n1681, n1489, n1519, n1588, n1508);
nand g1605 (n1617, n1528, n1576, n1517, n1590);
and  g1606 (n1651, n1484, n1542, n1521, n1483);
xor  g1607 (n1695, n1519, n1540, n1506, n1580);
and  g1608 (n1656, n1568, n1518, n1575, n1502);
nand g1609 (n1642, n1585, n1480, n1508, n1131);
nand g1610 (n1645, n1482, n1548, n1520, n1500);
nand g1611 (n1694, n1488, n1510, n1521, n1529);
and  g1612 (n1654, n1498, n1479, n1513, n1586);
nand g1613 (n1623, n1585, n1479, n1504, n1513);
or   g1614 (n1644, n1486, n1492, n1584, n1512);
or   g1615 (n1649, n1558, n1130, n1507, n1497);
and  g1616 (n1606, n1118, n1498, n1541, n1556);
nand g1617 (n1674, n1587, n1573, n1510, n1518);
nand g1618 (n1634, n1588, n1503, n1580, n1518);
xnor g1619 (n1698, n1481, n1583, n1523, n1120);
and  g1620 (n1605, n1498, n1489, n1516, n1124);
nand g1621 (n1616, n1127, n1128, n1487, n1582);
and  g1622 (n1671, n1495, n1535, n1516, n1577);
nor  g1623 (n1631, n1549, n1494, n1516, n1501);
xor  g1624 (n1648, n1486, n1485, n1588, n1581);
or   g1625 (n1613, n1552, n1504, n1510, n1500);
xnor g1626 (n1688, n1504, n1480, n1520, n1563);
nand g1627 (n1640, n1481, n1496, n1482, n1581);
nand g1628 (n1683, n1550, n1509, n1484, n1580);
and  g1629 (n1667, n1582, n1557, n1479, n1525);
xor  g1630 (n1630, n1520, n1483, n1125, n1583);
xnor g1631 (n1685, n1559, n1582, n1524, n1511);
nand g1632 (n1610, n1502, n1123, n1527, n1509);
and  g1633 (n1675, n1482, n1589, n1517, n1490);
xnor g1634 (n1641, n1489, n1514, n1519, n1505);
and  g1635 (n1620, n1525, n1547, n1565, n1488);
nand g1636 (n1650, n1529, n1506, n1527, n1119);
nand g1637 (n1615, n1537, n1526, n1578, n1528);
xor  g1638 (n1660, n1551, n1536, n1513, n1572);
or   g1639 (n1697, n1487, n1587, n1544, n1574);
nand g1640 (n1611, n1582, n1502, n1590, n1503);
xor  g1641 (n1670, n1579, n1494, n1515, n1507);
xor  g1642 (n1691, n1570, n1583, n1503, n1521);
nor  g1643 (n1664, n1488, n1589, n1501);
or   g1644 (n1625, n1579, n1483, n1485, n1588);
xor  g1645 (n1673, n1522, n1521, n1584, n1515);
xnor g1646 (n1692, n1533, n1497, n1553, n1539);
and  g1647 (n1666, n1525, n1491, n1513, n1515);
nor  g1648 (n1624, n1527, n1512, n1500, n1499);
nand g1649 (n1636, n1560, n1491, n1480, n1514);
nand g1650 (n1626, n1569, n1527, n1516, n1489);
nor  g1651 (n1665, n1587, n1511, n1585, n1495);
or   g1652 (n1633, n1499, n1505, n1522, n1538);
or   g1653 (n1655, n1522, n1586, n1523, n1562);
nor  g1654 (n1618, n1133, n1561, n1518, n1523);
and  g1655 (n1678, n1500, n1532, n1485, n1525);
and  g1656 (n1643, n1487, n1484, n1546, n1509);
xor  g1657 (n1647, n1578, n1493, n1484, n1515);
nand g1658 (n1657, n1488, n1526, n1590, n1478);
nor  g1659 (n1632, n1495, n1493, n1564, n1491);
xor  g1660 (n1682, n1506, n1517, n1590, n1528);
nand g1661 (n1661, n1498, n1486, n1497);
and  g1662 (n1619, n1585, n1495, n1493, n1581);
xor  g1663 (n1668, n1524, n1496, n1526, n1499);
nor  g1664 (n1612, n1504, n1497, n1502, n1543);
or   g1665 (n1621, n1490, n1508, n1506, n1528);
xor  g1666 (n1726, n1068, n1070);
and  g1667 (n1725, n1646, n1635, n1067, n1667);
and  g1668 (n1705, n1628, n1441, n1446);
nand g1669 (n1699, n1448, n1638, n1069, n1451);
xnor g1670 (n1733, n1608, n1451, n1449, n1606);
or   g1671 (n1701, n1448, n1444, n1140, n1445);
xnor g1672 (n1708, n1443, n1443, n1142, n1144);
or   g1673 (n1731, n1065, n1629, n1447, n1449);
nor  g1674 (n1721, n1449, n1150, n1149, n1447);
and  g1675 (n1719, n1611, n1066, n1446, n1445);
xor  g1676 (n1709, n1146, n1639, n1448, n1441);
and  g1677 (n1728, n1444, n1664, n1644, n1656);
or   g1678 (n1734, n1632, n1625, n1450, n1663);
xnor g1679 (n1732, n1607, n1440, n1647, n1652);
and  g1680 (n1713, n1451, n1444, n1634, n1605);
xnor g1681 (n1714, n1654, n1446, n1442, n1138);
xnor g1682 (n1704, n1657, n1630, n1151, n1614);
or   g1683 (n1735, n1669, n1665, n1445, n1640);
and  g1684 (n1729, n1137, n1441, n1620, n1135);
nor  g1685 (n1710, n1666, n1141, n1653, n1147);
xnor g1686 (n1711, n1623, n1450, n1661, n1442);
and  g1687 (n1707, n1670, n1626, n1659, n1627);
xnor g1688 (n1715, n1668, n1442, n1622);
nand g1689 (n1702, n1631, n1529, n1609, n1443);
xnor g1690 (n1722, n1443, n1649, n1530, n1134);
and  g1691 (n1716, n1671, n1148, n1645, n1651);
xor  g1692 (n1730, n1448, n1641, n1447, n1643);
or   g1693 (n1712, n1610, n1444, n1660, n1619);
nand g1694 (n1703, n1145, n1624, n1449, n1618);
nand g1695 (n1718, n1617, n1530, n1136, n1658);
and  g1696 (n1723, n1637, n1662, n1615, n1064);
nand g1697 (n1717, n1440, n1451, n1621, n1655);
nand g1698 (n1700, n1616, n1139, n1441, n1530);
xnor g1699 (n1706, n1445, n1633, n1450, n1447);
and  g1700 (n1727, n1612, n1440, n1143, n1650);
nand g1701 (n1720, n1636, n1530, n1450, n1613);
and  g1702 (n1724, n1440, n1642, n1648, n1531);
not  g1703 (n1739, n1706);
buf  g1704 (n1742, n1700);
not  g1705 (n1736, n1707);
not  g1706 (n1745, n1708);
not  g1707 (n1743, n1531);
buf  g1708 (n1738, n1703);
buf  g1709 (n1740, n1531);
buf  g1710 (n1741, n1701);
not  g1711 (n1744, n1705);
buf  g1712 (n1737, n1702);
or   g1713 (n1746, n1704, n1709, n1710, n1531);
xor  g1714 (n1774, n1156, n1742);
or   g1715 (n1775, n1598, n1680, n1591, n1741);
and  g1716 (n1772, n1739, n1600, n1591, n1602);
nor  g1717 (n1757, n1602, n1695, n1688, n1154);
xor  g1718 (n1760, n1596, n1693, n1601, n1597);
nand g1719 (n1752, n1683, n1602, n1593, n1597);
and  g1720 (n1750, n1685, n1673, n1594, n1743);
xor  g1721 (n1773, n1692, n1594, n1601, n1746);
nand g1722 (n1776, n1743, n1698, n1737, n1740);
and  g1723 (n1768, n1679, n1600, n1593, n1677);
xnor g1724 (n1762, n1746, n1596, n1745, n1744);
xnor g1725 (n1766, n1603, n1592, n1152, n1678);
nor  g1726 (n1765, n1744, n1742, n1675, n1592);
or   g1727 (n1767, n1601, n1596, n1604, n1595);
nand g1728 (n1749, n1593, n1744, n1691, n1736);
xor  g1729 (n1769, n1697, n1742, n1599, n1672);
xor  g1730 (n1754, n1598, n1597, n1599, n1600);
xnor g1731 (n1755, n1682, n1604, n1684, n1592);
xnor g1732 (n1758, n1743, n1741, n1599, n1745);
xnor g1733 (n1761, n1686, n1595, n1604, n1694);
and  g1734 (n1771, n1153, n1740, n1746, n1743);
and  g1735 (n1763, n1592, n1600, n1594, n1696);
xor  g1736 (n1770, n1604, n1687, n1745, n1598);
nand g1737 (n1753, n1597, n1738, n1599, n1603);
nor  g1738 (n1747, n1594, n1746, n1690, n1744);
nor  g1739 (n1764, n1681, n1603, n1595, n1742);
xor  g1740 (n1759, n1603, n1601, n1689, n1596);
nor  g1741 (n1748, n1591, n1741, n1595, n1674);
nand g1742 (n1751, n1593, n1155, n1676, n1745);
nand g1743 (n1756, n1591, n1598, n1741, n1602);
buf  g1744 (n1783, n1772);
not  g1745 (n1785, n1774);
not  g1746 (n1788, n1771);
not  g1747 (n1786, n1775);
not  g1748 (n1778, n1765);
buf  g1749 (n1782, n1767);
buf  g1750 (n1780, n1768);
buf  g1751 (n1777, n1766);
buf  g1752 (n1781, n1773);
buf  g1753 (n1779, n1769);
not  g1754 (n1787, n1770);
not  g1755 (n1784, n1776);
xor  g1756 (n1791, n1714, n1728, n1779, n1160);
xor  g1757 (n1794, n1785, n1720, n1163, n1158);
nor  g1758 (n1798, n1785, n1174, n1730, n1711);
or   g1759 (n1801, n1168, n1780, n1731, n1735);
and  g1760 (n1797, n1165, n1733, n1779, n1778);
xnor g1761 (n1808, n1780, n1785, n1167, n1172);
xnor g1762 (n1809, n1718, n1180, n1782, n1171);
or   g1763 (n1806, n1779, n1783, n1781, n1170);
xnor g1764 (n1792, n1159, n1782, n1726, n1713);
nand g1765 (n1807, n1785, n1169, n1175, n1777);
and  g1766 (n1804, n1780, n1725, n1178, n1781);
xnor g1767 (n1793, n1717, n1729, n1783, n1162);
xor  g1768 (n1803, n1179, n1778, n1157, n1782);
xor  g1769 (n1805, n1783, n1777, n1173, n1716);
nor  g1770 (n1790, n1712, n1721, n1166, n1161);
xor  g1771 (n1799, n1780, n1781, n1176, n1734);
nor  g1772 (n1796, n1783, n1715, n1784, n1778);
nor  g1773 (n1800, n1732, n1181, n1177, n1722);
nand g1774 (n1789, n1724, n1779, n1164, n1719);
nand g1775 (n1795, n1723, n1784, n1782);
or   g1776 (n1802, n1727, n1784, n1781, n1778);
buf  g1777 (n1813, n1798);
buf  g1778 (n1811, n1797);
buf  g1779 (n1812, n1796);
buf  g1780 (n1810, n1799);
buf  g1781 (n1825, n1801);
buf  g1782 (n1822, n1810);
buf  g1783 (n1827, n1811);
buf  g1784 (n1814, n1813);
not  g1785 (n1816, n1810);
not  g1786 (n1828, n1811);
not  g1787 (n1815, n1811);
not  g1788 (n1821, n1810);
buf  g1789 (n1824, n1800);
buf  g1790 (n1829, n1812);
buf  g1791 (n1826, n1813);
buf  g1792 (n1818, n1811);
not  g1793 (n1819, n1812);
not  g1794 (n1817, n1812);
buf  g1795 (n1820, n1812);
xnor g1796 (n1823, n1810, n1813);
xor  g1797 (n1847, n661, n1816, n647, n1819);
xor  g1798 (n1878, n665, n640, n662, n658);
xor  g1799 (n1842, n668, n646, n644, n633);
nand g1800 (n1877, n641, n1824, n1814, n1787);
xnor g1801 (n1869, n1817, n655, n1819, n663);
or   g1802 (n1890, n669, n644, n663, n656);
or   g1803 (n1848, n660, n639, n1809, n638);
xor  g1804 (n1882, n671, n658, n646, n631);
xnor g1805 (n1888, n1808, n1822, n1828, n670);
nand g1806 (n1830, n1828, n650, n639, n672);
xor  g1807 (n1854, n1827, n644, n646, n637);
or   g1808 (n1840, n670, n648, n1786, n643);
nor  g1809 (n1889, n1820, n1828, n643, n633);
xor  g1810 (n1850, n669, n631, n656, n671);
nor  g1811 (n1863, n1823, n1825, n1818, n641);
or   g1812 (n1872, n641, n1820, n1829);
and  g1813 (n1873, n1788, n640, n662, n1820);
xor  g1814 (n1838, n1827, n1825, n1816, n646);
or   g1815 (n1876, n665, n648, n636, n1823);
xnor g1816 (n1851, n1815, n647, n642, n658);
or   g1817 (n1875, n635, n637, n670, n1804);
or   g1818 (n1831, n1803, n666, n636, n1818);
xor  g1819 (n1846, n656, n645, n666, n651);
nor  g1820 (n1874, n645, n638, n658, n657);
nand g1821 (n1870, n1817, n637, n653, n659);
xor  g1822 (n1864, n652, n642, n639, n654);
xnor g1823 (n1880, n1829, n1788, n652);
xnor g1824 (n1867, n657, n1828, n638, n669);
xnor g1825 (n1865, n1815, n653, n636, n654);
or   g1826 (n1856, n647, n1787, n661, n668);
xnor g1827 (n1833, n634, n643, n640, n653);
xnor g1828 (n1855, n1826, n650, n1814, n1787);
and  g1829 (n1839, n648, n653, n637, n649);
xor  g1830 (n1860, n1820, n634, n664, n671);
nand g1831 (n1862, n640, n1802, n1827, n633);
and  g1832 (n1841, n651, n635, n1786, n1829);
nand g1833 (n1859, n651, n1786, n667, n660);
or   g1834 (n1879, n636, n1788, n668, n1817);
nand g1835 (n1852, n665, n655, n668, n1825);
or   g1836 (n1885, n635, n654, n632, n657);
xnor g1837 (n1845, n662, n1826, n651, n652);
and  g1838 (n1883, n1827, n1815, n635, n663);
or   g1839 (n1861, n663, n1822, n659);
xor  g1840 (n1837, n1819, n648, n666, n655);
xnor g1841 (n1881, n660, n649, n647, n1817);
nor  g1842 (n1849, n672, n645, n664, n671);
xnor g1843 (n1836, n1826, n1807, n650, n1821);
xnor g1844 (n1853, n664, n654, n662, n1787);
or   g1845 (n1868, n664, n667, n665);
xnor g1846 (n1834, n1825, n1821, n1824, n1816);
xor  g1847 (n1843, n1821, n643, n1805, n656);
or   g1848 (n1891, n659, n661, n1786, n633);
nor  g1849 (n1886, n649, n639, n1826, n672);
and  g1850 (n1832, n1824, n652, n1819, n661);
and  g1851 (n1866, n641, n642, n660, n1822);
nor  g1852 (n1857, n1823, n670, n1818, n634);
and  g1853 (n1884, n669, n657, n1824, n644);
and  g1854 (n1871, n667, n650, n1815, n666);
xor  g1855 (n1858, n638, n632, n659, n1806);
nand g1856 (n1835, n645, n1821, n632, n634);
nor  g1857 (n1844, n672, n632, n1823, n649);
and  g1858 (n1887, n1816, n642, n1818, n655);
not  g1859 (n1895, n1842);
buf  g1860 (n1908, n1846);
not  g1861 (n1911, n1832);
buf  g1862 (n1914, n1849);
buf  g1863 (n1907, n1833);
buf  g1864 (n1913, n1844);
not  g1865 (n1892, n1839);
buf  g1866 (n1906, n1853);
buf  g1867 (n1905, n1843);
buf  g1868 (n1893, n1838);
buf  g1869 (n1909, n1835);
not  g1870 (n1912, n1847);
buf  g1871 (n1904, n1845);
not  g1872 (n1900, n1834);
not  g1873 (n1902, n1830);
buf  g1874 (n1903, n1837);
not  g1875 (n1899, n1848);
buf  g1876 (n1901, n1852);
buf  g1877 (n1910, n1831);
not  g1878 (n1898, n1841);
buf  g1879 (n1897, n1851);
buf  g1880 (n1894, n1836);
buf  g1881 (n1915, n1840);
not  g1882 (n1896, n1850);
xor  g1883 (n1986, n1878, n1264, n1265, n1320);
xnor g1884 (n1964, n1194, n1203, n1865, n1915);
and  g1885 (n1960, n1899, n1912, n1895, n1906);
nor  g1886 (n1998, n1248, n1205, n1237, n1392);
nand g1887 (n1971, n1888, n1369, n1884, n1905);
and  g1888 (n1988, n1390, n1277, n1196, n1912);
xnor g1889 (n1990, n1221, n1879, n1882, n1210);
xor  g1890 (n1963, n1356, n1298, n1363, n1301);
nand g1891 (n1935, n1380, n1399, n1326, n1329);
nand g1892 (n1954, n1308, n1349, n1292, n1283);
nor  g1893 (n2003, n1281, n1244, n1198, n1314);
xor  g1894 (n1993, n1900, n1286, n1216, n1360);
or   g1895 (n1917, n1903, n1330, n1209, n1266);
nand g1896 (n1992, n1239, n1911, n1893, n1913);
nand g1897 (n1983, n1187, n1893, n1328, n1185);
nand g1898 (n1936, n1318, n1261, n1232, n1391);
xor  g1899 (n1942, n1895, n1206, n1212, n1910);
and  g1900 (n1922, n1347, n1897, n1406, n1309);
xnor g1901 (n1957, n1912, n1891, n1903, n1337);
xnor g1902 (n1965, n1395, n1348, n1355, n1350);
nor  g1903 (n2002, n1352, n1905, n1249, n1189);
nor  g1904 (n1920, n1370, n1302, n1898, n1268);
or   g1905 (n1969, n1195, n1873, n1907, n1361);
nor  g1906 (n1926, n1885, n1307, n1344, n1894);
nand g1907 (n1927, n1234, n1276, n1906, n1898);
xnor g1908 (n2004, n1304, n1902, n1910, n1345);
xor  g1909 (n1995, n1914, n1217, n1315, n1378);
nand g1910 (n1947, n1252, n1389, n1339, n1243);
and  g1911 (n1946, n1904, n1887, n1897, n1208);
xor  g1912 (n1974, n1306, n1250, n1338, n1229);
xor  g1913 (n1916, n1321, n1908, n1311, n1316);
nor  g1914 (n1938, n1880, n1898, n1859, n1335);
or   g1915 (n1945, n1071, n1227, n1883, n1379);
or   g1916 (n1961, n1364, n1377, n1904, n1257);
nor  g1917 (n1940, n1362, n1211, n1342, n1331);
and  g1918 (n1962, n1192, n1854, n1907, n1341);
xor  g1919 (n1996, n1263, n1228, n1327, n1199);
or   g1920 (n1932, n1224, n1313, n1894, n1274);
or   g1921 (n1978, n1897, n1905, n1384);
and  g1922 (n1979, n1855, n1319, n1365, n1915);
xor  g1923 (n1959, n1381, n1900, n1351, n1397);
xor  g1924 (n1976, n1317, n1402, n1374, n1219);
xor  g1925 (n1956, n1911, n1909, n1889, n1275);
xor  g1926 (n1999, n1220, n1282, n1393, n1353);
xor  g1927 (n1921, n1225, n1269, n1183, n1895);
nor  g1928 (n1968, n1182, n1914, n1201, n1901);
xnor g1929 (n1967, n1914, n1200, n1901, n1387);
nor  g1930 (n1985, n1407, n1408, n1354, n1291);
xor  g1931 (n1952, n1911, n1215, n1897, n1278);
and  g1932 (n1981, n1388, n1874, n1902, n1253);
nor  g1933 (n1966, n1197, n1207, n1403, n1204);
nor  g1934 (n1950, n1863, n1072, n1289, n1218);
nor  g1935 (n1918, n1396, n1190, n1913, n1231);
xor  g1936 (n1939, n1258, n1398, n1270, n1896);
xnor g1937 (n1955, n1272, n1366, n1322, n1906);
xnor g1938 (n1937, n1247, n1385, n1902, n1358);
xor  g1939 (n1941, n1235, n1903, n1236, n1909);
nand g1940 (n1949, n1899, n1899, n1284, n1188);
nor  g1941 (n2001, n1359, n1324, n1271, n1909);
or   g1942 (n1989, n1896, n1246, n1295, n1226);
nor  g1943 (n1933, n1186, n1273, n1202, n1871);
xor  g1944 (n1924, n1310, n1213, n1373, n1346);
nand g1945 (n2000, n1886, n1908, n1233);
and  g1946 (n1991, n1368, n1858, n1294, n1223);
xnor g1947 (n1951, n1312, n1193, n1372, n1915);
nor  g1948 (n1982, n1912, n1357, n1892, n1383);
nor  g1949 (n1997, n1241, n1296, n1267, n1903);
and  g1950 (n1973, n1861, n1881, n1256, n1191);
nand g1951 (n1994, n1240, n1242, n1222, n1890);
nand g1952 (n1929, n1259, n1899, n1913, n1904);
nand g1953 (n1987, n1367, n1305, n1376, n1299);
nor  g1954 (n1984, n1405, n1867, n1340, n1870);
nor  g1955 (n1980, n1303, n1857, n1287, n1913);
xor  g1956 (n1948, n1915, n1907, n1394, n1293);
xor  g1957 (n1953, n1914, n1375, n1901, n1251);
nand g1958 (n1928, n1868, n1872, n1386, n1895);
xnor g1959 (n1919, n1906, n1334, n1255, n1910);
or   g1960 (n1944, n1404, n1904, n1901, n1285);
or   g1961 (n1970, n1401, n1288, n1910, n1869);
xor  g1962 (n1975, n1238, n1254, n1184, n1896);
xnor g1963 (n1958, n1862, n1911, n1262, n1400);
xor  g1964 (n1925, n1900, n1214, n1290, n1902);
xnor g1965 (n1934, n1877, n1260, n1245, n1900);
or   g1966 (n1931, n1896, n1909, n1876, n1332);
or   g1967 (n1972, n1875, n1371, n1866, n1860);
xor  g1968 (n1930, n1297, n1908, n1280, n1856);
nor  g1969 (n1923, n1279, n1343, n1325, n1300);
xor  g1970 (n1943, n1336, n1898, n1382, n1333);
xnor g1971 (n1977, n1864, n1230, n1323, n1907);
or   g1972 (n2015, n1958, n1964, n1963, n1984);
xor  g1973 (n2008, n1955, n1981, n1973, n1934);
nor  g1974 (n2023, n1918, n1960, n1924, n1944);
xor  g1975 (n2005, n1994, n1940, n1971, n1916);
xnor g1976 (n2016, n1979, n1941, n1953, n1983);
xnor g1977 (n2026, n1956, n1990, n1967, n1945);
xor  g1978 (n2017, n1966, n1989, n1969, n1985);
nor  g1979 (n2013, n1937, n1954, n1949, n1977);
xor  g1980 (n2009, n1975, n1947, n1970, n1926);
nor  g1981 (n2024, n1929, n1939, n1957, n1972);
xnor g1982 (n2022, n1946, n1932, n1952, n1925);
and  g1983 (n2019, n1988, n1993, n1961, n1923);
nand g1984 (n2010, n1995, n1920, n1997, n1980);
and  g1985 (n2011, n1938, n1992, n1986, n1942);
nor  g1986 (n2007, n1919, n2002, n1943, n1930);
nor  g1987 (n2025, n1948, n1968, n1921, n1409);
nor  g1988 (n2020, n1965, n1976, n2000, n1987);
xor  g1989 (n2014, n1951, n1996, n1936, n2001);
nor  g1990 (n2012, n1928, n1982, n1922, n1950);
xnor g1991 (n2021, n1999, n1917, n1927, n1933);
or   g1992 (n2018, n1959, n1998, n1991, n1978);
nor  g1993 (n2006, n1962, n1974, n1931, n1935);
or   g1994 (n2031, n2023, n2017, n2021, n2025);
or   g1995 (n2032, n2015, n2019, n2003, n2010);
nor  g1996 (n2027, n2004, n2008, n2012, n2005);
nor  g1997 (n2030, n2007, n2013, n2024, n2026);
or   g1998 (n2028, n2022, n2009, n2016, n2020);
xor  g1999 (n2029, n2018, n2011, n2014, n2006);
endmodule
