

module Stat_100_53
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n100,
  n93,
  n80,
  n114,
  n99,
  n110,
  n107,
  n92,
  n84,
  n86,
  n79,
  n115,
  n91,
  n95,
  n88,
  n112,
  n117,
  n89,
  n132,
  n129,
  n120,
  n124,
  n128,
  n127,
  n125,
  n123,
  n119,
  n126,
  n122,
  n121,
  n131,
  n130
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n100;output n93;output n80;output n114;output n99;output n110;output n107;output n92;output n84;output n86;output n79;output n115;output n91;output n95;output n88;output n112;output n117;output n89;output n132;output n129;output n120;output n124;output n128;output n127;output n125;output n123;output n119;output n126;output n122;output n121;output n131;output n130;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n81;wire n82;wire n83;wire n85;wire n87;wire n90;wire n94;wire n96;wire n97;wire n98;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n108;wire n109;wire n111;wire n113;wire n116;wire n118;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;

  not
  g0
  (
    n41,
    n2
  );


  buf
  g1
  (
    n36,
    n2
  );


  not
  g2
  (
    KeyWire_0_15,
    n1
  );


  buf
  g3
  (
    KeyWire_0_5,
    n1
  );


  buf
  g4
  (
    n39,
    n2
  );


  buf
  g5
  (
    n34,
    n3
  );


  not
  g6
  (
    n42,
    n1
  );


  not
  g7
  (
    n38,
    n2
  );


  buf
  g8
  (
    n40,
    n3
  );


  not
  g9
  (
    n33,
    n1
  );


  not
  g10
  (
    n50,
    n33
  );


  not
  g11
  (
    n47,
    n34
  );


  buf
  g12
  (
    n48,
    n34
  );


  buf
  g13
  (
    KeyWire_0_14,
    n33
  );


  buf
  g14
  (
    n45,
    n33
  );


  buf
  g15
  (
    n49,
    n34
  );


  buf
  g16
  (
    n43,
    n34
  );


  buf
  g17
  (
    n44,
    n33
  );


  buf
  g18
  (
    n57,
    n45
  );


  buf
  g19
  (
    n67,
    n49
  );


  buf
  g20
  (
    n61,
    n43
  );


  buf
  g21
  (
    n51,
    n44
  );


  buf
  g22
  (
    n52,
    n46
  );


  buf
  g23
  (
    n55,
    n48
  );


  not
  g24
  (
    n53,
    n44
  );


  buf
  g25
  (
    n65,
    n35
  );


  not
  g26
  (
    n64,
    n47
  );


  buf
  g27
  (
    KeyWire_0_0,
    n44
  );


  not
  g28
  (
    n56,
    n45
  );


  buf
  g29
  (
    n63,
    n47
  );


  xor
  g30
  (
    n66,
    n44,
    n48
  );


  nor
  g31
  (
    n54,
    n46,
    n47
  );


  or
  g32
  (
    n59,
    n35,
    n35,
    n43,
    n48
  );


  nand
  g33
  (
    n62,
    n47,
    n45,
    n35,
    n46
  );


  nor
  g34
  (
    n68,
    n43,
    n43,
    n48,
    n49
  );


  xor
  g35
  (
    n60,
    n46,
    n36,
    n45
  );


  xor
  g36
  (
    n92,
    n62,
    n6
  );


  and
  g37
  (
    n94,
    n64,
    n29,
    n3,
    n32
  );


  nand
  g38
  (
    n70,
    n20,
    n67,
    n12,
    n32
  );


  xnor
  g39
  (
    n97,
    n67,
    n11,
    n30,
    n7
  );


  nor
  g40
  (
    n80,
    n15,
    n51,
    n29,
    n8
  );


  xnor
  g41
  (
    n91,
    n17,
    n61,
    n4
  );


  or
  g42
  (
    KeyWire_0_12,
    n51,
    n49,
    n18,
    n50
  );


  xor
  g43
  (
    n89,
    n56,
    n54,
    n27,
    n14
  );


  or
  g44
  (
    n109,
    n16,
    n36,
    n60,
    n15
  );


  nor
  g45
  (
    KeyWire_0_3,
    n59,
    n10,
    n54,
    n12
  );


  nor
  g46
  (
    KeyWire_0_4,
    n67,
    n50,
    n15,
    n55
  );


  xnor
  g47
  (
    KeyWire_0_7,
    n26,
    n16,
    n27,
    n20
  );


  and
  g48
  (
    KeyWire_0_8,
    n25,
    n64,
    n24,
    n58
  );


  or
  g49
  (
    n110,
    n63,
    n9,
    n22,
    n68
  );


  or
  g50
  (
    n99,
    n50,
    n6,
    n51,
    n8
  );


  xnor
  g51
  (
    n118,
    n68,
    n16,
    n14,
    n11
  );


  xor
  g52
  (
    n108,
    n10,
    n5,
    n66,
    n28
  );


  xnor
  g53
  (
    n82,
    n13,
    n57,
    n32,
    n7
  );


  nor
  g54
  (
    KeyWire_0_9,
    n10,
    n23,
    n63,
    n58
  );


  and
  g55
  (
    n77,
    n13,
    n64,
    n14,
    n62
  );


  nor
  g56
  (
    n93,
    n22,
    n24,
    n57,
    n66
  );


  or
  g57
  (
    n71,
    n23,
    n8,
    n18,
    n59
  );


  xnor
  g58
  (
    n105,
    n60,
    n64,
    n9,
    n4
  );


  nor
  g59
  (
    n69,
    n65,
    n26,
    n66,
    n21
  );


  and
  g60
  (
    n112,
    n25,
    n55,
    n59,
    n23
  );


  xnor
  g61
  (
    n98,
    n36,
    n49,
    n63,
    n8
  );


  xor
  g62
  (
    n88,
    n57,
    n12,
    n62,
    n18
  );


  and
  g63
  (
    n115,
    n52,
    n60,
    n25
  );


  xnor
  g64
  (
    n85,
    n18,
    n21,
    n50,
    n5
  );


  xnor
  g65
  (
    n102,
    n25,
    n7,
    n13,
    n26
  );


  or
  g66
  (
    n79,
    n61,
    n21,
    n27,
    n52
  );


  and
  g67
  (
    n96,
    n61,
    n55,
    n4,
    n30
  );


  nor
  g68
  (
    n74,
    n23,
    n59,
    n30
  );


  xor
  g69
  (
    KeyWire_0_6,
    n53,
    n62,
    n29,
    n10
  );


  and
  g70
  (
    n101,
    n21,
    n4,
    n58,
    n13
  );


  xnor
  g71
  (
    KeyWire_0_10,
    n54,
    n56,
    n31,
    n65
  );


  or
  g72
  (
    KeyWire_0_11,
    n52,
    n31,
    n54,
    n9
  );


  xor
  g73
  (
    n76,
    n22,
    n6,
    n67,
    n17
  );


  and
  g74
  (
    n73,
    n20,
    n15,
    n11,
    n19
  );


  or
  g75
  (
    n117,
    n65,
    n28,
    n5,
    n14
  );


  or
  g76
  (
    n114,
    n29,
    n31,
    n26,
    n68
  );


  and
  g77
  (
    n83,
    n17,
    n19,
    n58
  );


  nand
  g78
  (
    n104,
    n55,
    n5,
    n11,
    n53
  );


  or
  g79
  (
    n75,
    n17,
    n63,
    n22,
    n9
  );


  xnor
  g80
  (
    KeyWire_0_1,
    n56,
    n27,
    n28,
    n66
  );


  or
  g81
  (
    KeyWire_0_13,
    n56,
    n3,
    n53,
    n65
  );


  nor
  g82
  (
    n87,
    n32,
    n53,
    n68,
    n24
  );


  nor
  g83
  (
    n78,
    n57,
    n24,
    n31,
    n52
  );


  or
  g84
  (
    n90,
    n20,
    n7,
    n19,
    n6
  );


  nand
  g85
  (
    n81,
    n16,
    n51,
    n12,
    n28
  );


  nor
  g86
  (
    n129,
    n102,
    n41,
    n42
  );


  and
  g87
  (
    n127,
    n40,
    n106,
    n110,
    n88
  );


  nor
  g88
  (
    KeyWire_0_2,
    n91,
    n38,
    n101,
    n117
  );


  xor
  g89
  (
    n119,
    n94,
    n90,
    n92,
    n111
  );


  nand
  g90
  (
    n132,
    n98,
    n118,
    n37,
    n113
  );


  xor
  g91
  (
    n120,
    n95,
    n38,
    n87,
    n89
  );


  nor
  g92
  (
    n125,
    n93,
    n41,
    n42
  );


  and
  g93
  (
    n126,
    n103,
    n97,
    n38,
    n37
  );


  and
  g94
  (
    n128,
    n40,
    n37,
    n38,
    n115
  );


  xor
  g95
  (
    n131,
    n40,
    n41,
    n104,
    n109
  );


  xor
  g96
  (
    n121,
    n105,
    n41,
    n116,
    n114
  );


  and
  g97
  (
    n123,
    n39,
    n39,
    n107,
    n99
  );


  nor
  g98
  (
    n122,
    n112,
    n37,
    n108,
    n39
  );


  and
  g99
  (
    n130,
    n40,
    n39,
    n96,
    n100
  );


  xor
  KeyGate_0_0
  (
    n58,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n100,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n124,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n113,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n116,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n37,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n111,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n95,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n107,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n84,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n86,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n103,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n72,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n106,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n46,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n35,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


