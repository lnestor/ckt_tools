// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_226 written by SynthGen on 2021/04/05 11:23:26
module Stat_2000_226( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n739, n715, n1183, n1173, n1169, n1179, n1175, n1194,
 n1188, n1196, n1177, n1185, n1167, n1187, n1408, n1424,
 n1412, n1418, n1423, n1395, n1425, n1403, n1396, n1401,
 n1397, n1393, n1426, n1415, n1411, n1406, n2031, n2032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n739, n715, n1183, n1173, n1169, n1179, n1175, n1194,
 n1188, n1196, n1177, n1185, n1167, n1187, n1408, n1424,
 n1412, n1418, n1423, n1395, n1425, n1403, n1396, n1401,
 n1397, n1393, n1426, n1415, n1411, n1406, n2031, n2032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1168, n1170, n1171, n1172,
 n1174, n1176, n1178, n1180, n1181, n1182, n1184, n1186,
 n1189, n1190, n1191, n1192, n1193, n1195, n1197, n1198,
 n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
 n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
 n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
 n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
 n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
 n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
 n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
 n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
 n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
 n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
 n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
 n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
 n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
 n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
 n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
 n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
 n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
 n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
 n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
 n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
 n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
 n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
 n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
 n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
 n1391, n1392, n1394, n1398, n1399, n1400, n1402, n1404,
 n1405, n1407, n1409, n1410, n1413, n1414, n1416, n1417,
 n1419, n1420, n1421, n1422, n1427, n1428, n1429, n1430,
 n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
 n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
 n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
 n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
 n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
 n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
 n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
 n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
 n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
 n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
 n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
 n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
 n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
 n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
 n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
 n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
 n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
 n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
 n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
 n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
 n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
 n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
 n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
 n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
 n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
 n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
 n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
 n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
 n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
 n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
 n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
 n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
 n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
 n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
 n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
 n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
 n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
 n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
 n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
 n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
 n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
 n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
 n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
 n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
 n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
 n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
 n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
 n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
 n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
 n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
 n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
 n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
 n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
 n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
 n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
 n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
 n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
 n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
 n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
 n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
 n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
 n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
 n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
 n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
 n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
 n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
 n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
 n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
 n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
 n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
 n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
 n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
 n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
 n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
 n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030;

buf  g0 (n80, n32);
buf  g1 (n36, n4);
not  g2 (n35, n20);
not  g3 (n92, n28);
buf  g4 (n34, n15);
buf  g5 (n58, n23);
buf  g6 (n67, n7);
not  g7 (n123, n16);
not  g8 (n158, n1);
buf  g9 (n146, n6);
buf  g10 (n127, n32);
not  g11 (n82, n10);
not  g12 (n39, n12);
not  g13 (n62, n1);
not  g14 (n68, n8);
buf  g15 (n33, n22);
not  g16 (n156, n17);
not  g17 (n72, n10);
buf  g18 (n97, n24);
not  g19 (n77, n14);
buf  g20 (n154, n11);
buf  g21 (n87, n11);
buf  g22 (n139, n3);
not  g23 (n116, n2);
buf  g24 (n69, n19);
not  g25 (n151, n29);
not  g26 (n132, n16);
not  g27 (n101, n3);
buf  g28 (n88, n7);
buf  g29 (n38, n20);
buf  g30 (n118, n24);
not  g31 (n112, n3);
buf  g32 (n145, n25);
not  g33 (n100, n26);
buf  g34 (n138, n12);
not  g35 (n147, n20);
not  g36 (n81, n5);
buf  g37 (n129, n31);
buf  g38 (n160, n9);
not  g39 (n61, n14);
not  g40 (n109, n27);
buf  g41 (n78, n2);
buf  g42 (n65, n7);
buf  g43 (n89, n9);
not  g44 (n152, n8);
not  g45 (n55, n21);
not  g46 (n153, n10);
not  g47 (n108, n17);
buf  g48 (n90, n25);
not  g49 (n50, n23);
not  g50 (n121, n29);
buf  g51 (n111, n19);
not  g52 (n45, n17);
not  g53 (n110, n28);
buf  g54 (n122, n31);
not  g55 (n49, n9);
buf  g56 (n75, n31);
buf  g57 (n143, n25);
not  g58 (n119, n5);
not  g59 (n157, n26);
not  g60 (n128, n14);
not  g61 (n98, n22);
not  g62 (n148, n4);
not  g63 (n79, n24);
buf  g64 (n76, n15);
buf  g65 (n142, n18);
not  g66 (n43, n21);
not  g67 (n117, n10);
buf  g68 (n94, n22);
buf  g69 (n124, n28);
not  g70 (n113, n32);
buf  g71 (n74, n2);
not  g72 (n93, n24);
not  g73 (n115, n29);
buf  g74 (n137, n26);
not  g75 (n114, n14);
not  g76 (n63, n18);
not  g77 (n99, n13);
buf  g78 (n103, n26);
not  g79 (n107, n11);
not  g80 (n136, n5);
not  g81 (n125, n18);
not  g82 (n85, n4);
buf  g83 (n53, n29);
buf  g84 (n149, n9);
buf  g85 (n71, n4);
buf  g86 (n130, n6);
buf  g87 (n84, n23);
not  g88 (n54, n15);
buf  g89 (n150, n1);
buf  g90 (n83, n32);
buf  g91 (n140, n7);
buf  g92 (n70, n16);
buf  g93 (n41, n28);
not  g94 (n133, n12);
not  g95 (n59, n19);
not  g96 (n47, n13);
buf  g97 (n52, n11);
not  g98 (n56, n6);
buf  g99 (n51, n15);
not  g100 (n126, n30);
not  g101 (n106, n2);
not  g102 (n96, n21);
buf  g103 (n134, n19);
not  g104 (n46, n8);
buf  g105 (n44, n13);
not  g106 (n42, n30);
not  g107 (n104, n22);
not  g108 (n91, n5);
buf  g109 (n73, n1);
buf  g110 (n135, n3);
not  g111 (n64, n21);
not  g112 (n105, n25);
not  g113 (n48, n18);
not  g114 (n120, n16);
not  g115 (n141, n12);
buf  g116 (n131, n27);
not  g117 (n57, n30);
not  g118 (n37, n20);
not  g119 (n95, n30);
not  g120 (n60, n17);
buf  g121 (n40, n6);
buf  g122 (n144, n23);
buf  g123 (n159, n8);
buf  g124 (n66, n31);
buf  g125 (n155, n27);
buf  g126 (n102, n27);
not  g127 (n86, n13);
not  g128 (n292, n97);
not  g129 (n227, n143);
not  g130 (n652, n36);
not  g131 (n593, n46);
not  g132 (n226, n33);
buf  g133 (n286, n58);
buf  g134 (n208, n113);
not  g135 (n329, n39);
not  g136 (n231, n50);
buf  g137 (n243, n119);
buf  g138 (n238, n76);
buf  g139 (n449, n123);
buf  g140 (n589, n147);
buf  g141 (n366, n65);
not  g142 (n453, n66);
not  g143 (n300, n151);
not  g144 (n585, n33);
buf  g145 (n565, n153);
buf  g146 (n483, n77);
buf  g147 (n256, n159);
not  g148 (n628, n60);
buf  g149 (n202, n47);
not  g150 (n295, n37);
buf  g151 (n450, n114);
not  g152 (n595, n100);
not  g153 (n323, n101);
buf  g154 (n327, n113);
not  g155 (n291, n110);
not  g156 (n415, n126);
not  g157 (n284, n73);
buf  g158 (n165, n66);
buf  g159 (n599, n152);
not  g160 (n426, n124);
not  g161 (n511, n156);
not  g162 (n161, n146);
not  g163 (n663, n105);
not  g164 (n220, n157);
not  g165 (n367, n53);
buf  g166 (n425, n108);
buf  g167 (n169, n56);
not  g168 (n413, n95);
not  g169 (n167, n137);
buf  g170 (n640, n130);
not  g171 (n390, n131);
not  g172 (n513, n128);
not  g173 (n478, n126);
not  g174 (n424, n152);
buf  g175 (n171, n149);
not  g176 (n358, n44);
buf  g177 (n222, n50);
buf  g178 (n351, n70);
not  g179 (n214, n51);
buf  g180 (n297, n83);
buf  g181 (n491, n89);
not  g182 (n409, n45);
not  g183 (n439, n88);
not  g184 (n287, n94);
not  g185 (n645, n119);
not  g186 (n400, n118);
buf  g187 (n320, n120);
buf  g188 (n257, n47);
buf  g189 (n401, n154);
buf  g190 (n641, n100);
buf  g191 (n268, n146);
not  g192 (n212, n144);
not  g193 (n592, n130);
not  g194 (n606, n74);
not  g195 (n211, n93);
buf  g196 (n228, n72);
buf  g197 (n532, n72);
not  g198 (n411, n74);
buf  g199 (n482, n132);
buf  g200 (n240, n111);
not  g201 (n210, n84);
buf  g202 (n234, n36);
not  g203 (n190, n135);
not  g204 (n246, n79);
buf  g205 (n551, n44);
buf  g206 (n617, n97);
not  g207 (n388, n60);
buf  g208 (n659, n139);
not  g209 (n379, n154);
buf  g210 (n340, n74);
not  g211 (n625, n125);
buf  g212 (n492, n108);
buf  g213 (n163, n53);
buf  g214 (n229, n160);
buf  g215 (n441, n54);
buf  g216 (n455, n160);
not  g217 (n376, n80);
not  g218 (n354, n45);
not  g219 (n555, n106);
not  g220 (n255, n106);
buf  g221 (n578, n56);
buf  g222 (n557, n58);
not  g223 (n414, n42);
not  g224 (n462, n141);
buf  g225 (n536, n105);
not  g226 (n573, n115);
not  g227 (n479, n85);
not  g228 (n363, n135);
not  g229 (n259, n143);
not  g230 (n473, n99);
buf  g231 (n359, n72);
buf  g232 (n576, n131);
not  g233 (n647, n45);
not  g234 (n371, n41);
buf  g235 (n331, n114);
buf  g236 (n584, n70);
buf  g237 (n525, n157);
not  g238 (n362, n121);
buf  g239 (n270, n82);
not  g240 (n260, n92);
not  g241 (n446, n123);
not  g242 (n199, n122);
buf  g243 (n189, n64);
buf  g244 (n375, n101);
not  g245 (n484, n86);
buf  g246 (n445, n95);
buf  g247 (n644, n135);
not  g248 (n530, n100);
not  g249 (n187, n33);
buf  g250 (n466, n101);
not  g251 (n296, n117);
not  g252 (n254, n109);
not  g253 (n216, n54);
buf  g254 (n539, n36);
not  g255 (n407, n57);
buf  g256 (n468, n63);
not  g257 (n316, n61);
not  g258 (n274, n85);
buf  g259 (n639, n78);
buf  g260 (n381, n132);
buf  g261 (n281, n116);
buf  g262 (n408, n46);
not  g263 (n612, n54);
buf  g264 (n634, n120);
not  g265 (n494, n83);
buf  g266 (n197, n38);
buf  g267 (n633, n52);
not  g268 (n501, n81);
not  g269 (n609, n61);
not  g270 (n604, n49);
not  g271 (n384, n98);
not  g272 (n527, n42);
not  g273 (n572, n142);
not  g274 (n267, n121);
buf  g275 (n389, n133);
not  g276 (n334, n84);
not  g277 (n614, n158);
buf  g278 (n568, n155);
not  g279 (n613, n34);
not  g280 (n324, n156);
buf  g281 (n518, n46);
not  g282 (n338, n91);
buf  g283 (n514, n138);
not  g284 (n396, n98);
buf  g285 (n248, n110);
buf  g286 (n404, n56);
not  g287 (n262, n159);
not  g288 (n556, n40);
not  g289 (n610, n41);
not  g290 (n304, n102);
not  g291 (n350, n141);
not  g292 (n183, n123);
buf  g293 (n538, n127);
buf  g294 (n658, n121);
buf  g295 (n526, n41);
buf  g296 (n637, n55);
not  g297 (n280, n129);
not  g298 (n176, n114);
not  g299 (n269, n60);
buf  g300 (n651, n48);
buf  g301 (n193, n103);
not  g302 (n213, n144);
not  g303 (n397, n81);
not  g304 (n469, n150);
not  g305 (n326, n57);
buf  g306 (n600, n58);
buf  g307 (n310, n129);
buf  g308 (n422, n62);
buf  g309 (n219, n100);
not  g310 (n186, n97);
not  g311 (n205, n97);
not  g312 (n626, n49);
not  g313 (n447, n45);
buf  g314 (n412, n43);
buf  g315 (n416, n92);
not  g316 (n662, n59);
not  g317 (n464, n116);
buf  g318 (n622, n118);
not  g319 (n596, n95);
buf  g320 (n583, n75);
buf  g321 (n571, n131);
not  g322 (n488, n68);
buf  g323 (n548, n92);
not  g324 (n430, n82);
not  g325 (n343, n148);
buf  g326 (n545, n77);
not  g327 (n522, n34);
buf  g328 (n177, n133);
not  g329 (n303, n113);
buf  g330 (n348, n153);
not  g331 (n289, n52);
not  g332 (n239, n111);
buf  g333 (n458, n151);
not  g334 (n657, n65);
not  g335 (n448, n71);
buf  g336 (n503, n67);
buf  g337 (n519, n96);
buf  g338 (n523, n77);
not  g339 (n423, n109);
not  g340 (n386, n125);
not  g341 (n436, n74);
buf  g342 (n339, n75);
not  g343 (n504, n51);
not  g344 (n342, n34);
buf  g345 (n271, n93);
buf  g346 (n623, n39);
buf  g347 (n475, n88);
buf  g348 (n463, n114);
buf  g349 (n299, n147);
buf  g350 (n322, n111);
buf  g351 (n654, n35);
not  g352 (n452, n81);
not  g353 (n586, n94);
buf  g354 (n290, n69);
buf  g355 (n636, n63);
buf  g356 (n166, n57);
buf  g357 (n627, n38);
buf  g358 (n170, n109);
buf  g359 (n670, n115);
not  g360 (n440, n136);
buf  g361 (n629, n78);
buf  g362 (n650, n78);
buf  g363 (n476, n76);
not  g364 (n500, n64);
buf  g365 (n582, n63);
buf  g366 (n454, n89);
buf  g367 (n498, n87);
buf  g368 (n417, n90);
not  g369 (n508, n102);
buf  g370 (n383, n136);
not  g371 (n451, n117);
not  g372 (n369, n140);
buf  g373 (n567, n59);
not  g374 (n574, n70);
buf  g375 (n587, n104);
buf  g376 (n217, n86);
buf  g377 (n509, n124);
buf  g378 (n378, n71);
buf  g379 (n672, n148);
buf  g380 (n178, n36);
buf  g381 (n370, n64);
buf  g382 (n624, n144);
not  g383 (n631, n72);
not  g384 (n361, n106);
buf  g385 (n353, n53);
not  g386 (n546, n49);
buf  g387 (n278, n130);
not  g388 (n428, n150);
buf  g389 (n314, n133);
not  g390 (n225, n67);
not  g391 (n258, n108);
buf  g392 (n543, n89);
buf  g393 (n288, n88);
buf  g394 (n360, n110);
buf  g395 (n605, n119);
buf  g396 (n620, n91);
not  g397 (n632, n137);
not  g398 (n419, n107);
buf  g399 (n549, n159);
not  g400 (n434, n35);
not  g401 (n251, n94);
not  g402 (n164, n132);
not  g403 (n666, n67);
buf  g404 (n664, n121);
buf  g405 (n431, n149);
buf  g406 (n497, n104);
buf  g407 (n520, n124);
not  g408 (n279, n96);
not  g409 (n201, n145);
not  g410 (n465, n87);
buf  g411 (n250, n157);
buf  g412 (n328, n145);
buf  g413 (n560, n93);
buf  g414 (n275, n69);
buf  g415 (n437, n62);
not  g416 (n444, n71);
not  g417 (n649, n39);
not  g418 (n380, n84);
not  g419 (n377, n91);
buf  g420 (n182, n151);
not  g421 (n398, n107);
not  g422 (n364, n146);
buf  g423 (n619, n68);
buf  g424 (n427, n126);
buf  g425 (n387, n69);
not  g426 (n559, n80);
not  g427 (n318, n124);
not  g428 (n661, n101);
buf  g429 (n198, n112);
not  g430 (n655, n59);
not  g431 (n438, n83);
buf  g432 (n588, n55);
not  g433 (n341, n151);
not  g434 (n347, n134);
buf  g435 (n306, n90);
not  g436 (n276, n75);
buf  g437 (n204, n70);
not  g438 (n352, n96);
buf  g439 (n506, n145);
buf  g440 (n293, n35);
buf  g441 (n495, n87);
buf  g442 (n315, n34);
not  g443 (n597, n57);
buf  g444 (n537, n155);
buf  g445 (n496, n110);
buf  g446 (n313, n153);
not  g447 (n611, n140);
buf  g448 (n577, n85);
not  g449 (n528, n112);
buf  g450 (n552, n62);
buf  g451 (n547, n47);
not  g452 (n311, n128);
not  g453 (n391, n122);
not  g454 (n206, n55);
not  g455 (n283, n73);
not  g456 (n590, n103);
not  g457 (n481, n105);
not  g458 (n249, n119);
buf  g459 (n245, n145);
buf  g460 (n180, n132);
not  g461 (n667, n135);
not  g462 (n235, n102);
not  g463 (n515, n125);
not  g464 (n172, n128);
buf  g465 (n418, n50);
not  g466 (n173, n61);
buf  g467 (n194, n98);
not  g468 (n221, n75);
buf  g469 (n393, n152);
not  g470 (n233, n37);
not  g471 (n558, n83);
buf  g472 (n541, n80);
not  g473 (n207, n60);
not  g474 (n247, n42);
not  g475 (n472, n94);
not  g476 (n564, n86);
not  g477 (n325, n65);
not  g478 (n184, n76);
not  g479 (n531, n87);
buf  g480 (n507, n84);
buf  g481 (n365, n103);
buf  g482 (n668, n115);
not  g483 (n385, n40);
not  g484 (n242, n40);
buf  g485 (n540, n138);
not  g486 (n332, n159);
buf  g487 (n648, n155);
buf  g488 (n550, n56);
not  g489 (n357, n108);
buf  g490 (n218, n139);
not  g491 (n298, n106);
buf  g492 (n456, n157);
buf  g493 (n580, n143);
buf  g494 (n485, n107);
not  g495 (n554, n156);
not  g496 (n224, n150);
not  g497 (n669, n149);
buf  g498 (n253, n127);
buf  g499 (n534, n129);
not  g500 (n282, n120);
not  g501 (n294, n96);
not  g502 (n591, n141);
buf  g503 (n467, n141);
not  g504 (n368, n78);
not  g505 (n460, n128);
not  g506 (n330, n147);
buf  g507 (n374, n154);
not  g508 (n581, n133);
not  g509 (n312, n77);
not  g510 (n616, n149);
not  g511 (n337, n38);
not  g512 (n579, n109);
not  g513 (n191, n104);
buf  g514 (n575, n158);
buf  g515 (n471, n160);
buf  g516 (n356, n143);
buf  g517 (n470, n127);
not  g518 (n307, n93);
buf  g519 (n459, n61);
buf  g520 (n232, n137);
buf  g521 (n516, n118);
not  g522 (n236, n115);
not  g523 (n477, n127);
buf  g524 (n403, n66);
not  g525 (n244, n79);
buf  g526 (n521, n125);
not  g527 (n223, n140);
not  g528 (n429, n79);
buf  g529 (n480, n59);
not  g530 (n542, n134);
buf  g531 (n630, n44);
buf  g532 (n474, n91);
not  g533 (n336, n90);
buf  g534 (n569, n47);
buf  g535 (n486, n136);
buf  g536 (n175, n33);
not  g537 (n395, n160);
not  g538 (n435, n51);
not  g539 (n653, n82);
buf  g540 (n461, n118);
not  g541 (n443, n48);
buf  g542 (n344, n123);
not  g543 (n192, n44);
not  g544 (n349, n65);
buf  g545 (n535, n107);
buf  g546 (n372, n117);
not  g547 (n544, n92);
not  g548 (n671, n68);
not  g549 (n602, n85);
buf  g550 (n188, n136);
buf  g551 (n355, n142);
not  g552 (n502, n62);
not  g553 (n643, n81);
not  g554 (n512, n41);
not  g555 (n524, n131);
not  g556 (n493, n43);
not  g557 (n264, n49);
not  g558 (n392, n95);
not  g559 (n215, n52);
not  g560 (n301, n52);
not  g561 (n561, n88);
buf  g562 (n346, n39);
not  g563 (n570, n116);
not  g564 (n263, n73);
buf  g565 (n421, n148);
buf  g566 (n638, n105);
not  g567 (n162, n99);
not  g568 (n209, n154);
not  g569 (n406, n122);
buf  g570 (n457, n138);
not  g571 (n230, n158);
buf  g572 (n642, n35);
not  g573 (n308, n76);
not  g574 (n345, n102);
not  g575 (n399, n67);
buf  g576 (n252, n43);
buf  g577 (n394, n144);
buf  g578 (n487, n150);
buf  g579 (n319, n64);
not  g580 (n517, n46);
not  g581 (n553, n86);
not  g582 (n317, n153);
buf  g583 (n510, n148);
not  g584 (n373, n43);
buf  g585 (n665, n147);
not  g586 (n608, n82);
buf  g587 (n566, n58);
buf  g588 (n203, n142);
buf  g589 (n433, n69);
not  g590 (n272, n146);
buf  g591 (n174, n38);
not  g592 (n402, n139);
not  g593 (n200, n129);
not  g594 (n603, n99);
not  g595 (n533, n54);
buf  g596 (n181, n37);
not  g597 (n195, n48);
not  g598 (n405, n50);
buf  g599 (n185, n111);
not  g600 (n305, n152);
not  g601 (n382, n90);
buf  g602 (n179, n53);
buf  g603 (n273, n139);
buf  g604 (n333, n37);
buf  g605 (n285, n134);
buf  g606 (n266, n120);
not  g607 (n635, n155);
buf  g608 (n615, n112);
buf  g609 (n660, n103);
not  g610 (n499, n116);
buf  g611 (n420, n122);
buf  g612 (n410, n48);
not  g613 (n277, n113);
buf  g614 (n618, n55);
not  g615 (n594, n80);
not  g616 (n237, n40);
buf  g617 (n505, n63);
buf  g618 (n168, n73);
not  g619 (n563, n137);
not  g620 (n442, n142);
buf  g621 (n241, n138);
buf  g622 (n335, n130);
buf  g623 (n302, n140);
not  g624 (n656, n79);
buf  g625 (n321, n51);
not  g626 (n601, n66);
not  g627 (n265, n42);
buf  g628 (n432, n156);
buf  g629 (n607, n68);
buf  g630 (n621, n117);
buf  g631 (n489, n158);
not  g632 (n646, n112);
buf  g633 (n196, n104);
buf  g634 (n562, n99);
not  g635 (n309, n89);
not  g636 (n598, n71);
not  g637 (n490, n126);
buf  g638 (n261, n134);
not  g639 (n529, n98);
xnor g640 (n845, n430, n456, n333, n486);
nor  g641 (n685, n280, n461, n353, n357);
nand g642 (n814, n380, n332, n272, n378);
and  g643 (n851, n438, n407, n363, n423);
or   g644 (n903, n264, n484, n375, n369);
nand g645 (n726, n186, n319, n447, n303);
nand g646 (n746, n327, n233, n277, n426);
xor  g647 (n773, n167, n266, n442, n344);
xor  g648 (n843, n497, n459, n489, n417);
xor  g649 (n751, n348, n378, n398, n488);
nand g650 (n922, n367, n314, n269, n303);
xnor g651 (n800, n202, n282, n382, n266);
nand g652 (n863, n306, n344, n362, n229);
and  g653 (n693, n489, n386, n189, n480);
xor  g654 (n927, n165, n473, n287, n279);
nor  g655 (n912, n381, n322, n473, n428);
and  g656 (n749, n330, n244, n471, n478);
or   g657 (n870, n364, n381, n389, n383);
xor  g658 (n899, n409, n295, n274, n456);
or   g659 (n756, n446, n399, n313, n428);
nand g660 (n929, n387, n465, n406, n445);
and  g661 (n784, n452, n445, n314, n308);
or   g662 (n677, n348, n313, n300, n356);
xor  g663 (n824, n171, n410, n414, n369);
xnor g664 (n766, n297, n371, n434, n396);
and  g665 (n806, n230, n491, n351, n435);
and  g666 (n879, n334, n482, n312, n359);
nand g667 (n911, n255, n466, n352, n465);
or   g668 (n902, n416, n304, n450, n267);
xor  g669 (n859, n258, n311, n335, n461);
xor  g670 (n872, n385, n224, n377, n370);
or   g671 (n778, n422, n339, n408, n318);
xor  g672 (n865, n287, n260, n266, n269);
xnor g673 (n837, n445, n277, n205, n370);
or   g674 (n812, n425, n400, n417, n284);
nand g675 (n886, n274, n411, n290, n370);
and  g676 (n679, n345, n405, n421, n387);
nand g677 (n836, n309, n356, n444, n292);
nor  g678 (n890, n198, n372, n435);
and  g679 (n847, n330, n174, n380, n484);
nand g680 (n901, n423, n325, n289, n474);
xnor g681 (n690, n354, n446, n261, n176);
or   g682 (n793, n319, n338, n206, n342);
xor  g683 (n737, n490, n262, n449, n483);
xnor g684 (n834, n195, n355, n333, n484);
and  g685 (n842, n335, n460, n336, n326);
xor  g686 (n937, n398, n297, n481, n498);
xnor g687 (n909, n375, n315, n340, n390);
and  g688 (n700, n498, n307, n356, n455);
or   g689 (n704, n263, n361, n300, n420);
nand g690 (n829, n353, n259, n344, n245);
xnor g691 (n792, n390, n384, n161, n258);
and  g692 (n880, n295, n425, n163, n298);
or   g693 (n893, n367, n391, n458, n314);
xor  g694 (n817, n256, n493, n397, n360);
xnor g695 (n802, n472, n468, n414, n393);
xor  g696 (n908, n350, n178, n271, n427);
and  g697 (n830, n315, n187, n405, n376);
and  g698 (n915, n381, n359, n219, n291);
xnor g699 (n720, n434, n439, n416, n366);
nand g700 (n831, n475, n223, n409, n406);
and  g701 (n673, n379, n270, n448, n298);
xor  g702 (n796, n192, n265, n456, n293);
xor  g703 (n684, n427, n378, n443, n301);
xor  g704 (n926, n388, n373, n261, n291);
xnor g705 (n736, n331, n488, n411, n251);
and  g706 (n885, n292, n492, n455, n349);
nor  g707 (n846, n440, n336, n319, n307);
and  g708 (n923, n485, n418, n177, n326);
nand g709 (n730, n310, n388, n396, n458);
or   g710 (n891, n354, n375, n304, n267);
or   g711 (n686, n397, n469, n259, n472);
nand g712 (n921, n275, n299, n278);
or   g713 (n713, n431, n431, n443, n412);
nor  g714 (n876, n457, n166, n391, n276);
xor  g715 (n810, n489, n364, n493, n325);
or   g716 (n883, n388, n384, n261, n211);
and  g717 (n873, n359, n438, n296, n243);
xor  g718 (n848, n474, n276, n494, n280);
xor  g719 (n898, n342, n281, n370, n312);
xor  g720 (n887, n183, n465, n347, n381);
and  g721 (n930, n490, n448, n409, n469);
nand g722 (n764, n300, n345, n306, n318);
nor  g723 (n725, n466, n330, n394, n372);
nor  g724 (n884, n277, n419, n262, n497);
nor  g725 (n676, n321, n280, n413, n439);
xnor g726 (n680, n373, n424, n271, n391);
or   g727 (n900, n435, n497, n282, n321);
nor  g728 (n744, n284, n225, n464, n345);
xor  g729 (n743, n423, n216, n270, n353);
xor  g730 (n731, n291, n374, n433);
xor  g731 (n904, n308, n179, n313, n397);
nor  g732 (n894, n253, n494, n364, n487);
xnor g733 (n925, n326, n263, n324, n463);
xor  g734 (n933, n485, n320, n352, n309);
nand g735 (n809, n271, n459, n440, n443);
and  g736 (n758, n310, n287, n196, n355);
or   g737 (n936, n283, n279, n286, n449);
nand g738 (n869, n349, n386, n309, n318);
or   g739 (n807, n418, n348, n376, n337);
nor  g740 (n896, n297, n411, n435, n445);
xor  g741 (n708, n468, n252, n460, n422);
xnor g742 (n828, n356, n371, n485, n412);
and  g743 (n775, n317, n340, n305, n498);
or   g744 (n695, n403, n392, n408, n469);
xnor g745 (n740, n410, n263, n374, n349);
and  g746 (n729, n392, n376, n478, n258);
nand g747 (n808, n402, n348, n499, n281);
nand g748 (n741, n496, n301, n315, n324);
and  g749 (n748, n430, n443, n463, n254);
and  g750 (n785, n479, n295, n301, n382);
xnor g751 (n889, n184, n416, n349, n358);
and  g752 (n682, n441, n476, n492, n334);
and  g753 (n854, n282, n293, n241, n329);
nor  g754 (n783, n273, n362, n412, n299);
nor  g755 (n850, n494, n471, n221);
xor  g756 (n888, n302, n496, n374, n285);
xnor g757 (n935, n170, n427, n321, n473);
nand g758 (n739, n332, n437, n220, n260);
and  g759 (n841, n482, n457, n350, n360);
xnor g760 (n771, n315, n389, n199, n360);
nor  g761 (n916, n404, n368, n346, n292);
xnor g762 (n857, n320, n429, n188, n453);
nand g763 (n789, n289, n392, n433, n272);
nand g764 (n795, n465, n405, n375, n172);
nor  g765 (n815, n442, n391, n331, n288);
and  g766 (n849, n386, n493, n437, n477);
nand g767 (n840, n404, n401, n407, n384);
nor  g768 (n907, n397, n325, n327, n363);
or   g769 (n786, n246, n451, n311, n300);
or   g770 (n924, n294, n463, n407, n308);
xor  g771 (n747, n424, n351, n339, n438);
xor  g772 (n728, n386, n294, n353, n303);
xnor g773 (n701, n341, n477, n307, n476);
nand g774 (n691, n302, n434, n454, n476);
xor  g775 (n852, n331, n269, n413, n395);
nand g776 (n733, n310, n404, n342, n359);
xnor g777 (n860, n264, n478, n222, n447);
nor  g778 (n895, n268, n434, n487, n405);
nor  g779 (n750, n476, n290, n383, n436);
xor  g780 (n820, n265, n428, n292, n193);
xor  g781 (n727, n310, n483, n467, n323);
or   g782 (n787, n340, n257, n283, n273);
nand g783 (n913, n486, n411, n413, n340);
xnor g784 (n897, n347, n232, n432, n346);
and  g785 (n759, n417, n470, n446, n326);
xor  g786 (n735, n256, n460, n369, n164);
and  g787 (n791, n294, n361, n328, n362);
or   g788 (n801, n439, n472, n488, n461);
or   g789 (n772, n319, n485, n368, n395);
and  g790 (n892, n373, n406, n347, n366);
or   g791 (n878, n484, n431, n332, n317);
nand g792 (n774, n427, n453, n496, n328);
nand g793 (n753, n288, n328, n383, n217);
xor  g794 (n714, n346, n379, n248, n314);
nand g795 (n871, n255, n421, n268, n290);
xor  g796 (n855, n304, n238, n456, n479);
xnor g797 (n862, n384, n256, n415, n226);
nor  g798 (n813, n491, n471, n480, n369);
nor  g799 (n763, n394, n296, n444, n461);
xnor g800 (n853, n323, n210, n403, n285);
or   g801 (n767, n262, n267, n482, n338);
nand g802 (n805, n347, n422, n277, n256);
or   g803 (n719, n312, n185, n399, n306);
xor  g804 (n864, n394, n436, n459, n255);
nand g805 (n877, n316, n200, n288, n416);
nand g806 (n711, n367, n454, n285, n439);
or   g807 (n867, n260, n335, n323, n295);
and  g808 (n822, n467, n474, n379, n260);
xor  g809 (n868, n424, n237, n469, n406);
xor  g810 (n689, n488, n432, n451, n258);
xnor g811 (n705, n354, n377, n357, n432);
or   g812 (n914, n453, n190, n316, n419);
nand g813 (n882, n371, n395, n454, n472);
nand g814 (n825, n396, n440, n290, n419);
or   g815 (n939, n402, n351, n429, n274);
and  g816 (n917, n479, n312, n418, n452);
or   g817 (n938, n382, n388, n491, n430);
nor  g818 (n827, n392, n408, n478, n407);
nor  g819 (n832, n430, n380, n462, n343);
xnor g820 (n823, n257, n338, n400, n448);
nand g821 (n707, n389, n259, n417, n316);
xor  g822 (n715, n259, n242, n280, n376);
or   g823 (n782, n212, n420, n273, n352);
nand g824 (n724, n486, n483, n466, n283);
nand g825 (n717, n236, n180, n475, n234);
nor  g826 (n752, n361, n385, n366, n401);
xnor g827 (n770, n305, n299, n486, n425);
nand g828 (n797, n480, n284, n468, n350);
and  g829 (n838, n436, n325, n495, n366);
nand g830 (n745, n377, n449, n264, n477);
or   g831 (n780, n470, n304, n377, n331);
or   g832 (n702, n317, n448, n327, n399);
or   g833 (n755, n250, n308, n418, n487);
xnor g834 (n688, n313, n367, n181, n403);
nand g835 (n768, n473, n285, n275, n432);
nor  g836 (n732, n274, n169, n379, n477);
xnor g837 (n940, n311, n415, n235, n284);
and  g838 (n765, n362, n231, n303, n364);
nand g839 (n811, n335, n276, n299, n296);
nand g840 (n918, n344, n378, n341, n365);
or   g841 (n696, n329, n455, n343, n197);
xor  g842 (n716, n247, n336, n327, n447);
nor  g843 (n721, n426, n293, n492, n257);
nor  g844 (n826, n446, n428, n333, n429);
xnor g845 (n776, n275, n480, n475, n287);
nor  g846 (n881, n382, n227, n393, n279);
xor  g847 (n905, n400, n404, n263, n479);
and  g848 (n712, n426, n275, n361, n468);
and  g849 (n687, n270, n368, n398, n301);
nor  g850 (n866, n499, n393, n293, n289);
and  g851 (n803, n272, n462, n433, n239);
xnor g852 (n694, n398, n450, n481, n298);
nor  g853 (n760, n463, n306, n395, n339);
nor  g854 (n722, n341, n342, n286);
xor  g855 (n839, n288, n329, n441, n334);
xor  g856 (n761, n408, n459, n168, n401);
xnor g857 (n804, n324, n337, n368, n390);
xnor g858 (n920, n458, n266, n278, n457);
xnor g859 (n931, n447, n496, n466, n339);
nor  g860 (n906, n419, n423, n267, n318);
xor  g861 (n875, n414, n268, n352, n207);
nand g862 (n706, n302, n268, n357, n208);
or   g863 (n681, n402, n358, n265, n322);
and  g864 (n697, n271, n343, n283, n470);
and  g865 (n742, n452, n341, n444, n495);
or   g866 (n754, n457, n330, n354, n494);
or   g867 (n799, n355, n218, n422, n390);
and  g868 (n794, n426, n402, n444, n396);
nor  g869 (n819, n452, n328, n462, n357);
xnor g870 (n779, n297, n316, n450, n203);
nand g871 (n777, n191, n436, n294, n334);
and  g872 (n856, n333, n194, n403, n400);
xor  g873 (n757, n464, n482, n454, n249);
xor  g874 (n932, n305, n175, n324, n264);
nand g875 (n692, n449, n393, n498, n346);
xnor g876 (n861, n255, n410, n329, n495);
nor  g877 (n790, n336, n286, n414, n385);
or   g878 (n844, n358, n343, n491, n365);
xnor g879 (n821, n209, n279, n272, n438);
xnor g880 (n816, n481, n173, n490, n451);
or   g881 (n683, n464, n240, n273, n421);
or   g882 (n723, n317, n338, n497, n363);
or   g883 (n674, n453, n321, n311, n410);
nor  g884 (n734, n412, n276, n455, n467);
xnor g885 (n675, n495, n320, n214, n383);
and  g886 (n781, n490, n257, n302, n380);
xnor g887 (n703, n322, n365, n358, n269);
or   g888 (n718, n363, n481, n487, n442);
and  g889 (n798, n355, n182, n421, n270);
nor  g890 (n919, n483, n278, n281);
nor  g891 (n738, n429, n332, n467, n442);
nand g892 (n858, n373, n470, n282, n372);
and  g893 (n678, n415, n433, n460, n387);
nand g894 (n910, n493, n450, n320, n474);
xor  g895 (n769, n437, n424, n296, n289);
or   g896 (n818, n401, n213, n204, n420);
xnor g897 (n833, n489, n298, n441, n265);
xor  g898 (n788, n309, n399, n389, n323);
nand g899 (n709, n337, n440, n322, n351);
xor  g900 (n699, n492, n431, n387, n360);
xnor g901 (n762, n437, n420, n415, n215);
nand g902 (n710, n291, n307, n441, n458);
nor  g903 (n928, n451, n385, n337, n425);
or   g904 (n934, n464, n262, n462, n394);
xnor g905 (n698, n345, n371, n365, n261);
nand g906 (n874, n201, n409, n350, n228);
nand g907 (n835, n162, n475, n413, n305);
or   g908 (n1148, n640, n605, n569, n887);
nand g909 (n982, n638, n536, n515, n636);
xnor g910 (n1041, n592, n631, n500, n572);
xnor g911 (n1070, n704, n749, n620, n518);
nand g912 (n1149, n560, n529, n615, n587);
or   g913 (n1046, n502, n574, n659, n549);
xnor g914 (n1098, n630, n514, n622, n886);
and  g915 (n1133, n512, n641, n647, n607);
xor  g916 (n1107, n601, n659, n756, n658);
nand g917 (n1109, n534, n666, n632, n686);
or   g918 (n1152, n864, n551, n611, n733);
nor  g919 (n1075, n718, n654, n594, n633);
or   g920 (n963, n646, n503, n530, n578);
nand g921 (n1092, n593, n521, n586, n509);
xor  g922 (n1037, n577, n649, n595, n548);
and  g923 (n956, n600, n598, n627, n893);
nor  g924 (n1047, n667, n602, n800, n590);
or   g925 (n1159, n505, n649, n598, n645);
xor  g926 (n1134, n820, n668, n859, n727);
xnor g927 (n988, n506, n755, n678, n510);
xnor g928 (n977, n602, n603, n528, n648);
nand g929 (n1061, n639, n525, n837, n599);
and  g930 (n1150, n597, n843, n762, n620);
xnor g931 (n979, n879, n809, n556, n836);
xor  g932 (n1043, n806, n657, n882, n808);
xor  g933 (n1019, n878, n650, n831, n517);
and  g934 (n1027, n612, n518, n770, n594);
nand g935 (n1062, n615, n612, n601, n510);
xor  g936 (n1066, n509, n612, n703, n782);
nand g937 (n1079, n559, n580, n603, n554);
nor  g938 (n1108, n614, n547, n648, n661);
and  g939 (n1071, n559, n504, n766, n853);
and  g940 (n966, n538, n534, n740, n846);
xnor g941 (n1165, n544, n535, n790, n632);
and  g942 (n1063, n589, n659, n550, n665);
and  g943 (n1073, n535, n513, n574, n503);
xor  g944 (n1031, n714, n529, n516, n628);
xnor g945 (n1124, n657, n757, n812, n538);
xor  g946 (n1033, n538, n675, n735, n665);
xor  g947 (n952, n532, n590, n639, n585);
or   g948 (n1096, n610, n619, n581, n695);
xnor g949 (n1029, n642, n616, n537, n676);
nor  g950 (n980, n515, n765, n510, n728);
xnor g951 (n1086, n842, n521, n643, n701);
nor  g952 (n1099, n573, n604, n779, n521);
nor  g953 (n954, n577, n869, n618, n657);
nor  g954 (n984, n506, n594, n571, n513);
nand g955 (n1163, n553, n629, n562, n517);
nor  g956 (n969, n531, n691, n710, n620);
xor  g957 (n983, n635, n738, n645, n816);
or   g958 (n1128, n606, n900, n777, n797);
xor  g959 (n1007, n641, n507, n570, n523);
nor  g960 (n1009, n559, n776, n530, n641);
xor  g961 (n1156, n586, n668, n561, n522);
nor  g962 (n1054, n511, n606, n567, n637);
nor  g963 (n949, n538, n519, n540, n520);
and  g964 (n987, n665, n616, n888, n516);
nor  g965 (n1008, n519, n600, n612, n635);
xor  g966 (n955, n528, n590, n608, n663);
xor  g967 (n944, n659, n614, n767, n543);
xnor g968 (n1132, n744, n505, n646, n563);
xor  g969 (n1021, n663, n535, n504, n698);
xor  g970 (n989, n817, n634, n522, n615);
or   g971 (n981, n523, n562, n617, n582);
xor  g972 (n1042, n536, n699, n575, n500);
xor  g973 (n1144, n527, n608, n603, n563);
xnor g974 (n1069, n533, n655, n540, n568);
and  g975 (n959, n717, n605, n543, n683);
nor  g976 (n960, n720, n566, n531, n557);
nor  g977 (n994, n619, n752, n662, n898);
or   g978 (n1064, n589, n645, n581, n793);
xor  g979 (n1111, n653, n540, n833, n579);
or   g980 (n1091, n753, n617, n630, n524);
or   g981 (n1089, n880, n636, n628, n525);
or   g982 (n1038, n841, n845, n550);
xnor g983 (n1093, n537, n871, n571, n541);
xor  g984 (n1074, n618, n613, n614, n642);
nand g985 (n992, n828, n608, n537, n680);
and  g986 (n999, n515, n629, n599, n607);
xor  g987 (n942, n874, n811, n835, n677);
xnor g988 (n1115, n660, n656, n629, n534);
xor  g989 (n1100, n741, n666, n590, n622);
xor  g990 (n1157, n876, n570, n526, n865);
nand g991 (n1114, n583, n600, n601, n517);
or   g992 (n1013, n575, n604, n527, n715);
xor  g993 (n1000, n644, n507, n891, n557);
or   g994 (n1143, n568, n557, n664, n592);
and  g995 (n1095, n546, n613, n625, n595);
or   g996 (n1056, n520, n839, n791, n635);
or   g997 (n1105, n587, n524, n774, n775);
and  g998 (n976, n636, n652, n544, n586);
xor  g999 (n967, n539, n564, n730, n649);
nor  g1000 (n993, n586, n826, n642, n796);
and  g1001 (n1022, n854, n892, n631, n834);
nor  g1002 (n1080, n705, n618, n515, n801);
nand g1003 (n1025, n795, n579, n502, n522);
and  g1004 (n1094, n576, n589, n688, n747);
or   g1005 (n1118, n610, n638, n783, n643);
nand g1006 (n1024, n664, n549, n622, n588);
and  g1007 (n1001, n585, n499, n535, n639);
nor  g1008 (n1034, n870, n823, n521, n504);
or   g1009 (n1136, n550, n792, n598, n542);
xnor g1010 (n1116, n514, n637, n570, n739);
xor  g1011 (n1015, n519, n868, n615, n732);
nor  g1012 (n968, n555, n580, n664, n563);
nor  g1013 (n1050, n802, n501, n573, n863);
xnor g1014 (n1102, n611, n650, n531, n520);
xor  g1015 (n1123, n789, n697, n799, n584);
nor  g1016 (n1032, n662, n507, n501, n585);
xor  g1017 (n1028, n760, n544, n606, n661);
xor  g1018 (n1011, n584, n572, n518, n685);
xnor g1019 (n1018, n651, n707, n643, n655);
nand g1020 (n943, n528, n626, n623, n593);
or   g1021 (n1067, n696, n548, n651, n572);
nand g1022 (n1090, n556, n572, n566, n724);
and  g1023 (n974, n588, n647, n627, n591);
nor  g1024 (n1110, n508, n621, n526, n569);
or   g1025 (n1164, n523, n541, n609, n575);
xor  g1026 (n1087, n564, n646, n595, n848);
xor  g1027 (n1048, n667, n524, n608, n540);
and  g1028 (n1068, n784, n539, n578, n547);
xor  g1029 (n1057, n661, n617, n885, n507);
nand g1030 (n1077, n838, n743, n596, n543);
nor  g1031 (n1162, n682, n872, n599, n713);
xnor g1032 (n1076, n668, n509, n712, n532);
nand g1033 (n946, n579, n822, n561, n616);
xnor g1034 (n1160, n541, n821, n644, n624);
or   g1035 (n1101, n585, n751, n645, n623);
nand g1036 (n1053, n679, n617, n810, n737);
nand g1037 (n1142, n505, n895, n654, n638);
or   g1038 (n1131, n622, n580, n805, n537);
xor  g1039 (n985, n716, n827, n505, n551);
xor  g1040 (n1045, n544, n693, n546, n794);
or   g1041 (n948, n897, n589, n706, n815);
or   g1042 (n1005, n651, n639, n851, n502);
nor  g1043 (n971, n662, n655, n736, n648);
nor  g1044 (n986, n819, n640, n778, n502);
nand g1045 (n1039, n609, n554, n829, n624);
nand g1046 (n945, n654, n581, n588);
xnor g1047 (n947, n553, n519, n689, n652);
nand g1048 (n1121, n850, n875, n771, n619);
xor  g1049 (n1104, n630, n648, n511, n745);
and  g1050 (n1112, n576, n605, n656, n582);
nand g1051 (n1141, n577, n866, n553, n616);
or   g1052 (n1036, n621, n532, n511, n559);
xor  g1053 (n1072, n504, n514, n556, n552);
xnor g1054 (n1129, n877, n803, n595, n596);
xor  g1055 (n1153, n726, n646, n644, n541);
and  g1056 (n1154, n587, n536, n861, n746);
nor  g1057 (n951, n692, n596, n593, n506);
or   g1058 (n1017, n621, n856, n534, n840);
and  g1059 (n1044, n578, n609, n619, n527);
or   g1060 (n1055, n632, n641, n721, n552);
and  g1061 (n1020, n501, n547, n530, n602);
or   g1062 (n1125, n652, n526, n832, n633);
nor  g1063 (n1051, n661, n763, n729, n665);
xor  g1064 (n1016, n625, n798, n613, n830);
or   g1065 (n1059, n565, n533, n660, n722);
nand g1066 (n1126, n786, n583, n633, n587);
nor  g1067 (n1113, n542, n614, n658, n620);
nand g1068 (n995, n666, n857, n607, n564);
nor  g1069 (n1030, n600, n700, n862, n621);
xor  g1070 (n997, n558, n643, n690, n660);
xor  g1071 (n970, n593, n569, n561, n528);
nor  g1072 (n1085, n825, n525, n899, n663);
xnor g1073 (n961, n579, n558, n543);
nor  g1074 (n1127, n889, n884, n626, n630);
nand g1075 (n973, n582, n855, n568, n633);
xor  g1076 (n975, n570, n653, n545, n580);
nand g1077 (n1010, n552, n613, n631, n635);
nor  g1078 (n1146, n516, n571, n634, n847);
and  g1079 (n1103, n546, n560, n500, n708);
and  g1080 (n957, n522, n627, n601, n781);
xnor g1081 (n1012, n571, n629, n567, n563);
nand g1082 (n1122, n592, n561, n558, n565);
xor  g1083 (n991, n583, n551, n636, n759);
xor  g1084 (n1014, n574, n573, n638, n582);
xor  g1085 (n1151, n557, n512, n666, n576);
and  g1086 (n1097, n512, n533, n529, n642);
xor  g1087 (n1155, n725, n625, n592, n742);
and  g1088 (n1052, n653, n539, n511, n702);
nor  g1089 (n962, n577, n548, n723, n536);
nor  g1090 (n1166, n644, n560, n552, n525);
and  g1091 (n998, n598, n576, n768, n656);
nor  g1092 (n1023, n566, n565, n769, n508);
and  g1093 (n1065, n611, n547, n849, n605);
nor  g1094 (n958, n750, n780, n660, n664);
xnor g1095 (n1049, n551, n883, n628, n556);
xor  g1096 (n996, n637, n567, n658, n545);
xor  g1097 (n1083, n518, n647, n533, n549);
and  g1098 (n1006, n787, n567, n609, n542);
nor  g1099 (n1002, n632, n640, n748, n503);
nand g1100 (n1140, n555, n553, n554, n734);
or   g1101 (n1040, n896, n509, n584, n627);
nand g1102 (n990, n532, n510, n555, n512);
and  g1103 (n1139, n529, n565, n623, n596);
or   g1104 (n978, n545, n813, n890, n574);
xnor g1105 (n1078, n618, n731, n514, n761);
nand g1106 (n1119, n562, n852, n591, n773);
and  g1107 (n1145, n545, n807, n814, n662);
nor  g1108 (n1060, n555, n597, n566, n611);
xor  g1109 (n1120, n684, n594, n573, n531);
xor  g1110 (n953, n569, n772, n513, n719);
or   g1111 (n1082, n578, n597, n560, n658);
and  g1112 (n1003, n568, n562, n881, n709);
or   g1113 (n1161, n610, n575, n524, n694);
xnor g1114 (n1035, n526, n506, n508, n818);
nor  g1115 (n941, n804, n867, n824, n523);
and  g1116 (n1084, n501, n656, n764, n650);
and  g1117 (n964, n623, n626, n583);
and  g1118 (n1137, n548, n651, n508, n527);
or   g1119 (n1088, n711, n844, n637, n647);
xnor g1120 (n972, n591, n624, n681, n606);
xor  g1121 (n1130, n530, n663, n894, n599);
xor  g1122 (n1106, n858, n517, n754, n652);
xor  g1123 (n1117, n542, n650, n624, n667);
and  g1124 (n965, n657, n785, n520, n499);
and  g1125 (n1058, n539, n607, n549, n602);
nand g1126 (n1135, n634, n653, n655, n604);
nand g1127 (n1004, n581, n654, n610, n513);
and  g1128 (n1138, n667, n788, n500, n860);
nand g1129 (n1147, n516, n649, n640, n564);
xnor g1130 (n950, n634, n628, n604, n584);
or   g1131 (n1026, n687, n591, n668, n631);
nor  g1132 (n1081, n546, n873, n758, n503);
nand g1133 (n1158, n603, n625, n554, n597);
or   g1134 (n1194, n933, n1004, n960, n916);
xor  g1135 (n1168, n1015, n1049, n943, n1013);
xor  g1136 (n1171, n911, n932, n1063, n1068);
xor  g1137 (n1176, n907, n915, n1054, n957);
or   g1138 (n1172, n1023, n924, n920, n972);
xnor g1139 (n1202, n927, n1017, n1011, n1066);
nand g1140 (n1197, n1067, n903, n925, n975);
nor  g1141 (n1186, n948, n968, n1032, n1069);
and  g1142 (n1183, n1018, n1074, n909, n1061);
nor  g1143 (n1196, n934, n964, n990, n996);
nand g1144 (n1169, n1012, n984, n917, n1019);
nor  g1145 (n1195, n1031, n985, n904, n978);
nand g1146 (n1207, n1036, n1059, n918, n1041);
and  g1147 (n1187, n1008, n1046, n914, n1070);
xor  g1148 (n1184, n999, n1025, n912, n988);
nor  g1149 (n1191, n1053, n1035, n1052, n942);
nor  g1150 (n1204, n958, n1022, n928, n902);
or   g1151 (n1201, n1006, n908, n950, n997);
or   g1152 (n1181, n1062, n959, n966, n973);
or   g1153 (n1173, n1065, n923, n989, n1047);
or   g1154 (n1175, n986, n1021, n952, n969);
xor  g1155 (n1208, n1034, n1030, n1027, n955);
nand g1156 (n1189, n1003, n1029, n998, n1073);
and  g1157 (n1200, n944, n971, n1064, n1039);
xor  g1158 (n1180, n1048, n931, n947, n921);
or   g1159 (n1177, n981, n995, n1009, n976);
or   g1160 (n1182, n929, n919, n974, n953);
xnor g1161 (n1206, n930, n956, n946, n1055);
xnor g1162 (n1185, n901, n1057, n991, n1010);
or   g1163 (n1179, n1038, n1040, n951, n1028);
and  g1164 (n1167, n1005, n906, n1037, n1002);
xor  g1165 (n1190, n967, n970, n1051, n1020);
and  g1166 (n1192, n1000, n1043, n1058, n941);
or   g1167 (n1178, n1042, n1044, n949, n926);
xnor g1168 (n1193, n910, n1026, n980, n1016);
and  g1169 (n1203, n1007, n983, n945, n994);
nor  g1170 (n1174, n987, n913, n905, n922);
nand g1171 (n1188, n993, n1056, n1024, n1050);
xor  g1172 (n1170, n982, n992, n1071, n1014);
or   g1173 (n1198, n954, n979, n1001, n977);
or   g1174 (n1199, n1033, n1060, n961, n962);
xor  g1175 (n1205, n1072, n965, n1045, n963);
nand g1176 (n1222, n1079, n1145, n1195);
nand g1177 (n1214, n1098, n1119, n1189);
nor  g1178 (n1211, n1107, n1133, n1150, n1132);
xor  g1179 (n1212, n1105, n1193, n1115, n1096);
nor  g1180 (n1220, n1087, n1192, n1139, n1086);
nor  g1181 (n1226, n1116, n1190, n1184, n1185);
xnor g1182 (n1218, n1117, n1147, n1148, n1089);
and  g1183 (n1227, n1095, n1099, n1138, n1202);
xor  g1184 (n1217, n1142, n1084, n1194, n1088);
xnor g1185 (n1234, n1091, n1094, n1082, n1125);
xnor g1186 (n1230, n1141, n1118, n1093, n1108);
xor  g1187 (n1213, n1104, n1123, n1114, n1078);
xnor g1188 (n1219, n1129, n1201, n1090, n1134);
xor  g1189 (n1210, n1181, n1077, n1198, n1200);
or   g1190 (n1223, n1186, n1113, n1203, n1110);
nand g1191 (n1216, n1146, n1140, n1076, n1191);
nor  g1192 (n1232, n1135, n1130, n1122, n1187);
nor  g1193 (n1225, n1182, n1083, n1131, n1106);
and  g1194 (n1209, n1097, n1124, n1197, n1128);
nor  g1195 (n1228, n1112, n1188, n1137, n1111);
xnor g1196 (n1231, n1136, n1075, n1101, n1103);
and  g1197 (n1215, n1179, n1143, n1127, n1183);
and  g1198 (n1224, n1092, n1085, n1126, n1081);
xor  g1199 (n1221, n1180, n1120, n1199, n1121);
xor  g1200 (n1233, n1204, n1196, n1109, n1080);
nand g1201 (n1229, n1102, n1149, n1144, n1100);
not  g1202 (n1258, n1154);
not  g1203 (n1256, n1233);
buf  g1204 (n1240, n1225);
buf  g1205 (n1238, n1151);
not  g1206 (n1248, n1222);
not  g1207 (n1247, n1152);
not  g1208 (n1235, n1219);
not  g1209 (n1242, n1223);
buf  g1210 (n1237, n1210);
not  g1211 (n1236, n1215);
not  g1212 (n1252, n1226);
buf  g1213 (n1253, n1221);
buf  g1214 (n1260, n1212);
not  g1215 (n1239, n1214);
buf  g1216 (n1250, n1153);
buf  g1217 (n1254, n1216);
not  g1218 (n1241, n1227);
not  g1219 (n1246, n1234);
not  g1220 (n1245, n1211);
buf  g1221 (n1251, n1232);
not  g1222 (n1244, n1220);
not  g1223 (n1255, n1218);
nand g1224 (n1257, n1224, n1230);
and  g1225 (n1249, n1228, n1234);
and  g1226 (n1243, n1229, n1217);
nor  g1227 (n1259, n1209, n1155);
xnor g1228 (n1261, n1231, n1213);
not  g1229 (n1302, n1243);
not  g1230 (n1312, n1235);
not  g1231 (n1325, n1249);
buf  g1232 (n1262, n1250);
not  g1233 (n1275, n1242);
buf  g1234 (n1267, n1240);
not  g1235 (n1335, n1248);
not  g1236 (n1276, n1248);
not  g1237 (n1310, n1253);
not  g1238 (n1296, n1251);
not  g1239 (n1271, n1238);
not  g1240 (n1332, n1254);
not  g1241 (n1265, n1247);
buf  g1242 (n1334, n1240);
not  g1243 (n1329, n1254);
not  g1244 (n1294, n1248);
buf  g1245 (n1311, n1236);
buf  g1246 (n1322, n1242);
not  g1247 (n1326, n1235);
buf  g1248 (n1331, n1247);
not  g1249 (n1338, n1242);
buf  g1250 (n1297, n1252);
buf  g1251 (n1288, n1241);
buf  g1252 (n1336, n1237);
not  g1253 (n1289, n1239);
buf  g1254 (n1304, n1241);
not  g1255 (n1290, n1237);
not  g1256 (n1284, n1246);
not  g1257 (n1274, n1247);
buf  g1258 (n1317, n1243);
not  g1259 (n1330, n1241);
buf  g1260 (n1269, n1237);
buf  g1261 (n1318, n1237);
buf  g1262 (n1295, n1244);
not  g1263 (n1301, n1254);
not  g1264 (n1314, n1235);
not  g1265 (n1263, n1253);
not  g1266 (n1278, n1249);
not  g1267 (n1327, n1249);
buf  g1268 (n1292, n1243);
buf  g1269 (n1266, n1253);
not  g1270 (n1293, n1240);
not  g1271 (n1291, n1246);
not  g1272 (n1287, n1251);
buf  g1273 (n1303, n1236);
not  g1274 (n1300, n1252);
buf  g1275 (n1321, n1238);
buf  g1276 (n1299, n1246);
not  g1277 (n1283, n1244);
buf  g1278 (n1273, n1238);
buf  g1279 (n1340, n1249);
not  g1280 (n1333, n1241);
not  g1281 (n1268, n1250);
buf  g1282 (n1324, n1246);
buf  g1283 (n1308, n1254);
buf  g1284 (n1341, n1238);
buf  g1285 (n1313, n1239);
not  g1286 (n1315, n1245);
buf  g1287 (n1272, n1244);
buf  g1288 (n1279, n1240);
buf  g1289 (n1282, n1250);
buf  g1290 (n1264, n1253);
not  g1291 (n1316, n1242);
buf  g1292 (n1277, n1235);
not  g1293 (n1319, n1239);
not  g1294 (n1320, n1251);
not  g1295 (n1281, n1252);
buf  g1296 (n1339, n1239);
not  g1297 (n1309, n1251);
not  g1298 (n1328, n1245);
buf  g1299 (n1270, n1245);
not  g1300 (n1337, n1250);
buf  g1301 (n1280, n1248);
buf  g1302 (n1306, n1245);
not  g1303 (n1286, n1236);
not  g1304 (n1307, n1247);
buf  g1305 (n1305, n1244);
buf  g1306 (n1323, n1236);
not  g1307 (n1298, n1243);
not  g1308 (n1285, n1252);
xnor g1309 (n1353, n1255, n1261, n1288, n1272);
nand g1310 (n1376, n1284, n1273, n1298, n1264);
xnor g1311 (n1346, n1293, n1269, n1291, n1264);
nor  g1312 (n1364, n1290, n1276, n1299, n1257);
and  g1313 (n1350, n1288, n1272, n1259, n1290);
nand g1314 (n1382, n1292, n1263, n1287, n1268);
and  g1315 (n1361, n1284, n1301, n1265, n1283);
xnor g1316 (n1374, n1267, n1275, n1281, n1263);
xnor g1317 (n1383, n1262, n1270);
xnor g1318 (n1375, n1285, n1272, n1260, n1281);
or   g1319 (n1363, n1274, n1269, n1278, n1277);
and  g1320 (n1343, n1278, n1287, n1304, n1282);
xor  g1321 (n1344, n1281, n1290, n1292, n1274);
nand g1322 (n1351, n1279, n1260, n1289, n1286);
nand g1323 (n1372, n1264, n1294, n1265, n1295);
and  g1324 (n1370, n1276, n1275, n1289, n1260);
xor  g1325 (n1391, n1301, n1294, n1258, n1302);
or   g1326 (n1387, n1268, n1267, n1258, n1295);
or   g1327 (n1362, n1298, n1271, n1264, n1289);
or   g1328 (n1356, n1282, n1277, n1255, n1298);
nand g1329 (n1388, n1301, n1277, n1260, n1287);
xor  g1330 (n1373, n1289, n1257, n1297, n1274);
nor  g1331 (n1366, n1294, n1273, n1259, n1300);
nor  g1332 (n1354, n1293, n1276, n1302, n1280);
xnor g1333 (n1378, n1266, n1271, n1270);
nor  g1334 (n1347, n1303, n1295, n1262, n1256);
nand g1335 (n1385, n1285, n1276, n1274, n1265);
and  g1336 (n1359, n1303, n1266, n1283, n1286);
nand g1337 (n1380, n1297, n1300, n1257);
nor  g1338 (n1355, n1297, n1255, n1270, n1263);
xor  g1339 (n1371, n1293, n1303, n1298, n1256);
nand g1340 (n1367, n1275, n1257, n1285, n1286);
and  g1341 (n1384, n1256, n1266, n1285, n1296);
nand g1342 (n1357, n1299, n1303, n1258, n1291);
and  g1343 (n1358, n1268, n1259, n1301, n1299);
and  g1344 (n1368, n1255, n1280, n1279, n1261);
or   g1345 (n1348, n1279, n1291, n1283, n1272);
and  g1346 (n1379, n1282, n1290, n1267, n1291);
nand g1347 (n1381, n1273, n1271, n1302, n1284);
and  g1348 (n1345, n1278, n1299, n1261, n1296);
xor  g1349 (n1365, n1269, n1265, n1278, n1296);
or   g1350 (n1352, n1280, n1268, n1273, n1284);
xor  g1351 (n1386, n1288, n1287, n1304, n1261);
or   g1352 (n1349, n1293, n1294, n1256, n1277);
or   g1353 (n1369, n1258, n1269, n1292, n1295);
and  g1354 (n1342, n1304, n1292, n1266, n1283);
nor  g1355 (n1389, n1296, n1275, n1286, n1262);
nand g1356 (n1360, n1259, n1288, n1263, n1297);
nand g1357 (n1377, n1302, n1281, n1282, n1300);
xor  g1358 (n1390, n1304, n1267, n1279, n1280);
buf  g1359 (n1398, n1306);
buf  g1360 (n1412, n1311);
not  g1361 (n1414, n1305);
not  g1362 (n1419, n1308);
buf  g1363 (n1410, n1347);
not  g1364 (n1400, n1313);
buf  g1365 (n1406, n1312);
not  g1366 (n1417, n1365);
not  g1367 (n1422, n1358);
not  g1368 (n1404, n1343);
buf  g1369 (n1408, n1369);
not  g1370 (n1403, n1315);
buf  g1371 (n1423, n1313);
not  g1372 (n1415, n1367);
not  g1373 (n1394, n1346);
buf  g1374 (n1407, n1307);
buf  g1375 (n1418, n1315);
not  g1376 (n1401, n1313);
not  g1377 (n1420, n1310);
buf  g1378 (n1413, n1316);
xnor g1379 (n1393, n1352, n1307, n1362, n1305);
xor  g1380 (n1425, n1309, n1363, n1311, n1306);
nand g1381 (n1421, n1309, n1351, n1370, n1345);
nand g1382 (n1409, n1356, n1364, n1312, n1355);
xnor g1383 (n1405, n1308, n1305, n1376);
or   g1384 (n1411, n1361, n1312, n1315, n1307);
nor  g1385 (n1426, n1307, n1310, n1374, n1371);
xor  g1386 (n1399, n1350, n1308, n1306, n1314);
and  g1387 (n1416, n1344, n1309, n1357, n1375);
nand g1388 (n1397, n1349, n1308, n1314, n1372);
xnor g1389 (n1392, n1312, n1310, n1309);
xnor g1390 (n1424, n1315, n1314, n1313);
nor  g1391 (n1395, n1353, n1359, n1311, n1342);
xor  g1392 (n1396, n1373, n1311, n1354, n1348);
xor  g1393 (n1402, n1368, n1306, n1366, n1360);
not  g1394 (n1434, n1394);
not  g1395 (n1429, n1393);
not  g1396 (n1431, n1317);
buf  g1397 (n1427, n1397);
buf  g1398 (n1433, n1397);
buf  g1399 (n1436, n1398);
buf  g1400 (n1428, n1396);
buf  g1401 (n1437, n1316);
buf  g1402 (n1432, n1397);
xnor g1403 (n1430, n1398, n1317);
nand g1404 (n1435, n1395, n1398, n1316);
xnor g1405 (n1438, n1436, n1328, n1326, n1320);
or   g1406 (n1479, n1379, n1389, n1321, n1399);
nor  g1407 (n1461, n1435, n1427, n1329, n1431);
and  g1408 (n1452, n1436, n1378, n1389, n1433);
and  g1409 (n1476, n1381, n1431, n1325, n1388);
xnor g1410 (n1456, n1318, n1434, n1382, n1329);
nor  g1411 (n1450, n1401, n1332, n1382, n1387);
nand g1412 (n1444, n1390, n1386, n1431, n1327);
nor  g1413 (n1465, n1317, n1326, n1385, n1321);
nand g1414 (n1448, n1433, n1398, n1377, n1383);
and  g1415 (n1453, n1434, n1430, n1323, n1386);
and  g1416 (n1470, n1384, n1388, n1387, n1381);
or   g1417 (n1441, n1324, n1319, n1318, n1331);
and  g1418 (n1463, n1437, n1427, n1428, n1323);
or   g1419 (n1462, n1327, n1379, n1329, n1428);
xor  g1420 (n1478, n1432, n1391, n1325, n1427);
or   g1421 (n1471, n1320, n1428, n1387, n1324);
or   g1422 (n1455, n1391, n1400, n1434, n1331);
xor  g1423 (n1445, n1379, n1437, n1385, n1319);
nand g1424 (n1472, n1432, n1384, n1399, n1386);
nand g1425 (n1443, n1320, n1330, n1325, n1326);
xnor g1426 (n1440, n1328, n1434, n1321, n1317);
nor  g1427 (n1439, n1388, n1429, n1330);
nand g1428 (n1457, n1331, n1326, n1432, n1319);
nor  g1429 (n1449, n1430, n1383, n1323, n1321);
xnor g1430 (n1477, n1377, n1320, n1386, n1322);
xnor g1431 (n1469, n1400, n1389, n1430, n1380);
nand g1432 (n1468, n1390, n1437, n1436, n1378);
nor  g1433 (n1480, n1322, n1385, n1376, n1433);
nor  g1434 (n1474, n1330, n1322, n1325, n1327);
xnor g1435 (n1473, n1427, n1377, n1379, n1385);
and  g1436 (n1466, n1383, n1388, n1400, n1435);
or   g1437 (n1460, n1430, n1328, n1378);
xor  g1438 (n1442, n1428, n1431, n1389, n1429);
or   g1439 (n1451, n1436, n1384, n1327, n1399);
nor  g1440 (n1475, n1380, n1381, n1376);
xor  g1441 (n1454, n1323, n1390, n1380, n1382);
nor  g1442 (n1467, n1319, n1429, n1435, n1376);
or   g1443 (n1459, n1384, n1437, n1383, n1324);
nand g1444 (n1446, n1400, n1390, n1318, n1387);
or   g1445 (n1481, n1391, n1433, n1382, n1328);
or   g1446 (n1464, n1380, n1399, n1377, n1432);
xnor g1447 (n1447, n1329, n1429, n1391, n1318);
nor  g1448 (n1458, n1331, n1435, n1324, n1322);
not  g1449 (n1486, n1452);
not  g1450 (n1491, n1448);
buf  g1451 (n1484, n1450);
not  g1452 (n1485, n1439);
not  g1453 (n1496, n1449);
buf  g1454 (n1488, n1440);
buf  g1455 (n1492, n1438);
not  g1456 (n1483, n1446);
not  g1457 (n1482, n1444);
buf  g1458 (n1495, n1443);
buf  g1459 (n1490, n1442);
buf  g1460 (n1494, n1441);
not  g1461 (n1493, n1453);
not  g1462 (n1489, n1447);
not  g1463 (n1487, n1451);
not  g1464 (n1497, n1445);
or   g1465 (n1502, n1415, n1455, n1411, n1488);
nand g1466 (n1511, n1401, n1416, n1403, n1404);
xnor g1467 (n1528, n1490, n1404, n1418);
nor  g1468 (n1526, n1335, n1409, n1333, n1417);
xor  g1469 (n1514, n1413, n1489, n1409, n1421);
nor  g1470 (n1503, n1411, n1335, n1416, n1401);
xnor g1471 (n1504, n1410, n1408, n1418, n1484);
and  g1472 (n1523, n1418, n1334, n1485, n1409);
and  g1473 (n1529, n1413, n1411, n1409, n1484);
or   g1474 (n1507, n1421, n1406, n1412, n1414);
xnor g1475 (n1516, n1485, n1402, n1334, n1457);
nand g1476 (n1499, n1414, n1410, n1419, n1408);
and  g1477 (n1531, n1401, n1336, n1402, n1405);
nand g1478 (n1518, n1406, n1415, n1410, n1420);
and  g1479 (n1519, n1484, n1417, n1415, n1413);
nand g1480 (n1525, n1454, n1485, n1417, n1414);
xnor g1481 (n1532, n1417, n1404, n1403, n1407);
and  g1482 (n1501, n1407, n1490, n1333, n1484);
nor  g1483 (n1505, n1482, n1405, n1488, n1489);
xor  g1484 (n1521, n1487, n1482, n1411, n1332);
or   g1485 (n1522, n1487, n1482, n1334, n1485);
xor  g1486 (n1500, n1488, n1403, n1486, n1332);
xnor g1487 (n1513, n1489, n1419, n1416, n1487);
and  g1488 (n1509, n1483, n1420);
or   g1489 (n1510, n1334, n1482, n1406, n1413);
or   g1490 (n1506, n1490, n1408, n1488, n1483);
xor  g1491 (n1530, n1419, n1412, n1422, n1487);
and  g1492 (n1508, n1405, n1422, n1333);
xor  g1493 (n1512, n1414, n1406, n1486, n1420);
nand g1494 (n1524, n1419, n1489, n1335, n1402);
and  g1495 (n1520, n1486, n1405, n1402, n1416);
xnor g1496 (n1517, n1412, n1412, n1407, n1403);
xnor g1497 (n1515, n1421, n1418, n1332, n1486);
or   g1498 (n1498, n1483, n1407, n1410, n1421);
nand g1499 (n1527, n1408, n1456, n1335, n1415);
buf  g1500 (n1543, n1513);
not  g1501 (n1549, n1516);
buf  g1502 (n1546, n1504);
buf  g1503 (n1534, n1521);
not  g1504 (n1541, n1505);
buf  g1505 (n1545, n1515);
not  g1506 (n1560, n1509);
buf  g1507 (n1544, n1510);
not  g1508 (n1552, n1524);
not  g1509 (n1559, n1498);
not  g1510 (n1538, n1525);
not  g1511 (n1556, n1517);
not  g1512 (n1548, n1523);
not  g1513 (n1539, n1512);
not  g1514 (n1535, n1506);
not  g1515 (n1542, n1520);
buf  g1516 (n1540, n1522);
not  g1517 (n1557, n1503);
not  g1518 (n1537, n1499);
buf  g1519 (n1554, n1508);
not  g1520 (n1536, n1518);
buf  g1521 (n1547, n1514);
not  g1522 (n1553, n1511);
not  g1523 (n1551, n1507);
not  g1524 (n1533, n1519);
not  g1525 (n1558, n1500);
not  g1526 (n1550, n1502);
not  g1527 (n1555, n1501);
not  g1528 (n1587, n1534);
buf  g1529 (n1593, n1471);
buf  g1530 (n1632, n1475);
not  g1531 (n1597, n1543);
not  g1532 (n1608, n1492);
buf  g1533 (n1581, n1538);
not  g1534 (n1616, n1337);
not  g1535 (n1621, n1467);
not  g1536 (n1627, n1547);
not  g1537 (n1561, n1550);
buf  g1538 (n1572, n1546);
buf  g1539 (n1623, n1472);
not  g1540 (n1574, n1461);
buf  g1541 (n1595, n1475);
not  g1542 (n1626, n1538);
buf  g1543 (n1609, n1471);
buf  g1544 (n1594, n1474);
buf  g1545 (n1604, n1546);
not  g1546 (n1585, n1491);
buf  g1547 (n1619, n1495);
not  g1548 (n1598, n1544);
buf  g1549 (n1592, n1475);
buf  g1550 (n1566, n1468);
not  g1551 (n1596, n1462);
buf  g1552 (n1602, n1542);
not  g1553 (n1607, n1536);
buf  g1554 (n1611, n1541);
buf  g1555 (n1575, n1544);
buf  g1556 (n1631, n1544);
buf  g1557 (n1606, n1493);
not  g1558 (n1568, n1543);
buf  g1559 (n1599, n1465);
buf  g1560 (n1618, n1493);
not  g1561 (n1586, n1495);
not  g1562 (n1580, n1545);
not  g1563 (n1565, n1534);
not  g1564 (n1603, n1471);
buf  g1565 (n1590, n1459);
not  g1566 (n1630, n1535);
not  g1567 (n1576, n1541);
buf  g1568 (n1578, n1539);
buf  g1569 (n1615, n1536);
buf  g1570 (n1589, n1550);
not  g1571 (n1567, n1473);
buf  g1572 (n1613, n1464);
buf  g1573 (n1563, n1545);
buf  g1574 (n1617, n1161);
not  g1575 (n1583, n1470);
nand g1576 (n1569, n1469, n1472);
or   g1577 (n1573, n1494, n1460);
or   g1578 (n1610, n1472, n1540, n1539, n1474);
nand g1579 (n1564, n1492, n1156, n1160, n1336);
and  g1580 (n1625, n1548, n1538, n1533, n1549);
or   g1581 (n1612, n1550, n1548, n1541, n1492);
or   g1582 (n1628, n1472, n1458, n1473, n1542);
and  g1583 (n1571, n1537, n1491, n1549);
nand g1584 (n1562, n1159, n1158, n1539, n1543);
nand g1585 (n1570, n1539, n1537, n1336);
xnor g1586 (n1629, n1540, n1536, n1545, n1544);
xor  g1587 (n1588, n1474, n1547, n1491, n1538);
xnor g1588 (n1579, n1546, n1545, n1493, n1535);
nand g1589 (n1584, n1549, n1548, n1543, n1534);
or   g1590 (n1605, n1533, n1337, n1495, n1537);
and  g1591 (n1582, n1541, n1490, n1542, n1547);
and  g1592 (n1614, n1493, n1534, n1494);
or   g1593 (n1622, n1536, n1535, n1540, n1473);
nor  g1594 (n1591, n1336, n1337, n1474, n1495);
nor  g1595 (n1624, n1548, n1533, n1337, n1547);
xor  g1596 (n1620, n1533, n1494, n1471, n1546);
or   g1597 (n1577, n1492, n1542, n1473, n1491);
and  g1598 (n1601, n1475, n1535, n1550, n1466);
and  g1599 (n1600, n1157, n1463, n1540, n1496);
buf  g1600 (n1834, n1612);
not  g1601 (n1794, n1566);
not  g1602 (n1769, n1568);
buf  g1603 (n1793, n1582);
buf  g1604 (n1705, n1618);
buf  g1605 (n1844, n1555);
not  g1606 (n1784, n1593);
not  g1607 (n1648, n1621);
buf  g1608 (n1791, n1559);
not  g1609 (n1811, n1619);
not  g1610 (n1847, n1567);
not  g1611 (n1782, n1594);
not  g1612 (n1816, n1616);
buf  g1613 (n1693, n1341);
buf  g1614 (n1674, n1555);
not  g1615 (n1854, n1561);
buf  g1616 (n1742, n1579);
not  g1617 (n1747, n1573);
not  g1618 (n1745, n1594);
not  g1619 (n1827, n1602);
buf  g1620 (n1634, n1614);
not  g1621 (n1649, n669);
not  g1622 (n1800, n1586);
buf  g1623 (n1741, n1560);
not  g1624 (n1727, n1592);
not  g1625 (n1746, n1572);
not  g1626 (n1732, n1559);
buf  g1627 (n1828, n1603);
not  g1628 (n1724, n1611);
buf  g1629 (n1787, n1570);
not  g1630 (n1721, n1630);
buf  g1631 (n1848, n671);
not  g1632 (n1846, n1551);
buf  g1633 (n1754, n1589);
not  g1634 (n1717, n1592);
buf  g1635 (n1734, n1561);
not  g1636 (n1678, n1206);
buf  g1637 (n1756, n1584);
not  g1638 (n1819, n1621);
not  g1639 (n1656, n1608);
not  g1640 (n1707, n1565);
not  g1641 (n1663, n1558);
not  g1642 (n1807, n1608);
not  g1643 (n1825, n1606);
buf  g1644 (n1633, n1628);
not  g1645 (n1808, n1552);
buf  g1646 (n1760, n1604);
buf  g1647 (n1651, n1624);
not  g1648 (n1829, n1610);
buf  g1649 (n1691, n1588);
not  g1650 (n1711, n1615);
buf  g1651 (n1713, n1581);
not  g1652 (n1655, n1628);
buf  g1653 (n1753, n1584);
buf  g1654 (n1752, n1164);
buf  g1655 (n1809, n672);
not  g1656 (n1720, n1339);
buf  g1657 (n1641, n1626);
buf  g1658 (n1698, n1589);
not  g1659 (n1695, n1632);
buf  g1660 (n1817, n1601);
buf  g1661 (n1673, n1601);
not  g1662 (n1687, n1617);
buf  g1663 (n1843, n1586);
not  g1664 (n1798, n1602);
buf  g1665 (n1683, n1585);
buf  g1666 (n1778, n1480);
not  g1667 (n1661, n1165);
not  g1668 (n1676, n1625);
buf  g1669 (n1670, n1340);
not  g1670 (n1708, n1558);
not  g1671 (n1726, n1616);
buf  g1672 (n1772, n1593);
buf  g1673 (n1743, n1605);
not  g1674 (n1758, n1571);
not  g1675 (n1709, n1566);
not  g1676 (n1737, n1599);
buf  g1677 (n1842, n1426);
buf  g1678 (n1728, n1630);
not  g1679 (n1637, n1581);
not  g1680 (n1749, n1559);
buf  g1681 (n1820, n1340);
buf  g1682 (n1660, n1163);
buf  g1683 (n1821, n1607);
buf  g1684 (n1738, n1598);
not  g1685 (n1748, n1480);
buf  g1686 (n1849, n672);
not  g1687 (n1804, n1617);
not  g1688 (n1740, n1593);
not  g1689 (n1723, n1569);
buf  g1690 (n1658, n1477);
not  g1691 (n1725, n1628);
buf  g1692 (n1715, n1597);
not  g1693 (n1764, n1621);
buf  g1694 (n1735, n1560);
not  g1695 (n1642, n1574);
not  g1696 (n1763, n1562);
not  g1697 (n1675, n1588);
buf  g1698 (n1806, n1631);
buf  g1699 (n1671, n1587);
not  g1700 (n1704, n1612);
buf  g1701 (n1694, n1574);
not  g1702 (n1759, n1622);
not  g1703 (n1803, n1570);
buf  g1704 (n1799, n1162);
not  g1705 (n1666, n1579);
not  g1706 (n1700, n1584);
buf  g1707 (n1852, n1627);
buf  g1708 (n1767, n1424);
buf  g1709 (n1639, n1423);
not  g1710 (n1668, n1596);
buf  g1711 (n1647, n1592);
not  g1712 (n1680, n1611);
buf  g1713 (n1783, n1578);
not  g1714 (n1839, n1572);
buf  g1715 (n1835, n1605);
not  g1716 (n1719, n1565);
not  g1717 (n1654, n1478);
buf  g1718 (n1822, n1166);
not  g1719 (n1712, n1629);
buf  g1720 (n1686, n1166);
buf  g1721 (n1810, n1607);
not  g1722 (n1797, n1527);
buf  g1723 (n1688, n1600);
not  g1724 (n1792, n1426);
not  g1725 (n1702, n1562);
buf  g1726 (n1770, n1579);
buf  g1727 (n1774, n1529);
not  g1728 (n1850, n940);
not  g1729 (n1714, n1629);
buf  g1730 (n1853, n1586);
not  g1731 (n1801, n1425);
not  g1732 (n1729, n1551);
not  g1733 (n1766, n1596);
buf  g1734 (n1833, n1632);
buf  g1735 (n1730, n1599);
not  g1736 (n1744, n1605);
not  g1737 (n1771, n671);
buf  g1738 (n1699, n1564);
buf  g1739 (n1796, n1476);
not  g1740 (n1635, n1574);
not  g1741 (n1838, n1558);
buf  g1742 (n1775, n1594);
not  g1743 (n1837, n1581);
buf  g1744 (n1731, n1583);
buf  g1745 (n1773, n1424);
buf  g1746 (n1710, n1338);
not  g1747 (n1795, n1585);
buf  g1748 (n1823, n1562);
buf  g1749 (n1768, n1481);
and  g1750 (n1640, n1624, n1577, n1553);
and  g1751 (n1813, n1166, n1598, n1614, n1339);
xor  g1752 (n1659, n1599, n1565, n1617, n1556);
or   g1753 (n1677, n1557, n1592, n1496, n1607);
nor  g1754 (n1664, n1425, n1563, n1480, n1554);
xnor g1755 (n1669, n1557, n1426, n1621, n1423);
xor  g1756 (n1785, n1163, n1567, n1424, n1582);
xnor g1757 (n1718, n1164, n1479, n1531, n1555);
nor  g1758 (n1644, n1590, n1580, n1604, n1340);
xor  g1759 (n1780, n1165, n1341, n1563, n1616);
nor  g1760 (n1781, n1574, n1569, n1564, n1619);
or   g1761 (n1814, n1625, n1589, n1594, n1617);
nand g1762 (n1751, n1573, n1573, n1600, n1165);
or   g1763 (n1831, n1570, n1426, n1622, n1587);
nor  g1764 (n1681, n1532, n1568, n1497, n1612);
xnor g1765 (n1696, n1563, n1578, n1613, n1163);
xor  g1766 (n1697, n1570, n1568, n1575, n1609);
xnor g1767 (n1812, n1476, n1338, n1623, n1552);
or   g1768 (n1650, n1575, n1590, n1583, n1609);
xnor g1769 (n1706, n1576, n1618, n1554, n1591);
nand g1770 (n1845, n1595, n1575, n1615, n1497);
and  g1771 (n1638, n1632, n1207, n1477, n1580);
xnor g1772 (n1762, n1496, n1627, n670, n1618);
and  g1773 (n1750, n1564, n1580, n1551, n1582);
and  g1774 (n1739, n1620, n1627, n1586, n1619);
nand g1775 (n1851, n1611, n1476, n1571, n1596);
or   g1776 (n1777, n936, n670, n1163, n1554);
and  g1777 (n1805, n1620, n1571, n1607, n1557);
or   g1778 (n1645, n1591, n1563, n670, n1425);
nand g1779 (n1662, n1619, n1591, n1479, n1578);
and  g1780 (n1682, n1583, n1557, n1208, n1553);
or   g1781 (n1643, n1578, n1631, n1479, n1590);
nor  g1782 (n1840, n1165, n1559, n1604, n1576);
xor  g1783 (n1786, n1587, n1338, n1606, n1610);
and  g1784 (n1646, n1589, n1597, n1422, n1581);
xor  g1785 (n1689, n1614, n1613, n1477, n1424);
and  g1786 (n1701, n1590, n1596, n1624, n1601);
nand g1787 (n1672, n1600, n1553, n1588, n1625);
or   g1788 (n1755, n1591, n1579, n1477, n1595);
xnor g1789 (n1733, n670, n1497, n1599, n1587);
or   g1790 (n1790, n1609, n1624, n1585, n1628);
xor  g1791 (n1761, n1561, n1609, n669, n1564);
or   g1792 (n1665, n939, n1340, n1630, n1569);
xnor g1793 (n1636, n1608, n1476, n1598, n1595);
and  g1794 (n1779, n1580, n1595, n1603, n1481);
and  g1795 (n1832, n1603, n1571, n1584, n1588);
xnor g1796 (n1685, n935, n1602, n1629, n1577);
and  g1797 (n1855, n1569, n1585, n938, n1603);
nand g1798 (n1788, n671, n1478, n1597, n1630);
xnor g1799 (n1824, n1341, n1602, n1601, n1572);
or   g1800 (n1841, n1629, n1164, n1606, n1338);
nor  g1801 (n1692, n1593, n669, n1558, n1423);
xnor g1802 (n1703, n1481, n1166, n1339, n1613);
xnor g1803 (n1765, n1613, n1598, n1605, n1576);
xnor g1804 (n1836, n1610, n1626, n1631);
or   g1805 (n1818, n1615, n1425, n1556, n1528);
or   g1806 (n1716, n1339, n1422, n1572, n1555);
xnor g1807 (n1667, n1618, n1608, n1556, n1497);
and  g1808 (n1802, n1205, n1164, n1620, n1631);
and  g1809 (n1789, n1341, n1610, n1552, n1480);
nor  g1810 (n1815, n1479, n1623, n671, n669);
xor  g1811 (n1757, n1582, n1560, n1562, n1632);
nor  g1812 (n1830, n1627, n1481, n1614, n1478);
and  g1813 (n1657, n1600, n1626, n1576, n1622);
nor  g1814 (n1679, n1611, n1423, n1573, n1597);
or   g1815 (n1722, n1577, n1526, n1623, n1530);
and  g1816 (n1690, n1551, n1583, n1561, n1625);
xnor g1817 (n1684, n1554, n1567, n1568, n1604);
nor  g1818 (n1826, n1556, n1622, n1567, n1566);
nor  g1819 (n1776, n1612, n1552, n1566, n1553);
nand g1820 (n1736, n672, n1616, n1606, n1496);
xnor g1821 (n1653, n1623, n937, n1620, n1615);
xor  g1822 (n1652, n1478, n1575, n1560, n1565);
nor  g1823 (n1937, n1785, n1659, n1791, n1798);
xnor g1824 (n1857, n1769, n1749, n1846, n1817);
nand g1825 (n1875, n1817, n1800, n1734, n1827);
or   g1826 (n1960, n1683, n1823, n1810, n1674);
nand g1827 (n1963, n1818, n1850, n1783, n1777);
nand g1828 (n1982, n1773, n1708, n1770, n1836);
and  g1829 (n1914, n1715, n1778, n1795, n1757);
xnor g1830 (n1978, n1836, n1820, n1822, n1748);
xnor g1831 (n1905, n1707, n1824, n1852, n1780);
xnor g1832 (n1896, n1808, n1712, n1737, n1849);
nand g1833 (n1923, n1825, n1742, n1759, n1807);
xor  g1834 (n1931, n1749, n1790, n1838, n1762);
nand g1835 (n1908, n1842, n1810, n1831, n1837);
or   g1836 (n1885, n1797, n1832, n1660, n1779);
nor  g1837 (n1911, n1850, n1847, n1830, n1826);
xnor g1838 (n1915, n1817, n1842, n1652, n1725);
nor  g1839 (n1866, n1804, n1665, n1774, n1756);
nor  g1840 (n1930, n1781, n1648, n1798, n1760);
xnor g1841 (n1864, n1687, n1801, n1851, n1793);
nor  g1842 (n1925, n1785, n1761, n1830, n1788);
or   g1843 (n1918, n1816, n1705, n1719, n1855);
and  g1844 (n1901, n1826, n1664, n1776, n1787);
xor  g1845 (n1883, n1819, n1783, n1851, n1784);
xor  g1846 (n1909, n1853, n1788, n1699, n1786);
or   g1847 (n1917, n1841, n1789, n1851, n1744);
xnor g1848 (n1942, n1838, n1828, n1786, n1780);
xnor g1849 (n1859, n1807, n1662, n1789, n1803);
nand g1850 (n1916, n1783, n1827, n1677, n1705);
nand g1851 (n1939, n1824, n1852, n1771, n1818);
xor  g1852 (n1959, n1757, n1761, n1710, n1810);
and  g1853 (n1878, n1754, n1754, n1823, n1814);
nand g1854 (n1902, n1784, n1737, n1845, n1841);
xor  g1855 (n1904, n1713, n1821, n1779, n1800);
and  g1856 (n1961, n1736, n1739, n1786, n1721);
nor  g1857 (n1858, n1673, n1649, n1813, n1812);
nor  g1858 (n1899, n1773, n1684, n1730, n1780);
xor  g1859 (n1867, n1690, n1822, n1728, n1782);
nand g1860 (n1919, n1806, n1845, n1679, n1810);
and  g1861 (n1889, n1718, n1831, n1802, n1676);
nand g1862 (n1881, n1835, n1829, n1682, n1772);
nor  g1863 (n1862, n1655, n1650, n1852, n1809);
nor  g1864 (n1892, n1837, n1805, n1835, n1840);
or   g1865 (n1922, n1828, n1815, n1692);
xnor g1866 (n1967, n1829, n1709, n1818, n1775);
and  g1867 (n1893, n1803, n1846, n1755, n1784);
nand g1868 (n1983, n1747, n1724, n1833);
nor  g1869 (n1980, n1731, n1832, n1654, n1822);
nor  g1870 (n1962, n1796, n1732, n1731, n1704);
or   g1871 (n1928, n1694, n1789, n1779, n1806);
nor  g1872 (n1977, n1672, n1792, n1712, n1796);
or   g1873 (n1964, n1762, n1831, n1855, n1790);
and  g1874 (n1870, n1787, n1675, n1726, n1729);
xnor g1875 (n1953, n1847, n1719, n1803, n1741);
xnor g1876 (n1865, n1841, n1752, n1742, n1738);
xor  g1877 (n1884, n1793, n1748, n1693, n1667);
xnor g1878 (n1907, n1834, n1839, n1668);
nor  g1879 (n1880, n1835, n1815, n1799, n1670);
xnor g1880 (n1946, n1780, n1855, n1788, n1797);
and  g1881 (n1932, n1720, n1822, n1782, n1763);
nand g1882 (n1948, n1722, n672, n1814, n1807);
nand g1883 (n1936, n1854, n1771, n1849, n1697);
xor  g1884 (n1945, n1813, n1811, n1847, n1735);
or   g1885 (n1888, n1707, n1824, n1821, n1784);
or   g1886 (n1876, n1714, n1766, n1691, n1743);
or   g1887 (n1934, n1702, n1853, n1729, n1799);
xnor g1888 (n1981, n1808, n1826, n1829, n1811);
or   g1889 (n1951, n1750, n1767, n1755, n1723);
nand g1890 (n1920, n1788, n1850, n1710, n1686);
or   g1891 (n1898, n1815, n1803, n1769, n1844);
nor  g1892 (n1906, n1842, n1739, n1651, n1703);
nand g1893 (n1944, n1772, n1841, n1812, n1848);
xnor g1894 (n1974, n1658, n1838, n1805, n1745);
or   g1895 (n1968, n1701, n1794, n1795, n1793);
or   g1896 (n1900, n1801, n1730, n1716, n1802);
and  g1897 (n1891, n1718, n1753, n1818, n1775);
or   g1898 (n1860, n1843, n1816, n1758, n1751);
nand g1899 (n1926, n1740, n1819, n1760, n1720);
xnor g1900 (n1933, n1848, n1804, n1727, n1809);
and  g1901 (n1938, n1825, n1827, n1799, n1661);
and  g1902 (n1950, n1798, n1768, n1716, n1844);
nand g1903 (n1913, n1721, n1787, n1774, n1843);
xnor g1904 (n1975, n1656, n1826, n1767, n1795);
nor  g1905 (n1887, n1725, n1843, n1806, n1756);
nand g1906 (n1869, n1819, n1820, n1698, n1778);
or   g1907 (n1965, n1765, n1759, n1681, n1744);
xnor g1908 (n1856, n1800, n1834, n1835, n1746);
xnor g1909 (n1976, n1752, n1777, n1852, n1740);
or   g1910 (n1903, n1847, n1838, n1798, n1781);
xnor g1911 (n1895, n1824, n1845, n1827, n1792);
or   g1912 (n1873, n1823, n1669, n1854, n1829);
xnor g1913 (n1863, n1703, n1790, n1836, n1746);
and  g1914 (n1958, n1816, n1840, n1854, n1741);
xnor g1915 (n1890, n1808, n1783, n1776, n1657);
nand g1916 (n1971, n1817, n1821, n1695);
and  g1917 (n1868, n1723, n1671, n1764, n1728);
nor  g1918 (n1955, n1846, n1732, n1850, n1830);
xor  g1919 (n1877, n1706, n1825, n1805, n1804);
and  g1920 (n1979, n1794, n1834, n1704, n1848);
nor  g1921 (n1947, n1717, n1666, n1812, n1696);
xor  g1922 (n1966, n1711, n1766, n1724, n1688);
and  g1923 (n1897, n1796, n1751, n1753, n1781);
nand g1924 (n1874, n1765, n1782, n1853, n1792);
and  g1925 (n1935, n1812, n1828, n1685, n1813);
or   g1926 (n1910, n1809, n1787, n1792, n1848);
or   g1927 (n1894, n1770, n1709, n1830, n1717);
xor  g1928 (n1929, n1777, n1804, n1811, n1789);
or   g1929 (n1957, n1785, n1796, n1708, n1700);
xnor g1930 (n1984, n1745, n1747, n1791, n1823);
xor  g1931 (n1886, n1797, n1779, n1813, n1849);
xnor g1932 (n1924, n1734, n1736, n1786, n1842);
nor  g1933 (n1940, n1778, n1722, n1794, n1833);
nor  g1934 (n1969, n1689, n1836, n1840, n1839);
xor  g1935 (n1927, n1678, n1844, n1849, n1743);
nand g1936 (n1941, n1844, n1811, n1807, n1733);
or   g1937 (n1871, n1834, n1768, n1819, n1790);
and  g1938 (n1861, n1843, n1750, n1820, n1833);
nor  g1939 (n1912, n1663, n1738, n1714, n1764);
nor  g1940 (n1970, n1801, n1735, n1797, n1799);
nor  g1941 (n1985, n1832, n1837, n1733, n1706);
xnor g1942 (n1949, n1854, n1653, n1828, n1846);
xnor g1943 (n1879, n1777, n1713, n1781, n1839);
nor  g1944 (n1872, n1809, n1851, n1727, n1831);
or   g1945 (n1956, n1806, n1845, n1715, n1711);
and  g1946 (n1973, n1795, n1853, n1802, n1832);
nand g1947 (n1921, n1808, n1782, n1814, n1794);
or   g1948 (n1972, n1778, n1802, n1801, n1800);
xor  g1949 (n1882, n1840, n1758, n1814, n1805);
and  g1950 (n1954, n1785, n1816, n1680, n1820);
nor  g1951 (n1943, n1763, n1825, n1793, n1855);
nand g1952 (n1952, n1837, n1791, n1726);
xor  g1953 (n2013, n1896, n1912, n1931, n1902);
or   g1954 (n2004, n1978, n1939, n1895, n1893);
and  g1955 (n2007, n1944, n1905, n1900, n1907);
nor  g1956 (n2015, n1954, n1929, n1947, n1867);
nor  g1957 (n1998, n1903, n1878, n1924, n1964);
or   g1958 (n1996, n1973, n1914, n1983, n1962);
or   g1959 (n2012, n1937, n1943, n1934, n1857);
xor  g1960 (n1988, n1864, n1955, n1891, n1872);
or   g1961 (n2017, n1927, n1894, n1909, n1963);
xor  g1962 (n2016, n1925, n1911, n1877, n1887);
xnor g1963 (n2011, n1948, n1960, n1921, n1976);
xor  g1964 (n1994, n1908, n1886, n1979, n1951);
xnor g1965 (n2005, n1888, n1901, n1946, n1974);
nand g1966 (n1993, n1889, n1860, n1862, n1972);
nand g1967 (n1986, n1874, n1922, n1869, n1910);
or   g1968 (n2000, n1950, n1885, n1861, n1923);
xnor g1969 (n2006, n1980, n1898, n1906, n1875);
or   g1970 (n1991, n1913, n1904, n1949, n1940);
nor  g1971 (n2008, n1965, n1871, n1881, n1932);
xnor g1972 (n1989, n1868, n1956, n1942, n1866);
xnor g1973 (n1992, n1953, n1897, n1941, n1967);
nand g1974 (n1995, n1938, n1982, n1945, n1933);
or   g1975 (n2009, n1926, n1957, n1918, n1928);
or   g1976 (n2002, n1879, n1920, n1961, n1890);
nand g1977 (n2014, n1970, n1892, n1884, n1975);
nor  g1978 (n2010, n1880, n1856, n1968, n1916);
nand g1979 (n2001, n1876, n1873, n1959, n1883);
nand g1980 (n2003, n1935, n1958, n1882, n1870);
and  g1981 (n1997, n1952, n1930, n1859, n1971);
xor  g1982 (n1987, n1917, n1915, n1865, n1899);
xor  g1983 (n1999, n1981, n1919, n1977, n1863);
nand g1984 (n1990, n1969, n1936, n1966, n1858);
not  g1985 (n2020, n1988);
not  g1986 (n2018, n1993);
xnor g1987 (n2021, n1985, n1986);
xnor g1988 (n2022, n1990, n1984);
nor  g1989 (n2019, n1992, n1987, n1989, n1991);
nor  g1990 (n2025, n2022, n1999, n2010, n1998);
or   g1991 (n2026, n2001, n2017, n2011, n2003);
xnor g1992 (n2024, n2007, n2020, n2009, n2021);
xnor g1993 (n2027, n1996, n2004, n2022, n2019);
nand g1994 (n2029, n2016, n1997, n2014, n2006);
xnor g1995 (n2023, n2013, n2022, n2000, n2008);
nand g1996 (n2030, n2015, n2018, n2012, n1994);
and  g1997 (n2028, n2022, n1995, n2005, n2002);
nand g1998 (n2032, n2026, n2023, n2027, n2030);
xnor g1999 (n2031, n2028, n2029, n2024, n2025);
endmodule
