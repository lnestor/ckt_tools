// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_4000_362 written by SynthGen on 2021/04/05 11:24:27
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_4000_362 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n1141, n1144, n1227, n1235, n1230, n1228, n3849, n3850,
 n3855, n3848, n3851, n3856, n3854, n3847, n4020, n4025,
 n4021, n4026, n4018, n4027, n4031, n4024, n4016, n4032,
 n4029, n4017, n4028, n4015, n4030, n4022, n4023, n4019);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n1141, n1144, n1227, n1235, n1230, n1228, n3849, n3850,
 n3855, n3848, n3851, n3856, n3854, n3847, n4020, n4025,
 n4021, n4026, n4018, n4027, n4031, n4024, n4016, n4032,
 n4029, n4017, n4028, n4015, n4030, n4022, n4023, n4019;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1142, n1143, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1229, n1231, n1232, n1233, n1234, n1236, n1237, n1238,
 n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
 n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
 n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
 n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
 n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
 n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
 n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
 n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
 n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
 n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
 n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
 n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
 n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
 n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
 n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
 n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
 n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
 n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
 n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
 n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
 n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
 n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
 n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
 n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
 n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
 n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
 n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
 n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
 n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
 n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
 n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
 n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
 n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
 n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
 n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
 n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
 n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
 n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
 n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
 n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
 n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
 n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
 n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
 n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
 n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
 n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
 n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
 n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
 n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
 n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
 n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
 n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
 n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
 n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
 n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
 n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
 n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
 n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
 n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
 n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
 n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
 n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
 n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
 n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
 n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
 n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
 n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
 n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
 n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
 n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
 n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
 n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
 n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
 n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
 n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
 n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
 n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
 n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
 n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
 n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
 n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
 n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
 n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
 n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
 n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
 n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926,
 n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
 n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
 n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
 n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
 n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966,
 n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
 n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
 n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
 n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
 n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006,
 n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
 n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
 n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
 n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
 n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046,
 n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
 n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
 n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
 n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
 n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086,
 n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
 n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
 n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
 n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
 n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126,
 n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
 n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
 n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
 n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
 n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166,
 n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
 n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
 n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
 n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
 n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206,
 n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
 n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
 n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
 n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
 n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246,
 n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
 n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
 n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
 n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
 n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286,
 n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
 n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
 n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
 n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
 n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326,
 n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
 n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
 n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
 n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
 n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366,
 n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
 n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
 n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
 n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
 n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406,
 n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
 n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
 n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
 n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
 n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446,
 n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
 n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
 n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
 n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
 n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486,
 n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
 n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
 n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
 n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
 n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526,
 n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
 n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
 n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
 n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
 n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566,
 n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
 n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
 n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
 n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
 n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606,
 n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
 n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
 n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
 n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
 n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
 n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
 n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
 n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
 n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
 n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
 n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
 n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
 n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
 n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
 n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
 n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
 n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
 n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
 n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
 n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
 n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
 n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
 n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
 n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
 n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
 n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
 n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
 n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
 n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
 n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
 n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
 n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
 n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
 n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
 n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
 n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
 n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
 n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
 n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
 n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
 n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
 n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
 n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
 n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
 n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
 n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
 n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
 n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
 n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
 n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
 n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
 n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
 n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
 n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
 n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
 n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
 n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
 n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
 n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
 n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
 n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
 n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
 n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
 n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
 n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
 n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
 n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
 n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
 n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
 n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
 n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
 n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
 n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
 n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
 n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
 n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
 n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
 n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
 n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
 n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
 n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
 n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
 n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
 n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
 n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
 n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
 n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
 n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
 n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
 n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
 n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
 n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
 n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
 n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
 n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
 n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
 n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
 n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
 n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
 n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
 n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
 n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
 n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
 n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
 n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
 n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
 n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
 n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
 n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
 n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
 n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
 n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
 n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
 n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
 n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
 n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
 n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
 n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
 n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
 n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
 n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
 n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
 n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
 n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
 n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
 n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
 n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
 n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
 n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
 n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
 n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
 n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
 n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
 n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
 n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
 n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
 n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
 n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
 n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
 n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
 n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
 n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
 n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
 n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
 n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
 n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
 n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
 n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
 n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
 n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
 n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
 n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
 n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
 n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
 n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
 n3852, n3853, n3857, n3858, n3859, n3860, n3861, n3862,
 n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
 n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
 n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
 n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
 n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
 n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
 n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
 n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926,
 n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
 n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
 n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
 n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
 n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966,
 n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
 n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
 n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
 n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
 n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006,
 n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014;

buf  g0 (n127, n28);
not  g1 (n141, n27);
buf  g2 (n113, n8);
buf  g3 (n117, n16);
not  g4 (n47, n5);
not  g5 (n84, n19);
buf  g6 (n147, n6);
not  g7 (n115, n5);
buf  g8 (n49, n23);
buf  g9 (n62, n1);
not  g10 (n154, n4);
not  g11 (n121, n29);
buf  g12 (n157, n30);
buf  g13 (n64, n7);
not  g14 (n80, n31);
not  g15 (n158, n13);
buf  g16 (n107, n14);
buf  g17 (n79, n12);
buf  g18 (n52, n15);
not  g19 (n125, n28);
buf  g20 (n82, n16);
buf  g21 (n138, n24);
buf  g22 (n54, n17);
not  g23 (n37, n7);
buf  g24 (n71, n28);
buf  g25 (n57, n27);
not  g26 (n55, n18);
not  g27 (n122, n24);
not  g28 (n88, n3);
buf  g29 (n81, n11);
not  g30 (n143, n23);
not  g31 (n38, n20);
not  g32 (n61, n26);
buf  g33 (n36, n32);
not  g34 (n53, n15);
not  g35 (n68, n4);
buf  g36 (n41, n19);
buf  g37 (n108, n31);
buf  g38 (n102, n6);
buf  g39 (n95, n20);
buf  g40 (n46, n18);
buf  g41 (n150, n19);
buf  g42 (n51, n17);
buf  g43 (n59, n25);
buf  g44 (n50, n26);
not  g45 (n91, n4);
not  g46 (n69, n16);
not  g47 (n101, n8);
not  g48 (n151, n13);
not  g49 (n145, n1);
not  g50 (n146, n2);
not  g51 (n112, n9);
buf  g52 (n83, n30);
not  g53 (n120, n29);
not  g54 (n153, n22);
buf  g55 (n130, n11);
not  g56 (n74, n19);
buf  g57 (n40, n25);
not  g58 (n48, n2);
not  g59 (n44, n21);
not  g60 (n124, n22);
buf  g61 (n39, n25);
buf  g62 (n98, n29);
buf  g63 (n92, n8);
not  g64 (n137, n21);
buf  g65 (n72, n27);
buf  g66 (n65, n11);
buf  g67 (n100, n10);
not  g68 (n142, n22);
buf  g69 (n60, n18);
not  g70 (n152, n20);
buf  g71 (n110, n2);
buf  g72 (n86, n32);
buf  g73 (n104, n13);
not  g74 (n63, n27);
not  g75 (n77, n28);
buf  g76 (n136, n12);
buf  g77 (n135, n18);
not  g78 (n155, n30);
buf  g79 (n129, n9);
not  g80 (n149, n29);
not  g81 (n106, n17);
buf  g82 (n111, n6);
not  g83 (n33, n10);
buf  g84 (n43, n9);
not  g85 (n132, n25);
not  g86 (n109, n12);
not  g87 (n73, n3);
buf  g88 (n134, n11);
buf  g89 (n144, n5);
not  g90 (n118, n14);
buf  g91 (n128, n31);
not  g92 (n148, n6);
not  g93 (n105, n10);
not  g94 (n99, n1);
buf  g95 (n66, n9);
buf  g96 (n126, n15);
not  g97 (n96, n13);
not  g98 (n140, n14);
not  g99 (n133, n31);
buf  g100 (n42, n30);
buf  g101 (n34, n3);
buf  g102 (n45, n3);
buf  g103 (n156, n8);
buf  g104 (n67, n4);
not  g105 (n139, n10);
not  g106 (n76, n7);
not  g107 (n87, n24);
not  g108 (n94, n20);
buf  g109 (n90, n26);
not  g110 (n103, n15);
buf  g111 (n97, n22);
buf  g112 (n75, n26);
buf  g113 (n89, n12);
not  g114 (n119, n17);
not  g115 (n93, n16);
not  g116 (n114, n5);
buf  g117 (n78, n1);
buf  g118 (n56, n2);
buf  g119 (n35, n21);
buf  g120 (n85, n23);
buf  g121 (n131, n23);
not  g122 (n58, n21);
not  g123 (n70, n7);
not  g124 (n123, n24);
buf  g125 (n116, n14);
buf  g126 (n565, n94);
buf  g127 (n353, n74);
not  g128 (n372, n73);
not  g129 (n275, n85);
not  g130 (n197, n78);
buf  g131 (n534, n96);
not  g132 (n180, n66);
buf  g133 (n484, n95);
not  g134 (n216, n62);
not  g135 (n546, n36);
not  g136 (n417, n83);
not  g137 (n596, n93);
buf  g138 (n261, n79);
buf  g139 (n203, n77);
buf  g140 (n254, n106);
not  g141 (n271, n38);
buf  g142 (n475, n50);
buf  g143 (n260, n66);
buf  g144 (n218, n129);
not  g145 (n503, n108);
buf  g146 (n205, n47);
not  g147 (n226, n84);
not  g148 (n557, n123);
buf  g149 (n198, n117);
buf  g150 (n366, n108);
not  g151 (n194, n103);
not  g152 (n233, n44);
buf  g153 (n377, n94);
not  g154 (n617, n73);
buf  g155 (n295, n137);
buf  g156 (n424, n40);
buf  g157 (n431, n72);
not  g158 (n435, n61);
buf  g159 (n552, n93);
not  g160 (n612, n51);
buf  g161 (n515, n112);
buf  g162 (n455, n138);
not  g163 (n352, n83);
buf  g164 (n371, n127);
not  g165 (n615, n146);
buf  g166 (n597, n124);
buf  g167 (n419, n100);
not  g168 (n299, n97);
buf  g169 (n509, n96);
not  g170 (n441, n43);
buf  g171 (n554, n103);
not  g172 (n587, n136);
buf  g173 (n376, n79);
buf  g174 (n318, n39);
buf  g175 (n578, n103);
buf  g176 (n304, n110);
buf  g177 (n362, n126);
not  g178 (n330, n82);
buf  g179 (n526, n47);
buf  g180 (n355, n132);
buf  g181 (n429, n85);
buf  g182 (n327, n62);
buf  g183 (n363, n129);
not  g184 (n195, n146);
not  g185 (n505, n89);
not  g186 (n476, n107);
buf  g187 (n217, n35);
buf  g188 (n365, n49);
buf  g189 (n406, n77);
not  g190 (n234, n40);
not  g191 (n309, n103);
not  g192 (n305, n139);
not  g193 (n199, n65);
buf  g194 (n258, n124);
buf  g195 (n374, n122);
buf  g196 (n585, n87);
not  g197 (n164, n87);
buf  g198 (n408, n131);
buf  g199 (n346, n124);
buf  g200 (n522, n99);
not  g201 (n206, n62);
not  g202 (n191, n61);
buf  g203 (n277, n130);
buf  g204 (n265, n36);
buf  g205 (n564, n76);
buf  g206 (n321, n109);
not  g207 (n189, n65);
not  g208 (n286, n87);
not  g209 (n481, n100);
buf  g210 (n458, n115);
buf  g211 (n350, n70);
not  g212 (n369, n60);
not  g213 (n202, n63);
buf  g214 (n245, n149);
not  g215 (n457, n97);
not  g216 (n536, n130);
buf  g217 (n176, n110);
buf  g218 (n387, n53);
buf  g219 (n425, n106);
not  g220 (n323, n88);
not  g221 (n613, n114);
buf  g222 (n439, n133);
not  g223 (n568, n44);
not  g224 (n361, n92);
buf  g225 (n200, n71);
buf  g226 (n242, n50);
not  g227 (n506, n99);
not  g228 (n220, n136);
not  g229 (n231, n75);
not  g230 (n246, n34);
buf  g231 (n373, n68);
not  g232 (n300, n49);
buf  g233 (n567, n140);
not  g234 (n586, n81);
not  g235 (n268, n83);
buf  g236 (n338, n149);
not  g237 (n625, n130);
buf  g238 (n291, n121);
buf  g239 (n276, n53);
buf  g240 (n310, n143);
buf  g241 (n279, n129);
buf  g242 (n285, n86);
buf  g243 (n219, n87);
not  g244 (n456, n146);
buf  g245 (n436, n46);
buf  g246 (n328, n55);
buf  g247 (n336, n136);
not  g248 (n201, n45);
buf  g249 (n228, n69);
buf  g250 (n404, n56);
buf  g251 (n392, n41);
buf  g252 (n422, n130);
not  g253 (n620, n45);
buf  g254 (n434, n48);
not  g255 (n224, n125);
not  g256 (n560, n52);
not  g257 (n574, n69);
buf  g258 (n208, n51);
not  g259 (n614, n38);
buf  g260 (n595, n145);
not  g261 (n513, n117);
buf  g262 (n345, n116);
not  g263 (n561, n117);
not  g264 (n298, n98);
buf  g265 (n530, n70);
not  g266 (n500, n135);
not  g267 (n510, n141);
not  g268 (n379, n82);
not  g269 (n533, n122);
buf  g270 (n196, n65);
not  g271 (n524, n54);
buf  g272 (n284, n48);
buf  g273 (n253, n70);
buf  g274 (n339, n132);
buf  g275 (n581, n138);
not  g276 (n390, n78);
not  g277 (n433, n120);
buf  g278 (n239, n78);
buf  g279 (n320, n101);
not  g280 (n335, n122);
not  g281 (n440, n64);
buf  g282 (n263, n55);
buf  g283 (n472, n81);
not  g284 (n172, n60);
not  g285 (n532, n37);
buf  g286 (n237, n39);
not  g287 (n332, n47);
not  g288 (n187, n126);
buf  g289 (n572, n88);
not  g290 (n382, n128);
buf  g291 (n540, n33);
buf  g292 (n499, n107);
buf  g293 (n486, n126);
not  g294 (n492, n144);
buf  g295 (n368, n56);
buf  g296 (n415, n75);
buf  g297 (n529, n85);
not  g298 (n479, n101);
not  g299 (n531, n50);
not  g300 (n460, n33);
not  g301 (n541, n58);
not  g302 (n468, n142);
not  g303 (n311, n147);
buf  g304 (n504, n76);
not  g305 (n316, n42);
not  g306 (n412, n40);
not  g307 (n451, n37);
buf  g308 (n255, n58);
not  g309 (n488, n67);
buf  g310 (n495, n102);
buf  g311 (n493, n100);
not  g312 (n243, n98);
not  g313 (n293, n91);
buf  g314 (n525, n127);
not  g315 (n539, n99);
not  g316 (n396, n54);
not  g317 (n348, n147);
buf  g318 (n223, n91);
buf  g319 (n438, n59);
buf  g320 (n443, n51);
buf  g321 (n329, n65);
not  g322 (n409, n94);
not  g323 (n272, n48);
buf  g324 (n563, n144);
buf  g325 (n312, n118);
not  g326 (n256, n44);
buf  g327 (n393, n81);
not  g328 (n426, n51);
not  g329 (n494, n36);
buf  g330 (n463, n61);
buf  g331 (n559, n53);
buf  g332 (n236, n42);
not  g333 (n592, n81);
not  g334 (n183, n35);
not  g335 (n548, n108);
not  g336 (n259, n64);
buf  g337 (n502, n41);
not  g338 (n283, n69);
not  g339 (n221, n112);
not  g340 (n177, n62);
not  g341 (n623, n145);
not  g342 (n542, n148);
buf  g343 (n421, n93);
not  g344 (n163, n52);
buf  g345 (n577, n132);
buf  g346 (n580, n109);
buf  g347 (n303, n63);
not  g348 (n514, n118);
not  g349 (n364, n92);
buf  g350 (n257, n96);
not  g351 (n576, n148);
not  g352 (n167, n143);
not  g353 (n611, n123);
not  g354 (n621, n104);
buf  g355 (n528, n116);
buf  g356 (n354, n131);
buf  g357 (n401, n127);
not  g358 (n159, n77);
not  g359 (n566, n98);
buf  g360 (n241, n68);
not  g361 (n498, n91);
buf  g362 (n383, n147);
buf  g363 (n301, n80);
not  g364 (n604, n41);
buf  g365 (n414, n71);
buf  g366 (n170, n80);
buf  g367 (n386, n112);
not  g368 (n603, n76);
buf  g369 (n278, n141);
not  g370 (n508, n105);
buf  g371 (n477, n113);
not  g372 (n485, n66);
buf  g373 (n262, n101);
buf  g374 (n399, n43);
not  g375 (n518, n97);
buf  g376 (n297, n140);
not  g377 (n391, n68);
buf  g378 (n582, n95);
not  g379 (n606, n147);
not  g380 (n331, n39);
buf  g381 (n473, n139);
not  g382 (n192, n80);
not  g383 (n471, n133);
buf  g384 (n315, n117);
buf  g385 (n411, n140);
buf  g386 (n292, n115);
not  g387 (n445, n135);
not  g388 (n290, n72);
buf  g389 (n496, n53);
buf  g390 (n227, n102);
buf  g391 (n590, n143);
not  g392 (n161, n135);
buf  g393 (n388, n94);
not  g394 (n222, n92);
not  g395 (n470, n123);
buf  g396 (n340, n120);
not  g397 (n326, n142);
not  g398 (n232, n46);
buf  g399 (n521, n34);
buf  g400 (n235, n84);
buf  g401 (n249, n61);
buf  g402 (n584, n89);
buf  g403 (n593, n113);
not  g404 (n179, n104);
not  g405 (n359, n148);
not  g406 (n333, n134);
not  g407 (n594, n128);
buf  g408 (n357, n104);
not  g409 (n400, n96);
not  g410 (n190, n122);
buf  g411 (n535, n50);
buf  g412 (n413, n40);
buf  g413 (n307, n71);
not  g414 (n169, n119);
buf  g415 (n247, n71);
not  g416 (n405, n121);
buf  g417 (n461, n63);
not  g418 (n251, n38);
buf  g419 (n501, n58);
not  g420 (n394, n89);
not  g421 (n474, n73);
buf  g422 (n410, n83);
not  g423 (n193, n37);
not  g424 (n547, n121);
not  g425 (n543, n127);
buf  g426 (n314, n86);
buf  g427 (n238, n88);
not  g428 (n381, n35);
buf  g429 (n482, n107);
buf  g430 (n428, n60);
buf  g431 (n446, n134);
not  g432 (n287, n133);
not  g433 (n230, n134);
buf  g434 (n296, n60);
not  g435 (n448, n46);
buf  g436 (n356, n99);
buf  g437 (n512, n98);
buf  g438 (n166, n85);
not  g439 (n306, n125);
buf  g440 (n416, n116);
buf  g441 (n599, n86);
buf  g442 (n308, n140);
buf  g443 (n491, n143);
buf  g444 (n370, n138);
buf  g445 (n527, n110);
buf  g446 (n252, n102);
buf  g447 (n608, n112);
buf  g448 (n583, n131);
not  g449 (n325, n45);
buf  g450 (n489, n137);
not  g451 (n610, n74);
buf  g452 (n516, n90);
buf  g453 (n210, n120);
buf  g454 (n294, n145);
not  g455 (n168, n118);
not  g456 (n322, n114);
buf  g457 (n553, n90);
not  g458 (n403, n105);
buf  g459 (n380, n115);
not  g460 (n624, n56);
not  g461 (n453, n106);
buf  g462 (n579, n55);
buf  g463 (n215, n138);
buf  g464 (n267, n35);
not  g465 (n324, n48);
not  g466 (n437, n105);
buf  g467 (n464, n109);
not  g468 (n588, n59);
buf  g469 (n174, n120);
buf  g470 (n282, n131);
buf  g471 (n490, n146);
not  g472 (n337, n57);
not  g473 (n558, n33);
buf  g474 (n273, n107);
not  g475 (n537, n52);
not  g476 (n511, n44);
buf  g477 (n162, n135);
not  g478 (n447, n93);
buf  g479 (n619, n79);
buf  g480 (n367, n82);
buf  g481 (n598, n97);
not  g482 (n384, n86);
not  g483 (n545, n34);
buf  g484 (n589, n54);
buf  g485 (n186, n148);
not  g486 (n351, n82);
not  g487 (n274, n57);
buf  g488 (n555, n69);
buf  g489 (n622, n38);
not  g490 (n165, n45);
not  g491 (n469, n125);
not  g492 (n398, n123);
not  g493 (n181, n139);
not  g494 (n375, n58);
not  g495 (n289, n68);
buf  g496 (n212, n42);
buf  g497 (n211, n75);
not  g498 (n467, n88);
buf  g499 (n569, n90);
buf  g500 (n317, n41);
buf  g501 (n517, n116);
buf  g502 (n160, n89);
buf  g503 (n188, n37);
not  g504 (n250, n137);
not  g505 (n378, n64);
buf  g506 (n430, n74);
buf  g507 (n319, n64);
not  g508 (n618, n141);
not  g509 (n523, n33);
buf  g510 (n550, n57);
not  g511 (n402, n70);
buf  g512 (n483, n136);
buf  g513 (n480, n72);
buf  g514 (n538, n114);
buf  g515 (n344, n139);
buf  g516 (n601, n57);
buf  g517 (n389, n109);
buf  g518 (n450, n101);
not  g519 (n449, n128);
not  g520 (n213, n92);
buf  g521 (n184, n137);
not  g522 (n605, n132);
not  g523 (n459, n118);
buf  g524 (n171, n76);
buf  g525 (n178, n39);
not  g526 (n360, n113);
buf  g527 (n280, n66);
not  g528 (n288, n100);
buf  g529 (n616, n126);
buf  g530 (n432, n104);
not  g531 (n385, n114);
buf  g532 (n407, n144);
buf  g533 (n607, n119);
buf  g534 (n266, n108);
not  g535 (n544, n63);
buf  g536 (n209, n95);
not  g537 (n556, n111);
not  g538 (n427, n77);
not  g539 (n444, n34);
not  g540 (n204, n80);
not  g541 (n397, n124);
not  g542 (n573, n67);
buf  g543 (n487, n56);
buf  g544 (n225, n73);
buf  g545 (n519, n128);
buf  g546 (n347, n59);
not  g547 (n575, n79);
not  g548 (n571, n105);
not  g549 (n462, n145);
buf  g550 (n343, n102);
buf  g551 (n229, n84);
not  g552 (n240, n141);
not  g553 (n570, n142);
not  g554 (n466, n47);
not  g555 (n349, n55);
not  g556 (n602, n49);
buf  g557 (n442, n113);
not  g558 (n423, n42);
buf  g559 (n549, n106);
buf  g560 (n395, n119);
buf  g561 (n334, n46);
not  g562 (n600, n144);
not  g563 (n562, n84);
not  g564 (n452, n90);
not  g565 (n185, n133);
buf  g566 (n420, n129);
buf  g567 (n207, n67);
not  g568 (n281, n119);
not  g569 (n269, n115);
buf  g570 (n465, n59);
not  g571 (n507, n149);
buf  g572 (n341, n95);
not  g573 (n244, n52);
not  g574 (n418, n110);
not  g575 (n478, n43);
not  g576 (n497, n91);
buf  g577 (n342, n134);
buf  g578 (n520, n43);
not  g579 (n302, n111);
not  g580 (n609, n78);
buf  g581 (n173, n72);
not  g582 (n313, n111);
buf  g583 (n358, n74);
buf  g584 (n182, n67);
buf  g585 (n551, n36);
not  g586 (n248, n75);
not  g587 (n175, n54);
buf  g588 (n214, n49);
buf  g589 (n270, n142);
buf  g590 (n454, n121);
buf  g591 (n591, n111);
buf  g592 (n264, n125);
buf  g593 (n705, n527);
buf  g594 (n699, n332);
buf  g595 (n636, n340);
buf  g596 (n1020, n424);
buf  g597 (n731, n592);
buf  g598 (n628, n229);
not  g599 (n854, n248);
not  g600 (n929, n577);
buf  g601 (n693, n342);
buf  g602 (n856, n502);
buf  g603 (n914, n340);
not  g604 (n1048, n544);
buf  g605 (n665, n287);
not  g606 (n1090, n610);
buf  g607 (n772, n185);
buf  g608 (n938, n538);
buf  g609 (n751, n329);
buf  g610 (n804, n497);
buf  g611 (n1110, n204);
buf  g612 (n1052, n344);
buf  g613 (n1008, n328);
not  g614 (n631, n226);
not  g615 (n808, n420);
buf  g616 (n944, n378);
not  g617 (n737, n623);
not  g618 (n775, n549);
not  g619 (n1105, n277);
not  g620 (n1095, n573);
not  g621 (n956, n187);
buf  g622 (n717, n504);
not  g623 (n695, n245);
buf  g624 (n662, n588);
buf  g625 (n1039, n270);
not  g626 (n960, n364);
not  g627 (n786, n250);
buf  g628 (n849, n294);
nor  g629 (n1078, n503, n335, n372, n442);
nor  g630 (n839, n533, n272, n432, n244);
nor  g631 (n677, n398, n553, n166, n365);
nand g632 (n1050, n503, n520, n190, n555);
xor  g633 (n824, n576, n308, n269, n619);
and  g634 (n716, n382, n550, n177, n482);
xor  g635 (n1031, n178, n274, n303, n270);
nor  g636 (n904, n397, n204, n175, n336);
xor  g637 (n656, n162, n349, n262, n310);
and  g638 (n889, n511, n421, n229, n233);
and  g639 (n947, n207, n381, n185, n521);
nor  g640 (n919, n416, n263, n196, n172);
nand g641 (n638, n583, n206, n445, n441);
and  g642 (n753, n555, n188, n334, n210);
xnor g643 (n723, n506, n607, n246, n416);
or   g644 (n846, n546, n243, n349, n162);
or   g645 (n762, n413, n401, n415, n503);
xor  g646 (n711, n273, n547, n388, n305);
nor  g647 (n1072, n328, n603, n248, n494);
and  g648 (n1003, n585, n488, n283, n264);
or   g649 (n814, n344, n567, n622, n279);
xnor g650 (n822, n266, n405, n472, n327);
nand g651 (n684, n391, n616, n522, n169);
or   g652 (n853, n179, n427, n437, n291);
nor  g653 (n1044, n460, n180, n340, n547);
xnor g654 (n785, n443, n224, n235, n298);
nand g655 (n881, n496, n473, n358, n318);
nand g656 (n877, n383, n367, n365, n488);
and  g657 (n958, n591, n513, n236, n304);
nand g658 (n727, n623, n616, n585, n170);
or   g659 (n626, n534, n388, n605, n198);
xnor g660 (n851, n409, n556, n278, n289);
nand g661 (n870, n199, n591, n551, n183);
or   g662 (n812, n558, n423, n599, n550);
xnor g663 (n663, n371, n526, n305, n198);
nand g664 (n734, n586, n448, n453, n366);
or   g665 (n689, n223, n621, n438, n389);
xnor g666 (n992, n608, n588, n182, n169);
and  g667 (n967, n289, n430, n557, n398);
or   g668 (n761, n311, n508, n537, n545);
nand g669 (n726, n512, n418, n218, n610);
nor  g670 (n1042, n456, n540, n195, n220);
and  g671 (n707, n300, n342, n619, n452);
nand g672 (n879, n168, n460, n335, n344);
nand g673 (n791, n454, n431, n261, n205);
nor  g674 (n900, n375, n571, n621, n196);
nor  g675 (n680, n552, n398, n558, n602);
nor  g676 (n650, n468, n306, n204, n584);
and  g677 (n923, n320, n284, n324, n269);
or   g678 (n941, n300, n552, n569, n159);
xor  g679 (n1053, n582, n213, n336, n500);
nor  g680 (n1066, n591, n449, n519, n604);
nor  g681 (n925, n348, n283, n378, n449);
and  g682 (n997, n327, n483, n496, n401);
or   g683 (n752, n557, n349, n468, n535);
nand g684 (n976, n424, n256, n345, n261);
and  g685 (n940, n267, n280, n455, n510);
xnor g686 (n664, n433, n354, n502, n577);
xor  g687 (n776, n355, n333, n612, n286);
and  g688 (n893, n355, n381, n467, n527);
nand g689 (n950, n267, n260, n169, n539);
xnor g690 (n810, n174, n542, n453, n297);
and  g691 (n708, n377, n431, n290, n295);
or   g692 (n780, n208, n232, n436, n527);
and  g693 (n895, n508, n537, n433, n369);
nand g694 (n872, n488, n323, n184, n379);
nor  g695 (n660, n502, n533, n255, n189);
xor  g696 (n719, n526, n441, n574, n339);
or   g697 (n1017, n226, n387, n364, n334);
xor  g698 (n1064, n425, n593, n612, n401);
xor  g699 (n1023, n192, n383, n530, n565);
or   g700 (n735, n469, n410, n399, n475);
xnor g701 (n1012, n277, n380, n429, n341);
xnor g702 (n649, n561, n275, n478, n623);
or   g703 (n779, n274, n273, n611, n587);
xor  g704 (n1104, n569, n572, n556, n247);
or   g705 (n1098, n396, n325, n434, n215);
and  g706 (n789, n295, n227, n539, n222);
nor  g707 (n683, n313, n412, n245, n494);
nand g708 (n888, n163, n377, n455, n563);
and  g709 (n953, n209, n220, n460, n168);
nand g710 (n1111, n250, n254, n568, n541);
or   g711 (n722, n565, n563, n264, n609);
xor  g712 (n1086, n517, n501, n166, n562);
and  g713 (n927, n290, n211, n536, n466);
and  g714 (n829, n439, n271, n406, n548);
nand g715 (n729, n179, n603, n314, n449);
nor  g716 (n1085, n483, n579, n291, n395);
xor  g717 (n797, n229, n407, n194, n404);
and  g718 (n685, n287, n176, n620, n382);
nor  g719 (n876, n437, n252, n209, n481);
and  g720 (n818, n351, n440, n519, n578);
or   g721 (n1054, n315, n181, n485, n203);
or   g722 (n811, n261, n577, n532, n499);
nor  g723 (n955, n206, n456, n408, n212);
xnor g724 (n1024, n263, n507, n236, n605);
xor  g725 (n1071, n575, n479, n235, n319);
xor  g726 (n821, n197, n622, n453, n378);
xnor g727 (n1002, n389, n516, n587, n215);
nor  g728 (n743, n450, n218, n467, n422);
xnor g729 (n970, n525, n279, n376, n304);
nand g730 (n945, n251, n541, n445, n319);
xnor g731 (n741, n442, n511, n516, n360);
nor  g732 (n667, n445, n580, n492, n308);
nand g733 (n1035, n499, n397, n552, n350);
xor  g734 (n1025, n177, n235, n214, n614);
nor  g735 (n1088, n336, n447, n333, n305);
or   g736 (n725, n356, n446, n214, n318);
nor  g737 (n1089, n305, n208, n459, n440);
xnor g738 (n847, n186, n480, n368, n241);
or   g739 (n1056, n281, n599, n592, n374);
nor  g740 (n783, n331, n590, n620, n485);
and  g741 (n864, n162, n362, n603, n262);
and  g742 (n777, n436, n334, n229, n575);
and  g743 (n1058, n326, n381, n195, n366);
nor  g744 (n977, n584, n522, n480, n532);
nand g745 (n718, n301, n597, n433, n271);
xor  g746 (n644, n342, n603, n483, n329);
xor  g747 (n989, n514, n271, n242, n390);
nor  g748 (n912, n436, n495, n513, n198);
nor  g749 (n740, n339, n431, n396, n569);
xnor g750 (n988, n608, n475, n612, n404);
xnor g751 (n1018, n400, n356, n176, n601);
nand g752 (n790, n523, n296, n492, n191);
nor  g753 (n819, n320, n215, n188, n609);
xor  g754 (n848, n595, n590, n231, n423);
xor  g755 (n873, n213, n412, n544, n207);
nand g756 (n800, n479, n473, n345, n457);
xor  g757 (n984, n166, n313, n186, n341);
xnor g758 (n1026, n435, n411, n457, n461);
nor  g759 (n987, n463, n522, n370, n540);
or   g760 (n1080, n173, n562, n471, n574);
xor  g761 (n1059, n531, n206, n197, n568);
nor  g762 (n713, n466, n194, n258, n201);
xor  g763 (n763, n470, n281, n443, n271);
xnor g764 (n961, n533, n529, n213, n487);
nor  g765 (n1021, n190, n364, n201, n333);
and  g766 (n805, n190, n478, n523, n241);
nand g767 (n855, n454, n484, n273, n448);
nor  g768 (n714, n459, n596, n606, n234);
nor  g769 (n978, n551, n462, n506, n585);
xor  g770 (n896, n422, n373, n348, n534);
xnor g771 (n653, n219, n327, n440, n590);
xor  g772 (n1049, n599, n216, n353, n370);
and  g773 (n887, n232, n390, n385, n564);
nand g774 (n959, n445, n393, n171, n595);
nor  g775 (n646, n379, n518, n322, n287);
nor  g776 (n841, n387, n163, n467, n490);
and  g777 (n968, n186, n458, n323, n335);
and  g778 (n796, n430, n439, n570, n386);
xor  g779 (n993, n407, n504, n233, n415);
or   g780 (n632, n212, n282, n230, n302);
nand g781 (n774, n619, n546, n485, n347);
nand g782 (n830, n543, n285, n406, n435);
and  g783 (n652, n415, n437, n361, n458);
nand g784 (n964, n417, n518, n403, n180);
or   g785 (n756, n339, n270, n402, n365);
nor  g786 (n857, n521, n384, n509, n414);
xnor g787 (n837, n419, n572, n598, n329);
nand g788 (n629, n298, n308, n524, n456);
nand g789 (n702, n284, n324, n350, n406);
and  g790 (n911, n356, n312, n330, n570);
nor  g791 (n736, n346, n441, n179, n289);
and  g792 (n907, n463, n208, n379, n368);
and  g793 (n971, n251, n586, n541, n252);
nor  g794 (n1014, n484, n377, n223, n400);
and  g795 (n715, n338, n191, n257, n370);
xor  g796 (n894, n266, n374, n415, n220);
nand g797 (n630, n439, n266, n189, n325);
xnor g798 (n745, n600, n194, n386, n589);
nor  g799 (n669, n358, n346, n600, n528);
or   g800 (n1114, n295, n212, n588, n175);
and  g801 (n1091, n618, n538, n482, n255);
and  g802 (n996, n367, n559, n560, n575);
xnor g803 (n673, n411, n294, n358, n372);
xnor g804 (n831, n518, n172, n586, n314);
and  g805 (n1103, n274, n604, n399, n228);
and  g806 (n882, n418, n515, n182, n589);
xor  g807 (n1043, n539, n211, n525, n286);
nor  g808 (n645, n193, n432, n358, n312);
and  g809 (n771, n554, n393, n582, n326);
and  g810 (n738, n311, n412, n328, n387);
and  g811 (n778, n535, n477, n593, n253);
xnor g812 (n637, n337, n277, n353, n549);
xor  g813 (n982, n532, n497, n227, n407);
nor  g814 (n840, n324, n256, n436, n495);
xor  g815 (n1062, n510, n509, n474, n609);
nand g816 (n991, n248, n371, n264, n296);
or   g817 (n952, n403, n596, n163, n567);
xor  g818 (n850, n353, n593, n387, n614);
xor  g819 (n1004, n225, n604, n388, n459);
and  g820 (n692, n216, n240, n268, n429);
xor  g821 (n749, n243, n345, n361, n456);
xnor g822 (n875, n581, n451, n558, n321);
or   g823 (n901, n192, n420, n428, n294);
nand g824 (n874, n488, n164, n435, n623);
nand g825 (n681, n512, n489, n317, n591);
and  g826 (n948, n425, n465, n285, n349);
nor  g827 (n1087, n602, n360, n438, n611);
or   g828 (n747, n597, n410, n493, n173);
xnor g829 (n954, n239, n473, n570, n372);
or   g830 (n886, n239, n338, n224, n513);
and  g831 (n1001, n582, n304, n468, n594);
xnor g832 (n815, n618, n386, n474, n171);
nand g833 (n668, n509, n517, n272, n564);
or   g834 (n1038, n231, n533, n354, n167);
nand g835 (n983, n579, n583, n275, n617);
or   g836 (n1107, n617, n471, n571, n281);
nand g837 (n994, n380, n500, n171, n393);
xnor g838 (n1005, n464, n452, n189, n539);
nand g839 (n817, n359, n457, n555, n385);
xor  g840 (n1069, n586, n529, n350, n550);
nand g841 (n802, n594, n275, n389, n391);
and  g842 (n869, n417, n434, n228, n315);
nand g843 (n635, n246, n496, n434, n222);
or   g844 (n899, n481, n383, n405, n554);
nor  g845 (n750, n544, n476, n529, n223);
nor  g846 (n679, n609, n523, n310, n287);
xor  g847 (n917, n160, n260, n372, n583);
nor  g848 (n794, n579, n298, n499, n606);
xnor g849 (n792, n525, n453, n398, n385);
and  g850 (n1096, n278, n249, n414, n462);
and  g851 (n981, n359, n309, n251, n390);
nand g852 (n892, n180, n205, n159, n520);
xnor g853 (n671, n337, n232, n249, n193);
and  g854 (n1007, n394, n580, n288, n413);
nand g855 (n807, n351, n510, n452, n542);
nor  g856 (n728, n540, n475, n530, n318);
nand g857 (n935, n330, n369, n601);
nand g858 (n765, n190, n326, n607, n421);
xor  g859 (n845, n531, n203, n506, n312);
or   g860 (n710, n329, n182, n382, n313);
or   g861 (n1076, n243, n307, n560, n228);
nor  g862 (n1100, n430, n485, n331, n268);
or   g863 (n1028, n392, n215, n547, n167);
or   g864 (n682, n238, n308, n185, n302);
nor  g865 (n1084, n244, n484, n205, n494);
nor  g866 (n744, n208, n176, n242, n487);
nand g867 (n1083, n306, n399, n341, n554);
nand g868 (n926, n578, n216, n498, n379);
nor  g869 (n1063, n435, n569, n514, n490);
nand g870 (n773, n218, n202, n259, n319);
and  g871 (n654, n513, n391, n491, n199);
xor  g872 (n969, n368, n465, n505, n200);
and  g873 (n1033, n252, n438, n281, n564);
and  g874 (n868, n470, n481, n293, n427);
xor  g875 (n721, n250, n265, n278, n442);
nor  g876 (n827, n363, n274, n548, n245);
and  g877 (n1057, n592, n350, n391, n385);
nand g878 (n1082, n447, n542, n175, n236);
xor  g879 (n659, n161, n606, n217, n417);
or   g880 (n746, n253, n576, n343, n519);
or   g881 (n921, n608, n339, n254, n443);
xor  g882 (n764, n460, n524, n432, n303);
xor  g883 (n724, n594, n276, n402, n515);
xor  g884 (n897, n505, n553, n486, n472);
or   g885 (n769, n509, n384, n390, n618);
nor  g886 (n703, n501, n454, n232, n173);
xnor g887 (n742, n314, n617, n354, n341);
or   g888 (n787, n535, n446, n237, n346);
nand g889 (n627, n263, n200, n262, n174);
nor  g890 (n834, n159, n483, n285, n562);
and  g891 (n890, n380, n330, n363, n165);
xnor g892 (n998, n550, n535, n273, n170);
and  g893 (n674, n306, n322, n470, n371);
nor  g894 (n643, n479, n269, n231, n245);
nand g895 (n980, n301, n241, n418, n227);
nor  g896 (n825, n332, n570, n250, n321);
or   g897 (n906, n444, n621, n234, n258);
nand g898 (n666, n226, n411, n292, n280);
nor  g899 (n670, n343, n160, n510, n360);
and  g900 (n1093, n521, n201, n292, n353);
or   g901 (n844, n595, n451, n161, n455);
xnor g902 (n866, n237, n386, n225, n484);
nor  g903 (n803, n289, n374, n348, n573);
nor  g904 (n833, n219, n337, n288, n195);
xor  g905 (n861, n567, n301, n587, n508);
xnor g906 (n1070, n470, n448, n337, n307);
xor  g907 (n865, n584, n284, n552, n589);
and  g908 (n852, n294, n314, n467, n515);
nand g909 (n957, n331, n538, n585, n347);
xor  g910 (n1027, n531, n421, n514, n519);
or   g911 (n1067, n184, n482, n366, n486);
xnor g912 (n1010, n463, n174, n493, n607);
nand g913 (n1116, n517, n202, n438, n322);
xnor g914 (n1040, n439, n446, n381, n384);
or   g915 (n909, n580, n221, n352, n482);
xor  g916 (n863, n530, n581, n203, n458);
nand g917 (n946, n278, n400, n414, n310);
and  g918 (n720, n426, n410, n181, n594);
nor  g919 (n784, n621, n502, n237, n557);
xnor g920 (n920, n583, n600, n522, n319);
nor  g921 (n647, n425, n620, n419, n322);
xor  g922 (n891, n551, n489, n469, n471);
xnor g923 (n908, n619, n428, n534, n299);
nor  g924 (n816, n255, n589, n297, n618);
and  g925 (n1022, n536, n440, n597, n507);
nor  g926 (n902, n272, n293, n276, n375);
xnor g927 (n930, n450, n429, n352, n421);
nor  g928 (n823, n545, n590, n283, n280);
nor  g929 (n905, n374, n204, n409, n317);
xor  g930 (n697, n181, n224, n409, n265);
nand g931 (n759, n575, n617, n501, n574);
xnor g932 (n1051, n181, n561, n492, n196);
and  g933 (n1030, n355, n556, n455, n324);
or   g934 (n965, n333, n572, n516, n174);
xnor g935 (n1109, n237, n362, n612, n556);
or   g936 (n973, n345, n394, n447, n321);
or   g937 (n986, n325, n432, n416, n357);
nor  g938 (n862, n486, n359, n179, n476);
and  g939 (n690, n184, n545, n613, n230);
nor  g940 (n1075, n469, n236, n361, n163);
nand g941 (n966, n269, n551, n606, n286);
xnor g942 (n1077, n498, n520, n231, n560);
xnor g943 (n1047, n442, n206, n363, n615);
or   g944 (n962, n234, n178, n295, n524);
and  g945 (n1032, n182, n316, n369, n392);
nor  g946 (n634, n357, n234, n516, n607);
nor  g947 (n932, n263, n567, n394, n226);
xor  g948 (n1094, n481, n224, n448, n183);
and  g949 (n910, n450, n253, n506, n211);
and  g950 (n1106, n543, n466, n266, n265);
and  g951 (n859, n193, n169, n464, n392);
xor  g952 (n884, n430, n414, n473, n327);
or   g953 (n937, n461, n284, n200, n178);
and  g954 (n1000, n409, n161, n199, n419);
nand g955 (n1034, n614, n404, n564, n297);
nand g956 (n1074, n602, n290, n498, n328);
xor  g957 (n995, n316, n203, n230, n541);
xor  g958 (n795, n423, n177, n217, n615);
xnor g959 (n838, n238, n395, n402, n286);
and  g960 (n661, n176, n581, n260, n487);
and  g961 (n639, n476, n165, n172, n598);
nand g962 (n782, n288, n542, n558, n545);
or   g963 (n655, n282, n444, n366, n310);
nor  g964 (n943, n242, n219, n402, n301);
or   g965 (n951, n173, n600, n318, n244);
or   g966 (n836, n357, n422, n240, n159);
nor  g967 (n642, n601, n240, n466, n511);
nand g968 (n640, n303, n247, n428, n511);
nor  g969 (n676, n423, n251, n346, n548);
or   g970 (n806, n543, n620, n192, n413);
xnor g971 (n758, n315, n427, n197, n451);
nand g972 (n1036, n573, n480, n187, n596);
xnor g973 (n860, n383, n193, n408, n260);
nand g974 (n1019, n614, n446, n447, n478);
xor  g975 (n933, n323, n429, n464, n164);
xor  g976 (n913, n491, n160, n405, n501);
or   g977 (n1113, n209, n220, n425, n256);
xor  g978 (n754, n243, n497, n494, n426);
nor  g979 (n691, n261, n189, n526, n299);
or   g980 (n1055, n370, n471, n397, n309);
nor  g981 (n1073, n450, n362, n468, n526);
nor  g982 (n1081, n394, n209, n180, n168);
xnor g983 (n696, n475, n375, n472, n161);
or   g984 (n922, n582, n321, n431, n413);
nand g985 (n733, n547, n428, n240, n512);
nand g986 (n781, n486, n320, n291, n449);
nand g987 (n704, n530, n257, n525, n307);
xor  g988 (n706, n427, n380, n272, n300);
nor  g989 (n766, n557, n499, n491, n373);
nand g990 (n835, n565, n315, n571, n196);
nand g991 (n820, n587, n419, n317, n187);
xor  g992 (n931, n312, n167, n221);
nand g993 (n1108, n343, n200, n316, n406);
nand g994 (n832, n469, n565, n611, n170);
and  g995 (n732, n579, n309, n230, n443);
nor  g996 (n730, n242, n246, n593, n171);
and  g997 (n694, n233, n508, n363, n210);
xor  g998 (n701, n566, n360, n543, n537);
xnor g999 (n949, n257, n265, n392, n546);
nand g1000 (n801, n524, n241, n490, n496);
nand g1001 (n1029, n389, n610, n202, n401);
xnor g1002 (n979, n400, n311, n205, n538);
or   g1003 (n1102, n338, n605, n462, n536);
or   g1004 (n700, n367, n214, n457, n247);
xnor g1005 (n898, n228, n577, n225, n325);
nor  g1006 (n972, n572, n426, n555, n396);
nand g1007 (n739, n595, n598, n267, n498);
or   g1008 (n1112, n191, n323, n183, n162);
nor  g1009 (n1068, n262, n505, n290, n233);
xor  g1010 (n903, n566, n299, n219, n317);
nor  g1011 (n858, n477, n597, n424, n336);
or   g1012 (n942, n177, n395, n167, n188);
xor  g1013 (n799, n497, n330, n175, n331);
nand g1014 (n1079, n573, n554, n164, n500);
or   g1015 (n1009, n514, n246, n529, n186);
nand g1016 (n1101, n505, n347, n292, n248);
nor  g1017 (n885, n357, n571, n568, n292);
and  g1018 (n1115, n420, n187, n388, n303);
nor  g1019 (n928, n351, n393, n352, n239);
nand g1020 (n809, n528, n216, n444, n581);
or   g1021 (n1011, n214, n198, n610, n207);
or   g1022 (n1046, n285, n580, n395, n576);
and  g1023 (n1016, n459, n218, n549, n252);
xnor g1024 (n641, n254, n184, n507, n377);
or   g1025 (n878, n382, n259, n601, n254);
nand g1026 (n1099, n531, n172, n194, n364);
or   g1027 (n867, n528, n464, n343, n536);
or   g1028 (n651, n288, n613, n441, n412);
xnor g1029 (n657, n417, n217, n355, n563);
nand g1030 (n788, n615, n433, n563, n375);
nor  g1031 (n768, n320, n222, n249, n221);
nand g1032 (n1015, n235, n348, n212, n562);
and  g1033 (n813, n452, n500, n185, n309);
nand g1034 (n918, n523, n326, n371, n493);
nand g1035 (n974, n210, n559, n165, n367);
xnor g1036 (n658, n222, n277, n534, n276);
xnor g1037 (n963, n368, n296, n279, n293);
and  g1038 (n1041, n407, n465, n521, n578);
xnor g1039 (n672, n418, n376, n168, n561);
nor  g1040 (n748, n165, n462, n622, n559);
and  g1041 (n880, n507, n302, n282, n275);
nor  g1042 (n843, n378, n477, n183, n313);
and  g1043 (n915, n299, n279, n306, n512);
xor  g1044 (n924, n338, n568, n537, n316);
xnor g1045 (n1045, n239, n340, n576, n424);
nor  g1046 (n760, n602, n259, n160, n444);
nand g1047 (n633, n559, n307, n302, n478);
xor  g1048 (n1065, n613, n411, n334, n461);
or   g1049 (n1013, n408, n296, n504, n546);
or   g1050 (n934, n405, n347, n622, n283);
xnor g1051 (n1117, n247, n332, n267, n426);
xor  g1052 (n767, n332, n403, n258, n487);
xnor g1053 (n755, n354, n416, n365, n335);
xnor g1054 (n675, n504, n170, n495, n311);
xor  g1055 (n990, n373, n227, n434, n540);
nand g1056 (n1092, n561, n566, n352, n276);
and  g1057 (n975, n495, n300, n164, n249);
nor  g1058 (n828, n605, n397, n259, n293);
nor  g1059 (n648, n297, n422, n207, n238);
or   g1060 (n688, n344, n304, n477, n298);
xor  g1061 (n826, n270, n282, n615, n598);
xor  g1062 (n798, n578, n342, n465, n553);
nand g1063 (n842, n396, n566, n616, n604);
nand g1064 (n1061, n199, n223, n493, n258);
xnor g1065 (n793, n384, n244, n192, n515);
nor  g1066 (n871, n201, n404, n480, n359);
nor  g1067 (n985, n210, n280, n361, n553);
nand g1068 (n1037, n489, n613, n238, n451);
and  g1069 (n709, n454, n373, n596, n264);
and  g1070 (n999, n520, n410, n574, n479);
xor  g1071 (n1006, n476, n458, n408, n202);
nand g1072 (n936, n490, n213, n256, n351);
xnor g1073 (n687, n291, n403, n217, n592);
or   g1074 (n770, n544, n255, n420, n191);
nand g1075 (n883, n548, n527, n356, n178);
nand g1076 (n1060, n461, n195, n437, n472);
xor  g1077 (n686, n599, n257, n532, n376);
nand g1078 (n698, n489, n474, n528, n463);
or   g1079 (n939, n474, n611, n362, n518);
xnor g1080 (n712, n560, n616, n549, n503);
and  g1081 (n757, n268, n517, n588, n399);
xnor g1082 (n678, n492, n225, n211, n197);
xnor g1083 (n1097, n268, n188, n584, n491);
xor  g1084 (n916, n376, n253, n608, n166);
buf  g1085 (n1118, n653);
not  g1086 (n1139, n632);
buf  g1087 (n1122, n645);
buf  g1088 (n1135, n634);
not  g1089 (n1136, n640);
not  g1090 (n1137, n637);
not  g1091 (n1119, n638);
buf  g1092 (n1121, n636);
not  g1093 (n1134, n626);
not  g1094 (n1120, n641);
not  g1095 (n1133, n643);
buf  g1096 (n1124, n642);
buf  g1097 (n1129, n630);
buf  g1098 (n1130, n649);
buf  g1099 (n1123, n646);
buf  g1100 (n1125, n644);
buf  g1101 (n1126, n635);
buf  g1102 (n1138, n627);
buf  g1103 (n1128, n631);
not  g1104 (n1131, n628);
xor  g1105 (n1132, n639, n633, n650, n651);
and  g1106 (n1127, n629, n648, n647, n652);
and  g1107 (n1146, n1126, n677, n663, n685);
nor  g1108 (n1142, n687, n674, n655, n689);
xor  g1109 (n1140, n675, n688, n1122, n670);
xor  g1110 (n1151, n656, n658, n662, n676);
xor  g1111 (n1143, n668, n681, n683, n684);
xor  g1112 (n1147, n669, n686, n664, n1125);
or   g1113 (n1149, n667, n1127, n654, n673);
nand g1114 (n1150, n665, n682, n661, n1120);
xor  g1115 (n1144, n671, n657, n1121, n1124);
xnor g1116 (n1148, n1123, n659, n1119, n660);
xnor g1117 (n1145, n1118, n680, n678, n679);
and  g1118 (n1141, n1128, n1129, n672, n666);
not  g1119 (n1152, n1144);
buf  g1120 (n1161, n1145);
buf  g1121 (n1154, n1146);
buf  g1122 (n1155, n1147);
buf  g1123 (n1156, n1149);
not  g1124 (n1153, n1142);
buf  g1125 (n1159, n1148);
buf  g1126 (n1158, n1150);
buf  g1127 (n1157, n1143);
buf  g1128 (n1160, n1151);
buf  g1129 (n1162, n1161);
buf  g1130 (n1163, n153);
nand g1131 (n1169, n150, n151);
xnor g1132 (n1167, n1158, n149, n1160, n150);
or   g1133 (n1168, n1155, n150, n153, n154);
xnor g1134 (n1170, n1159, n153, n152, n1157);
and  g1135 (n1166, n152, n152, n154, n151);
xor  g1136 (n1171, n1152, n153, n154);
nor  g1137 (n1165, n150, n151, n1153);
or   g1138 (n1164, n1154, n155, n1156, n152);
buf  g1139 (n1172, n1165);
buf  g1140 (n1190, n1165);
not  g1141 (n1179, n1162);
not  g1142 (n1176, n1166);
buf  g1143 (n1185, n1165);
buf  g1144 (n1188, n1166);
not  g1145 (n1186, n1163);
not  g1146 (n1182, n1162);
not  g1147 (n1189, n1164);
buf  g1148 (n1184, n1165);
not  g1149 (n1174, n1166);
buf  g1150 (n1187, n1162);
buf  g1151 (n1191, n1163);
not  g1152 (n1173, n1163);
not  g1153 (n1178, n1164);
buf  g1154 (n1175, n1166);
not  g1155 (n1177, n1162);
not  g1156 (n1180, n1164);
buf  g1157 (n1181, n1163);
not  g1158 (n1183, n1164);
not  g1159 (n1197, n701);
xor  g1160 (n1194, n699, n703, n1172);
xor  g1161 (n1198, n694, n690, n706, n1173);
xor  g1162 (n1196, n693, n700, n697, n1173);
xnor g1163 (n1195, n705, n698, n702, n695);
or   g1164 (n1192, n1173, n1172, n696);
xor  g1165 (n1193, n704, n691, n692, n1172);
not  g1166 (n1201, n1196);
not  g1167 (n1207, n1183);
nor  g1168 (n1199, n1183, n1187);
xnor g1169 (n1226, n709, n715, n1175, n1181);
xnor g1170 (n1200, n1176, n1192, n1186);
and  g1171 (n1224, n708, n1198, n1184, n1179);
nand g1172 (n1204, n1194, n713, n1182, n1181);
xnor g1173 (n1221, n1178, n1185, n1197, n1194);
nor  g1174 (n1217, n721, n1195, n1178, n1192);
xnor g1175 (n1208, n1186, n720, n1184, n1180);
nand g1176 (n1223, n1178, n1196, n1197, n1187);
xor  g1177 (n1203, n1177, n1179, n1176);
xnor g1178 (n1211, n1195, n1174, n724, n1193);
xor  g1179 (n1214, n1177, n714, n1194, n1193);
xnor g1180 (n1225, n1181, n1198, n1173, n1187);
xnor g1181 (n1218, n710, n1174, n1178, n711);
and  g1182 (n1220, n1196, n624, n722, n718);
nand g1183 (n1216, n712, n1184, n1177, n1174);
nor  g1184 (n1209, n1182, n1198, n1183, n1186);
and  g1185 (n1210, n1184, n1183, n1180, n719);
nor  g1186 (n1202, n1174, n1175, n1195, n717);
nand g1187 (n1205, n1177, n707, n1175, n1193);
or   g1188 (n1222, n1179, n1176, n1182, n1197);
xor  g1189 (n1215, n1181, n1195, n1194, n1196);
xor  g1190 (n1206, n1193, n1192, n1179, n1198);
and  g1191 (n1213, n1180, n1186, n1182, n1185);
nor  g1192 (n1212, n1180, n1185, n1175);
and  g1193 (n1219, n716, n1187, n1197, n723);
xnor g1194 (n1230, n728, n1207, n1203);
nand g1195 (n1227, n1207, n1199);
xnor g1196 (n1234, n1200, n729, n1208, n1204);
xor  g1197 (n1229, n624, n1208, n1205, n725);
xnor g1198 (n1232, n1205, n1202, n1201);
or   g1199 (n1231, n1203, n1207, n1202);
nand g1200 (n1235, n730, n1200, n1204);
nand g1201 (n1236, n1206, n1200, n1205, n1204);
xnor g1202 (n1237, n727, n1201, n1206, n1200);
xnor g1203 (n1228, n1206, n1208, n1201, n1203);
xnor g1204 (n1233, n1201, n1208, n1205, n1199);
nor  g1205 (n1238, n726, n1207, n1203, n1206);
buf  g1206 (n1241, n1236);
not  g1207 (n1243, n1238);
not  g1208 (n1242, n1237);
not  g1209 (n1246, n1232);
buf  g1210 (n1244, n1231);
buf  g1211 (n1240, n1233);
buf  g1212 (n1245, n1234);
buf  g1213 (n1239, n1235);
not  g1214 (n1248, n1246);
buf  g1215 (n1272, n1210);
not  g1216 (n1271, n1132);
nand g1217 (n1269, n156, n1240, n1168);
and  g1218 (n1262, n1167, n1240, n1188, n1190);
or   g1219 (n1252, n624, n1167, n1168, n158);
xnor g1220 (n1267, n625, n1167, n1239, n1189);
or   g1221 (n1261, n1245, n1211, n731, n156);
or   g1222 (n1256, n1241, n1243, n733);
and  g1223 (n1255, n1167, n1246, n157, n1209);
nor  g1224 (n1270, n158, n1171, n735, n155);
xnor g1225 (n1274, n1191, n1243, n155, n1170);
nor  g1226 (n1265, n1133, n155, n1188);
or   g1227 (n1278, n1137, n1130, n736, n1242);
xor  g1228 (n1263, n1239, n1242, n1246, n1171);
or   g1229 (n1275, n1188, n1239, n1245, n1131);
nand g1230 (n1247, n1212, n158, n1191, n624);
nor  g1231 (n1266, n1209, n1134, n1211, n1245);
xor  g1232 (n1253, n1243, n1240, n1171);
nand g1233 (n1276, n1136, n157, n156, n1240);
and  g1234 (n1250, n1242, n1190, n1245, n1210);
and  g1235 (n1254, n1169, n1244, n158);
xnor g1236 (n1264, n1191, n1244, n1170, n732);
or   g1237 (n1257, n1246, n1189, n1211, n157);
xor  g1238 (n1273, n625, n1139, n1189, n1239);
nor  g1239 (n1249, n156, n1169, n1168, n32);
and  g1240 (n1277, n1168, n1210, n1169, n1244);
xnor g1241 (n1268, n1190, n1210, n1242, n1241);
xor  g1242 (n1251, n1191, n734, n1135, n1170);
nor  g1243 (n1259, n1241, n1189, n1190, n1209);
nand g1244 (n1258, n1209, n32, n157, n1170);
nand g1245 (n1260, n1211, n1169, n1138, n1241);
not  g1246 (n1290, n1267);
not  g1247 (n1331, n1250);
not  g1248 (n1285, n1272);
buf  g1249 (n1307, n1261);
buf  g1250 (n1313, n1254);
buf  g1251 (n1324, n1257);
buf  g1252 (n1311, n1264);
not  g1253 (n1299, n1266);
not  g1254 (n1302, n1254);
buf  g1255 (n1297, n1250);
not  g1256 (n1287, n1268);
buf  g1257 (n1280, n1264);
buf  g1258 (n1295, n1276);
buf  g1259 (n1294, n1257);
buf  g1260 (n1337, n1248);
not  g1261 (n1322, n1249);
buf  g1262 (n1305, n1255);
not  g1263 (n1286, n1257);
buf  g1264 (n1328, n1262);
buf  g1265 (n1304, n1252);
not  g1266 (n1283, n1264);
not  g1267 (n1296, n1271);
not  g1268 (n1323, n1270);
not  g1269 (n1293, n1254);
not  g1270 (n1303, n1274);
not  g1271 (n1308, n1275);
not  g1272 (n1316, n1265);
buf  g1273 (n1281, n1263);
buf  g1274 (n1292, n1275);
not  g1275 (n1318, n1260);
not  g1276 (n1335, n1256);
buf  g1277 (n1330, n1255);
buf  g1278 (n1301, n1269);
buf  g1279 (n1310, n1266);
buf  g1280 (n1312, n1266);
buf  g1281 (n1319, n1255);
buf  g1282 (n1317, n1271);
buf  g1283 (n1325, n1248);
not  g1284 (n1288, n1265);
buf  g1285 (n1298, n1261);
nor  g1286 (n1291, n1273, n1249);
and  g1287 (n1289, n1251, n1273, n1259, n1268);
nand g1288 (n1333, n1259, n1254, n1260, n1276);
xnor g1289 (n1300, n1275, n1256, n1271, n1273);
xor  g1290 (n1338, n1253, n1274, n1249);
nand g1291 (n1279, n1258, n1251, n1267);
nor  g1292 (n1306, n1273, n1252, n1248, n1268);
nand g1293 (n1320, n1258, n1249, n1272, n1264);
or   g1294 (n1315, n1270, n1272, n1271, n1276);
xnor g1295 (n1326, n1260, n1263, n1269, n1268);
xnor g1296 (n1309, n1263, n1275, n1269, n1276);
xor  g1297 (n1327, n1266, n1259, n1247);
nor  g1298 (n1332, n1255, n1256, n1260, n1270);
xor  g1299 (n1334, n1261, n1263, n1257, n1250);
xnor g1300 (n1329, n1250, n1252, n1274, n1267);
xor  g1301 (n1336, n1247, n1258, n1269, n1253);
xnor g1302 (n1321, n1262, n1258, n1267, n1253);
xor  g1303 (n1282, n1272, n1270, n1253, n1261);
nor  g1304 (n1284, n1262, n1251, n1252, n1265);
xnor g1305 (n1314, n1248, n1265, n1256, n1262);
not  g1306 (n1340, n1283);
not  g1307 (n1344, n1282);
not  g1308 (n1345, n1280);
not  g1309 (n1341, n1281);
not  g1310 (n1346, n1279);
buf  g1311 (n1342, n1286);
buf  g1312 (n1339, n1285);
not  g1313 (n1343, n1284);
nor  g1314 (n1348, n1301, n1222, n1317, n1214);
nor  g1315 (n1364, n1312, n1339, n1217);
nand g1316 (n1369, n1298, n1345, n1213, n1222);
and  g1317 (n1347, n1340, n1316, n1223, n1341);
and  g1318 (n1371, n1220, n1218, n1339, n1342);
nand g1319 (n1353, n1216, n1217, n1221, n1293);
and  g1320 (n1370, n1302, n1294, n1341, n1310);
nor  g1321 (n1373, n1311, n1223, n1304, n1342);
and  g1322 (n1362, n737, n1346, n1289);
nor  g1323 (n1354, n1346, n1218, n1213, n1219);
nand g1324 (n1360, n1215, n1339, n1224, n1212);
xnor g1325 (n1358, n1215, n1300, n1313, n1344);
xor  g1326 (n1363, n1345, n1218, n1215, n1290);
xnor g1327 (n1352, n1222, n1340, n1212, n1305);
xnor g1328 (n1359, n1218, n1217, n1345, n1340);
and  g1329 (n1365, n1221, n1216, n1303, n1344);
xnor g1330 (n1349, n1343, n1220, n1314, n1307);
or   g1331 (n1361, n1295, n1296, n1344, n1342);
xor  g1332 (n1350, n1288, n1221, n1224, n1341);
and  g1333 (n1356, n1213, n1343, n1219);
and  g1334 (n1368, n1287, n1220, n1343, n1346);
nand g1335 (n1357, n1212, n1216, n1308, n1222);
and  g1336 (n1351, n1309, n1292, n1219, n1297);
and  g1337 (n1372, n1214, n1214, n1299, n1306);
nor  g1338 (n1367, n1344, n1223, n1213);
nor  g1339 (n1355, n1214, n1215, n1216, n1221);
or   g1340 (n1366, n1345, n1315, n1291, n1220);
buf  g1341 (n1376, n1358);
nand g1342 (n1378, n1348, n1349, n1357);
nand g1343 (n1375, n1354, n1353, n1355, n1362);
nor  g1344 (n1377, n1347, n1351, n1361, n1352);
xor  g1345 (n1374, n1356, n1350, n1359, n1360);
and  g1346 (n1380, n1365, n1364, n1363, n738);
nand g1347 (n1379, n1375, n1366, n1374, n739);
buf  g1348 (n1382, n740);
buf  g1349 (n1383, n1379);
and  g1350 (n1381, n1379, n1380, n742, n741);
buf  g1351 (n1386, n1382);
not  g1352 (n1387, n746);
or   g1353 (n1385, n743, n1381, n1383, n745);
xnor g1354 (n1384, n748, n1383, n747, n744);
buf  g1355 (n1389, n1384);
buf  g1356 (n1390, n1387);
not  g1357 (n1394, n1386);
not  g1358 (n1392, n749);
not  g1359 (n1388, n1387);
not  g1360 (n1393, n1385);
or   g1361 (n1391, n1386, n1385);
not  g1362 (n1399, n758);
not  g1363 (n1405, n1392);
not  g1364 (n1398, n761);
buf  g1365 (n1401, n1390);
buf  g1366 (n1395, n1389);
not  g1367 (n1400, n757);
not  g1368 (n1403, n756);
not  g1369 (n1409, n1391);
buf  g1370 (n1397, n1391);
buf  g1371 (n1404, n754);
nor  g1372 (n1402, n1388, n1392, n1391);
and  g1373 (n1406, n763, n1390, n1392, n755);
nand g1374 (n1396, n751, n760, n1389, n753);
nor  g1375 (n1407, n764, n1390, n1391, n762);
or   g1376 (n1408, n750, n752, n759, n1388);
not  g1377 (n1437, n1398);
buf  g1378 (n1415, n1397);
not  g1379 (n1433, n1396);
buf  g1380 (n1422, n1395);
not  g1381 (n1427, n1401);
buf  g1382 (n1426, n1400);
not  g1383 (n1423, n1401);
not  g1384 (n1428, n1395);
buf  g1385 (n1432, n1401);
not  g1386 (n1425, n1400);
buf  g1387 (n1416, n1399);
buf  g1388 (n1436, n1396);
not  g1389 (n1417, n1397);
not  g1390 (n1430, n1397);
buf  g1391 (n1424, n1401);
buf  g1392 (n1414, n1395);
not  g1393 (n1434, n1398);
buf  g1394 (n1421, n1399);
not  g1395 (n1410, n1400);
buf  g1396 (n1419, n1398);
not  g1397 (n1435, n1396);
buf  g1398 (n1431, n1397);
not  g1399 (n1418, n1396);
not  g1400 (n1429, n1399);
not  g1401 (n1413, n1399);
buf  g1402 (n1420, n1400);
not  g1403 (n1411, n1395);
buf  g1404 (n1412, n1398);
nand g1405 (n1480, n932, n1020, n882, n888);
nor  g1406 (n1473, n1046, n1412, n1018, n1437);
xor  g1407 (n1467, n956, n1058, n839, n902);
and  g1408 (n1488, n906, n987, n785, n977);
nand g1409 (n1451, n1007, n1099, n815, n789);
nand g1410 (n1527, n983, n1431, n865, n1012);
and  g1411 (n1541, n939, n1072, n1040, n823);
nand g1412 (n1539, n825, n836, n1426, n961);
xnor g1413 (n1511, n842, n801, n1014, n1090);
nor  g1414 (n1535, n1085, n872, n811, n997);
nor  g1415 (n1509, n1424, n1418, n1435);
nand g1416 (n1470, n926, n879, n1414, n876);
xor  g1417 (n1452, n1415, n1434, n978);
nor  g1418 (n1510, n1414, n1041, n870, n1079);
xnor g1419 (n1514, n1436, n949, n974, n1083);
nand g1420 (n1482, n1019, n930, n883, n810);
xor  g1421 (n1528, n1412, n1427, n994, n792);
xor  g1422 (n1462, n807, n847, n1418, n1092);
nand g1423 (n1502, n1021, n1037, n1425, n775);
and  g1424 (n1495, n862, n942, n915, n958);
nor  g1425 (n1524, n1000, n765, n1057, n880);
or   g1426 (n1474, n890, n1434, n934, n768);
nor  g1427 (n1464, n874, n984, n885, n875);
nand g1428 (n1477, n821, n777, n1002, n1437);
or   g1429 (n1441, n793, n1028, n1420, n944);
or   g1430 (n1494, n820, n848, n922, n979);
xor  g1431 (n1515, n1042, n972, n1424, n791);
nand g1432 (n1486, n854, n1418, n1009, n867);
or   g1433 (n1442, n1004, n771, n1036, n925);
nand g1434 (n1504, n931, n914, n849, n877);
xor  g1435 (n1461, n892, n1027, n1017, n1421);
xnor g1436 (n1481, n953, n1088, n1414, n1074);
and  g1437 (n1538, n951, n917, n1076, n803);
xor  g1438 (n1542, n866, n918, n1034, n1432);
and  g1439 (n1438, n1437, n941, n1432, n1429);
and  g1440 (n1508, n857, n1431, n995, n779);
xnor g1441 (n1526, n959, n1428, n1100, n829);
xor  g1442 (n1478, n774, n843, n860, n967);
xor  g1443 (n1453, n816, n1084, n884, n905);
and  g1444 (n1479, n921, n1424, n1087, n895);
xor  g1445 (n1498, n993, n1436, n878, n1421);
nor  g1446 (n1497, n1430, n1081, n1078, n1416);
nand g1447 (n1484, n991, n809, n1051, n955);
and  g1448 (n1448, n936, n827, n858, n1026);
or   g1449 (n1546, n1431, n973, n800, n844);
and  g1450 (n1457, n996, n896, n1420, n1410);
nor  g1451 (n1499, n1435, n1097, n1047, n963);
nor  g1452 (n1447, n1048, n1412, n1064, n1428);
nor  g1453 (n1444, n773, n1035, n1421, n1032);
or   g1454 (n1503, n784, n841, n1417, n835);
and  g1455 (n1476, n869, n1414, n1432, n971);
xor  g1456 (n1449, n935, n975, n1422, n903);
xnor g1457 (n1483, n1098, n999, n986, n873);
xor  g1458 (n1501, n889, n990, n893, n1433);
nand g1459 (n1459, n1411, n1003, n1082, n1077);
nor  g1460 (n1458, n1436, n1413, n798, n913);
xnor g1461 (n1492, n769, n1420, n1433, n1428);
or   g1462 (n1540, n1006, n928, n1435, n1030);
nor  g1463 (n1516, n813, n1023, n1015, n1418);
xnor g1464 (n1471, n1029, n945, n891, n916);
nor  g1465 (n1530, n933, n794, n1417, n1430);
xnor g1466 (n1521, n969, n907, n1049, n1086);
xor  g1467 (n1450, n859, n1423, n992, n776);
or   g1468 (n1446, n846, n797, n1080, n899);
nor  g1469 (n1465, n1411, n834, n1415, n1063);
or   g1470 (n1490, n911, n1005, n1070, n833);
or   g1471 (n1544, n795, n871, n1054, n950);
or   g1472 (n1512, n988, n1053, n802, n1416);
nor  g1473 (n1455, n861, n1425, n1428, n1431);
nor  g1474 (n1520, n923, n1096, n910, n1427);
xnor g1475 (n1456, n1071, n1038, n929, n863);
xor  g1476 (n1445, n1067, n1425, n1089, n1437);
nor  g1477 (n1547, n1062, n780, n1069, n805);
xnor g1478 (n1519, n799, n817, n957, n1429);
and  g1479 (n1463, n822, n1415, n919, n852);
and  g1480 (n1534, n864, n1420, n1422, n788);
nand g1481 (n1533, n1043, n1419, n1093, n868);
xnor g1482 (n1472, n920, n840, n981, n818);
or   g1483 (n1440, n898, n960, n786, n1091);
and  g1484 (n1525, n787, n1065, n1410, n908);
and  g1485 (n1475, n900, n1426, n909, n946);
xor  g1486 (n1529, n830, n964, n772, n1056);
nor  g1487 (n1468, n804, n943, n832, n770);
nor  g1488 (n1439, n1022, n998, n924, n1044);
nor  g1489 (n1505, n1024, n1001, n1424, n778);
or   g1490 (n1548, n952, n968, n940, n1413);
or   g1491 (n1487, n856, n1066, n1033, n1025);
xnor g1492 (n1523, n966, n1059, n1417, n1421);
xor  g1493 (n1536, n947, n1423, n783, n1095);
or   g1494 (n1469, n912, n1422, n1075, n855);
nor  g1495 (n1489, n819, n1419, n850, n1427);
nand g1496 (n1466, n904, n814, n894, n901);
xor  g1497 (n1549, n1426, n1413, n985, n1417);
xor  g1498 (n1537, n1425, n1423, n782, n927);
xor  g1499 (n1543, n1011, n948, n980, n806);
xor  g1500 (n1513, n1432, n790, n1008, n1412);
xor  g1501 (n1496, n1427, n1416, n1039, n1410);
xnor g1502 (n1531, n1434, n1430, n1422, n1031);
and  g1503 (n1507, n826, n808, n1050, n1413);
and  g1504 (n1493, n1433, n881, n965, n1423);
nand g1505 (n1517, n1429, n976, n1055, n796);
nand g1506 (n1545, n1411, n1013, n1052, n1016);
nor  g1507 (n1506, n831, n812, n1433, n853);
xor  g1508 (n1491, n1429, n824, n1436, n1045);
xor  g1509 (n1485, n970, n1010, n851, n767);
xnor g1510 (n1518, n954, n1419, n766, n989);
xnor g1511 (n1532, n1073, n1419, n1061, n1430);
xor  g1512 (n1454, n1094, n982, n1415, n897);
or   g1513 (n1500, n838, n1410, n887, n781);
nand g1514 (n1460, n1068, n837, n828, n938);
xnor g1515 (n1443, n937, n962, n1060, n1426);
nor  g1516 (n1522, n886, n1416, n1411, n845);
buf  g1517 (n1560, n1447);
not  g1518 (n1571, n1444);
buf  g1519 (n1585, n1448);
not  g1520 (n1555, n1440);
buf  g1521 (n1554, n1439);
not  g1522 (n1570, n1441);
not  g1523 (n1573, n1442);
buf  g1524 (n1578, n1444);
buf  g1525 (n1584, n1442);
not  g1526 (n1566, n1443);
not  g1527 (n1579, n1445);
not  g1528 (n1583, n1446);
not  g1529 (n1574, n1448);
buf  g1530 (n1567, n1446);
not  g1531 (n1568, n1449);
buf  g1532 (n1557, n1438);
buf  g1533 (n1576, n1447);
buf  g1534 (n1572, n1444);
not  g1535 (n1550, n1440);
buf  g1536 (n1582, n1449);
buf  g1537 (n1580, n1446);
not  g1538 (n1553, n1439);
not  g1539 (n1561, n1442);
buf  g1540 (n1551, n1448);
not  g1541 (n1564, n1447);
not  g1542 (n1563, n1438);
buf  g1543 (n1552, n1439);
not  g1544 (n1559, n1441);
buf  g1545 (n1575, n1449);
buf  g1546 (n1581, n1440);
buf  g1547 (n1556, n1445);
not  g1548 (n1569, n1443);
not  g1549 (n1558, n1441);
buf  g1550 (n1565, n1438);
not  g1551 (n1562, n1443);
buf  g1552 (n1577, n1445);
buf  g1553 (n1696, n1498);
not  g1554 (n1624, n1497);
buf  g1555 (n1622, n1478);
buf  g1556 (n1658, n1517);
not  g1557 (n1685, n1493);
not  g1558 (n1729, n1452);
buf  g1559 (n1633, n1581);
not  g1560 (n1641, n1538);
buf  g1561 (n1712, n1527);
buf  g1562 (n1589, n1498);
buf  g1563 (n1605, n1532);
buf  g1564 (n1596, n1511);
not  g1565 (n1705, n1534);
buf  g1566 (n1695, n1547);
buf  g1567 (n1599, n1524);
not  g1568 (n1647, n1523);
not  g1569 (n1688, n1503);
not  g1570 (n1704, n1554);
nand g1571 (n1694, n1578, n1484, n1523, n1566);
nor  g1572 (n1699, n1527, n1466, n1529, n1482);
xnor g1573 (n1675, n1473, n1473, n1451, n1547);
and  g1574 (n1621, n1487, n1526, n1559, n1468);
or   g1575 (n1648, n1460, n1565, n1551, n1530);
or   g1576 (n1714, n1495, n1489, n1473, n1377);
xnor g1577 (n1623, n1465, n1487, n1574, n1585);
and  g1578 (n1607, n1524, n1452, n1458, n1499);
nand g1579 (n1681, n1461, n1548, n1552, n1484);
and  g1580 (n1635, n1474, n1557, n1525, n1545);
or   g1581 (n1703, n1544, n1481, n1525, n1535);
xnor g1582 (n1593, n1553, n1501, n1570, n1511);
and  g1583 (n1654, n1539, n1462, n1512, n1576);
xnor g1584 (n1717, n1505, n1554, n1490, n1504);
nand g1585 (n1668, n1577, n1491, n1557, n1506);
nand g1586 (n1682, n1555, n1551, n1487, n1572);
nand g1587 (n1592, n1516, n1517, n1485, n1499);
or   g1588 (n1728, n1554, n1520, n1570, n1538);
nand g1589 (n1630, n1581, n1581, n1573, n1541);
nand g1590 (n1700, n1481, n1486, n1509, n1531);
xnor g1591 (n1595, n1573, n1562, n1533, n1510);
or   g1592 (n1697, n1513, n1581, n1527, n1532);
nor  g1593 (n1662, n1463, n1492, n1535, n1458);
xor  g1594 (n1660, n1512, n1553, n1461, n1508);
xnor g1595 (n1659, n1567, n1478, n1585, n1540);
and  g1596 (n1598, n1485, n1490, n1504, n1543);
nor  g1597 (n1614, n1552, n1503, n1561, n1516);
or   g1598 (n1590, n1543, n1507, n1550, n1573);
xor  g1599 (n1676, n1508, n1471, n1495, n1557);
or   g1600 (n1613, n1460, n1521, n1450, n1545);
xor  g1601 (n1646, n1583, n1510, n1528, n1522);
or   g1602 (n1632, n1501, n1543, n1535, n1556);
nand g1603 (n1628, n1476, n1528, n1465, n1492);
xnor g1604 (n1693, n1463, n1479, n1576, n1571);
xor  g1605 (n1612, n1580, n1500, n1545, n1555);
or   g1606 (n1719, n1546, n1514, n1468, n1495);
nor  g1607 (n1603, n1531, n1519, n1584, n1534);
and  g1608 (n1606, n1378, n1539, n1568, n1475);
and  g1609 (n1610, n1489, n1469, n1570, n1524);
and  g1610 (n1670, n1489, n1482, n1520, n1542);
xnor g1611 (n1643, n1482, n1543, n1457, n1515);
xor  g1612 (n1698, n1477, n1470, n1515, n1494);
xnor g1613 (n1726, n1479, n1504, n1567, n1464);
nor  g1614 (n1608, n1498, n1564, n1467, n1509);
xnor g1615 (n1645, n1496, n1464, n1451, n1556);
nand g1616 (n1587, n1480, n1462, n1530, n1537);
nand g1617 (n1651, n1504, n1486, n1502);
nor  g1618 (n1627, n1517, n1522, n1487, n1474);
nor  g1619 (n1721, n1578, n1575, n1559, n1493);
xnor g1620 (n1720, n1479, n1538, n1488, n1525);
nor  g1621 (n1680, n1578, n1520, n1452, n1515);
and  g1622 (n1609, n1450, n1476, n1507, n1579);
nor  g1623 (n1640, n1495, n1528, n1525, n1505);
xnor g1624 (n1689, n1556, n1464, n1450, n1474);
xnor g1625 (n1725, n1454, n1467, n1575, n1576);
and  g1626 (n1683, n1514, n1524, n1488, n1578);
or   g1627 (n1642, n1519, n1477, n1583, n1499);
nor  g1628 (n1619, n1563, n1536, n1559, n1476);
xor  g1629 (n1650, n1563, n1472, n1512, n1515);
and  g1630 (n1639, n1473, n1555, n1534, n1541);
xor  g1631 (n1637, n1500, n1523, n1563, n1522);
nor  g1632 (n1709, n1559, n1558, n1506, n1496);
and  g1633 (n1600, n1470, n1551, n1544, n1519);
nand g1634 (n1701, n1552, n1514, n1455, n1489);
and  g1635 (n1664, n1490, n1570, n1472, n1497);
nand g1636 (n1690, n1584, n1556, n1577, n1485);
nand g1637 (n1636, n1469, n1475, n1513, n1471);
nand g1638 (n1702, n1458, n1513, n1486, n1469);
xnor g1639 (n1597, n1554, n1516, n1541, n1560);
and  g1640 (n1652, n1459, n1496, n1483, n1567);
nand g1641 (n1644, n1529, n1518, n1542, n1566);
xor  g1642 (n1667, n1520, n1486, n1585, n1547);
or   g1643 (n1687, n1572, n1584, n1492, n1523);
or   g1644 (n1588, n1571, n1499, n1533, n1575);
and  g1645 (n1707, n1492, n1552, n1583, n1479);
and  g1646 (n1711, n1569, n1582, n1453, n1511);
nand g1647 (n1708, n1468, n1568, n1569, n1567);
nor  g1648 (n1656, n1560, n1472, n1566, n1475);
or   g1649 (n1679, n1521, n1485, n1562, n1582);
nor  g1650 (n1657, n1517, n1546, n1457, n1553);
xnor g1651 (n1692, n1574, n1566, n1579, n1580);
and  g1652 (n1617, n1490, n1505, n1546, n1522);
xnor g1653 (n1629, n1535, n1491, n1526, n1503);
nor  g1654 (n1678, n1501, n1475, n1548, n1494);
nand g1655 (n1611, n1536, n1530, n1488, n1583);
nand g1656 (n1723, n1483, n1503, n1481, n1459);
or   g1657 (n1671, n1531, n1557, n1453, n1561);
xnor g1658 (n1672, n1530, n1502, n1565, n1457);
or   g1659 (n1615, n1505, n1512, n1456, n1526);
and  g1660 (n1722, n1480, n1558, n1494, n1476);
or   g1661 (n1655, n1533, n1573, n1477, n1455);
nor  g1662 (n1653, n1580, n1550, n1474, n1496);
xnor g1663 (n1715, n1534, n1572, n1506, n1538);
nor  g1664 (n1718, n1542, n1529, n1574, n1501);
xnor g1665 (n1594, n1508, n1510, n1536, n1471);
and  g1666 (n1661, n1572, n1507, n1544, n1528);
xnor g1667 (n1674, n1478, n1558, n1536, n1471);
and  g1668 (n1673, n1462, n1571, n1521, n1506);
nor  g1669 (n1677, n1531, n1519, n1521, n1579);
xor  g1670 (n1620, n1569, n1565, n1467, n1527);
or   g1671 (n1686, n1539, n1483, n1513, n1537);
nand g1672 (n1649, n1545, n1455, n1491, n1540);
nand g1673 (n1665, n1574, n1532, n1502, n1456);
nand g1674 (n1669, n1463, n1537, n1466, n1493);
nand g1675 (n1625, n1544, n1582, n1484, n1526);
xnor g1676 (n1586, n1454, n1480, n1470, n1465);
xor  g1677 (n1601, n1550, n1548, n1560, n1564);
nand g1678 (n1638, n1537, n1470, n1565, n1497);
xor  g1679 (n1604, n1500, n1577, n1509, n1466);
nand g1680 (n1684, n1514, n1550, n1497, n1456);
and  g1681 (n1663, n1560, n1518, n1542, n1569);
xor  g1682 (n1724, n1453, n1494, n1508, n1553);
xor  g1683 (n1626, n1488, n1575, n1518, n1562);
nor  g1684 (n1616, n1568, n1511, n1493, n1540);
and  g1685 (n1716, n1558, n1481, n1480, n1562);
or   g1686 (n1691, n1564, n1491, n1498, n1478);
xnor g1687 (n1618, n1460, n1376, n1518, n1540);
and  g1688 (n1634, n1532, n1571, n1509, n1547);
or   g1689 (n1666, n1582, n1484, n1561);
nor  g1690 (n1727, n1482, n1529, n1539, n1454);
nor  g1691 (n1602, n1461, n1584, n1579, n1510);
xnor g1692 (n1713, n1564, n1555, n1516, n1577);
nor  g1693 (n1631, n1563, n1472, n1507, n1551);
nor  g1694 (n1591, n1459, n1576, n1533, n1451);
xnor g1695 (n1706, n1546, n1483, n1541, n1568);
or   g1696 (n1710, n1580, n1500, n1585, n1477);
not  g1697 (n2149, n1594);
not  g1698 (n2069, n1592);
buf  g1699 (n1818, n1694);
buf  g1700 (n2295, n1690);
buf  g1701 (n2055, n1631);
buf  g1702 (n1893, n1674);
buf  g1703 (n2105, n1613);
buf  g1704 (n1936, n1655);
not  g1705 (n1899, n1641);
not  g1706 (n1851, n1667);
buf  g1707 (n2288, n1671);
buf  g1708 (n1872, n1714);
buf  g1709 (n2050, n1721);
buf  g1710 (n1831, n1727);
buf  g1711 (n1875, n1607);
not  g1712 (n2134, n1706);
buf  g1713 (n2218, n1634);
not  g1714 (n1780, n1594);
not  g1715 (n2094, n1692);
not  g1716 (n1981, n1592);
buf  g1717 (n1920, n1608);
not  g1718 (n1951, n1670);
not  g1719 (n1871, n1662);
buf  g1720 (n1988, n1105);
not  g1721 (n2184, n1587);
buf  g1722 (n1783, n1624);
not  g1723 (n2238, n1616);
buf  g1724 (n1976, n1597);
buf  g1725 (n2067, n1710);
buf  g1726 (n2128, n1714);
buf  g1727 (n2084, n1689);
not  g1728 (n1907, n1640);
buf  g1729 (n2133, n1603);
not  g1730 (n1992, n1601);
buf  g1731 (n2029, n1670);
buf  g1732 (n2173, n1716);
not  g1733 (n1958, n1724);
buf  g1734 (n1770, n1693);
not  g1735 (n1828, n1675);
not  g1736 (n1793, n1716);
not  g1737 (n2066, n1701);
not  g1738 (n1748, n1710);
buf  g1739 (n1733, n1626);
buf  g1740 (n2042, n1632);
buf  g1741 (n1952, n1636);
not  g1742 (n1888, n1588);
buf  g1743 (n2145, n1647);
not  g1744 (n2228, n1666);
buf  g1745 (n1977, n1599);
not  g1746 (n2119, n1620);
not  g1747 (n2085, n1638);
buf  g1748 (n1879, n1715);
buf  g1749 (n1815, n1694);
buf  g1750 (n2167, n1588);
not  g1751 (n2232, n1674);
buf  g1752 (n2110, n1661);
not  g1753 (n1751, n1656);
buf  g1754 (n1971, n1590);
buf  g1755 (n2198, n1394);
buf  g1756 (n2292, n1650);
not  g1757 (n1759, n1643);
buf  g1758 (n2070, n1640);
not  g1759 (n1795, n1655);
buf  g1760 (n1821, n1653);
buf  g1761 (n1959, n1708);
not  g1762 (n2108, n1714);
buf  g1763 (n1985, n1654);
buf  g1764 (n2098, n1677);
not  g1765 (n1973, n1652);
buf  g1766 (n2284, n1644);
buf  g1767 (n2111, n1652);
not  g1768 (n2188, n1103);
not  g1769 (n2081, n1655);
buf  g1770 (n1832, n1686);
not  g1771 (n2201, n1632);
not  g1772 (n1999, n1699);
not  g1773 (n2087, n1678);
not  g1774 (n1867, n1719);
buf  g1775 (n1752, n1659);
buf  g1776 (n1826, n1718);
buf  g1777 (n1891, n1606);
buf  g1778 (n2044, n1685);
buf  g1779 (n1801, n1617);
not  g1780 (n2025, n1703);
buf  g1781 (n2005, n1672);
buf  g1782 (n2073, n1643);
not  g1783 (n1924, n1702);
buf  g1784 (n2250, n1675);
buf  g1785 (n1775, n1711);
buf  g1786 (n2199, n1594);
not  g1787 (n2291, n1610);
not  g1788 (n2010, n1596);
not  g1789 (n1843, n1597);
buf  g1790 (n2285, n1726);
not  g1791 (n1796, n1608);
not  g1792 (n2008, n1646);
buf  g1793 (n1850, n1608);
not  g1794 (n2019, n1598);
not  g1795 (n2273, n1589);
not  g1796 (n2101, n1711);
buf  g1797 (n1838, n1676);
not  g1798 (n2013, n1668);
buf  g1799 (n1797, n1637);
not  g1800 (n1822, n1612);
not  g1801 (n1906, n1605);
buf  g1802 (n2182, n1652);
not  g1803 (n2107, n1635);
buf  g1804 (n1814, n1714);
not  g1805 (n1987, n1688);
not  g1806 (n2086, n1693);
not  g1807 (n2132, n1630);
buf  g1808 (n2220, n1393);
not  g1809 (n2233, n1615);
buf  g1810 (n2117, n1594);
buf  g1811 (n1945, n1600);
buf  g1812 (n2287, n1104);
not  g1813 (n2155, n1589);
not  g1814 (n2022, n1716);
buf  g1815 (n1877, n1642);
not  g1816 (n2118, n1720);
buf  g1817 (n1873, n1671);
not  g1818 (n2046, n1599);
buf  g1819 (n1842, n1648);
buf  g1820 (n2102, n1632);
buf  g1821 (n1950, n1595);
buf  g1822 (n2264, n1688);
buf  g1823 (n2270, n1698);
buf  g1824 (n2282, n1619);
not  g1825 (n2205, n1697);
buf  g1826 (n2003, n1713);
buf  g1827 (n1840, n1697);
not  g1828 (n2209, n1640);
buf  g1829 (n2126, n1654);
not  g1830 (n2063, n1680);
not  g1831 (n2278, n1597);
buf  g1832 (n2179, n1649);
not  g1833 (n2169, n1653);
buf  g1834 (n1889, n1618);
buf  g1835 (n1844, n1619);
not  g1836 (n1990, n1586);
buf  g1837 (n1972, n1693);
not  g1838 (n2141, n1702);
not  g1839 (n2164, n1647);
buf  g1840 (n2100, n1627);
buf  g1841 (n1753, n1706);
buf  g1842 (n1943, n1705);
not  g1843 (n2300, n1705);
buf  g1844 (n1970, n1675);
buf  g1845 (n2196, n1625);
not  g1846 (n2213, n1669);
buf  g1847 (n2052, n1592);
buf  g1848 (n2243, n1393);
not  g1849 (n2174, n1614);
buf  g1850 (n1955, n1604);
buf  g1851 (n1912, n1698);
not  g1852 (n1964, n1682);
buf  g1853 (n2131, n1661);
not  g1854 (n1868, n1662);
not  g1855 (n1803, n1621);
not  g1856 (n2170, n1624);
not  g1857 (n1993, n1614);
not  g1858 (n2048, n1611);
not  g1859 (n2212, n1722);
not  g1860 (n2263, n1101);
buf  g1861 (n1997, n1660);
buf  g1862 (n1755, n1713);
buf  g1863 (n1865, n1687);
buf  g1864 (n2033, n1642);
buf  g1865 (n2047, n1593);
not  g1866 (n1789, n1681);
not  g1867 (n2020, n1651);
not  g1868 (n2142, n1600);
not  g1869 (n2299, n1626);
buf  g1870 (n1781, n1694);
buf  g1871 (n1807, n1663);
not  g1872 (n2241, n1634);
not  g1873 (n1904, n1661);
not  g1874 (n1967, n1729);
buf  g1875 (n1863, n1667);
buf  g1876 (n2137, n1631);
buf  g1877 (n1954, n1659);
buf  g1878 (n2258, n1641);
buf  g1879 (n1806, n1622);
not  g1880 (n1817, n1602);
not  g1881 (n2214, n1601);
not  g1882 (n2023, n1680);
not  g1883 (n2227, n1709);
buf  g1884 (n1827, n1631);
not  g1885 (n2115, n1698);
not  g1886 (n2181, n1682);
buf  g1887 (n2056, n1606);
buf  g1888 (n2014, n1644);
buf  g1889 (n1901, n1664);
not  g1890 (n2125, n1623);
buf  g1891 (n2071, n1593);
buf  g1892 (n2301, n1691);
not  g1893 (n1880, n1645);
buf  g1894 (n2224, n1699);
buf  g1895 (n2231, n1717);
not  g1896 (n1834, n1704);
not  g1897 (n2193, n1613);
not  g1898 (n2266, n1707);
not  g1899 (n1922, n1639);
not  g1900 (n2180, n1710);
not  g1901 (n2172, n1637);
not  g1902 (n1737, n1728);
buf  g1903 (n2146, n1658);
not  g1904 (n2016, n1614);
buf  g1905 (n2060, n1692);
buf  g1906 (n1749, n1721);
buf  g1907 (n1866, n1588);
buf  g1908 (n1932, n1612);
buf  g1909 (n2153, n1691);
buf  g1910 (n1984, n1612);
buf  g1911 (n1809, n1635);
buf  g1912 (n1812, n1718);
buf  g1913 (n2058, n1626);
buf  g1914 (n2150, n1106);
not  g1915 (n2267, n1641);
not  g1916 (n2253, n1623);
buf  g1917 (n2247, n1606);
buf  g1918 (n2161, n1646);
buf  g1919 (n2234, n1604);
not  g1920 (n1942, n1633);
buf  g1921 (n1849, n1642);
not  g1922 (n1915, n1663);
not  g1923 (n2035, n1678);
not  g1924 (n2135, n1607);
not  g1925 (n2176, n1606);
not  g1926 (n1963, n1635);
buf  g1927 (n2075, n1613);
buf  g1928 (n1900, n1625);
not  g1929 (n2039, n1707);
not  g1930 (n1882, n1622);
not  g1931 (n1769, n1665);
not  g1932 (n2203, n1609);
buf  g1933 (n1919, n1644);
buf  g1934 (n2144, n1612);
buf  g1935 (n2026, n1703);
buf  g1936 (n2297, n1589);
not  g1937 (n1799, n1588);
not  g1938 (n2024, n1715);
not  g1939 (n2254, n1679);
not  g1940 (n1895, n1692);
not  g1941 (n2239, n1610);
buf  g1942 (n2077, n1697);
buf  g1943 (n1833, n1628);
buf  g1944 (n1824, n1727);
buf  g1945 (n2240, n1677);
buf  g1946 (n1830, n1719);
not  g1947 (n1961, n1661);
not  g1948 (n2268, n1684);
not  g1949 (n1836, n1707);
not  g1950 (n2225, n1721);
not  g1951 (n2261, n1695);
buf  g1952 (n1876, n1724);
not  g1953 (n1946, n1684);
buf  g1954 (n2293, n1590);
not  g1955 (n2124, n1723);
buf  g1956 (n2256, n1642);
not  g1957 (n2252, n1682);
not  g1958 (n1772, n1659);
buf  g1959 (n1734, n1673);
buf  g1960 (n2040, n1703);
buf  g1961 (n2021, n1713);
not  g1962 (n1837, n1683);
buf  g1963 (n1750, n1698);
buf  g1964 (n1760, n1705);
buf  g1965 (n1825, n1628);
not  g1966 (n1966, n1645);
buf  g1967 (n1839, n1596);
not  g1968 (n1841, n1669);
buf  g1969 (n1918, n1727);
buf  g1970 (n1858, n1623);
not  g1971 (n2078, n1605);
buf  g1972 (n1897, n1628);
not  g1973 (n1940, n1725);
not  g1974 (n1884, n1630);
not  g1975 (n2211, n1629);
not  g1976 (n2269, n1641);
buf  g1977 (n1887, n1621);
buf  g1978 (n1823, n1648);
buf  g1979 (n1948, n1670);
buf  g1980 (n2244, n1715);
buf  g1981 (n2001, n1652);
buf  g1982 (n2186, n1656);
buf  g1983 (n2158, n1587);
not  g1984 (n1757, n1674);
not  g1985 (n1938, n1648);
not  g1986 (n2030, n1723);
buf  g1987 (n1785, n1713);
buf  g1988 (n1881, n1677);
not  g1989 (n1996, n1636);
not  g1990 (n2157, n1681);
buf  g1991 (n2009, n1595);
buf  g1992 (n2064, n1658);
not  g1993 (n1957, n1710);
not  g1994 (n2206, n1701);
buf  g1995 (n2147, n1615);
buf  g1996 (n2177, n1621);
not  g1997 (n2248, n1689);
not  g1998 (n2304, n1603);
not  g1999 (n1917, n1687);
buf  g2000 (n2091, n1704);
not  g2001 (n2138, n1638);
not  g2002 (n2208, n1673);
buf  g2003 (n1965, n1715);
not  g2004 (n2305, n1599);
buf  g2005 (n2187, n1625);
not  g2006 (n1732, n1684);
not  g2007 (n1991, n1685);
buf  g2008 (n1896, n1645);
not  g2009 (n1929, n1660);
buf  g2010 (n2251, n1609);
not  g2011 (n1947, n1650);
not  g2012 (n2204, n1718);
not  g2013 (n2221, n1627);
not  g2014 (n2230, n1729);
buf  g2015 (n2127, n1631);
buf  g2016 (n1845, n1657);
not  g2017 (n1835, n1637);
not  g2018 (n2162, n1668);
not  g2019 (n2272, n1687);
buf  g2020 (n1805, n1672);
buf  g2021 (n2004, n1610);
not  g2022 (n2089, n1688);
buf  g2023 (n1935, n1636);
not  g2024 (n1949, n1676);
not  g2025 (n2045, n1690);
buf  g2026 (n1986, n1717);
buf  g2027 (n2109, n1394);
buf  g2028 (n2302, n1687);
not  g2029 (n1808, n1620);
buf  g2030 (n1846, n1634);
buf  g2031 (n2189, n1628);
buf  g2032 (n2274, n1394);
buf  g2033 (n1730, n1650);
buf  g2034 (n2160, n1678);
not  g2035 (n1994, n1666);
buf  g2036 (n2151, n1616);
not  g2037 (n1898, n1647);
not  g2038 (n1995, n1664);
not  g2039 (n2219, n1632);
not  g2040 (n1862, n1703);
not  g2041 (n2116, n1726);
buf  g2042 (n1790, n1665);
buf  g2043 (n2074, n1720);
buf  g2044 (n2088, n1598);
not  g2045 (n2143, n1666);
buf  g2046 (n2027, n1673);
not  g2047 (n2303, n1665);
not  g2048 (n2242, n1638);
not  g2049 (n1735, n1721);
not  g2050 (n1738, n1640);
buf  g2051 (n2166, n1651);
buf  g2052 (n1869, n1649);
buf  g2053 (n2034, n1596);
buf  g2054 (n1739, n1636);
buf  g2055 (n1933, n1720);
buf  g2056 (n1848, n1394);
buf  g2057 (n2129, n1700);
not  g2058 (n1763, n1593);
buf  g2059 (n2168, n1622);
buf  g2060 (n1746, n1644);
not  g2061 (n1736, n1627);
not  g2062 (n2018, n1699);
not  g2063 (n2096, n1672);
buf  g2064 (n1883, n1664);
buf  g2065 (n1892, n1719);
not  g2066 (n1860, n1622);
not  g2067 (n2103, n1712);
buf  g2068 (n2015, n1728);
buf  g2069 (n2194, n1586);
buf  g2070 (n2290, n1614);
not  g2071 (n1782, n1591);
not  g2072 (n1926, n1723);
buf  g2073 (n1820, n1648);
buf  g2074 (n1989, n1693);
buf  g2075 (n2043, n1681);
not  g2076 (n1804, n1718);
buf  g2077 (n2106, n1711);
buf  g2078 (n2215, n1587);
not  g2079 (n1861, n1618);
not  g2080 (n2236, n1691);
buf  g2081 (n1794, n1591);
buf  g2082 (n1921, n1611);
not  g2083 (n2006, n1607);
not  g2084 (n2294, n1646);
buf  g2085 (n1962, n1618);
buf  g2086 (n1786, n1102);
not  g2087 (n2061, n1728);
not  g2088 (n2217, n1602);
not  g2089 (n1914, n1673);
buf  g2090 (n2082, n1627);
buf  g2091 (n2051, n1607);
buf  g2092 (n1878, n1604);
buf  g2093 (n2097, n1668);
buf  g2094 (n2099, n1702);
not  g2095 (n1811, n1680);
not  g2096 (n1791, n1654);
not  g2097 (n1743, n1600);
not  g2098 (n2265, n1656);
buf  g2099 (n1885, n1601);
not  g2100 (n2216, n1616);
buf  g2101 (n2190, n1686);
not  g2102 (n1756, n1655);
buf  g2103 (n2036, n1708);
not  g2104 (n1905, n1695);
not  g2105 (n2235, n1646);
not  g2106 (n2148, n1726);
not  g2107 (n2154, n1393);
not  g2108 (n2156, n1591);
buf  g2109 (n2260, n1608);
buf  g2110 (n1944, n1651);
not  g2111 (n1853, n1663);
buf  g2112 (n1784, n1621);
not  g2113 (n1975, n1701);
not  g2114 (n1930, n1658);
not  g2115 (n2281, n1672);
buf  g2116 (n1956, n1616);
not  g2117 (n1934, n1725);
not  g2118 (n2053, n1605);
not  g2119 (n2002, n1657);
buf  g2120 (n2112, n1700);
buf  g2121 (n1776, n1696);
not  g2122 (n2104, n1586);
buf  g2123 (n2120, n1708);
buf  g2124 (n2031, n1624);
buf  g2125 (n2113, n1722);
buf  g2126 (n1802, n1596);
buf  g2127 (n1902, n1589);
not  g2128 (n1911, n1666);
buf  g2129 (n1980, n1692);
buf  g2130 (n2065, n1602);
buf  g2131 (n1927, n1617);
not  g2132 (n2076, n1679);
buf  g2133 (n2000, n1707);
buf  g2134 (n2276, n1635);
not  g2135 (n1974, n1590);
buf  g2136 (n1754, n1639);
not  g2137 (n2095, n1592);
buf  g2138 (n1747, n1601);
not  g2139 (n2192, n1706);
not  g2140 (n2197, n1630);
buf  g2141 (n1798, n1728);
buf  g2142 (n2185, n1729);
buf  g2143 (n2202, n1712);
buf  g2144 (n1890, n1682);
buf  g2145 (n2195, n1676);
buf  g2146 (n2271, n1603);
buf  g2147 (n2011, n1702);
not  g2148 (n1778, n1618);
buf  g2149 (n1998, n1619);
not  g2150 (n2007, n1681);
buf  g2151 (n2255, n1662);
buf  g2152 (n1744, n1643);
buf  g2153 (n1788, n1711);
buf  g2154 (n2059, n1697);
not  g2155 (n2093, n1651);
not  g2156 (n1766, n1689);
not  g2157 (n1765, n1609);
buf  g2158 (n1764, n1656);
buf  g2159 (n1909, n1657);
not  g2160 (n1731, n1669);
buf  g2161 (n1816, n1680);
buf  g2162 (n1742, n1684);
buf  g2163 (n1913, n1695);
buf  g2164 (n2165, n1654);
not  g2165 (n1741, n1620);
buf  g2166 (n1855, n1657);
buf  g2167 (n2171, n1708);
buf  g2168 (n2136, n1688);
not  g2169 (n1773, n1686);
not  g2170 (n2092, n1623);
buf  g2171 (n2191, n1694);
not  g2172 (n1908, n1630);
buf  g2173 (n1968, n1709);
not  g2174 (n2226, n1639);
not  g2175 (n2012, n1676);
buf  g2176 (n2139, n1685);
buf  g2177 (n2121, n1611);
not  g2178 (n2090, n1704);
not  g2179 (n2283, n1696);
buf  g2180 (n1978, n1586);
buf  g2181 (n1777, n1619);
buf  g2182 (n2028, n1643);
not  g2183 (n1903, n1683);
buf  g2184 (n1771, n1720);
buf  g2185 (n2183, n1645);
buf  g2186 (n2080, n1633);
not  g2187 (n2289, n1653);
buf  g2188 (n1983, n1649);
not  g2189 (n2114, n1706);
buf  g2190 (n1857, n1729);
not  g2191 (n2259, n1671);
buf  g2192 (n2123, n1658);
buf  g2193 (n2072, n1393);
buf  g2194 (n1910, n1590);
buf  g2195 (n1800, n1600);
buf  g2196 (n2245, n1699);
not  g2197 (n2237, n1683);
buf  g2198 (n1923, n1701);
buf  g2199 (n2140, n1679);
buf  g2200 (n2130, n1597);
not  g2201 (n1937, n1653);
buf  g2202 (n2286, n1700);
not  g2203 (n2249, n1725);
not  g2204 (n1939, n1717);
not  g2205 (n1740, n1690);
buf  g2206 (n1916, n1664);
buf  g2207 (n1819, n1649);
buf  g2208 (n2210, n1634);
not  g2209 (n2037, n1696);
not  g2210 (n1792, n1678);
not  g2211 (n2054, n1671);
not  g2212 (n1852, n1696);
not  g2213 (n2159, n1722);
not  g2214 (n1925, n1605);
not  g2215 (n2229, n1689);
buf  g2216 (n1941, n1725);
buf  g2217 (n2083, n1380);
buf  g2218 (n1856, n1669);
not  g2219 (n2175, n1668);
not  g2220 (n1886, n1609);
buf  g2221 (n2122, n1598);
buf  g2222 (n2277, n1610);
not  g2223 (n1874, n1639);
buf  g2224 (n2280, n1717);
buf  g2225 (n2275, n1633);
not  g2226 (n1829, n1624);
not  g2227 (n1761, n1723);
not  g2228 (n2068, n1686);
buf  g2229 (n1982, n1637);
not  g2230 (n2057, n1633);
buf  g2231 (n1859, n1611);
buf  g2232 (n2257, n1695);
not  g2233 (n2262, n1712);
not  g2234 (n1969, n1620);
buf  g2235 (n1953, n1691);
buf  g2236 (n1810, n1626);
buf  g2237 (n2041, n1722);
not  g2238 (n1787, n1667);
buf  g2239 (n1854, n1595);
buf  g2240 (n2246, n1629);
buf  g2241 (n1758, n1107);
buf  g2242 (n2038, n1617);
not  g2243 (n2296, n1683);
not  g2244 (n2223, n1647);
not  g2245 (n1847, n1638);
not  g2246 (n1864, n1716);
buf  g2247 (n1979, n1615);
not  g2248 (n2163, n1724);
buf  g2249 (n2298, n1629);
buf  g2250 (n1774, n1704);
buf  g2251 (n2017, n1598);
not  g2252 (n1931, n1613);
buf  g2253 (n2222, n1625);
not  g2254 (n2049, n1604);
not  g2255 (n2079, n1709);
buf  g2256 (n1768, n1685);
buf  g2257 (n1767, n1674);
buf  g2258 (n1762, n1712);
not  g2259 (n1894, n1705);
buf  g2260 (n2279, n1670);
not  g2261 (n1779, n1719);
buf  g2262 (n2200, n1700);
buf  g2263 (n2207, n1677);
buf  g2264 (n1870, n1724);
buf  g2265 (n1928, n1617);
not  g2266 (n2032, n1615);
and  g2267 (n1813, n1667, n1603);
xnor g2268 (n2178, n1591, n1660, n1659, n1602);
or   g2269 (n2062, n1726, n1587, n1665, n1663);
xor  g2270 (n2152, n1595, n1599, n1690, n1709);
nand g2271 (n1960, n1662, n1727, n1593, n1660);
nand g2272 (n1745, n1629, n1650, n1679, n1675);
not  g2273 (n2428, n1990);
buf  g2274 (n3438, n2039);
not  g2275 (n2860, n2159);
buf  g2276 (n3250, n1931);
buf  g2277 (n3570, n1750);
not  g2278 (n2533, n2263);
not  g2279 (n3154, n1944);
not  g2280 (n3451, n2124);
not  g2281 (n3041, n1827);
buf  g2282 (n2575, n2003);
buf  g2283 (n3104, n2126);
not  g2284 (n2981, n2128);
buf  g2285 (n3442, n1838);
not  g2286 (n2799, n2220);
not  g2287 (n2711, n1793);
not  g2288 (n3299, n1931);
buf  g2289 (n2891, n2222);
not  g2290 (n2426, n1867);
buf  g2291 (n3336, n2036);
not  g2292 (n3487, n2053);
not  g2293 (n2918, n1843);
not  g2294 (n3381, n1899);
buf  g2295 (n2693, n2059);
buf  g2296 (n2613, n2193);
buf  g2297 (n2703, n1988);
buf  g2298 (n2994, n2127);
buf  g2299 (n2848, n2184);
buf  g2300 (n2657, n2015);
not  g2301 (n2805, n2082);
buf  g2302 (n2774, n1933);
buf  g2303 (n2489, n1944);
not  g2304 (n2556, n1988);
buf  g2305 (n2697, n1407);
buf  g2306 (n3082, n2266);
buf  g2307 (n3345, n2093);
buf  g2308 (n3449, n2155);
buf  g2309 (n3358, n1802);
not  g2310 (n3198, n2107);
not  g2311 (n3244, n1887);
not  g2312 (n3492, n2032);
not  g2313 (n2551, n1792);
not  g2314 (n2892, n2082);
buf  g2315 (n3223, n2148);
not  g2316 (n2895, n1869);
buf  g2317 (n3084, n2127);
not  g2318 (n3501, n1915);
not  g2319 (n3016, n2133);
not  g2320 (n3480, n1992);
not  g2321 (n3183, n2215);
buf  g2322 (n2319, n2267);
buf  g2323 (n3535, n1787);
not  g2324 (n2769, n2189);
not  g2325 (n2737, n2130);
not  g2326 (n2328, n1960);
buf  g2327 (n2659, n1965);
not  g2328 (n2338, n2055);
buf  g2329 (n3165, n2029);
buf  g2330 (n3404, n1769);
not  g2331 (n3114, n2004);
buf  g2332 (n3204, n1826);
not  g2333 (n2803, n2067);
buf  g2334 (n2735, n1755);
not  g2335 (n2558, n1914);
not  g2336 (n3057, n1402);
buf  g2337 (n2496, n1818);
not  g2338 (n2924, n2096);
not  g2339 (n3465, n1832);
buf  g2340 (n2450, n1939);
not  g2341 (n2595, n2114);
buf  g2342 (n2755, n1927);
not  g2343 (n3567, n2264);
buf  g2344 (n3382, n1901);
buf  g2345 (n3145, n2031);
not  g2346 (n2451, n1915);
not  g2347 (n3253, n2024);
not  g2348 (n3488, n2245);
buf  g2349 (n2869, n2213);
buf  g2350 (n2427, n2073);
buf  g2351 (n3008, n1407);
not  g2352 (n2654, n2199);
not  g2353 (n2567, n2257);
buf  g2354 (n2806, n1959);
buf  g2355 (n2494, n2072);
buf  g2356 (n2968, n2019);
buf  g2357 (n3290, n1883);
buf  g2358 (n3519, n2163);
buf  g2359 (n3127, n2253);
not  g2360 (n2749, n2170);
buf  g2361 (n2813, n1896);
buf  g2362 (n3254, n1990);
buf  g2363 (n2868, n1886);
not  g2364 (n2384, n2224);
buf  g2365 (n3237, n2290);
not  g2366 (n2701, n1878);
not  g2367 (n2316, n1937);
not  g2368 (n2762, n2303);
buf  g2369 (n2761, n2099);
buf  g2370 (n2359, n1829);
not  g2371 (n3096, n2136);
not  g2372 (n3302, n2123);
buf  g2373 (n3272, n1864);
not  g2374 (n2962, n2125);
not  g2375 (n2344, n2294);
buf  g2376 (n2557, n1877);
not  g2377 (n2442, n1776);
not  g2378 (n2925, n1924);
not  g2379 (n2829, n1816);
buf  g2380 (n2497, n1944);
buf  g2381 (n3426, n1404);
not  g2382 (n2624, n2000);
buf  g2383 (n2910, n1787);
buf  g2384 (n3394, n2225);
buf  g2385 (n2974, n1987);
not  g2386 (n3396, n2272);
buf  g2387 (n2626, n1408);
not  g2388 (n3533, n1871);
buf  g2389 (n3243, n1971);
not  g2390 (n2424, n2030);
not  g2391 (n2437, n2000);
buf  g2392 (n3474, n2169);
buf  g2393 (n2771, n1790);
buf  g2394 (n2398, n2023);
buf  g2395 (n3398, n2297);
buf  g2396 (n3142, n1917);
not  g2397 (n3115, n1851);
buf  g2398 (n2425, n2195);
not  g2399 (n3326, n2225);
buf  g2400 (n2719, n1111);
not  g2401 (n3322, n2269);
buf  g2402 (n2388, n2023);
buf  g2403 (n2789, n1908);
not  g2404 (n3123, n2249);
not  g2405 (n3403, n2141);
buf  g2406 (n2678, n1876);
buf  g2407 (n3386, n1880);
buf  g2408 (n2381, n2179);
not  g2409 (n2760, n1901);
buf  g2410 (n3370, n1967);
not  g2411 (n2589, n2046);
buf  g2412 (n3318, n2075);
not  g2413 (n2430, n1757);
buf  g2414 (n2941, n2097);
buf  g2415 (n3051, n2117);
buf  g2416 (n2397, n2108);
not  g2417 (n3425, n2146);
not  g2418 (n2683, n2066);
buf  g2419 (n2696, n2206);
not  g2420 (n3528, n1961);
not  g2421 (n2562, n2256);
buf  g2422 (n3282, n2134);
buf  g2423 (n3062, n1882);
buf  g2424 (n3077, n1912);
buf  g2425 (n2436, n1899);
buf  g2426 (n3561, n1848);
buf  g2427 (n3087, n2204);
buf  g2428 (n3085, n2144);
not  g2429 (n3242, n2111);
not  g2430 (n2480, n2121);
not  g2431 (n3280, n2186);
not  g2432 (n2842, n1995);
buf  g2433 (n2585, n1821);
buf  g2434 (n2509, n1848);
not  g2435 (n3140, n2249);
buf  g2436 (n3066, n2229);
buf  g2437 (n2690, n1853);
not  g2438 (n3011, n2101);
not  g2439 (n2700, n2152);
buf  g2440 (n2725, n1730);
not  g2441 (n2523, n2282);
buf  g2442 (n2993, n2149);
not  g2443 (n3543, n2159);
buf  g2444 (n2541, n2185);
not  g2445 (n2444, n1739);
not  g2446 (n2965, n2121);
not  g2447 (n3541, n1894);
buf  g2448 (n2705, n2196);
buf  g2449 (n3021, n2004);
buf  g2450 (n3342, n2167);
buf  g2451 (n2874, n2280);
not  g2452 (n2420, n2228);
not  g2453 (n3484, n1860);
not  g2454 (n3010, n1732);
not  g2455 (n2311, n2016);
not  g2456 (n3030, n1929);
buf  g2457 (n2720, n1404);
not  g2458 (n2904, n2270);
buf  g2459 (n2669, n2043);
buf  g2460 (n2505, n2096);
buf  g2461 (n2315, n2014);
not  g2462 (n2521, n2180);
not  g2463 (n3300, n2095);
buf  g2464 (n2409, n2189);
not  g2465 (n3070, n2120);
buf  g2466 (n3267, n2192);
buf  g2467 (n2449, n1828);
buf  g2468 (n3549, n2158);
not  g2469 (n2591, n1923);
not  g2470 (n3189, n2195);
not  g2471 (n2491, n1802);
buf  g2472 (n2759, n2008);
not  g2473 (n2744, n2019);
buf  g2474 (n2845, n1961);
not  g2475 (n2676, n2284);
not  g2476 (n2743, n1796);
buf  g2477 (n2630, n1813);
not  g2478 (n3159, n2167);
buf  g2479 (n2840, n1875);
not  g2480 (n3368, n1894);
buf  g2481 (n2615, n2271);
not  g2482 (n2861, n1995);
not  g2483 (n2940, n1805);
buf  g2484 (n2673, n1848);
not  g2485 (n2818, n1403);
buf  g2486 (n2461, n2013);
buf  g2487 (n3294, n1740);
buf  g2488 (n2317, n1898);
buf  g2489 (n2643, n2148);
not  g2490 (n3330, n1920);
buf  g2491 (n2423, n2203);
buf  g2492 (n2609, n1983);
not  g2493 (n3291, n2274);
not  g2494 (n2622, n1906);
buf  g2495 (n3390, n2212);
buf  g2496 (n3285, n2069);
buf  g2497 (n2881, n1995);
not  g2498 (n3222, n1940);
not  g2499 (n2825, n1408);
buf  g2500 (n2441, n1988);
not  g2501 (n3035, n2160);
buf  g2502 (n3428, n2238);
not  g2503 (n2400, n2077);
buf  g2504 (n2837, n1942);
buf  g2505 (n2960, n2090);
not  g2506 (n2752, n1945);
buf  g2507 (n2472, n1745);
buf  g2508 (n3040, n2254);
not  g2509 (n3281, n1889);
buf  g2510 (n3516, n2300);
not  g2511 (n2808, n2048);
not  g2512 (n2379, n2232);
not  g2513 (n3172, n2121);
buf  g2514 (n3439, n2096);
not  g2515 (n3053, n1948);
not  g2516 (n2466, n2031);
buf  g2517 (n3468, n1918);
buf  g2518 (n2517, n2130);
buf  g2519 (n3113, n2068);
not  g2520 (n2353, n1977);
not  g2521 (n2973, n1972);
buf  g2522 (n3103, n2017);
buf  g2523 (n2607, n1974);
buf  g2524 (n2366, n1810);
not  g2525 (n2688, n2018);
not  g2526 (n3216, n1907);
buf  g2527 (n2531, n1944);
not  g2528 (n2715, n1409);
not  g2529 (n2470, n2189);
not  g2530 (n3555, n2215);
not  g2531 (n2951, n2063);
not  g2532 (n2686, n2297);
buf  g2533 (n2432, n1951);
buf  g2534 (n2897, n1866);
not  g2535 (n2367, n1972);
buf  g2536 (n3546, n2089);
not  g2537 (n3068, n2042);
not  g2538 (n3235, n2301);
not  g2539 (n2545, n1933);
buf  g2540 (n3099, n2242);
buf  g2541 (n2820, n1967);
not  g2542 (n3392, n2270);
buf  g2543 (n2456, n2139);
buf  g2544 (n2792, n2188);
buf  g2545 (n3080, n2114);
not  g2546 (n2401, n2181);
buf  g2547 (n3109, n1830);
not  g2548 (n2515, n1950);
buf  g2549 (n3153, n2003);
not  g2550 (n3043, n1926);
buf  g2551 (n3185, n2181);
not  g2552 (n3264, n2124);
not  g2553 (n3262, n1812);
buf  g2554 (n3412, n1225);
not  g2555 (n2342, n1926);
not  g2556 (n2952, n2098);
buf  g2557 (n2922, n1402);
not  g2558 (n3045, n2028);
buf  g2559 (n3058, n2135);
not  g2560 (n3469, n2298);
not  g2561 (n3167, n1819);
buf  g2562 (n2620, n1871);
buf  g2563 (n2991, n1761);
buf  g2564 (n3323, n2208);
not  g2565 (n2856, n1977);
buf  g2566 (n2581, n2029);
not  g2567 (n2791, n2057);
not  g2568 (n3246, n1911);
buf  g2569 (n3436, n2231);
buf  g2570 (n2467, n1856);
not  g2571 (n2525, n2080);
not  g2572 (n2816, n2278);
not  g2573 (n3102, n1981);
not  g2574 (n2957, n2244);
not  g2575 (n2390, n2140);
not  g2576 (n3268, n2002);
buf  g2577 (n2386, n2219);
buf  g2578 (n2888, n2141);
buf  g2579 (n3462, n1961);
not  g2580 (n3117, n2208);
buf  g2581 (n2361, n1987);
buf  g2582 (n3489, n1954);
buf  g2583 (n2695, n2300);
not  g2584 (n2309, n2293);
not  g2585 (n2590, n1972);
buf  g2586 (n2872, n2063);
not  g2587 (n3328, n1941);
not  g2588 (n2464, n2169);
buf  g2589 (n3341, n2184);
not  g2590 (n3182, n1804);
not  g2591 (n3337, n1908);
not  g2592 (n2513, n1940);
not  g2593 (n3174, n2049);
not  g2594 (n3233, n1956);
buf  g2595 (n2689, n2082);
not  g2596 (n2641, n1733);
not  g2597 (n2768, n2210);
buf  g2598 (n3470, n1818);
not  g2599 (n3572, n2258);
not  g2600 (n3201, n1787);
buf  g2601 (n3359, n1879);
buf  g2602 (n2666, n2111);
not  g2603 (n3307, n1895);
buf  g2604 (n3269, n1805);
buf  g2605 (n2445, n2004);
buf  g2606 (n3176, n2132);
buf  g2607 (n2510, n2129);
buf  g2608 (n2375, n1829);
not  g2609 (n3437, n2136);
buf  g2610 (n2336, n2059);
not  g2611 (n3418, n1992);
buf  g2612 (n3406, n1915);
buf  g2613 (n3479, n2221);
not  g2614 (n3357, n1885);
not  g2615 (n3255, n1849);
buf  g2616 (n2605, n1920);
buf  g2617 (n3052, n1970);
buf  g2618 (n3106, n2265);
buf  g2619 (n2618, n1902);
buf  g2620 (n3321, n2060);
buf  g2621 (n2950, n2077);
buf  g2622 (n2429, n1796);
not  g2623 (n2572, n1921);
not  g2624 (n2739, n2024);
buf  g2625 (n2753, n1967);
buf  g2626 (n3547, n2246);
buf  g2627 (n2422, n1829);
not  g2628 (n2870, n2305);
not  g2629 (n2930, n2224);
buf  g2630 (n2937, n1989);
not  g2631 (n2644, n1850);
buf  g2632 (n2604, n1225);
not  g2633 (n3097, n1912);
buf  g2634 (n2529, n1903);
buf  g2635 (n3150, n1993);
buf  g2636 (n3213, n2278);
not  g2637 (n2652, n2015);
buf  g2638 (n3151, n1802);
buf  g2639 (n2549, n2154);
buf  g2640 (n3017, n2274);
not  g2641 (n2625, n1800);
not  g2642 (n2483, n1731);
buf  g2643 (n3383, n1736);
not  g2644 (n2959, n1836);
buf  g2645 (n3111, n2202);
buf  g2646 (n3419, n2046);
buf  g2647 (n2844, n1904);
not  g2648 (n2944, n2157);
not  g2649 (n2826, n2301);
buf  g2650 (n3554, n1226);
not  g2651 (n2898, n1916);
not  g2652 (n3033, n1790);
buf  g2653 (n2402, n2223);
buf  g2654 (n2849, n2092);
not  g2655 (n2518, n1934);
not  g2656 (n3160, n1990);
buf  g2657 (n3378, n2296);
buf  g2658 (n3491, n1850);
buf  g2659 (n2824, n2304);
not  g2660 (n3132, n1984);
buf  g2661 (n3197, n2105);
buf  g2662 (n3289, n2044);
not  g2663 (n3525, n1851);
not  g2664 (n2969, n1812);
not  g2665 (n2351, n2131);
not  g2666 (n3372, n2284);
not  g2667 (n3050, n2033);
buf  g2668 (n3138, n2174);
not  g2669 (n2569, n2043);
not  g2670 (n3196, n2199);
not  g2671 (n2487, n1854);
buf  g2672 (n2378, n1997);
buf  g2673 (n2349, n2076);
not  g2674 (n2582, n2098);
not  g2675 (n3037, n2143);
buf  g2676 (n3485, n1835);
not  g2677 (n3497, n1761);
not  g2678 (n2335, n2197);
not  g2679 (n2783, n1818);
buf  g2680 (n3120, n1856);
not  g2681 (n2987, n2150);
not  g2682 (n3518, n2024);
not  g2683 (n2574, n2216);
buf  g2684 (n3251, n1984);
buf  g2685 (n2859, n2231);
not  g2686 (n2851, n1966);
buf  g2687 (n3144, n1828);
buf  g2688 (n3331, n2039);
buf  g2689 (n3047, n1926);
not  g2690 (n3149, n1915);
buf  g2691 (n2628, n1895);
buf  g2692 (n3108, n1978);
not  g2693 (n2520, n2281);
buf  g2694 (n3121, n2210);
not  g2695 (n2867, n1758);
not  g2696 (n2677, n2016);
not  g2697 (n2866, n2167);
not  g2698 (n2320, n1955);
not  g2699 (n2337, n1874);
not  g2700 (n2503, n2120);
buf  g2701 (n3352, n2190);
not  g2702 (n2306, n1965);
not  g2703 (n3514, n1919);
buf  g2704 (n2920, n2253);
buf  g2705 (n3188, n2021);
not  g2706 (n3229, n1798);
not  g2707 (n3483, n2155);
not  g2708 (n2307, n1916);
buf  g2709 (n2637, n1852);
not  g2710 (n3275, n1797);
buf  g2711 (n2971, n2270);
buf  g2712 (n3441, n2128);
not  g2713 (n2889, n1847);
not  g2714 (n2712, n2079);
buf  g2715 (n2499, n2211);
buf  g2716 (n2901, n2298);
buf  g2717 (n2742, n2168);
buf  g2718 (n2632, n2105);
buf  g2719 (n2612, n2170);
not  g2720 (n3100, n1900);
buf  g2721 (n3531, n1785);
not  g2722 (n2563, n1744);
buf  g2723 (n2846, n2267);
buf  g2724 (n3329, n2026);
buf  g2725 (n2958, n2028);
not  g2726 (n2333, n2206);
not  g2727 (n2784, n1747);
not  g2728 (n2787, n2089);
buf  g2729 (n3402, n2056);
not  g2730 (n2926, n2293);
buf  g2731 (n3141, n1766);
buf  g2732 (n3498, n1798);
buf  g2733 (n3542, n1872);
buf  g2734 (n2838, n2115);
not  g2735 (n2722, n2034);
not  g2736 (n3356, n1948);
not  g2737 (n3376, n2227);
buf  g2738 (n3308, n1913);
not  g2739 (n2490, n2206);
buf  g2740 (n2916, n2071);
not  g2741 (n3458, n2156);
not  g2742 (n3334, n1843);
not  g2743 (n2362, n1892);
not  g2744 (n2747, n2055);
buf  g2745 (n2741, n1946);
buf  g2746 (n2757, n2057);
not  g2747 (n3094, n2064);
buf  g2748 (n2418, n1919);
not  g2749 (n3293, n2266);
not  g2750 (n3472, n2223);
not  g2751 (n3346, n2164);
not  g2752 (n3367, n1858);
not  g2753 (n3076, n1755);
not  g2754 (n2392, n2280);
not  g2755 (n2797, n2120);
not  g2756 (n2972, n1843);
not  g2757 (n3504, n2240);
not  g2758 (n2358, n2291);
not  g2759 (n2372, n2008);
not  g2760 (n2404, n2282);
not  g2761 (n2945, n1998);
not  g2762 (n2751, n2009);
buf  g2763 (n2833, n2007);
buf  g2764 (n2639, n1939);
buf  g2765 (n2479, n1891);
buf  g2766 (n3315, n1963);
buf  g2767 (n3059, n2097);
buf  g2768 (n3227, n1929);
buf  g2769 (n2501, n2158);
buf  g2770 (n2540, n1896);
buf  g2771 (n3309, n2009);
buf  g2772 (n2999, n2003);
buf  g2773 (n2790, n2168);
not  g2774 (n2433, n1890);
buf  g2775 (n2936, n1985);
buf  g2776 (n2614, n1946);
not  g2777 (n3475, n1946);
buf  g2778 (n3416, n2010);
not  g2779 (n2627, n1804);
not  g2780 (n2502, n1983);
not  g2781 (n2566, n1911);
buf  g2782 (n3266, n1908);
buf  g2783 (n3028, n2131);
not  g2784 (n2929, n2126);
buf  g2785 (n2875, n2299);
not  g2786 (n3417, n1957);
not  g2787 (n2360, n1889);
not  g2788 (n3556, n1993);
buf  g2789 (n3249, n2179);
buf  g2790 (n2890, n1927);
buf  g2791 (n2393, n2281);
not  g2792 (n3093, n1980);
buf  g2793 (n2435, n2005);
buf  g2794 (n2530, n2009);
not  g2795 (n3360, n1947);
not  g2796 (n3320, n1803);
buf  g2797 (n2635, n1964);
not  g2798 (n2453, n2241);
not  g2799 (n3507, n1921);
buf  g2800 (n2347, n2252);
not  g2801 (n2915, n1952);
buf  g2802 (n3105, n2243);
buf  g2803 (n2727, n2211);
not  g2804 (n2616, n1738);
buf  g2805 (n2619, n2101);
not  g2806 (n2853, n1833);
buf  g2807 (n3375, n2170);
not  g2808 (n2650, n2302);
not  g2809 (n3283, n2083);
not  g2810 (n2671, n2222);
not  g2811 (n2564, n1849);
buf  g2812 (n3125, n2213);
not  g2813 (n3078, n2278);
not  g2814 (n3310, n2087);
not  g2815 (n2956, n1834);
not  g2816 (n3231, n2129);
buf  g2817 (n3092, n2171);
not  g2818 (n2447, n2036);
not  g2819 (n3044, n2239);
buf  g2820 (n3453, n2046);
buf  g2821 (n2446, n2249);
not  g2822 (n2687, n2215);
not  g2823 (n2642, n2286);
buf  g2824 (n3245, n2179);
buf  g2825 (n2610, n1999);
not  g2826 (n3232, n2067);
buf  g2827 (n2764, n2163);
not  g2828 (n3239, n2165);
not  g2829 (n2341, n2186);
not  g2830 (n2876, n2155);
buf  g2831 (n2454, n2063);
buf  g2832 (n2417, n2085);
not  g2833 (n3536, n2060);
not  g2834 (n3377, n1791);
not  g2835 (n3036, n2066);
not  g2836 (n3348, n1927);
buf  g2837 (n2863, n2302);
buf  g2838 (n2692, n1804);
not  g2839 (n3202, n2079);
buf  g2840 (n2570, n2027);
not  g2841 (n3456, n2191);
not  g2842 (n3317, n1797);
buf  g2843 (n2405, n2154);
not  g2844 (n3020, n2091);
buf  g2845 (n3147, n2233);
not  g2846 (n3075, n2208);
buf  g2847 (n3327, n2161);
not  g2848 (n3301, n2161);
buf  g2849 (n2346, n1830);
buf  g2850 (n2656, n2221);
not  g2851 (n2421, n1906);
buf  g2852 (n2345, n1770);
not  g2853 (n2781, n2214);
not  g2854 (n2592, n1914);
buf  g2855 (n3569, n2251);
not  g2856 (n2584, n2048);
not  g2857 (n2810, n2033);
not  g2858 (n3284, n2056);
not  g2859 (n2323, n1964);
buf  g2860 (n2596, n1821);
not  g2861 (n3486, n1754);
not  g2862 (n2526, n1884);
not  g2863 (n3064, n2169);
not  g2864 (n3199, n2163);
not  g2865 (n2679, n2228);
buf  g2866 (n3313, n1799);
not  g2867 (n2395, n1792);
not  g2868 (n3072, n1409);
not  g2869 (n2508, n2080);
buf  g2870 (n3316, n2238);
buf  g2871 (n2933, n1892);
buf  g2872 (n2460, n2044);
buf  g2873 (n2312, n2205);
buf  g2874 (n2455, n1864);
buf  g2875 (n2814, n2047);
not  g2876 (n3400, n2254);
buf  g2877 (n2996, n2042);
buf  g2878 (n3529, n2142);
buf  g2879 (n3476, n2240);
not  g2880 (n3081, n1854);
buf  g2881 (n2647, n1918);
buf  g2882 (n3210, n1997);
buf  g2883 (n2662, n2017);
not  g2884 (n3004, n2151);
buf  g2885 (n3179, n1801);
buf  g2886 (n3225, n2012);
not  g2887 (n2914, n1921);
not  g2888 (n3420, n2305);
buf  g2889 (n3540, n2043);
not  g2890 (n2823, n2053);
not  g2891 (n2667, n2012);
buf  g2892 (n3157, n1963);
buf  g2893 (n2736, n2129);
buf  g2894 (n2416, n1972);
not  g2895 (n3550, n1872);
not  g2896 (n2631, n2117);
buf  g2897 (n2324, n1815);
not  g2898 (n3450, n2117);
buf  g2899 (n3224, n1868);
not  g2900 (n3091, n2017);
buf  g2901 (n2629, n1925);
not  g2902 (n3466, n2300);
buf  g2903 (n2385, n2207);
not  g2904 (n2537, n2111);
not  g2905 (n3461, n1950);
not  g2906 (n2796, n2117);
buf  g2907 (n3380, n2078);
buf  g2908 (n2758, n2263);
not  g2909 (n2408, n2074);
buf  g2910 (n3305, n2072);
buf  g2911 (n3431, n2129);
buf  g2912 (n3169, n1990);
buf  g2913 (n3090, n1783);
buf  g2914 (n3513, n2256);
buf  g2915 (n2963, n2178);
not  g2916 (n3560, n1742);
not  g2917 (n3156, n1842);
not  g2918 (n2365, n2027);
buf  g2919 (n2670, n2011);
not  g2920 (n3517, n1939);
buf  g2921 (n2550, n2285);
buf  g2922 (n2989, n1751);
not  g2923 (n2655, n1909);
not  g2924 (n3074, n1224);
buf  g2925 (n3391, n2291);
not  g2926 (n2495, n2018);
not  g2927 (n2410, n1858);
not  g2928 (n2331, n1407);
buf  g2929 (n3347, n2118);
not  g2930 (n2583, n2001);
buf  g2931 (n3515, n2113);
not  g2932 (n2640, n1840);
not  g2933 (n2913, n1752);
buf  g2934 (n2522, n1780);
buf  g2935 (n3112, n1823);
buf  g2936 (n3110, n1968);
not  g2937 (n3071, n1962);
not  g2938 (n3083, n1975);
buf  g2939 (n2462, n1937);
buf  g2940 (n3527, n2192);
buf  g2941 (n2507, n2262);
buf  g2942 (n2732, n1855);
buf  g2943 (n3195, n1943);
not  g2944 (n3343, n2146);
buf  g2945 (n2717, n1763);
buf  g2946 (n2912, n2083);
not  g2947 (n2419, n2283);
not  g2948 (n3564, n1910);
not  g2949 (n3209, n1798);
not  g2950 (n3065, n2027);
not  g2951 (n2606, n2112);
buf  g2952 (n2862, n2227);
not  g2953 (n2954, n2245);
not  g2954 (n3166, n1981);
not  g2955 (n2726, n2204);
buf  g2956 (n2754, n2233);
buf  g2957 (n3226, n2228);
buf  g2958 (n3203, n2290);
buf  g2959 (n2376, n1759);
buf  g2960 (n3385, n1803);
not  g2961 (n2779, n1973);
not  g2962 (n2932, n2153);
not  g2963 (n2413, n2076);
buf  g2964 (n2988, n1910);
not  g2965 (n3173, n2283);
buf  g2966 (n3349, n2198);
buf  g2967 (n3354, n2067);
buf  g2968 (n3502, n2299);
buf  g2969 (n3006, n2007);
buf  g2970 (n3055, n2303);
buf  g2971 (n3369, n2241);
not  g2972 (n3207, n2178);
not  g2973 (n2439, n2253);
buf  g2974 (n3340, n1935);
buf  g2975 (n2661, n2150);
not  g2976 (n2982, n1837);
buf  g2977 (n2802, n2078);
buf  g2978 (n2370, n2272);
not  g2979 (n2415, n2085);
not  g2980 (n3311, n2109);
not  g2981 (n3355, n2235);
not  g2982 (n2469, n2192);
buf  g2983 (n3562, n2226);
not  g2984 (n3271, n2260);
not  g2985 (n2985, n1839);
not  g2986 (n2873, n1957);
not  g2987 (n3170, n2295);
not  g2988 (n2553, n1806);
buf  g2989 (n2778, n2047);
not  g2990 (n2638, n1941);
buf  g2991 (n2903, n2036);
buf  g2992 (n2330, n2064);
not  g2993 (n3493, n1977);
not  g2994 (n2383, n2035);
buf  g2995 (n2852, n1917);
buf  g2996 (n3049, n1939);
not  g2997 (n3228, n1948);
buf  g2998 (n2369, n1984);
not  g2999 (n2434, n1861);
buf  g3000 (n2544, n2104);
not  g3001 (n3494, n1801);
buf  g3002 (n3332, n2212);
buf  g3003 (n2352, n1893);
buf  g3004 (n2308, n1841);
buf  g3005 (n2947, n2198);
buf  g3006 (n3101, n1996);
buf  g3007 (n3126, n2138);
not  g3008 (n2334, n1804);
buf  g3009 (n2939, n1999);
buf  g3010 (n2902, n2024);
not  g3011 (n3374, n2044);
buf  g3012 (n2684, n2083);
not  g3013 (n2593, n2247);
not  g3014 (n3481, n2246);
buf  g3015 (n3303, n1892);
buf  g3016 (n2391, n2122);
buf  g3017 (n3338, n1965);
buf  g3018 (n2776, n1909);
buf  g3019 (n3363, n2201);
buf  g3020 (n2680, n2156);
buf  g3021 (n3031, n1929);
not  g3022 (n2407, n1814);
buf  g3023 (n3429, n1936);
not  g3024 (n2716, n2167);
not  g3025 (n3175, n2265);
not  g3026 (n3163, n1969);
buf  g3027 (n2827, n2288);
not  g3028 (n3522, n1859);
buf  g3029 (n2554, n2146);
not  g3030 (n2399, n1789);
buf  g3031 (n2380, n1991);
buf  g3032 (n3373, n2025);
not  g3033 (n3365, n1738);
buf  g3034 (n2807, n1850);
buf  g3035 (n2528, n1861);
buf  g3036 (n2746, n2201);
buf  g3037 (n2906, n1940);
not  g3038 (n2547, n2055);
buf  g3039 (n2675, n1952);
buf  g3040 (n2368, n1791);
buf  g3041 (n2560, n2163);
buf  g3042 (n3136, n1910);
not  g3043 (n2819, n1895);
not  g3044 (n3413, n2214);
not  g3045 (n2382, n2286);
buf  g3046 (n3273, n1937);
buf  g3047 (n2339, n2068);
not  g3048 (n3261, n2065);
not  g3049 (n2782, n1753);
buf  g3050 (n2493, n2073);
not  g3051 (n3260, n1899);
not  g3052 (n2355, n2080);
not  g3053 (n2542, n2050);
buf  g3054 (n3448, n1806);
buf  g3055 (n3473, n2084);
buf  g3056 (n3019, n1824);
not  g3057 (n2310, n1943);
buf  g3058 (n2793, n2294);
buf  g3059 (n2514, n2174);
buf  g3060 (n2406, n1844);
not  g3061 (n3131, n1881);
buf  g3062 (n3545, n1935);
buf  g3063 (n3164, n1874);
buf  g3064 (n3205, n2159);
buf  g3065 (n3452, n1834);
not  g3066 (n3433, n1788);
not  g3067 (n3025, n2269);
buf  g3068 (n2934, n1875);
buf  g3069 (n2579, n1782);
buf  g3070 (n2621, n2162);
buf  g3071 (n2363, n2177);
not  g3072 (n3424, n2108);
not  g3073 (n3325, n2025);
not  g3074 (n2734, n2107);
not  g3075 (n3333, n1977);
buf  g3076 (n3395, n2175);
buf  g3077 (n2927, n2176);
not  g3078 (n3551, n2116);
not  g3079 (n3060, n1919);
buf  g3080 (n3061, n1743);
not  g3081 (n2685, n2089);
buf  g3082 (n2371, n2243);
buf  g3083 (n3364, n1815);
buf  g3084 (n2577, n2279);
not  g3085 (n3234, n2284);
buf  g3086 (n3295, n2259);
not  g3087 (n2475, n1994);
not  g3088 (n2953, n2225);
not  g3089 (n2598, n2111);
buf  g3090 (n2740, n2039);
buf  g3091 (n2917, n1920);
buf  g3092 (n2681, n2278);
not  g3093 (n3177, n1866);
buf  g3094 (n2811, n2116);
not  g3095 (n2651, n2103);
buf  g3096 (n2552, n1907);
not  g3097 (n3384, n2195);
not  g3098 (n3537, n2257);
buf  g3099 (n3018, n2110);
buf  g3100 (n2387, n2223);
not  g3101 (n2763, n1812);
not  g3102 (n3252, n2184);
not  g3103 (n3220, n1875);
buf  g3104 (n3276, n2296);
not  g3105 (n2975, n1913);
buf  g3106 (n2835, n2181);
buf  g3107 (n2649, n1808);
not  g3108 (n2729, n2235);
not  g3109 (n2477, n1822);
buf  g3110 (n2886, n1405);
buf  g3111 (n2458, n2101);
not  g3112 (n2543, n2242);
not  g3113 (n2702, n1811);
not  g3114 (n3435, n2060);
buf  g3115 (n3371, n1828);
buf  g3116 (n3443, n2038);
not  g3117 (n2938, n1815);
not  g3118 (n3005, n2128);
buf  g3119 (n3000, n2059);
buf  g3120 (n3559, n1843);
not  g3121 (n2834, n2285);
buf  g3122 (n3471, n2234);
not  g3123 (n2847, n2093);
not  g3124 (n2883, n2037);
buf  g3125 (n3506, n2289);
buf  g3126 (n3388, n2069);
buf  g3127 (n2473, n1909);
buf  g3128 (n3069, n2175);
not  g3129 (n3027, n2144);
not  g3130 (n3503, n2068);
buf  g3131 (n2403, n1979);
buf  g3132 (n3319, n2143);
buf  g3133 (n2885, n1934);
buf  g3134 (n2942, n1885);
not  g3135 (n3259, n2261);
buf  g3136 (n2322, n1981);
not  g3137 (n3482, n1773);
not  g3138 (n3247, n2177);
not  g3139 (n2682, n2196);
not  g3140 (n3161, n1949);
buf  g3141 (n3135, n1794);
buf  g3142 (n3098, n2086);
not  g3143 (n3079, n1903);
buf  g3144 (n2983, n1775);
not  g3145 (n2723, n2186);
buf  g3146 (n3558, n1864);
buf  g3147 (n2694, n2273);
buf  g3148 (n2484, n2276);
buf  g3149 (n3029, n1854);
buf  g3150 (n3511, n2075);
not  g3151 (n2519, n1797);
buf  g3152 (n3490, n2181);
not  g3153 (n2794, n1920);
not  g3154 (n3265, n2247);
buf  g3155 (n2377, n2141);
not  g3156 (n3563, n1765);
buf  g3157 (n3128, n2033);
not  g3158 (n2986, n2087);
buf  g3159 (n2831, n1836);
buf  g3160 (n2485, n1110);
not  g3161 (n2894, n2158);
not  g3162 (n2713, n1932);
not  g3163 (n2998, n1806);
buf  g3164 (n3230, n2038);
buf  g3165 (n2327, n2197);
buf  g3166 (n3200, n2119);
not  g3167 (n2884, n2070);
not  g3168 (n3510, n2216);
buf  g3169 (n2786, n2277);
not  g3170 (n2858, n2197);
not  g3171 (n2772, n1888);
buf  g3172 (n2646, n2268);
not  g3173 (n3178, n1785);
not  g3174 (n3422, n2244);
not  g3175 (n2357, n1966);
not  g3176 (n2580, n2230);
buf  g3177 (n3236, n2180);
buf  g3178 (n3211, n2260);
buf  g3179 (n3393, n2250);
not  g3180 (n2992, n2234);
buf  g3181 (n2830, n2200);
not  g3182 (n3206, n1955);
not  g3183 (n3107, n1747);
buf  g3184 (n3500, n1793);
not  g3185 (n3389, n1793);
not  g3186 (n2587, n2250);
not  g3187 (n2600, n1796);
buf  g3188 (n2465, n1837);
buf  g3189 (n3530, n2140);
buf  g3190 (n2770, n2122);
not  g3191 (n3526, n2102);
not  g3192 (n2724, n2289);
not  g3193 (n2850, n2138);
buf  g3194 (n3012, n2201);
buf  g3195 (n3571, n1947);
not  g3196 (n2935, n2153);
buf  g3197 (n3067, n2061);
buf  g3198 (n2459, n2088);
not  g3199 (n2788, n1989);
not  g3200 (n3421, n1403);
buf  g3201 (n2800, n1845);
buf  g3202 (n3495, n1841);
buf  g3203 (n3089, n1855);
not  g3204 (n3180, n1900);
buf  g3205 (n3122, n1956);
buf  g3206 (n2970, n2214);
buf  g3207 (n2532, n2282);
buf  g3208 (n2506, n1860);
buf  g3209 (n2516, n2303);
not  g3210 (n3015, n2172);
buf  g3211 (n3278, n1807);
not  g3212 (n3192, n1839);
buf  g3213 (n2911, n2203);
buf  g3214 (n3557, n1799);
buf  g3215 (n2966, n1935);
not  g3216 (n2909, n1963);
buf  g3217 (n3241, n2106);
not  g3218 (n3405, n2023);
buf  g3219 (n3039, n2013);
xnor g3220 (n3379, n1835, n1861, n2133);
or   g3221 (n3133, n1783, n2165, n2118, n1986);
xor  g3222 (n2854, n1826, n2019, n2087, n2103);
xor  g3223 (n2855, n1857, n1985, n1867, n1742);
and  g3224 (n3534, n1936, n2296, n2239, n2266);
nand g3225 (n2864, n1979, n1873, n2045, n1823);
and  g3226 (n2313, n2102, n2096, n2126, n2189);
nand g3227 (n2396, n2010, n2247, n2287, n2286);
xnor g3228 (n3366, n1917, n1771, n1851, n2259);
nor  g3229 (n3162, n1820, n1918, n2166, n1799);
nand g3230 (n2350, n2079, n1817, n1875, n1800);
and  g3231 (n3568, n1957, n2112, n1953, n1822);
nor  g3232 (n2980, n1976, n1945, n2288, n2135);
and  g3233 (n2597, n1837, n2240, n2261, n2022);
or   g3234 (n3478, n1994, n2275, n2095, n2078);
and  g3235 (n2617, n1896, n2211, n1941, n1993);
nor  g3236 (n2534, n2125, n2097, n2052, n2288);
nand g3237 (n2452, n2258, n2209, n1968, n2235);
xnor g3238 (n2414, n1406, n1823, n1979, n2180);
xnor g3239 (n3544, n1784, n2017, n1842, n1730);
xor  g3240 (n2871, n1966, n1856, n2300, n2065);
xor  g3241 (n3194, n2149, n1816, n1901, n1786);
and  g3242 (n3095, n2217, n2042, n1914, n2273);
nor  g3243 (n2887, n2018, n2216, n2176, n2232);
and  g3244 (n3240, n2175, n1734, n2088, n1994);
xor  g3245 (n3086, n1962, n2072, n2021, n2304);
or   g3246 (n3296, n1869, n2265, n2025, n2258);
and  g3247 (n2573, n2246, n2248, n2138, n1935);
or   g3248 (n2561, n1905, n1785, n1918, n2028);
xor  g3249 (n2775, n2102, n2002, n2139, n1958);
nor  g3250 (n2809, n1809, n1743, n2280, n2248);
and  g3251 (n2511, n1406, n1954, n1797, n2221);
nand g3252 (n3499, n2138, n1970, n2136, n2124);
xnor g3253 (n3361, n2072, n2239, n2162, n1895);
nand g3254 (n2733, n2151, n2247, n2176, n2118);
nor  g3255 (n3286, n1998, n1786, n2043, n2074);
and  g3256 (n2821, n2082, n1853, n2194, n2145);
nor  g3257 (n3184, n1225, n2037, n2154, n1880);
nand g3258 (n3046, n2145, n2149, n1840, n1996);
or   g3259 (n3042, n2064, n1948, n2103, n1953);
xor  g3260 (n2603, n2110, n2153, n1942, n2016);
nor  g3261 (n3088, n2236, n1862, n1902, n2021);
nor  g3262 (n3351, n1992, n1822, n2142, n2173);
nor  g3263 (n3277, n1969, n2110, n1985, n1825);
and  g3264 (n3168, n2196, n2194, n1810, n2127);
and  g3265 (n3003, n1919, n2287, n1735, n1903);
xnor g3266 (n3038, n2039, n2023, n2299, n2099);
nor  g3267 (n3148, n2143, n2236, n2125, n2203);
and  g3268 (n2504, n2114, n2273, n2280, n2294);
or   g3269 (n3446, n2027, n2100, n2302, n2172);
nand g3270 (n3054, n1860, n1760, n2268, n1788);
xor  g3271 (n2314, n2217, n1973, n2220, n1931);
xor  g3272 (n2714, n1741, n1754, n2224, n1971);
and  g3273 (n2785, n2092, n2062, n1855, n1980);
or   g3274 (n3350, n2053, n1838, n1845, n1882);
xor  g3275 (n3401, n1986, n2218, n2150, n1817);
nor  g3276 (n2524, n1938, n1979, n2118, n1768);
nand g3277 (n2706, n1782, n1764, n2086, n2112);
nand g3278 (n2653, n2188, n1813, n1832, n2094);
nor  g3279 (n3274, n2001, n1982, n1762, n2291);
and  g3280 (n3218, n2276, n2137, n2151, n2054);
and  g3281 (n3455, n1923, n2254, n1904, n1112);
xor  g3282 (n2321, n1794, n1733, n2213, n1846);
and  g3283 (n2691, n1889, n2037, n2196, n2256);
nor  g3284 (n2412, n1933, n1993, n1862, n2016);
and  g3285 (n2546, n1768, n1986, n1745, n2275);
nor  g3286 (n3459, n2286, n1930, n1789, n1886);
and  g3287 (n3565, n1933, n2219, n2304, n2276);
nor  g3288 (n2708, n2054, n2095, n2064, n1834);
nor  g3289 (n2839, n1952, n2239, n2106, n1898);
xor  g3290 (n2481, n2075, n2103, n1876, n2070);
xnor g3291 (n2329, n1819, n1894, n1780, n1845);
nor  g3292 (n3026, n2022, n2101, n2140, n1880);
or   g3293 (n2900, n2092, n1813, n2200, n2255);
nor  g3294 (n2801, n2164, n2051, n1931, n2074);
nand g3295 (n2601, n2085, n2252, n2257, n2148);
nor  g3296 (n3193, n1930, n2061, n2026, n2250);
xnor g3297 (n3181, n2245, n1787, n1833, n2065);
xor  g3298 (n3190, n1865, n1752, n1868, n1890);
xor  g3299 (n3256, n2014, n2299, n2244, n2100);
xor  g3300 (n2431, n2179, n1801, n2227, n1904);
nand g3301 (n3573, n1808, n1776, n2301, n2060);
or   g3302 (n2536, n2001, n1807, n2305, n2298);
or   g3303 (n2948, n1408, n1841, n1912, n1991);
or   g3304 (n2332, n1951, n2209, n2028, n2171);
nand g3305 (n2599, n1891, n1871, n2105, n1975);
nand g3306 (n2857, n2059, n1872, n2173, n2174);
nor  g3307 (n3238, n1402, n1949, n2265, n2185);
xor  g3308 (n2535, n2066, n1921, n1913, n2049);
xor  g3309 (n3460, n2000, n2219, n1827, n2031);
nand g3310 (n2976, n2210, n2035, n2071, n1405);
nand g3311 (n2602, n1809, n2269, n1881, n2073);
xnor g3312 (n2893, n1849, n2202, n2068, n2073);
nand g3313 (n2880, n2221, n1978, n2295, n2282);
xnor g3314 (n2663, n1820, n2295, n2045, n1922);
xnor g3315 (n2750, n1924, n2105, n2035, n2206);
xnor g3316 (n2539, n2246, n1964, n1841, n1959);
and  g3317 (n3335, n1748, n1842, n2081, n2020);
or   g3318 (n3463, n2134, n1996, n1811, n1971);
or   g3319 (n2905, n2157, n2050, n2259, n1923);
xnor g3320 (n2411, n1734, n1942, n1878, n1867);
or   g3321 (n3208, n2157, n2093, n1906, n2095);
and  g3322 (n3014, n2113, n2249, n2251, n2261);
xnor g3323 (n3434, n1891, n2084, n2141, n2230);
and  g3324 (n2955, n1922, n1889, n2225, n1746);
xnor g3325 (n3279, n2076, n1878, n1846, n2144);
nand g3326 (n3009, n2275, n2131, n2005, n2033);
xnor g3327 (n3324, n2070, n1792, n1958, n2200);
xor  g3328 (n3304, n2125, n2065, n1838, n2240);
or   g3329 (n2931, n2098, n2114, n1774, n1894);
xor  g3330 (n3248, n1809, n2271, n2295, n2030);
nand g3331 (n3454, n2137, n2149, n2147, n1942);
and  g3332 (n3143, n1951, n1911, n2188, n2069);
or   g3333 (n3023, n2229, n1888, n1795, n1862);
and  g3334 (n2995, n1879, n2070, n1405, n1898);
or   g3335 (n3073, n1825, n2119, n2271, n2005);
or   g3336 (n2457, n1749, n1817, n1947, n2267);
nor  g3337 (n2389, n1969, n1834, n1795, n2277);
or   g3338 (n2765, n1938, n2116, n2183, n2207);
nor  g3339 (n3509, n2049, n1839, n1884, n1823);
nor  g3340 (n3523, n2237, n1873, n2215, n1949);
nor  g3341 (n2964, n1949, n1963, n1859, n1956);
or   g3342 (n2674, n2207, n2092, n2108, n2021);
nor  g3343 (n3263, n2255, n2178, n1877, n1893);
or   g3344 (n2780, n2022, n1932, n2287, n1891);
nand g3345 (n2879, n1978, n1778, n2056, n1857);
xnor g3346 (n2730, n1924, n2187, n2183, n1981);
xnor g3347 (n2822, n1830, n1886, n2006, n1887);
nor  g3348 (n3001, n2235, n2279, n2137, n2224);
xnor g3349 (n2877, n2292, n2020, n1897, n2113);
xnor g3350 (n2777, n1842, n2099, n1960, n2054);
nand g3351 (n3344, n2212, n1903, n2087, n2277);
nor  g3352 (n2658, n1941, n1900, n1753, n1402);
nor  g3353 (n3574, n1870, n1848, n2015, n2298);
xor  g3354 (n3139, n1735, n2048, n2126, n1975);
xnor g3355 (n3553, n2199, n1962, n1885, n2182);
or   g3356 (n3415, n2123, n1960, n2289, n1869);
xor  g3357 (n2721, n1970, n2171, n1790, n2182);
nand g3358 (n3444, n1767, n2032, n1884, n2256);
xnor g3359 (n3399, n1825, n2132, n1984, n1882);
nand g3360 (n2665, n2088, n2275, n1767, n1998);
xor  g3361 (n2967, n2258, n2201, n1868, n2290);
nor  g3362 (n2586, n2154, n2041, n2243, n1983);
xor  g3363 (n3287, n1853, n1786, n2090, n2009);
xnor g3364 (n2946, n2109, n2143, n1409, n1896);
xor  g3365 (n3496, n2226, n1858, n2243, n2231);
xnor g3366 (n2611, n2130, n1885, n1873, n2045);
or   g3367 (n3292, n2140, n2230, n2099, n1976);
or   g3368 (n3118, n1805, n2030, n1748, n2214);
xnor g3369 (n2923, n2165, n1407, n1838, n2198);
and  g3370 (n2340, n1863, n2128, n2044, n2199);
nand g3371 (n2664, n2242, n1936, n2175, n2279);
and  g3372 (n3212, n1757, n2058, n2202, n2229);
nand g3373 (n3407, n2077, n1822, n2293, n1859);
xnor g3374 (n2756, n1870, n2287, n1925, n1937);
xor  g3375 (n3397, n2304, n2190, n1999, n2177);
xor  g3376 (n2660, n1406, n2002, n2283, n2058);
xnor g3377 (n3130, n2161, n1923, n2109, n1751);
and  g3378 (n2648, n2152, n1962, n1910, n2135);
or   g3379 (n2354, n2057, n2204, n1890, n2205);
nand g3380 (n2766, n1906, n1900, n2091, n1816);
and  g3381 (n2565, n1995, n2052, n2260, n2255);
xnor g3382 (n2548, n2209, n2007, n1965, n1409);
and  g3383 (n3152, n2090, n1762, n2220, n1961);
and  g3384 (n2977, n1976, n1905, n1866, n2292);
or   g3385 (n2921, n2190, n1858, n2002, n1844);
xor  g3386 (n2471, n2041, n1784, n1865, n1790);
xnor g3387 (n3411, n2230, n1873, n1879, n2165);
or   g3388 (n2356, n2185, n2172, n1802, n2203);
nor  g3389 (n2961, n1840, n1801, n2209, n2166);
xnor g3390 (n3539, n2259, n1901, n2051, n1982);
and  g3391 (n3158, n2241, n1934, n1786, n1874);
or   g3392 (n2348, n1908, n1890, n1827, n2268);
xnor g3393 (n2718, n1953, n2147, n1850, n2262);
nand g3394 (n3566, n2104, n1865, n2234, n2272);
xor  g3395 (n2907, n2119, n1225, n1955, n1731);
nand g3396 (n2804, n2270, n2008, n1840, n2164);
xor  g3397 (n2645, n1771, n2019, n1781, n2218);
xor  g3398 (n2908, n2160, n2055, n1970, n1997);
xnor g3399 (n2841, n2250, n2155, n1960, n1795);
xor  g3400 (n2623, n1892, n2015, n2185, n1820);
and  g3401 (n2448, n2168, n2127, n2013, n2077);
or   g3402 (n3521, n2232, n2227, n2156, n1897);
nor  g3403 (n3124, n2046, n1958, n1980, n1798);
and  g3404 (n2795, n2008, n2232, n2124, n1860);
nand g3405 (n3187, n2292, n2158, n2197, n1826);
xor  g3406 (n3387, n1959, n1870, n1749, n1852);
xnor g3407 (n2828, n1770, n1807, n1763, n2078);
xor  g3408 (n3137, n2257, n1867, n1732, n2104);
xor  g3409 (n3520, n2071, n2174, n1932, n1987);
and  g3410 (n2896, n2093, n2248, n2226, n2200);
xnor g3411 (n3447, n1943, n2146, n1862, n1811);
nor  g3412 (n2698, n1777, n1983, n2047, n2036);
nor  g3413 (n2943, n1404, n1952, n1991, n1759);
xor  g3414 (n2578, n2193, n2191, n2058, n2079);
xnor g3415 (n2843, n2234, n1817, n1803, n2268);
xor  g3416 (n3146, n1773, n2115, n2054, n2123);
or   g3417 (n2738, n1907, n1930, n1792, n1405);
nand g3418 (n2634, n2172, n2020, n1997, n1824);
and  g3419 (n3134, n1746, n1224, n1805, n1884);
xor  g3420 (n2709, n1956, n1904, n2038, n2292);
xor  g3421 (n3524, n2218, n1813, n2131, n2130);
nor  g3422 (n2555, n2040, n2219, n2025, n1876);
xor  g3423 (n2699, n1859, n2006, n2058, n1789);
xnor g3424 (n3297, n1847, n1902, n1812, n1998);
xor  g3425 (n2773, n2195, n1846, n2063, n2134);
xor  g3426 (n2949, n2303, n1831, n1807, n2122);
xnor g3427 (n2588, n1883, n1980, n2134, n2109);
or   g3428 (n2899, n2297, n2011, n2022, n1835);
nor  g3429 (n2527, n2106, n2075, n1844, n2301);
xor  g3430 (n2559, n2045, n1932, n2110, n2262);
and  g3431 (n2500, n2264, n2011, n1897, n2226);
or   g3432 (n2343, n2081, n1954, n2191, n2139);
and  g3433 (n2571, n1880, n2263, n1796, n2056);
or   g3434 (n3048, n1737, n1969, n2285, n2162);
xor  g3435 (n3548, n1928, n1820, n1886, n2236);
nor  g3436 (n3214, n1911, n1883, n1758, n2291);
nor  g3437 (n3171, n2133, n1816, n2288, n2217);
xnor g3438 (n2882, n2145, n2242, n2061, n1861);
xor  g3439 (n2394, n1766, n1964, n1864, n1877);
and  g3440 (n2979, n2183, n1866, n2094, n1916);
xnor g3441 (n2476, n1814, n1934, n1854, n1955);
and  g3442 (n3410, n2089, n2013, n1853, n1926);
nor  g3443 (n3306, n2289, n1772, n1789, n1781);
or   g3444 (n2767, n1788, n2187, n1945, n1957);
xor  g3445 (n3034, n2091, n2216, n1832, n2040);
xor  g3446 (n2498, n2107, n1810, n1806, n2030);
xnor g3447 (n3002, n1818, n2097, n1999, n2198);
or   g3448 (n3056, n2171, n2007, n2001, n2184);
nor  g3449 (n2836, n2223, n1855, n1814, n2251);
xnor g3450 (n2865, n2052, n1774, n2062, n1403);
and  g3451 (n2704, n2053, n1958, n1945, n2202);
nor  g3452 (n3538, n2156, n2081, n2260, n1825);
xor  g3453 (n3219, n1791, n2047, n2293, n2094);
nor  g3454 (n2710, n1874, n2261, n2208, n2147);
xor  g3455 (n3427, n2211, n1847, n1925, n1927);
xor  g3456 (n3298, n1856, n2168, n1865, n2137);
nor  g3457 (n3032, n1800, n1868, n1794, n1814);
or   g3458 (n3423, n1845, n1739, n1877, n1936);
nand g3459 (n2748, n2241, n2285, n2237, n2104);
or   g3460 (n2325, n2091, n1893, n1950, n2106);
xnor g3461 (n3409, n1851, n2086, n2228, n2183);
xnor g3462 (n2978, n2253, n1795, n2194, n1839);
nor  g3463 (n3312, n2081, n1772, n2164, n1837);
xnor g3464 (n2984, n1829, n2076, n1869, n1887);
xor  g3465 (n2373, n1808, n1847, n1905, n1951);
nand g3466 (n2878, n2051, n2182, n1974, n2166);
and  g3467 (n3116, n1779, n2192, n1872, n2115);
nor  g3468 (n2492, n2267, n2100, n2176, n1898);
nor  g3469 (n2318, n1902, n1912, n2032, n1971);
xor  g3470 (n2482, n2108, n2083, n2034, n2150);
and  g3471 (n3508, n1737, n2132, n2255, n2264);
nor  g3472 (n2745, n1740, n2272, n1810, n2153);
and  g3473 (n2478, n1888, n1881, n2220, n1938);
and  g3474 (n2488, n2014, n2237, n1819, n1876);
nand g3475 (n2990, n2052, n2061, n2190, n1777);
and  g3476 (n2474, n2088, n1947, n2237, n2193);
xor  g3477 (n3186, n2116, n1986, n1809, n1764);
xnor g3478 (n3575, n1778, n1922, n2048, n2252);
xor  g3479 (n2594, n1821, n1967, n1808, n2193);
xor  g3480 (n3430, n2276, n1828, n2212, n1987);
nand g3481 (n2633, n2157, n2100, n2142, n2102);
xnor g3482 (n2608, n2032, n2182, n2264, n1836);
or   g3483 (n3257, n2279, n1857, n1883, n1989);
or   g3484 (n3288, n2004, n1741, n2026, n2229);
nand g3485 (n2486, n1811, n2274, n2107, n1881);
xnor g3486 (n3477, n2086, n2284, n2218, n1835);
nand g3487 (n2672, n2038, n2266, n2098, n2122);
and  g3488 (n2728, n1922, n1863, n1815, n1973);
and  g3489 (n2668, n2269, n1760, n1800, n2010);
nor  g3490 (n3119, n2020, n1905, n2191, n1968);
nor  g3491 (n3155, n1989, n2069, n2037, n1849);
nor  g3492 (n3457, n1953, n1976, n2034, n2244);
or   g3493 (n2798, n1924, n2113, n2012, n1907);
nor  g3494 (n3270, n2231, n2050, n1836, n2049);
nor  g3495 (n2364, n2294, n1893, n1879, n2090);
and  g3496 (n2440, n1959, n1888, n1821, n2217);
nand g3497 (n2468, n1824, n2011, n2034, n2263);
xor  g3498 (n2538, n1978, n2042, n1831, n2085);
and  g3499 (n3314, n1406, n2297, n1968, n2066);
and  g3500 (n2512, n2180, n2115, n1928, n2135);
nand g3501 (n2443, n1988, n1852, n2005, n1857);
xnor g3502 (n3362, n2112, n2062, n2035, n2204);
xnor g3503 (n3007, n2120, n2136, n2029, n1756);
nor  g3504 (n3217, n1882, n1982, n2139, n2283);
nor  g3505 (n3339, n2071, n2254, n1846, n1109);
xor  g3506 (n3013, n1938, n1785, n1966, n2251);
xor  g3507 (n3408, n2281, n1991, n2173, n2151);
nand g3508 (n3445, n2233, n2041, n2062, n1830);
nor  g3509 (n2576, n2210, n1928, n2161, n1404);
xnor g3510 (n3221, n1940, n2152, n2123, n2006);
xor  g3511 (n2438, n2205, n1943, n1929, n2148);
xnor g3512 (n2997, n2222, n2188, n1769, n1994);
nand g3513 (n3215, n1793, n2040, n2029, n1803);
xor  g3514 (n2817, n2187, n1819, n2018, n1870);
nor  g3515 (n3532, n2277, n2057, n2177, n2160);
xnor g3516 (n2812, n1909, n2169, n2273, n2084);
xnor g3517 (n3024, n1928, n1794, n2205, n2050);
or   g3518 (n2568, n1832, n2094, n2290, n1913);
xor  g3519 (n2636, n2162, n2051, n1844, n1779);
nand g3520 (n3432, n2010, n2274, n2133, n2305);
xnor g3521 (n2326, n1852, n1744, n1831, n2159);
nand g3522 (n2832, n2006, n2067, n2012, n1750);
or   g3523 (n3512, n1950, n1108, n1975, n2084);
xor  g3524 (n3505, n1826, n1863, n2271, n2119);
xnor g3525 (n2919, n1799, n2040, n2166, n2238);
or   g3526 (n2463, n1824, n2281, n2026, n2173);
xor  g3527 (n3022, n1765, n1914, n2170, n2194);
xnor g3528 (n3129, n2207, n1973, n2245, n1897);
xor  g3529 (n3258, n2080, n2238, n2041, n2213);
nor  g3530 (n3191, n1403, n1974, n2222, n2014);
xnor g3531 (n2731, n1827, n1788, n1736, n2152);
xor  g3532 (n2928, n2132, n2296, n2236, n2000);
nand g3533 (n2815, n1833, n2186, n1899, n1946);
xor  g3534 (n3353, n2003, n2252, n1775, n1863);
xnor g3535 (n3464, n1878, n1887, n1871, n1917);
or   g3536 (n2374, n1831, n2142, n1992, n2248);
xnor g3537 (n3063, n2178, n2074, n1756, n2160);
xnor g3538 (n3552, n1985, n1833, n2144, n2121);
nor  g3539 (n3440, n2262, n2187, n1954, n1930);
and  g3540 (n3467, n2302, n1925, n1982, n2145);
xnor g3541 (n2707, n1916, n1996, n2233, n2031);
xor  g3542 (n3414, n2147, n1791, n1974, n1408);
xnor g3543 (n3715, n3374, n3218, n2711, n2646);
and  g3544 (n3652, n2957, n3192, n3152, n2576);
nor  g3545 (n3825, n3029, n2455, n3131, n2444);
nor  g3546 (n3802, n3187, n3115, n2969, n3012);
xor  g3547 (n3824, n3276, n3318, n3081, n3288);
xnor g3548 (n3601, n2530, n2650, n2440, n2602);
nand g3549 (n3650, n2840, n2490, n2565, n2975);
nand g3550 (n3744, n2731, n2500, n2984, n2314);
xnor g3551 (n3737, n2591, n3369, n3051, n3170);
or   g3552 (n3816, n2473, n2360, n2666, n3172);
or   g3553 (n3663, n625, n2846, n3100, n2637);
or   g3554 (n3752, n3281, n3353, n2985, n3196);
xnor g3555 (n3591, n3212, n2799, n2729, n2364);
xor  g3556 (n3749, n2395, n2325, n3213, n2393);
xnor g3557 (n3603, n2789, n2959, n3362, n2371);
xor  g3558 (n3739, n2970, n2811, n3347, n3105);
and  g3559 (n3581, n2622, n2806, n2588, n2605);
or   g3560 (n3777, n3193, n3195, n3252, n3366);
nor  g3561 (n3803, n3054, n2404, n2768, n2735);
nor  g3562 (n3799, n2887, n3207, n2410, n2706);
xnor g3563 (n3643, n2869, n2829, n2815, n2408);
and  g3564 (n3639, n2837, n2313, n2720, n3214);
or   g3565 (n3645, n2770, n2485, n2931, n2457);
xor  g3566 (n3771, n2425, n3200, n3136, n2403);
and  g3567 (n3784, n2898, n3215, n3056, n3246);
xor  g3568 (n3583, n2648, n2849, n3120, n2863);
nor  g3569 (n3659, n3117, n2709, n2871, n2551);
nor  g3570 (n3822, n2361, n2600, n2934, n2704);
nor  g3571 (n3634, n2651, n3098, n2665, n2780);
and  g3572 (n3655, n2385, n2357, n3072, n2818);
and  g3573 (n3718, n2702, n2306, n2868, n3166);
or   g3574 (n3719, n2794, n3021, n2430, n3287);
xor  g3575 (n3750, n3150, n2564, n2582, n3317);
or   g3576 (n3665, n2899, n2906, n2921, n3080);
xor  g3577 (n3690, n2628, n3335, n2426, n2762);
xor  g3578 (n3658, n2427, n2642, n3352, n3043);
or   g3579 (n3769, n3359, n2981, n625, n2675);
or   g3580 (n3689, n2351, n2459, n2561, n3239);
or   g3581 (n3606, n3241, n3129, n3074, n3387);
and  g3582 (n3697, n2534, n2420, n3206, n2539);
and  g3583 (n3654, n3046, n2626, n2330, n2381);
nor  g3584 (n3732, n2315, n2874, n2634, n3154);
nand g3585 (n3811, n2765, n2388, n2496, n3248);
or   g3586 (n3790, n2980, n3173, n3107, n3175);
nand g3587 (n3660, n2544, n3000, n2912, n2323);
and  g3588 (n3832, n2986, n2919, n2320, n2932);
and  g3589 (n3806, n3020, n3044, n2476, n2669);
xor  g3590 (n3704, n3119, n2629, n3284, n2880);
nor  g3591 (n3836, n2453, n2469, n3083, n3132);
xor  g3592 (n3743, n3004, n2813, n2715, n2807);
nand g3593 (n3599, n2690, n2826, n3094, n3176);
xnor g3594 (n3683, n2830, n2960, n3073, n3373);
xor  g3595 (n3741, n3314, n2595, n2992, n3025);
and  g3596 (n3835, n2358, n3121, n2758, n3104);
and  g3597 (n3681, n2858, n2487, n2533, n3033);
or   g3598 (n3696, n2432, n3270, n3112, n2713);
xnor g3599 (n3782, n2434, n2667, n2621, n3199);
xor  g3600 (n3623, n3090, n2525, n3310, n2707);
or   g3601 (n3585, n2643, n2925, n2601, n3194);
xor  g3602 (n3600, n3035, n3363, n2892, n3086);
nand g3603 (n3612, n2394, n2499, n2831, n3222);
and  g3604 (n3805, n2865, n3165, n2955, n2538);
and  g3605 (n3778, n2732, n2619, n2982, n2311);
xor  g3606 (n3589, n2705, n3266, n3267, n2749);
xor  g3607 (n3667, n3065, n2573, n3336, n2333);
nor  g3608 (n3789, n2687, n3343, n2821, n2583);
or   g3609 (n3843, n2350, n3296, n2479, n3082);
nor  g3610 (n3598, n2372, n3042, n2618, n3227);
and  g3611 (n3796, n2436, n2861, n3377, n2775);
or   g3612 (n3605, n3245, n2703, n3340, n2719);
nor  g3613 (n3578, n2519, n2673, n2378, n3014);
or   g3614 (n3619, n3240, n2342, n3174, n3124);
xnor g3615 (n3620, n3303, n2961, n3308, n2545);
xnor g3616 (n3726, n2805, n2498, n2615, n3371);
nand g3617 (n3767, n3251, n2438, n2741, n3208);
nand g3618 (n3635, n3226, n2407, n3069, n3143);
nand g3619 (n3730, n3280, n3095, n2839, n2700);
or   g3620 (n3691, n2645, n2461, n2978, n3238);
nor  g3621 (n3703, n2418, n3253, n3367, n2733);
and  g3622 (n3819, n2578, n3139, n3289, n3109);
nor  g3623 (n3609, n3102, n2492, n3186, n2764);
xnor g3624 (n3580, n2718, n3024, n2493, n2750);
or   g3625 (n3631, n2389, n3356, n3316, n3164);
xnor g3626 (n3670, n3191, n3002, n3268, n2902);
xor  g3627 (n3729, n3262, n2725, n2827, n3167);
and  g3628 (n3842, n2716, n3277, n2918, n2581);
and  g3629 (n3773, n2512, n3063, n3106, n2922);
xnor g3630 (n3651, n3315, n2446, n2515, n2606);
xor  g3631 (n3801, n2474, n2930, n2965, n2397);
xor  g3632 (n3821, n3198, n3005, n3327, n2537);
or   g3633 (n3838, n2421, n3326, n3321, n3032);
xor  g3634 (n3734, n3030, n2708, n3091, n2488);
and  g3635 (n3761, n2613, n2557, n3089, n3342);
and  g3636 (n3675, n2696, n2950, n2543, n3354);
nor  g3637 (n3624, n2437, n3261, n2774, n3008);
nor  g3638 (n3786, n3163, n2456, n2940, n2689);
xor  g3639 (n3616, n2318, n2604, n3145, n2558);
and  g3640 (n3793, n2470, n2416, n2611, n2693);
xor  g3641 (n3679, n3275, n2392, n3062, n2793);
nand g3642 (n3577, n2995, n2363, n2938, n2677);
xnor g3643 (n3710, n2562, n2359, n3379, n3299);
xnor g3644 (n3694, n2550, n3231, n2656, n2738);
xnor g3645 (n3831, n2998, n3023, n2607, n3197);
xnor g3646 (n3757, n2527, n3350, n2356, n2897);
xnor g3647 (n3638, n2464, n3161, n2948, n3211);
nand g3648 (n3829, n2993, n3092, n2460, n2941);
and  g3649 (n3637, n2745, n3228, n2483, n3304);
and  g3650 (n3765, n3169, n3085, n3237, n3225);
nand g3651 (n3834, n2324, n3149, n3339, n2326);
xnor g3652 (n3837, n2623, n3077, n3037, n2592);
and  g3653 (n3785, n2343, n2792, n3123, n2855);
nor  g3654 (n3632, n2463, n2570, n3027, n2327);
xor  g3655 (n3731, n2532, n2736, n2510, n2658);
xnor g3656 (n3705, n3305, n3130, n3156, n2767);
xnor g3657 (n3671, n2809, n2382, n3018, n3031);
nand g3658 (n3846, n2953, n3378, n3257, n3177);
or   g3659 (n3677, n2663, n2726, n2317, n2872);
xnor g3660 (n3717, n3148, n3135, n3244, n2877);
nand g3661 (n3775, n2526, n3122, n2489, n2312);
nor  g3662 (n3745, n2698, n2795, n2585, n3385);
or   g3663 (n3695, n2340, n2891, n3272, n2390);
or   g3664 (n3827, n2820, n3205, n2516, n3203);
xor  g3665 (n3640, n2332, n2402, n2610, n2654);
xnor g3666 (n3613, n2579, n2901, n2783, n3348);
nand g3667 (n3685, n3220, n3221, n2670, n2505);
and  g3668 (n3629, n3313, n3357, n2518, n3380);
and  g3669 (n3617, n3210, n2724, n3181, n3151);
xnor g3670 (n3666, n2817, n2710, n2743, n2433);
xor  g3671 (n3587, n2836, n2668, n2942, n2979);
and  g3672 (n3676, n2882, n2697, n2857, n2797);
or   g3673 (n3725, n2308, n2355, n2954, n2835);
xnor g3674 (n3708, n2554, n2913, n2369, n3328);
xnor g3675 (n3608, n3278, n3057, n2522, n2679);
or   g3676 (n3810, n2467, n3153, n3125, n2688);
nor  g3677 (n3714, n2400, n3016, n2883, n2547);
xor  g3678 (n3693, n2419, n2660, n2958, n3217);
xnor g3679 (n3633, n2454, n2563, n2852, n3292);
xor  g3680 (n3661, n3223, n3264, n2338, n2435);
and  g3681 (n3788, n3061, n2681, n3028, n3079);
nand g3682 (n3584, n3345, n3301, n2782, n2334);
or   g3683 (n3783, n2401, n2541, n3118, n2683);
or   g3684 (n3597, n2633, n2365, n2814, n2640);
xor  g3685 (n3688, n2399, n3338, n2928, n2442);
nor  g3686 (n3807, n2672, n2652, n2380, n3110);
or   g3687 (n3748, n2577, n2406, n2747, n2347);
xnor g3688 (n3678, n3370, n2445, n2923, n2354);
nor  g3689 (n3582, n2495, n3040, n2462, n3279);
and  g3690 (n3812, n3179, n3015, n3282, n2674);
or   g3691 (n3830, n2411, n2692, n2335, n2963);
xnor g3692 (n3664, n2662, n2988, n3097, n3160);
xor  g3693 (n3701, n3265, n3320, n2739, n2486);
xnor g3694 (n3747, n2497, n2721, n2911, n3093);
xnor g3695 (n3622, n3114, n2329, n3344, n3361);
and  g3696 (n3673, n2447, n3157, n2480, n3047);
xor  g3697 (n3763, n2916, n2310, n2566, n3201);
xor  g3698 (n3576, n2804, n3302, n3141, n2501);
or   g3699 (n3716, n2370, n2450, n2834, n2309);
nor  g3700 (n3653, n2568, n2990, n2991, n3127);
xor  g3701 (n3610, n3243, n2744, n2374, n2346);
nand g3702 (n3594, n2653, n3319, n2517, n2307);
nor  g3703 (n3668, n2755, n3283, n2860, n2603);
or   g3704 (n3682, n2757, n3133, n3162, n2412);
nand g3705 (n3808, n2742, n2614, n2344, n3116);
xnor g3706 (n3709, n2812, n3383, n2422, n2552);
or   g3707 (n3740, n2348, n3066, n2376, n2494);
nand g3708 (n3795, n3067, n2722, n2695, n2760);
nand g3709 (n3592, n2885, n2714, n3140, n3180);
nor  g3710 (n3641, n2838, n2952, n3096, n3332);
nor  g3711 (n3707, n2567, n3182, n2366, n2754);
or   g3712 (n3833, n2417, n2889, n2321, n2572);
nand g3713 (n3590, n2478, n3293, n3060, n3155);
and  g3714 (n3674, n2472, n2638, n2484, n2802);
xor  g3715 (n3792, n2686, n2723, n2691, n2856);
nand g3716 (n3800, n2477, n2584, n2535, n3070);
xor  g3717 (n3776, n2769, n2798, n2468, n2502);
xor  g3718 (n3712, n3111, n3147, n2386, n2594);
nand g3719 (n3669, n2933, n3307, n2593, n2659);
xor  g3720 (n3736, n2778, n3324, n2509, n2717);
nor  g3721 (n3699, n2513, n3011, n3224, n2909);
xnor g3722 (n3815, n2630, n2842, n3019, n3346);
nor  g3723 (n3713, n2597, n2475, n2546, n3146);
nand g3724 (n3720, n2977, n2641, n2560, n2983);
or   g3725 (n3735, n3075, n3009, n3360, n3045);
or   g3726 (n3579, n3269, n2694, n2974, n2947);
or   g3727 (n3813, n2824, n2949, n2413, n2661);
or   g3728 (n3630, n2383, n2590, n2878, n3048);
xnor g3729 (n3649, n2808, n3190, n2803, n3329);
nor  g3730 (n3711, n2520, n2571, n2893, n3055);
xor  g3731 (n3794, n2375, n2748, n3236, n3108);
xor  g3732 (n3780, n3312, n3189, n2625, n3219);
xor  g3733 (n3754, n2586, n3087, n3295, n2671);
nand g3734 (n3706, n2349, n2853, n2377, n2841);
xor  g3735 (n3636, n2449, n2927, n2773, n3188);
xnor g3736 (n3628, n2448, n2753, n2458, n2612);
xor  g3737 (n3781, n2685, n2951, n2999, n2439);
nand g3738 (n3723, n2647, n3050, n2845, n2989);
and  g3739 (n3755, n2859, n2756, n3041, n2908);
xnor g3740 (n3602, n3006, n3365, n3099, n3138);
xnor g3741 (n3727, n3290, n3036, n2945, n3311);
xor  g3742 (n3607, n2763, n2785, n2790, n2553);
xor  g3743 (n3604, n3171, n2542, n2636, n2854);
xor  g3744 (n3839, n2373, n2336, n2903, n3209);
nand g3745 (n3627, n2844, n2465, n2339, n3247);
nand g3746 (n3596, n3026, n2781, n3159, n2548);
nand g3747 (n3595, n3084, n2825, n2482, n2491);
nand g3748 (n3845, n2631, n2876, n2900, n2730);
and  g3749 (n3738, n2828, n2779, n3325, n2776);
and  g3750 (n3823, n2740, n2362, n2786, n2924);
xnor g3751 (n3684, n2664, n2620, n2728, n2962);
and  g3752 (n3648, n3168, n2443, n2810, n2796);
nor  g3753 (n3762, n2387, n2529, n3274, n3078);
or   g3754 (n3841, n2384, n2452, n3298, n3113);
nor  g3755 (n3759, n2507, n3184, n3142, n3234);
and  g3756 (n3768, n2644, n3128, n2678, n2639);
xnor g3757 (n3687, n2540, n2655, n2341, n2914);
or   g3758 (n3764, n2431, n3263, n2971, n2956);
xnor g3759 (n3692, n2935, n3233, n3330, n3384);
and  g3760 (n3698, n2396, n2879, n2368, n3103);
and  g3761 (n3844, n3255, n2379, n2441, n3049);
xor  g3762 (n3797, n2599, n2864, n2866, n2352);
or   g3763 (n3593, n2967, n2964, n3242, n2676);
and  g3764 (n3787, n3088, n2609, n2920, n2890);
nand g3765 (n3647, n2451, n2398, n3376, n2737);
nor  g3766 (n3618, n2617, n3017, n2910, n2886);
nor  g3767 (n3804, n2996, n2632, n2580, n2589);
xnor g3768 (n3626, n2508, n3306, n2784, n3101);
or   g3769 (n3672, n2816, n2466, n3386, n2896);
and  g3770 (n3680, n2504, n3022, n2331, n2699);
nor  g3771 (n3758, n2875, n3178, n2800, n2549);
nor  g3772 (n3840, n3368, n3349, n3271, n2832);
nor  g3773 (n3770, n2772, n2531, n3358, n2587);
and  g3774 (n3772, n2319, n2787, n2414, n3202);
nor  g3775 (n3728, n2569, n2471, n3134, n2759);
or   g3776 (n3614, n2712, n3059, n3294, n2939);
and  g3777 (n3779, n3229, n2976, n2746, n2946);
nand g3778 (n3809, n3232, n2405, n2833, n3058);
xor  g3779 (n3646, n2867, n3309, n2409, n3256);
or   g3780 (n3798, n2503, n2761, n3158, n3331);
nor  g3781 (n3642, n3258, n2524, n2624, n3183);
xnor g3782 (n3817, n2337, n2429, n2966, n3039);
or   g3783 (n3621, n2701, n2917, n3053, n2823);
nand g3784 (n3611, n2751, n3068, n2870, n2766);
or   g3785 (n3818, n2847, n2843, n2929, n2353);
xor  g3786 (n3586, n3381, n3038, n3076, n2575);
xnor g3787 (n3733, n2680, n2506, n2367, n2734);
xnor g3788 (n3644, n2423, n2555, n2727, n2345);
nor  g3789 (n3702, n2862, n3334, n2523, n2514);
or   g3790 (n3746, n3204, n2322, n2936, n3285);
nor  g3791 (n3657, n2973, n2881, n2850, n2848);
xnor g3792 (n3721, n2428, n2635, n2791, n2328);
or   g3793 (n3700, n3297, n2997, n2987, n2556);
xnor g3794 (n3791, n3351, n2616, n2528, n2944);
nor  g3795 (n3820, n2536, n2819, n2904, n3001);
xnor g3796 (n3686, n2801, n2994, n2391, n2511);
xnor g3797 (n3625, n3144, n3010, n2481, n2649);
nor  g3798 (n3751, n3249, n3337, n2574, n3052);
nor  g3799 (n3724, n2943, n3291, n3375, n3064);
xnor g3800 (n3753, n2559, n3323, n3013, n2888);
xnor g3801 (n3588, n3230, n3382, n2627, n3185);
nand g3802 (n3742, n3254, n2937, n2684, n2657);
nor  g3803 (n3662, n2752, n3372, n3235, n2682);
xor  g3804 (n3756, n3126, n2415, n3333, n2905);
xnor g3805 (n3766, n2521, n2972, n3137, n3273);
nor  g3806 (n3826, n3250, n3341, n2907, n2895);
or   g3807 (n3615, n2608, n3286, n3007, n2915);
and  g3808 (n3814, n2968, n2822, n3322, n3071);
nor  g3809 (n3760, n3260, n2788, n3364, n2873);
xor  g3810 (n3722, n3003, n3355, n3216, n2884);
nand g3811 (n3828, n2316, n2598, n2851, n2777);
nand g3812 (n3774, n2771, n2596, n3259, n2926);
and  g3813 (n3656, n2894, n3034, n3300, n2424);
nand g3814 (n3847, n3577, n3615, n3597, n3580);
nand g3815 (n3856, n3579, n3606, n3602, n3599);
xnor g3816 (n3851, n3605, n3593, n3613, n3607);
or   g3817 (n3848, n3601, n3610, n3598, n3584);
xnor g3818 (n3855, n3595, n3614, n3596, n3600);
and  g3819 (n3852, n3583, n3611, n3586, n3589);
nand g3820 (n3854, n3582, n3591, n3578, n3576);
or   g3821 (n3850, n3594, n3608, n3590, n3581);
or   g3822 (n3853, n3612, n3587, n3585, n3609);
nor  g3823 (n3849, n3603, n3592, n3604, n3588);
xor  g3824 (n3857, n3855, n3617, n3856, n3619);
or   g3825 (n3858, n3616, n3618, n3620, n3621);
buf  g3826 (n3859, n3857);
or   g3827 (n3860, n1369, n1367, n3857, n1371);
nand g3828 (n3862, n1370, n1226, n1368, n3858);
nand g3829 (n3861, n3858, n1113, n1226);
not  g3830 (n3877, n3624);
xnor g3831 (n3873, n3859, n1319, n3860, n1278);
xnor g3832 (n3875, n1278, n1325, n1323, n1372);
xor  g3833 (n3878, n3623, n3862, n3622, n1333);
nand g3834 (n3872, n1321, n3629, n1278, n1549);
and  g3835 (n3876, n1329, n3628, n3860, n1327);
nand g3836 (n3866, n1549, n3861, n1332, n3860);
or   g3837 (n3865, n3630, n3859, n1549, n3860);
nor  g3838 (n3868, n1331, n1326, n1548, n3861);
and  g3839 (n3863, n1324, n3625, n1337, n1320);
or   g3840 (n3864, n1278, n1330, n1373, n1318);
xor  g3841 (n3871, n3859, n1335, n3862, n1336);
nor  g3842 (n3867, n1328, n1338, n1277);
xnor g3843 (n3869, n3859, n3861, n1322, n1334);
xor  g3844 (n3870, n1277, n3861, n3627, n3862);
or   g3845 (n3874, n1549, n3862, n1277, n3626);
nand g3846 (n3904, n3481, n3874, n1117, n3456);
or   g3847 (n3923, n3865, n3505, n3437, n3543);
and  g3848 (n3920, n3413, n3876, n3399, n3520);
xnor g3849 (n3885, n3870, n3561, n3470, n3445);
xor  g3850 (n3913, n3540, n3433, n3864, n3868);
xor  g3851 (n3900, n3562, n3865, n3553, n3417);
and  g3852 (n3909, n3556, n3439, n3874, n3432);
or   g3853 (n3908, n3557, n3421, n3513, n3541);
and  g3854 (n3910, n3504, n3575, n3877, n3441);
xor  g3855 (n3895, n3572, n3555, n3479, n3528);
xor  g3856 (n3942, n3868, n3878, n3539, n3873);
xnor g3857 (n3921, n3863, n3482, n3865, n3406);
xnor g3858 (n3917, n3524, n3480, n3868, n3418);
xor  g3859 (n3929, n3395, n3442, n3431, n3483);
xnor g3860 (n3925, n3875, n3409, n3874, n3451);
nor  g3861 (n3927, n3865, n3554, n3497, n3877);
nor  g3862 (n3931, n3452, n3546, n3465, n3533);
xnor g3863 (n3907, n3872, n3870, n3569, n3869);
or   g3864 (n3937, n3478, n3570, n3400, n3878);
nand g3865 (n3912, n3494, n1114, n3873, n3551);
nor  g3866 (n3930, n3467, n3566, n3550, n3429);
and  g3867 (n3897, n3453, n3402, n3863, n3872);
xnor g3868 (n3890, n3527, n3488, n3866, n3450);
and  g3869 (n3896, n3863, n3427, n3872, n3573);
nand g3870 (n3889, n3871, n3475, n3869, n3501);
xor  g3871 (n3936, n3537, n3508, n3870, n3873);
xnor g3872 (n3881, n3466, n3515, n3510, n3491);
nor  g3873 (n3898, n3871, n3552, n3391, n3536);
nor  g3874 (n3893, n1115, n3518, n3542, n3864);
or   g3875 (n3883, n3517, n3878, n3499, n3875);
or   g3876 (n3903, n3398, n3411, n3876, n3871);
and  g3877 (n3911, n3485, n3455, n3463, n3435);
nor  g3878 (n3906, n3531, n3404, n3509, n3490);
and  g3879 (n3888, n3492, n3571, n3459, n3867);
xnor g3880 (n3924, n3477, n3388, n3568, n3436);
or   g3881 (n3884, n3548, n3397, n3476, n3454);
and  g3882 (n3894, n3472, n3506, n3872, n3512);
or   g3883 (n3880, n3449, n3877, n3428, n3538);
xnor g3884 (n3938, n3521, n3567, n1116, n3870);
or   g3885 (n3887, n3549, n3498, n3560, n3493);
nor  g3886 (n3916, n3522, n3530, n3396, n3460);
and  g3887 (n3926, n3864, n3486, n3496, n3464);
nor  g3888 (n3922, n3519, n3484, n3868, n3438);
nor  g3889 (n3928, n3444, n3407, n3430, n3869);
nand g3890 (n3892, n3425, n3878, n3877, n3403);
xor  g3891 (n3941, n3500, n3408, n3866, n3867);
and  g3892 (n3891, n3468, n3394, n3523, n3871);
and  g3893 (n3901, n3390, n3461, n3876, n3434);
or   g3894 (n3886, n3526, n3559, n3866, n3448);
or   g3895 (n3932, n3516, n3863, n3412, n3876);
xnor g3896 (n3919, n3864, n3426, n3392, n3544);
nor  g3897 (n3939, n3866, n3447, n3405, n3547);
and  g3898 (n3933, n3457, n3574, n3873, n3420);
and  g3899 (n3918, n3875, n3867, n3495, n3458);
or   g3900 (n3934, n3422, n3525, n3502, n3443);
xor  g3901 (n3902, n3867, n3446, n3565, n3545);
xnor g3902 (n3915, n3410, n3416, n3414, n3471);
xor  g3903 (n3914, n3462, n3558, n3473, n3487);
and  g3904 (n3899, n3424, n3563, n3529, n3564);
xor  g3905 (n3905, n3875, n3440, n3869, n3423);
or   g3906 (n3882, n3534, n3419, n3511, n3393);
nand g3907 (n3935, n3489, n3535, n3401, n3874);
xnor g3908 (n3940, n3469, n3389, n3532, n3503);
nand g3909 (n3879, n3474, n3415, n3507, n3514);
nor  g3910 (n3988, n3704, n3841, n3743, n3715);
or   g3911 (n3974, n3754, n3779, n3664, n3687);
and  g3912 (n3984, n3925, n3773, n3711, n3902);
nand g3913 (n3980, n3836, n3832, n3924, n3918);
xnor g3914 (n3963, n3776, n3768, n3818, n3914);
nand g3915 (n3972, n3908, n3785, n3751, n3699);
nor  g3916 (n4010, n3937, n3730, n3766, n3634);
nand g3917 (n3943, n3938, n3815, n3939, n3679);
or   g3918 (n3981, n3895, n3915, n3659, n3791);
nor  g3919 (n4002, n3710, n3845, n3834, n3680);
and  g3920 (n3987, n3926, n3705, n3642, n3896);
nand g3921 (n3964, n3676, n3805, n3712, n3667);
and  g3922 (n3951, n3792, n3767, n3631, n3894);
xor  g3923 (n3989, n3787, n3700, n3665, n3723);
nor  g3924 (n3993, n3770, n3758, n3720, n3652);
and  g3925 (n3971, n3753, n3752, n3930, n3736);
or   g3926 (n4009, n3802, n3934, n3635, n3729);
xor  g3927 (n3954, n3820, n3782, n3674, n3786);
nand g3928 (n4004, n3844, n3681, n3798, n3727);
xnor g3929 (n3986, n3839, n3647, n3813, n3812);
nor  g3930 (n3947, n3677, n3718, n3826, n3735);
and  g3931 (n3944, n3660, n3817, n3808, n3821);
xnor g3932 (n3994, n3935, n3835, n3684, n3886);
xnor g3933 (n3977, n3666, n3749, n3748, n3673);
nand g3934 (n3991, n3788, n3790, n3693, n3900);
xnor g3935 (n3955, n3940, n3734, n3827, n3824);
nor  g3936 (n4005, n3807, n3672, n3784, n3745);
and  g3937 (n3978, n3881, n3638, n3883, n3759);
and  g3938 (n3995, n3891, n3724, n3655, n3939);
nor  g3939 (n3982, n3662, n3632, n3901, n3695);
xor  g3940 (n3950, n3757, n3933, n3903, n3898);
or   g3941 (n4000, n3941, n3889, n3899, n3940);
xor  g3942 (n3998, n3942, n3649, n3651, n3640);
and  g3943 (n3965, n3880, n3694, n3838, n3733);
nor  g3944 (n3953, n3761, n3641, n3721, n3750);
or   g3945 (n3985, n3739, n3897, n3708, n3714);
xnor g3946 (n3948, n3690, n3911, n3707, n3936);
xor  g3947 (n3945, n3904, n3816, n3756, n3804);
or   g3948 (n3983, n3794, n3747, n3726, n3656);
nor  g3949 (n3959, n3709, n3837, n3774, n3842);
nand g3950 (n4012, n3795, n3917, n3728, n3738);
nand g3951 (n3956, n3731, n3741, n3703, n3799);
nor  g3952 (n3967, n3906, n3780, n3829, n3801);
and  g3953 (n3966, n3658, n3670, n3645, n3920);
nor  g3954 (n4008, n3760, n3814, n3907, n3650);
xor  g3955 (n4011, n3769, n3919, n3840, n3669);
xor  g3956 (n3946, n3633, n3686, n3942, n3809);
xnor g3957 (n3968, n3936, n3732, n3698, n3719);
or   g3958 (n3949, n3697, n3639, n3909, n3764);
and  g3959 (n3957, n3843, n3646, n3921, n3654);
nand g3960 (n3961, n3806, n3713, n3884, n3746);
nand g3961 (n3962, n3830, n3913, n3689, n3828);
xnor g3962 (n3973, n3912, n3923, n3783, n3882);
xnor g3963 (n4001, n3661, n3668, n3893, n3777);
nor  g3964 (n3958, n3825, n3701, n3755, n3916);
nor  g3965 (n3999, n3778, n3725, n3928, n3717);
nand g3966 (n3992, n3796, n3823, n3744, n3722);
nor  g3967 (n3952, n3763, n3932, n3683, n3803);
xor  g3968 (n4014, n3888, n3833, n3929, n3742);
and  g3969 (n3990, n3682, n3831, n3922, n3685);
xnor g3970 (n4003, n3887, n3653, n3775, n3797);
xor  g3971 (n3996, n3636, n3793, n3737, n3762);
and  g3972 (n3960, n3879, n3811, n3937, n3771);
xnor g3973 (n4006, n3927, n3941, n3931, n3671);
and  g3974 (n3979, n3765, n3692, n3716, n3800);
and  g3975 (n3970, n3935, n3740, n3706, n3643);
and  g3976 (n3997, n3637, n3789, n3781, n3938);
xnor g3977 (n4007, n3810, n3678, n3910, n3663);
nand g3978 (n3976, n3905, n3822, n3846, n3819);
or   g3979 (n3975, n3702, n3696, n3892, n3657);
xnor g3980 (n4013, n3644, n3885, n3688, n3675);
nor  g3981 (n3969, n3648, n3691, n3772, n3890);
nand g3982 (n4015, n3951, n3956, n3993, n3972);
or   g3983 (n4031, n3958, n3980, n3995, n3960);
or   g3984 (n4026, n3962, n4003, n3999, n3952);
and  g3985 (n4018, n4004, n3944, n3990, n4011);
nor  g3986 (n4028, n3965, n3982, n3961, n4007);
and  g3987 (n4019, n3998, n3953, n4000, n4010);
or   g3988 (n4022, n3970, n3984, n3992, n3985);
xnor g3989 (n4023, n3968, n3971, n3946, n4005);
or   g3990 (n4017, n3966, n3994, n3986, n3983);
and  g3991 (n4020, n4008, n3974, n3978, n3989);
xnor g3992 (n4029, n4001, n3981, n3976, n4014);
or   g3993 (n4025, n3979, n3955, n4009, n3975);
and  g3994 (n4016, n3948, n3964, n3991, n3987);
nor  g3995 (n4021, n3977, n3947, n4006, n3959);
nand g3996 (n4024, n3949, n3996, n3967, n4002);
nand g3997 (n4027, n4013, n3945, n3957, n3963);
xor  g3998 (n4030, n3997, n3988, n3954, n3943);
or   g3999 (n4032, n4012, n3950, n3969, n3973);
endmodule
