

module Stat_3000_432
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n82,
  n74,
  n57,
  n41,
  n114,
  n61,
  n70,
  n121,
  n112,
  n85,
  n104,
  n124,
  n67,
  n132,
  n117,
  n76,
  n1107,
  n1108,
  n1113,
  n1116,
  n3011,
  n3015,
  n3014,
  n3010,
  n3009,
  n3013,
  n3008,
  n3022,
  n3024,
  n3030,
  n3031,
  n3032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n82;
  output n74;
  output n57;
  output n41;
  output n114;
  output n61;
  output n70;
  output n121;
  output n112;
  output n85;
  output n104;
  output n124;
  output n67;
  output n132;
  output n117;
  output n76;
  output n1107;
  output n1108;
  output n1113;
  output n1116;
  output n3011;
  output n3015;
  output n3014;
  output n3010;
  output n3009;
  output n3013;
  output n3008;
  output n3022;
  output n3024;
  output n3030;
  output n3031;
  output n3032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n58;
  wire n59;
  wire n60;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n68;
  wire n69;
  wire n71;
  wire n72;
  wire n73;
  wire n75;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n83;
  wire n84;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n113;
  wire n115;
  wire n116;
  wire n118;
  wire n119;
  wire n120;
  wire n122;
  wire n123;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1114;
  wire n1115;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3012;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3023;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n80,
    n27
  );


  not
  g1
  (
    n59,
    n16
  );


  not
  g2
  (
    n127,
    n3
  );


  buf
  g3
  (
    n60,
    n8
  );


  buf
  g4
  (
    n52,
    n21
  );


  buf
  g5
  (
    n36,
    n20
  );


  buf
  g6
  (
    n132,
    n16
  );


  buf
  g7
  (
    KeyWire_0_29,
    n21
  );


  not
  g8
  (
    n71,
    n26
  );


  not
  g9
  (
    n97,
    n25
  );


  buf
  g10
  (
    n102,
    n15
  );


  not
  g11
  (
    n114,
    n11
  );


  not
  g12
  (
    n87,
    n26
  );


  not
  g13
  (
    n84,
    n18
  );


  buf
  g14
  (
    n110,
    n31
  );


  buf
  g15
  (
    n103,
    n14
  );


  buf
  g16
  (
    n124,
    n25
  );


  not
  g17
  (
    n118,
    n18
  );


  not
  g18
  (
    n40,
    n19
  );


  not
  g19
  (
    n56,
    n1
  );


  buf
  g20
  (
    n90,
    n27
  );


  buf
  g21
  (
    n38,
    n3
  );


  buf
  g22
  (
    n61,
    n6
  );


  buf
  g23
  (
    n119,
    n20
  );


  not
  g24
  (
    n77,
    n19
  );


  not
  g25
  (
    n39,
    n12
  );


  buf
  g26
  (
    n86,
    n22
  );


  buf
  g27
  (
    n106,
    n8
  );


  not
  g28
  (
    n116,
    n26
  );


  buf
  g29
  (
    n54,
    n15
  );


  not
  g30
  (
    n120,
    n17
  );


  not
  g31
  (
    n46,
    n6
  );


  not
  g32
  (
    n101,
    n24
  );


  buf
  g33
  (
    n108,
    n2
  );


  buf
  g34
  (
    n70,
    n26
  );


  buf
  g35
  (
    n104,
    n9
  );


  not
  g36
  (
    n55,
    n5
  );


  buf
  g37
  (
    n58,
    n10
  );


  not
  g38
  (
    n65,
    n13
  );


  not
  g39
  (
    n126,
    n23
  );


  not
  g40
  (
    n68,
    n24
  );


  buf
  g41
  (
    n123,
    n11
  );


  not
  g42
  (
    n48,
    n22
  );


  buf
  g43
  (
    n111,
    n14
  );


  not
  g44
  (
    KeyWire_0_22,
    n19
  );


  not
  g45
  (
    n45,
    n20
  );


  not
  g46
  (
    n81,
    n23
  );


  not
  g47
  (
    n78,
    n3
  );


  buf
  g48
  (
    n100,
    n9
  );


  buf
  g49
  (
    n34,
    n28
  );


  not
  g50
  (
    n41,
    n29
  );


  not
  g51
  (
    n66,
    n27
  );


  not
  g52
  (
    n113,
    n13
  );


  buf
  g53
  (
    n112,
    n7
  );


  not
  g54
  (
    n37,
    n13
  );


  not
  g55
  (
    KeyWire_0_6,
    n30
  );


  buf
  g56
  (
    n69,
    n30
  );


  buf
  g57
  (
    n121,
    n23
  );


  not
  g58
  (
    n42,
    n12
  );


  not
  g59
  (
    n72,
    n28
  );


  not
  g60
  (
    n47,
    n5
  );


  not
  g61
  (
    n122,
    n28
  );


  not
  g62
  (
    n107,
    n6
  );


  buf
  g63
  (
    n115,
    n22
  );


  buf
  g64
  (
    n35,
    n27
  );


  buf
  g65
  (
    n79,
    n4
  );


  not
  g66
  (
    n128,
    n11
  );


  not
  g67
  (
    n74,
    n10
  );


  buf
  g68
  (
    n91,
    n7
  );


  not
  g69
  (
    n53,
    n30
  );


  not
  g70
  (
    n83,
    n31
  );


  not
  g71
  (
    n98,
    n17
  );


  buf
  g72
  (
    n67,
    n2
  );


  not
  g73
  (
    n57,
    n25
  );


  buf
  g74
  (
    n64,
    n18
  );


  buf
  g75
  (
    n76,
    n17
  );


  buf
  g76
  (
    n125,
    n29
  );


  buf
  g77
  (
    n130,
    n29
  );


  not
  g78
  (
    n82,
    n4
  );


  not
  g79
  (
    n50,
    n29
  );


  buf
  g80
  (
    n96,
    n1
  );


  not
  g81
  (
    n95,
    n25
  );


  not
  g82
  (
    n89,
    n15
  );


  not
  g83
  (
    n94,
    n5
  );


  buf
  g84
  (
    n85,
    n12
  );


  buf
  g85
  (
    n105,
    n30
  );


  buf
  g86
  (
    n88,
    n4
  );


  not
  g87
  (
    n51,
    n14
  );


  not
  g88
  (
    n63,
    n16
  );


  buf
  g89
  (
    n117,
    n9
  );


  not
  g90
  (
    n49,
    n7
  );


  buf
  g91
  (
    n109,
    n28
  );


  not
  g92
  (
    n44,
    n8
  );


  buf
  g93
  (
    n33,
    n24
  );


  not
  g94
  (
    n129,
    n2
  );


  not
  g95
  (
    n99,
    n1
  );


  not
  g96
  (
    n43,
    n31
  );


  buf
  g97
  (
    n75,
    n31
  );


  buf
  g98
  (
    n73,
    n10
  );


  not
  g99
  (
    n62,
    n21
  );


  buf
  g100
  (
    n332,
    n120
  );


  buf
  g101
  (
    n374,
    n61
  );


  not
  g102
  (
    n203,
    n38
  );


  not
  g103
  (
    n473,
    n91
  );


  buf
  g104
  (
    n407,
    n71
  );


  not
  g105
  (
    n158,
    n68
  );


  not
  g106
  (
    n471,
    n128
  );


  not
  g107
  (
    n272,
    n87
  );


  buf
  g108
  (
    n313,
    n104
  );


  not
  g109
  (
    n134,
    n66
  );


  not
  g110
  (
    n392,
    n65
  );


  buf
  g111
  (
    n323,
    n56
  );


  buf
  g112
  (
    n213,
    n121
  );


  buf
  g113
  (
    n315,
    n122
  );


  not
  g114
  (
    n464,
    n56
  );


  buf
  g115
  (
    n152,
    n78
  );


  not
  g116
  (
    n389,
    n93
  );


  not
  g117
  (
    n502,
    n63
  );


  buf
  g118
  (
    n357,
    n115
  );


  buf
  g119
  (
    n308,
    n126
  );


  buf
  g120
  (
    n229,
    n34
  );


  buf
  g121
  (
    n133,
    n107
  );


  not
  g122
  (
    n230,
    n79
  );


  not
  g123
  (
    n404,
    n96
  );


  not
  g124
  (
    n336,
    n124
  );


  buf
  g125
  (
    n261,
    n110
  );


  buf
  g126
  (
    n453,
    n91
  );


  buf
  g127
  (
    n439,
    n58
  );


  buf
  g128
  (
    n376,
    n108
  );


  buf
  g129
  (
    n183,
    n79
  );


  not
  g130
  (
    n296,
    n105
  );


  not
  g131
  (
    n472,
    n48
  );


  buf
  g132
  (
    KeyWire_0_31,
    n123
  );


  not
  g133
  (
    KeyWire_0_15,
    n62
  );


  not
  g134
  (
    n335,
    n73
  );


  not
  g135
  (
    n483,
    n50
  );


  buf
  g136
  (
    n454,
    n97
  );


  not
  g137
  (
    n321,
    n58
  );


  not
  g138
  (
    n177,
    n106
  );


  not
  g139
  (
    n197,
    n34
  );


  buf
  g140
  (
    n388,
    n118
  );


  buf
  g141
  (
    n157,
    n111
  );


  buf
  g142
  (
    n316,
    n92
  );


  not
  g143
  (
    n419,
    n123
  );


  not
  g144
  (
    n284,
    n103
  );


  not
  g145
  (
    n244,
    n92
  );


  not
  g146
  (
    n222,
    n73
  );


  buf
  g147
  (
    n493,
    n79
  );


  buf
  g148
  (
    n383,
    n38
  );


  not
  g149
  (
    n145,
    n39
  );


  buf
  g150
  (
    n173,
    n132
  );


  not
  g151
  (
    n504,
    n46
  );


  buf
  g152
  (
    n167,
    n88
  );


  not
  g153
  (
    n142,
    n117
  );


  buf
  g154
  (
    n154,
    n47
  );


  not
  g155
  (
    n136,
    n62
  );


  buf
  g156
  (
    n162,
    n51
  );


  buf
  g157
  (
    n148,
    n70
  );


  not
  g158
  (
    n266,
    n57
  );


  not
  g159
  (
    KeyWire_0_28,
    n85
  );


  buf
  g160
  (
    n372,
    n130
  );


  not
  g161
  (
    n487,
    n124
  );


  buf
  g162
  (
    n475,
    n115
  );


  not
  g163
  (
    n243,
    n110
  );


  not
  g164
  (
    n438,
    n117
  );


  buf
  g165
  (
    n351,
    n114
  );


  not
  g166
  (
    n458,
    n128
  );


  not
  g167
  (
    n385,
    n83
  );


  not
  g168
  (
    n288,
    n106
  );


  not
  g169
  (
    n141,
    n90
  );


  not
  g170
  (
    n248,
    n35
  );


  not
  g171
  (
    n364,
    n126
  );


  not
  g172
  (
    n302,
    n112
  );


  buf
  g173
  (
    n146,
    n107
  );


  buf
  g174
  (
    n344,
    n99
  );


  buf
  g175
  (
    n137,
    n118
  );


  buf
  g176
  (
    n184,
    n45
  );


  not
  g177
  (
    n198,
    n128
  );


  not
  g178
  (
    n211,
    n60
  );


  buf
  g179
  (
    n452,
    n54
  );


  buf
  g180
  (
    n415,
    n131
  );


  buf
  g181
  (
    n495,
    n117
  );


  not
  g182
  (
    n492,
    n110
  );


  buf
  g183
  (
    n330,
    n70
  );


  not
  g184
  (
    n373,
    n82
  );


  buf
  g185
  (
    n401,
    n37
  );


  buf
  g186
  (
    n189,
    n131
  );


  buf
  g187
  (
    n235,
    n109
  );


  buf
  g188
  (
    n236,
    n119
  );


  buf
  g189
  (
    n247,
    n101
  );


  not
  g190
  (
    n496,
    n127
  );


  not
  g191
  (
    n138,
    n67
  );


  not
  g192
  (
    n371,
    n72
  );


  not
  g193
  (
    n500,
    n66
  );


  not
  g194
  (
    n216,
    n54
  );


  not
  g195
  (
    n449,
    n125
  );


  not
  g196
  (
    n366,
    n74
  );


  buf
  g197
  (
    n176,
    n71
  );


  buf
  g198
  (
    n411,
    n53
  );


  not
  g199
  (
    n349,
    n62
  );


  not
  g200
  (
    n512,
    n68
  );


  not
  g201
  (
    n207,
    n93
  );


  not
  g202
  (
    n422,
    n47
  );


  buf
  g203
  (
    n461,
    n69
  );


  buf
  g204
  (
    n513,
    n39
  );


  buf
  g205
  (
    n305,
    n81
  );


  not
  g206
  (
    n283,
    n77
  );


  buf
  g207
  (
    n242,
    n67
  );


  not
  g208
  (
    n187,
    n112
  );


  buf
  g209
  (
    n246,
    n90
  );


  not
  g210
  (
    n440,
    n47
  );


  not
  g211
  (
    n150,
    n89
  );


  buf
  g212
  (
    n204,
    n71
  );


  buf
  g213
  (
    n466,
    n42
  );


  not
  g214
  (
    n338,
    n41
  );


  buf
  g215
  (
    n292,
    n49
  );


  buf
  g216
  (
    n277,
    n55
  );


  buf
  g217
  (
    n274,
    n98
  );


  not
  g218
  (
    n180,
    n91
  );


  buf
  g219
  (
    n149,
    n116
  );


  buf
  g220
  (
    n486,
    n35
  );


  buf
  g221
  (
    n267,
    n82
  );


  buf
  g222
  (
    n185,
    n102
  );


  not
  g223
  (
    n463,
    n125
  );


  buf
  g224
  (
    n363,
    n89
  );


  not
  g225
  (
    n484,
    n59
  );


  buf
  g226
  (
    n360,
    n77
  );


  not
  g227
  (
    n468,
    n54
  );


  not
  g228
  (
    n358,
    n86
  );


  not
  g229
  (
    n205,
    n75
  );


  not
  g230
  (
    n359,
    n60
  );


  buf
  g231
  (
    n278,
    n57
  );


  not
  g232
  (
    n498,
    n39
  );


  buf
  g233
  (
    n379,
    n115
  );


  buf
  g234
  (
    n161,
    n119
  );


  not
  g235
  (
    n225,
    n113
  );


  buf
  g236
  (
    n437,
    n89
  );


  not
  g237
  (
    n408,
    n53
  );


  buf
  g238
  (
    n442,
    n107
  );


  buf
  g239
  (
    n218,
    n102
  );


  buf
  g240
  (
    n514,
    n113
  );


  not
  g241
  (
    n465,
    n93
  );


  buf
  g242
  (
    n506,
    n114
  );


  not
  g243
  (
    n319,
    n98
  );


  not
  g244
  (
    n390,
    n49
  );


  not
  g245
  (
    n451,
    n70
  );


  buf
  g246
  (
    n345,
    n74
  );


  not
  g247
  (
    n171,
    n111
  );


  not
  g248
  (
    n253,
    n86
  );


  not
  g249
  (
    n251,
    n78
  );


  not
  g250
  (
    n159,
    n63
  );


  buf
  g251
  (
    n318,
    n72
  );


  buf
  g252
  (
    n329,
    n95
  );


  not
  g253
  (
    n325,
    n81
  );


  buf
  g254
  (
    n234,
    n95
  );


  not
  g255
  (
    n356,
    n59
  );


  not
  g256
  (
    n233,
    n101
  );


  buf
  g257
  (
    n343,
    n105
  );


  buf
  g258
  (
    n350,
    n37
  );


  buf
  g259
  (
    n348,
    n109
  );


  buf
  g260
  (
    n300,
    n80
  );


  buf
  g261
  (
    n309,
    n76
  );


  buf
  g262
  (
    n239,
    n42
  );


  buf
  g263
  (
    n402,
    n46
  );


  buf
  g264
  (
    n260,
    n91
  );


  buf
  g265
  (
    n250,
    n120
  );


  not
  g266
  (
    n231,
    n80
  );


  not
  g267
  (
    n431,
    n100
  );


  buf
  g268
  (
    n447,
    n77
  );


  buf
  g269
  (
    n462,
    n84
  );


  buf
  g270
  (
    n306,
    n88
  );


  not
  g271
  (
    n507,
    n77
  );


  not
  g272
  (
    n286,
    n92
  );


  buf
  g273
  (
    n400,
    n132
  );


  not
  g274
  (
    n215,
    n111
  );


  buf
  g275
  (
    n287,
    n112
  );


  not
  g276
  (
    n485,
    n40
  );


  not
  g277
  (
    n221,
    n63
  );


  not
  g278
  (
    n280,
    n116
  );


  buf
  g279
  (
    n327,
    n63
  );


  buf
  g280
  (
    n474,
    n44
  );


  buf
  g281
  (
    n144,
    n64
  );


  not
  g282
  (
    n254,
    n66
  );


  buf
  g283
  (
    n258,
    n53
  );


  buf
  g284
  (
    n151,
    n111
  );


  buf
  g285
  (
    n499,
    n108
  );


  not
  g286
  (
    n303,
    n105
  );


  buf
  g287
  (
    n378,
    n35
  );


  buf
  g288
  (
    n270,
    n113
  );


  buf
  g289
  (
    n224,
    n98
  );


  not
  g290
  (
    n301,
    n100
  );


  not
  g291
  (
    n294,
    n92
  );


  buf
  g292
  (
    n489,
    n129
  );


  not
  g293
  (
    n240,
    n103
  );


  buf
  g294
  (
    n456,
    n86
  );


  not
  g295
  (
    n426,
    n98
  );


  buf
  g296
  (
    n428,
    n118
  );


  not
  g297
  (
    n397,
    n102
  );


  buf
  g298
  (
    n467,
    n69
  );


  not
  g299
  (
    n409,
    n52
  );


  not
  g300
  (
    n307,
    n109
  );


  not
  g301
  (
    n460,
    n82
  );


  not
  g302
  (
    n135,
    n129
  );


  not
  g303
  (
    n252,
    n88
  );


  not
  g304
  (
    n334,
    n127
  );


  buf
  g305
  (
    n314,
    n97
  );


  not
  g306
  (
    n181,
    n62
  );


  buf
  g307
  (
    n339,
    n100
  );


  buf
  g308
  (
    n347,
    n120
  );


  buf
  g309
  (
    n435,
    n131
  );


  not
  g310
  (
    n368,
    n72
  );


  not
  g311
  (
    n219,
    n106
  );


  not
  g312
  (
    n380,
    n61
  );


  not
  g313
  (
    n174,
    n84
  );


  buf
  g314
  (
    n433,
    n104
  );


  not
  g315
  (
    n361,
    n95
  );


  buf
  g316
  (
    n398,
    n78
  );


  buf
  g317
  (
    n191,
    n104
  );


  not
  g318
  (
    n156,
    n108
  );


  not
  g319
  (
    n153,
    n94
  );


  buf
  g320
  (
    n370,
    n49
  );


  not
  g321
  (
    n436,
    n80
  );


  buf
  g322
  (
    n386,
    n34
  );


  buf
  g323
  (
    n209,
    n42
  );


  buf
  g324
  (
    n241,
    n103
  );


  not
  g325
  (
    n226,
    n119
  );


  not
  g326
  (
    n194,
    n36
  );


  not
  g327
  (
    n263,
    n114
  );


  buf
  g328
  (
    n228,
    n45
  );


  not
  g329
  (
    n424,
    n107
  );


  buf
  g330
  (
    n396,
    n59
  );


  buf
  g331
  (
    n320,
    n60
  );


  not
  g332
  (
    n455,
    n81
  );


  not
  g333
  (
    n480,
    n130
  );


  not
  g334
  (
    n477,
    n97
  );


  not
  g335
  (
    n342,
    n131
  );


  buf
  g336
  (
    n238,
    n116
  );


  buf
  g337
  (
    n354,
    n76
  );


  buf
  g338
  (
    KeyWire_0_43,
    n76
  );


  not
  g339
  (
    n289,
    n88
  );


  not
  g340
  (
    n432,
    n101
  );


  buf
  g341
  (
    n394,
    n41
  );


  buf
  g342
  (
    n175,
    n56
  );


  buf
  g343
  (
    n291,
    n73
  );


  not
  g344
  (
    n365,
    n61
  );


  buf
  g345
  (
    n515,
    n102
  );


  not
  g346
  (
    n423,
    n114
  );


  not
  g347
  (
    n281,
    n64
  );


  buf
  g348
  (
    n418,
    n64
  );


  buf
  g349
  (
    n481,
    n110
  );


  buf
  g350
  (
    n410,
    n94
  );


  not
  g351
  (
    n482,
    n52
  );


  not
  g352
  (
    n469,
    n65
  );


  buf
  g353
  (
    n256,
    n99
  );


  not
  g354
  (
    n501,
    n64
  );


  buf
  g355
  (
    n193,
    n68
  );


  buf
  g356
  (
    n279,
    n112
  );


  not
  g357
  (
    n237,
    n55
  );


  buf
  g358
  (
    n446,
    n59
  );


  buf
  g359
  (
    n430,
    n66
  );


  buf
  g360
  (
    n417,
    n95
  );


  not
  g361
  (
    n160,
    n75
  );


  not
  g362
  (
    n367,
    n43
  );


  buf
  g363
  (
    n412,
    n83
  );


  buf
  g364
  (
    n212,
    n55
  );


  not
  g365
  (
    n494,
    n113
  );


  not
  g366
  (
    n304,
    n57
  );


  not
  g367
  (
    n271,
    n83
  );


  buf
  g368
  (
    n352,
    n125
  );


  not
  g369
  (
    n429,
    n74
  );


  not
  g370
  (
    n182,
    n115
  );


  buf
  g371
  (
    n444,
    n69
  );


  not
  g372
  (
    n387,
    n126
  );


  buf
  g373
  (
    n168,
    n52
  );


  not
  g374
  (
    n337,
    n103
  );


  buf
  g375
  (
    n406,
    n51
  );


  buf
  g376
  (
    n268,
    n129
  );


  buf
  g377
  (
    n297,
    n87
  );


  not
  g378
  (
    n322,
    n67
  );


  buf
  g379
  (
    n457,
    n89
  );


  not
  g380
  (
    n503,
    n125
  );


  buf
  g381
  (
    n164,
    n56
  );


  not
  g382
  (
    n355,
    n122
  );


  buf
  g383
  (
    n165,
    n76
  );


  not
  g384
  (
    n190,
    n99
  );


  not
  g385
  (
    n285,
    n96
  );


  buf
  g386
  (
    n196,
    n117
  );


  not
  g387
  (
    n490,
    n108
  );


  buf
  g388
  (
    n331,
    n106
  );


  buf
  g389
  (
    n405,
    n61
  );


  buf
  g390
  (
    n511,
    n40
  );


  buf
  g391
  (
    n140,
    n94
  );


  buf
  g392
  (
    n208,
    n127
  );


  not
  g393
  (
    n179,
    n118
  );


  buf
  g394
  (
    n399,
    n121
  );


  buf
  g395
  (
    n245,
    n87
  );


  buf
  g396
  (
    n166,
    n123
  );


  buf
  g397
  (
    n445,
    n101
  );


  not
  g398
  (
    n312,
    n96
  );


  buf
  g399
  (
    n377,
    n50
  );


  not
  g400
  (
    n172,
    n126
  );


  not
  g401
  (
    n163,
    n46
  );


  buf
  g402
  (
    KeyWire_0_9,
    n87
  );


  not
  g403
  (
    n202,
    n82
  );


  buf
  g404
  (
    n147,
    n122
  );


  buf
  g405
  (
    n249,
    n40
  );


  not
  g406
  (
    n420,
    n122
  );


  not
  g407
  (
    n333,
    n49
  );


  not
  g408
  (
    n491,
    n124
  );


  not
  g409
  (
    n478,
    n132
  );


  buf
  g410
  (
    n259,
    n129
  );


  buf
  g411
  (
    KeyWire_0_19,
    n58
  );


  not
  g412
  (
    n326,
    n70
  );


  not
  g413
  (
    n362,
    n84
  );


  buf
  g414
  (
    n298,
    n121
  );


  not
  g415
  (
    n290,
    n37
  );


  not
  g416
  (
    n293,
    n43
  );


  buf
  g417
  (
    n273,
    n93
  );


  buf
  g418
  (
    n232,
    n41
  );


  not
  g419
  (
    n416,
    n79
  );


  not
  g420
  (
    n200,
    n123
  );


  buf
  g421
  (
    n317,
    n94
  );


  buf
  g422
  (
    n311,
    n97
  );


  not
  g423
  (
    n265,
    n104
  );


  buf
  g424
  (
    n340,
    n55
  );


  not
  g425
  (
    n299,
    n65
  );


  not
  g426
  (
    n220,
    n109
  );


  not
  g427
  (
    n413,
    n90
  );


  buf
  g428
  (
    n403,
    n85
  );


  not
  g429
  (
    n223,
    n58
  );


  not
  g430
  (
    n170,
    n83
  );


  buf
  g431
  (
    n476,
    n50
  );


  not
  g432
  (
    KeyWire_0_34,
    n85
  );


  not
  g433
  (
    n217,
    n44
  );


  buf
  g434
  (
    n441,
    n48
  );


  buf
  g435
  (
    n206,
    n33
  );


  buf
  g436
  (
    n421,
    n44
  );


  buf
  g437
  (
    n178,
    n33
  );


  buf
  g438
  (
    n295,
    n60
  );


  not
  g439
  (
    n450,
    n85
  );


  not
  g440
  (
    n282,
    n81
  );


  buf
  g441
  (
    n276,
    n74
  );


  buf
  g442
  (
    n510,
    n53
  );


  buf
  g443
  (
    n341,
    n120
  );


  buf
  g444
  (
    n509,
    n100
  );


  buf
  g445
  (
    n199,
    n119
  );


  buf
  g446
  (
    n214,
    n45
  );


  not
  g447
  (
    n434,
    n130
  );


  not
  g448
  (
    n346,
    n72
  );


  not
  g449
  (
    n169,
    n124
  );


  not
  g450
  (
    n395,
    n78
  );


  buf
  g451
  (
    n479,
    n116
  );


  buf
  g452
  (
    n375,
    n38
  );


  not
  g453
  (
    n275,
    n71
  );


  not
  g454
  (
    n470,
    n36
  );


  not
  g455
  (
    n188,
    n43
  );


  buf
  g456
  (
    n186,
    n68
  );


  not
  g457
  (
    n310,
    n73
  );


  buf
  g458
  (
    n139,
    n54
  );


  not
  g459
  (
    n391,
    n86
  );


  not
  g460
  (
    n384,
    n90
  );


  buf
  g461
  (
    n505,
    n69
  );


  not
  g462
  (
    n508,
    n48
  );


  buf
  g463
  (
    n155,
    n65
  );


  buf
  g464
  (
    n393,
    n96
  );


  not
  g465
  (
    n353,
    n51
  );


  buf
  g466
  (
    n324,
    n99
  );


  buf
  g467
  (
    n427,
    n57
  );


  not
  g468
  (
    n459,
    n36
  );


  not
  g469
  (
    n195,
    n75
  );


  not
  g470
  (
    n262,
    n51
  );


  not
  g471
  (
    KeyWire_0_8,
    n52
  );


  buf
  g472
  (
    n269,
    n33
  );


  not
  g473
  (
    n369,
    n84
  );


  buf
  g474
  (
    n488,
    n128
  );


  buf
  g475
  (
    n497,
    n127
  );


  not
  g476
  (
    n227,
    n130
  );


  not
  g477
  (
    n143,
    n121
  );


  not
  g478
  (
    n210,
    n80
  );


  not
  g479
  (
    n201,
    n75
  );


  not
  g480
  (
    n192,
    n105
  );


  buf
  g481
  (
    n425,
    n67
  );


  buf
  g482
  (
    n414,
    n50
  );


  and
  g483
  (
    n744,
    n349,
    n405,
    n420,
    n137
  );


  xnor
  g484
  (
    n845,
    n465,
    n475,
    n427,
    n432
  );


  or
  g485
  (
    n607,
    n262,
    n371,
    n295,
    n473
  );


  xnor
  g486
  (
    n584,
    n464,
    n486,
    n281,
    n473
  );


  xnor
  g487
  (
    n673,
    n175,
    n151,
    n283,
    n453
  );


  and
  g488
  (
    n769,
    n32,
    n398,
    n396,
    n254
  );


  and
  g489
  (
    n752,
    n234,
    n32,
    n485,
    n253
  );


  xor
  g490
  (
    n608,
    n486,
    n434,
    n502,
    n409
  );


  and
  g491
  (
    n681,
    n430,
    n431,
    n465,
    n370
  );


  xor
  g492
  (
    n863,
    n481,
    n401,
    n461,
    n483
  );


  xor
  g493
  (
    n756,
    n156,
    n287,
    n351,
    n338
  );


  and
  g494
  (
    n799,
    n305,
    n285,
    n395,
    n295
  );


  or
  g495
  (
    n663,
    n491,
    n487,
    n368,
    n346
  );


  or
  g496
  (
    n619,
    n335,
    n498,
    n200,
    n161
  );


  xor
  g497
  (
    n711,
    n250,
    n291,
    n408,
    n350
  );


  and
  g498
  (
    n525,
    n219,
    n413,
    n358,
    n199
  );


  or
  g499
  (
    n755,
    n258,
    n252,
    n427,
    n407
  );


  xor
  g500
  (
    n821,
    n215,
    n349,
    n288,
    n144
  );


  or
  g501
  (
    n874,
    n132,
    n393,
    n312,
    n353
  );


  nand
  g502
  (
    n658,
    n484,
    n231,
    n338,
    n171
  );


  xor
  g503
  (
    n792,
    n165,
    n217,
    n234,
    n466
  );


  xor
  g504
  (
    n568,
    n323,
    n454,
    n306,
    n313
  );


  and
  g505
  (
    n677,
    n248,
    n329,
    n449,
    n241
  );


  xor
  g506
  (
    KeyWire_0_26,
    n136,
    n181,
    n330,
    n501
  );


  xor
  g507
  (
    n871,
    n386,
    n456,
    n275,
    n241
  );


  xor
  g508
  (
    n807,
    n491,
    n216,
    n218,
    n484
  );


  nor
  g509
  (
    n870,
    n209,
    n438,
    n161,
    n328
  );


  nor
  g510
  (
    n665,
    n422,
    n296,
    n419,
    n186
  );


  or
  g511
  (
    n879,
    n427,
    n193,
    n212,
    n505
  );


  or
  g512
  (
    n586,
    n255,
    n343,
    n379,
    n384
  );


  nor
  g513
  (
    n782,
    n176,
    n355,
    n429,
    n172
  );


  and
  g514
  (
    n827,
    n319,
    n433,
    n475,
    n268
  );


  xor
  g515
  (
    n788,
    n413,
    n464,
    n426,
    n390
  );


  nand
  g516
  (
    n594,
    n170,
    n259,
    n381,
    n178
  );


  nor
  g517
  (
    n614,
    n296,
    n441,
    n247,
    n142
  );


  nor
  g518
  (
    n732,
    n501,
    n382,
    n446,
    n435
  );


  and
  g519
  (
    n790,
    n384,
    n457,
    n352,
    n250
  );


  nand
  g520
  (
    n723,
    n421,
    n290,
    n344,
    n141
  );


  xor
  g521
  (
    n580,
    n389,
    n332,
    n274,
    n170
  );


  nor
  g522
  (
    n552,
    n246,
    n319,
    n261,
    n150
  );


  xnor
  g523
  (
    n604,
    n230,
    n354,
    n399,
    n398
  );


  nor
  g524
  (
    n569,
    n301,
    n476,
    n287,
    n438
  );


  xor
  g525
  (
    n796,
    n389,
    n190,
    n484,
    n184
  );


  and
  g526
  (
    n704,
    n141,
    n205,
    n262,
    n460
  );


  and
  g527
  (
    n545,
    n273,
    n221,
    n392,
    n475
  );


  nor
  g528
  (
    n589,
    n264,
    n479,
    n457,
    n207
  );


  or
  g529
  (
    n612,
    n225,
    n214,
    n277,
    n323
  );


  nand
  g530
  (
    n777,
    n242,
    n259,
    n186,
    n314
  );


  or
  g531
  (
    n726,
    n306,
    n134,
    n316,
    n392
  );


  and
  g532
  (
    n578,
    n415,
    n209,
    n240,
    n136
  );


  nor
  g533
  (
    n798,
    n208,
    n439,
    n165,
    n251
  );


  and
  g534
  (
    n536,
    n296,
    n368,
    n250,
    n315
  );


  nor
  g535
  (
    n558,
    n412,
    n396,
    n496,
    n439
  );


  xnor
  g536
  (
    n676,
    n238,
    n426,
    n234,
    n265
  );


  or
  g537
  (
    n808,
    n423,
    n308,
    n244,
    n220
  );


  xor
  g538
  (
    n795,
    n242,
    n339,
    n239,
    n188
  );


  nand
  g539
  (
    n715,
    n492,
    n266,
    n135,
    n197
  );


  nand
  g540
  (
    n877,
    n364,
    n440,
    n495,
    n150
  );


  or
  g541
  (
    n735,
    n337,
    n193,
    n244,
    n411
  );


  xor
  g542
  (
    n564,
    n329,
    n494,
    n291,
    n194
  );


  nand
  g543
  (
    n836,
    n437,
    n279,
    n195,
    n429
  );


  xnor
  g544
  (
    n518,
    n315,
    n276,
    n159,
    n389
  );


  xnor
  g545
  (
    n844,
    n385,
    n192,
    n365,
    n403
  );


  nor
  g546
  (
    n856,
    n299,
    n391,
    n212,
    n312
  );


  nor
  g547
  (
    n738,
    n491,
    n276,
    n376,
    n315
  );


  xor
  g548
  (
    n534,
    n459,
    n239,
    n341,
    n222
  );


  xor
  g549
  (
    n826,
    n461,
    n412,
    n321,
    n353
  );


  xnor
  g550
  (
    n590,
    n324,
    n456,
    n274,
    n487
  );


  xnor
  g551
  (
    n760,
    n154,
    n374,
    n357,
    n421
  );


  nand
  g552
  (
    n764,
    n320,
    n323,
    n423,
    n395
  );


  xnor
  g553
  (
    n631,
    n481,
    n441,
    n478,
    n424
  );


  nand
  g554
  (
    n862,
    n140,
    n291,
    n295,
    n134
  );


  nor
  g555
  (
    n779,
    n278,
    n145,
    n361,
    n294
  );


  xnor
  g556
  (
    n532,
    n180,
    n206,
    n317,
    n416
  );


  nand
  g557
  (
    n717,
    n448,
    n442,
    n284,
    n193
  );


  nor
  g558
  (
    n630,
    n474,
    n298,
    n428,
    n354
  );


  or
  g559
  (
    n579,
    n156,
    n281,
    n190,
    n299
  );


  xnor
  g560
  (
    n588,
    n135,
    n210,
    n318,
    n495
  );


  nor
  g561
  (
    n739,
    n266,
    n294,
    n350,
    n311
  );


  nor
  g562
  (
    n875,
    n211,
    n493,
    n452,
    n181
  );


  nand
  g563
  (
    n794,
    n320,
    n248,
    n274,
    n451
  );


  xnor
  g564
  (
    n650,
    n282,
    n257,
    n353,
    n154
  );


  xnor
  g565
  (
    n621,
    n431,
    n162,
    n209,
    n253
  );


  xnor
  g566
  (
    n867,
    n201,
    n422,
    n181,
    n478
  );


  or
  g567
  (
    n637,
    n290,
    n204,
    n394,
    n200
  );


  and
  g568
  (
    n694,
    n198,
    n442,
    n499
  );


  nand
  g569
  (
    n617,
    n416,
    n492,
    n154,
    n399
  );


  nor
  g570
  (
    n709,
    n424,
    n359,
    n275,
    n218
  );


  xor
  g571
  (
    n664,
    n280,
    n179,
    n467,
    n171
  );


  xnor
  g572
  (
    n696,
    n450,
    n294,
    n233,
    n286
  );


  and
  g573
  (
    n705,
    n260,
    n177,
    n402,
    n221
  );


  or
  g574
  (
    n698,
    n400,
    n305,
    n295,
    n169
  );


  xor
  g575
  (
    n841,
    n288,
    n357,
    n369,
    n381
  );


  and
  g576
  (
    n817,
    n501,
    n397,
    n250,
    n358
  );


  xnor
  g577
  (
    n753,
    n329,
    n394,
    n504,
    n373
  );


  nor
  g578
  (
    n859,
    n139,
    n147,
    n427,
    n356
  );


  nand
  g579
  (
    n659,
    n228,
    n310,
    n374,
    n251
  );


  nand
  g580
  (
    n649,
    n190,
    n140,
    n161,
    n325
  );


  xnor
  g581
  (
    n749,
    n193,
    n206,
    n225,
    n273
  );


  xor
  g582
  (
    n866,
    n419,
    n187,
    n416,
    n417
  );


  xnor
  g583
  (
    KeyWire_0_17,
    n367,
    n380,
    n192,
    n254
  );


  or
  g584
  (
    n600,
    n505,
    n175,
    n439,
    n445
  );


  nor
  g585
  (
    n577,
    n257,
    n199,
    n363,
    n160
  );


  nand
  g586
  (
    n574,
    n159,
    n196,
    n178,
    n333
  );


  nor
  g587
  (
    n759,
    n202,
    n374,
    n381,
    n383
  );


  or
  g588
  (
    n561,
    n269,
    n447,
    n489,
    n371
  );


  nand
  g589
  (
    n666,
    n366,
    n421,
    n349,
    n372
  );


  xor
  g590
  (
    n731,
    n500,
    n406,
    n229,
    n147
  );


  and
  g591
  (
    n791,
    n247,
    n267,
    n322,
    n157
  );


  and
  g592
  (
    KeyWire_0_40,
    n313,
    n453,
    n149,
    n190
  );


  xnor
  g593
  (
    n567,
    n300,
    n454,
    n468,
    n333
  );


  and
  g594
  (
    n685,
    n226,
    n505,
    n367,
    n366
  );


  nand
  g595
  (
    n529,
    n332,
    n311,
    n499,
    n360
  );


  xnor
  g596
  (
    n776,
    n211,
    n169,
    n349,
    n449
  );


  nor
  g597
  (
    n849,
    n189,
    n430,
    n146,
    n488
  );


  or
  g598
  (
    n623,
    n486,
    n248,
    n341,
    n348
  );


  nor
  g599
  (
    n797,
    n340,
    n138,
    n169,
    n436
  );


  nand
  g600
  (
    n846,
    n242,
    n207,
    n362,
    n479
  );


  or
  g601
  (
    n830,
    n471,
    n245,
    n463,
    n203
  );


  xor
  g602
  (
    n720,
    n151,
    n461,
    n394,
    n285
  );


  nor
  g603
  (
    n691,
    n203,
    n503,
    n277,
    n463
  );


  or
  g604
  (
    n716,
    n286,
    n298,
    n191,
    n443
  );


  nor
  g605
  (
    n842,
    n263,
    n182,
    n335,
    n314
  );


  xor
  g606
  (
    n713,
    n304,
    n365,
    n271,
    n236
  );


  or
  g607
  (
    n642,
    n376,
    n346,
    n275,
    n496
  );


  xor
  g608
  (
    n810,
    n497,
    n339,
    n463,
    n180
  );


  xor
  g609
  (
    n686,
    n183,
    n153,
    n148,
    n502
  );


  xor
  g610
  (
    n550,
    n470,
    n173,
    n167,
    n251
  );


  nand
  g611
  (
    n628,
    n379,
    n358,
    n285,
    n377
  );


  nand
  g612
  (
    n747,
    n398,
    n343,
    n267,
    n484
  );


  xnor
  g613
  (
    n850,
    n330,
    n303,
    n222,
    n208
  );


  xor
  g614
  (
    n876,
    n195,
    n153,
    n423
  );


  and
  g615
  (
    n662,
    n297,
    n266,
    n476,
    n284
  );


  or
  g616
  (
    n690,
    n339,
    n478,
    n459,
    n441
  );


  xor
  g617
  (
    n783,
    n246,
    n290,
    n346,
    n277
  );


  and
  g618
  (
    n554,
    n493,
    n405,
    n375,
    n155
  );


  and
  g619
  (
    n603,
    n502,
    n217,
    n198,
    n254
  );


  or
  g620
  (
    n657,
    n213,
    n362,
    n229,
    n233
  );


  nand
  g621
  (
    n766,
    n179,
    n372,
    n292,
    n237
  );


  xor
  g622
  (
    n743,
    n191,
    n437,
    n404,
    n236
  );


  or
  g623
  (
    n718,
    n462,
    n448,
    n378,
    n418
  );


  xnor
  g624
  (
    n632,
    n401,
    n150,
    n213,
    n142
  );


  or
  g625
  (
    n535,
    n353,
    n224,
    n481,
    n319
  );


  xor
  g626
  (
    n660,
    n287,
    n292,
    n324,
    n326
  );


  and
  g627
  (
    n672,
    n264,
    n282,
    n394,
    n246
  );


  nor
  g628
  (
    n805,
    n407,
    n405,
    n380,
    n474
  );


  and
  g629
  (
    n814,
    n359,
    n306,
    n246,
    n155
  );


  and
  g630
  (
    n671,
    n280,
    n435,
    n376,
    n344
  );


  and
  g631
  (
    n888,
    n430,
    n356,
    n379,
    n210
  );


  nand
  g632
  (
    KeyWire_0_37,
    n205,
    n328,
    n399
  );


  or
  g633
  (
    n884,
    n342,
    n278,
    n195,
    n317
  );


  or
  g634
  (
    n835,
    n406,
    n335,
    n348
  );


  nand
  g635
  (
    n889,
    n406,
    n256,
    n320,
    n196
  );


  nand
  g636
  (
    n670,
    n139,
    n194,
    n503,
    n153
  );


  xnor
  g637
  (
    n724,
    n407,
    n312,
    n163,
    n152
  );


  nand
  g638
  (
    n573,
    n171,
    n396,
    n176,
    n488
  );


  nand
  g639
  (
    n523,
    n334,
    n479,
    n492,
    n368
  );


  xor
  g640
  (
    n640,
    n339,
    n377,
    n361,
    n408
  );


  nor
  g641
  (
    n627,
    n386,
    n228,
    n216,
    n185
  );


  or
  g642
  (
    n736,
    n462,
    n219,
    n362,
    n387
  );


  and
  g643
  (
    n887,
    n223,
    n241,
    n254,
    n466
  );


  and
  g644
  (
    n750,
    n418,
    n274,
    n428,
    n443
  );


  or
  g645
  (
    n643,
    n160,
    n331,
    n375,
    n366
  );


  xor
  g646
  (
    n598,
    n336,
    n308,
    n229,
    n480
  );


  xnor
  g647
  (
    n881,
    n471,
    n312,
    n245,
    n300
  );


  or
  g648
  (
    n800,
    n456,
    n184,
    n351,
    n379
  );


  nor
  g649
  (
    n772,
    n204,
    n414,
    n373,
    n393
  );


  xor
  g650
  (
    n634,
    n257,
    n420,
    n504,
    n302
  );


  and
  g651
  (
    n644,
    n331,
    n337,
    n304,
    n260
  );


  or
  g652
  (
    n745,
    n249,
    n397,
    n448,
    n227
  );


  nor
  g653
  (
    n572,
    n206,
    n336,
    n277,
    n320
  );


  xnor
  g654
  (
    n785,
    n223,
    n347,
    n364,
    n345
  );


  and
  g655
  (
    KeyWire_0_61,
    n404,
    n241,
    n467,
    n410
  );


  and
  g656
  (
    n857,
    n478,
    n326,
    n294,
    n380
  );


  xor
  g657
  (
    n780,
    n460,
    n450,
    n360,
    n233
  );


  nand
  g658
  (
    n751,
    n133,
    n158,
    n428,
    n259
  );


  or
  g659
  (
    n865,
    n201,
    n408,
    n252,
    n504
  );


  and
  g660
  (
    n539,
    n436,
    n386,
    n382
  );


  xor
  g661
  (
    n609,
    n480,
    n482,
    n227,
    n269
  );


  nand
  g662
  (
    n565,
    n403,
    n367,
    n146,
    n497
  );


  and
  g663
  (
    n563,
    n281,
    n474,
    n191,
    n258
  );


  xnor
  g664
  (
    n748,
    n454,
    n388,
    n148,
    n472
  );


  xnor
  g665
  (
    n812,
    n181,
    n350,
    n301,
    n497
  );


  and
  g666
  (
    n542,
    n166,
    n143,
    n223,
    n468
  );


  and
  g667
  (
    n730,
    n222,
    n414,
    n365,
    n483
  );


  and
  g668
  (
    n530,
    n186,
    n140,
    n235,
    n411
  );


  or
  g669
  (
    n754,
    n302,
    n458,
    n423,
    n232
  );


  and
  g670
  (
    n597,
    n268,
    n372,
    n226,
    n391
  );


  xor
  g671
  (
    KeyWire_0_36,
    n228,
    n170,
    n402,
    n152
  );


  or
  g672
  (
    n543,
    n315,
    n227,
    n201,
    n162
  );


  or
  g673
  (
    n585,
    n272,
    n362,
    n437,
    n239
  );


  and
  g674
  (
    n703,
    n213,
    n455,
    n318,
    n397
  );


  xnor
  g675
  (
    n576,
    n166,
    n269,
    n228,
    n462
  );


  or
  g676
  (
    n684,
    n276,
    n243,
    n472,
    n385
  );


  nand
  g677
  (
    n773,
    n223,
    n187,
    n196,
    n341
  );


  or
  g678
  (
    n864,
    n231,
    n305,
    n377,
    n327
  );


  nor
  g679
  (
    n707,
    n372,
    n404,
    n426,
    n432
  );


  and
  g680
  (
    n652,
    n174,
    n331,
    n224,
    n436
  );


  and
  g681
  (
    n700,
    n165,
    n477,
    n331,
    n345
  );


  xnor
  g682
  (
    n728,
    n316,
    n413,
    n200,
    n210
  );


  nand
  g683
  (
    n555,
    n163,
    n470,
    n137,
    n468
  );


  nand
  g684
  (
    n633,
    n185,
    n264,
    n143,
    n446
  );


  or
  g685
  (
    n626,
    n425,
    n249,
    n240,
    n279
  );


  xor
  g686
  (
    n768,
    n270,
    n400,
    n252,
    n260
  );


  and
  g687
  (
    n823,
    n197,
    n347,
    n490,
    n307
  );


  xor
  g688
  (
    n647,
    n168,
    n297,
    n261,
    n350
  );


  nor
  g689
  (
    n522,
    n238,
    n502,
    n290,
    n235
  );


  and
  g690
  (
    n692,
    n425,
    n488,
    n400,
    n480
  );


  and
  g691
  (
    n714,
    n158,
    n152,
    n332,
    n392
  );


  xnor
  g692
  (
    n837,
    n160,
    n177,
    n265,
    n383
  );


  xnor
  g693
  (
    n721,
    n206,
    n272,
    n238,
    n235
  );


  and
  g694
  (
    n787,
    n326,
    n214,
    n225,
    n215
  );


  nand
  g695
  (
    n667,
    n413,
    n377,
    n470,
    n163
  );


  xor
  g696
  (
    n547,
    n437,
    n205,
    n279,
    n433
  );


  xor
  g697
  (
    n834,
    n305,
    n32,
    n224,
    n146
  );


  xor
  g698
  (
    n591,
    n336,
    n134,
    n297,
    n286
  );


  xnor
  g699
  (
    n702,
    n370,
    n319,
    n189,
    n308
  );


  and
  g700
  (
    n806,
    n230,
    n187,
    n383,
    n174
  );


  and
  g701
  (
    n734,
    n232,
    n325,
    n279,
    n169
  );


  and
  g702
  (
    n813,
    n485,
    n141,
    n395,
    n182
  );


  nand
  g703
  (
    n757,
    n168,
    n179,
    n393,
    n201
  );


  nor
  g704
  (
    n582,
    n402,
    n355,
    n195,
    n203
  );


  and
  g705
  (
    n854,
    n433,
    n221,
    n219,
    n261
  );


  xnor
  g706
  (
    n521,
    n161,
    n432,
    n449,
    n462
  );


  xnor
  g707
  (
    n740,
    n445,
    n340,
    n272,
    n156
  );


  and
  g708
  (
    n688,
    n405,
    n282,
    n293,
    n429
  );


  xor
  g709
  (
    n669,
    n386,
    n168,
    n327,
    n335
  );


  and
  g710
  (
    n562,
    n454,
    n301,
    n155,
    n184
  );


  nand
  g711
  (
    n595,
    n184,
    n288,
    n232,
    n442
  );


  nor
  g712
  (
    n638,
    n457,
    n260,
    n409,
    n450
  );


  xnor
  g713
  (
    n706,
    n378,
    n135,
    n343,
    n271
  );


  nand
  g714
  (
    n741,
    n417,
    n474,
    n218,
    n316
  );


  xnor
  g715
  (
    n725,
    n337,
    n273,
    n412,
    n258
  );


  and
  g716
  (
    n828,
    n493,
    n482,
    n267,
    n301
  );


  nor
  g717
  (
    n775,
    n435,
    n450,
    n496,
    n348
  );


  nand
  g718
  (
    n699,
    n194,
    n180,
    n328,
    n284
  );


  xnor
  g719
  (
    n839,
    n152,
    n197,
    n480,
    n194
  );


  and
  g720
  (
    n538,
    n451,
    n180,
    n466,
    n200
  );


  nor
  g721
  (
    n528,
    n286,
    n472,
    n459,
    n420
  );


  nor
  g722
  (
    KeyWire_0_0,
    n455,
    n154,
    n485,
    n148
  );


  xor
  g723
  (
    n802,
    n489,
    n183,
    n266,
    n495
  );


  xnor
  g724
  (
    n646,
    n207,
    n475,
    n236,
    n342
  );


  and
  g725
  (
    KeyWire_0_46,
    n162,
    n483,
    n247,
    n292
  );


  nand
  g726
  (
    n654,
    n136,
    n258,
    n343,
    n188
  );


  xnor
  g727
  (
    n520,
    n453,
    n280,
    n473,
    n177
  );


  xnor
  g728
  (
    n548,
    n396,
    n333,
    n498,
    n291
  );


  xor
  g729
  (
    n765,
    n464,
    n458,
    n360,
    n355
  );


  xnor
  g730
  (
    n804,
    n270,
    n345,
    n492,
    n313
  );


  xor
  g731
  (
    n639,
    n408,
    n230,
    n164,
    n363
  );


  or
  g732
  (
    n687,
    n136,
    n324,
    n476,
    n431
  );


  and
  g733
  (
    n678,
    n469,
    n202,
    n263,
    n415
  );


  or
  g734
  (
    n853,
    n418,
    n387,
    n308,
    n442
  );


  or
  g735
  (
    n722,
    n278,
    n445,
    n148,
    n321
  );


  xnor
  g736
  (
    n596,
    n321,
    n346,
    n340,
    n378
  );


  nor
  g737
  (
    n625,
    n139,
    n160,
    n392,
    n493
  );


  xnor
  g738
  (
    n829,
    n333,
    n202,
    n429,
    n256
  );


  nand
  g739
  (
    n803,
    n164,
    n483,
    n296,
    n459
  );


  nand
  g740
  (
    n601,
    n375,
    n357,
    n411,
    n222
  );


  xnor
  g741
  (
    n832,
    n334,
    n163,
    n397,
    n133
  );


  nand
  g742
  (
    n712,
    n330,
    n342,
    n133,
    n419
  );


  or
  g743
  (
    n855,
    n310,
    n192,
    n173,
    n457
  );


  xnor
  g744
  (
    n742,
    n440,
    n204,
    n167,
    n182
  );


  nand
  g745
  (
    n575,
    n303,
    n391,
    n311,
    n262
  );


  and
  g746
  (
    n682,
    n232,
    n470,
    n500,
    n272
  );


  xnor
  g747
  (
    n524,
    n307,
    n385,
    n354,
    n426
  );


  or
  g748
  (
    n587,
    n382,
    n401,
    n151,
    n300
  );


  and
  g749
  (
    n843,
    n289,
    n226,
    n142,
    n425
  );


  xor
  g750
  (
    n820,
    n448,
    n309,
    n271
  );


  xor
  g751
  (
    n533,
    n456,
    n468,
    n488,
    n498
  );


  xnor
  g752
  (
    n519,
    n336,
    n490,
    n210,
    n371
  );


  or
  g753
  (
    n549,
    n225,
    n187,
    n302,
    n469
  );


  nand
  g754
  (
    n570,
    n310,
    n438,
    n482,
    n220
  );


  nor
  g755
  (
    n541,
    n477,
    n421,
    n257,
    n352
  );


  nand
  g756
  (
    n761,
    n175,
    n216,
    n356,
    n245
  );


  or
  g757
  (
    n620,
    n255,
    n32,
    n388,
    n422
  );


  nor
  g758
  (
    n559,
    n419,
    n189,
    n402,
    n309
  );


  xor
  g759
  (
    n635,
    n217,
    n434,
    n487,
    n139
  );


  and
  g760
  (
    n833,
    n142,
    n143,
    n316,
    n255
  );


  xor
  g761
  (
    n708,
    n440,
    n158,
    n289,
    n354
  );


  nor
  g762
  (
    n885,
    n269,
    n494,
    n293,
    n455
  );


  xor
  g763
  (
    n544,
    n157,
    n176,
    n159,
    n303
  );


  nor
  g764
  (
    n873,
    n446,
    n412,
    n164,
    n414
  );


  xor
  g765
  (
    n815,
    n496,
    n283,
    n149,
    n268
  );


  nand
  g766
  (
    n824,
    n172,
    n326,
    n170,
    n183
  );


  nor
  g767
  (
    n697,
    n275,
    n133,
    n145,
    n398
  );


  nand
  g768
  (
    n701,
    n376,
    n174,
    n229,
    n334
  );


  or
  g769
  (
    n551,
    n431,
    n461,
    n345,
    n263
  );


  nand
  g770
  (
    n872,
    n436,
    n297,
    n146,
    n391
  );


  xnor
  g771
  (
    n571,
    n490,
    n317,
    n451,
    n282
  );


  and
  g772
  (
    n583,
    n243,
    n449,
    n158,
    n417
  );


  nand
  g773
  (
    n848,
    n247,
    n439,
    n490,
    n216
  );


  and
  g774
  (
    n847,
    n197,
    n381,
    n435,
    n504
  );


  nor
  g775
  (
    n683,
    n466,
    n341,
    n473,
    n443
  );


  xor
  g776
  (
    n852,
    n366,
    n447,
    n293,
    n298
  );


  nor
  g777
  (
    n546,
    n471,
    n157,
    n185,
    n368
  );


  nor
  g778
  (
    n786,
    n369,
    n378,
    n351,
    n310
  );


  xnor
  g779
  (
    n653,
    n441,
    n159,
    n263,
    n401
  );


  and
  g780
  (
    n605,
    n481,
    n179,
    n298,
    n140
  );


  and
  g781
  (
    n858,
    n347,
    n231,
    n218,
    n409
  );


  nand
  g782
  (
    n606,
    n403,
    n245,
    n156,
    n469
  );


  xor
  g783
  (
    n599,
    n444,
    n302,
    n268,
    n318
  );


  nand
  g784
  (
    n793,
    n292,
    n178,
    n410,
    n342
  );


  nor
  g785
  (
    n641,
    n213,
    n207,
    n344,
    n162
  );


  and
  g786
  (
    n655,
    n145,
    n371,
    n271,
    n249
  );


  and
  g787
  (
    n733,
    n264,
    n214,
    n338,
    n485
  );


  or
  g788
  (
    n622,
    n325,
    n498,
    n464,
    n373
  );


  xor
  g789
  (
    n811,
    n172,
    n211,
    n373,
    n198
  );


  xor
  g790
  (
    n616,
    n329,
    n463,
    n243,
    n198
  );


  and
  g791
  (
    n729,
    n414,
    n425,
    n355,
    n303
  );


  nand
  g792
  (
    n615,
    n205,
    n265,
    n239,
    n472
  );


  or
  g793
  (
    n557,
    n237,
    n220,
    n221,
    n240
  );


  nand
  g794
  (
    n758,
    n400,
    n364,
    n233,
    n325
  );


  and
  g795
  (
    n851,
    n288,
    n452,
    n361,
    n167
  );


  or
  g796
  (
    n593,
    n384,
    n293,
    n388,
    n467
  );


  xnor
  g797
  (
    n556,
    n224,
    n357,
    n327,
    n183
  );


  nand
  g798
  (
    n727,
    n500,
    n383,
    n270,
    n489
  );


  xnor
  g799
  (
    n679,
    n323,
    n359,
    n452,
    n157
  );


  or
  g800
  (
    n868,
    n141,
    n307,
    n188,
    n235
  );


  or
  g801
  (
    n801,
    n166,
    n192,
    n309,
    n395
  );


  xor
  g802
  (
    n560,
    n501,
    n410,
    n446,
    n447
  );


  nand
  g803
  (
    n693,
    n300,
    n191,
    n465,
    n428
  );


  xor
  g804
  (
    n674,
    n407,
    n208,
    n137,
    n167
  );


  xnor
  g805
  (
    n695,
    n262,
    n166,
    n199,
    n253
  );


  nand
  g806
  (
    n822,
    n243,
    n432,
    n322,
    n231
  );


  nor
  g807
  (
    n613,
    n403,
    n332,
    n491,
    n418
  );


  xor
  g808
  (
    n516,
    n318,
    n214,
    n365,
    n212
  );


  xnor
  g809
  (
    n763,
    n208,
    n363,
    n196,
    n138
  );


  nand
  g810
  (
    n689,
    n317,
    n364,
    n367,
    n255
  );


  and
  g811
  (
    n880,
    n283,
    n424,
    n202,
    n338
  );


  nand
  g812
  (
    n831,
    n287,
    n253,
    n477,
    n352
  );


  nand
  g813
  (
    n818,
    n322,
    n322,
    n334,
    n434
  );


  xnor
  g814
  (
    n668,
    n495,
    n227,
    n289,
    n280
  );


  nor
  g815
  (
    n592,
    n299,
    n145,
    n237,
    n234
  );


  nor
  g816
  (
    n636,
    n445,
    n244,
    n138,
    n369
  );


  or
  g817
  (
    n767,
    n203,
    n344,
    n416,
    n330
  );


  nor
  g818
  (
    n789,
    n285,
    n447,
    n240,
    n410
  );


  xor
  g819
  (
    n675,
    n256,
    n209,
    n307,
    n143
  );


  or
  g820
  (
    n566,
    n393,
    n503,
    n420,
    n390
  );


  and
  g821
  (
    n656,
    n409,
    n176,
    n321,
    n173
  );


  xnor
  g822
  (
    n770,
    n164,
    n134,
    n273,
    n144
  );


  xnor
  g823
  (
    n526,
    n369,
    n211,
    n415,
    n311
  );


  xnor
  g824
  (
    n840,
    n304,
    n283,
    n351,
    n487
  );


  xor
  g825
  (
    n553,
    n284,
    n174,
    n261,
    n144
  );


  xor
  g826
  (
    n774,
    n237,
    n389,
    n199,
    n173
  );


  xnor
  g827
  (
    n710,
    n168,
    n324,
    n380,
    n177
  );


  and
  g828
  (
    n537,
    n147,
    n188,
    n259,
    n370
  );


  or
  g829
  (
    n602,
    n149,
    n385,
    n172,
    n443
  );


  and
  g830
  (
    n618,
    n444,
    n276,
    n217,
    n278
  );


  and
  g831
  (
    n771,
    n455,
    n438,
    n149,
    n453
  );


  nor
  g832
  (
    n838,
    n359,
    n186,
    n444,
    n352
  );


  xor
  g833
  (
    n624,
    n433,
    n249,
    n356,
    n189
  );


  xnor
  g834
  (
    n882,
    n390,
    n256,
    n304,
    n503
  );


  nand
  g835
  (
    n611,
    n458,
    n251,
    n361,
    n252
  );


  or
  g836
  (
    n746,
    n137,
    n226,
    n151,
    n185
  );


  xnor
  g837
  (
    n861,
    n314,
    n248,
    n363,
    n390
  );


  and
  g838
  (
    n581,
    n165,
    n360,
    n424,
    n451
  );


  xor
  g839
  (
    n762,
    n494,
    n458,
    n465,
    n135
  );


  or
  g840
  (
    n878,
    n155,
    n242,
    n471,
    n387
  );


  xor
  g841
  (
    n531,
    n500,
    n406,
    n265,
    n489
  );


  nand
  g842
  (
    n645,
    n444,
    n452,
    n182,
    n486
  );


  nor
  g843
  (
    n629,
    n494,
    n399,
    n215,
    n270
  );


  xnor
  g844
  (
    n825,
    n404,
    n138,
    n175,
    n476
  );


  nor
  g845
  (
    n784,
    n430,
    n314,
    n440,
    n220
  );


  and
  g846
  (
    n648,
    n384,
    n299,
    n358,
    n469
  );


  xor
  g847
  (
    n661,
    n244,
    n479,
    n215,
    n236
  );


  xor
  g848
  (
    n869,
    n477,
    n499,
    n387,
    n417
  );


  xnor
  g849
  (
    n860,
    n467,
    n204,
    n347,
    n411
  );


  xor
  g850
  (
    n680,
    n374,
    n212,
    n375,
    n313
  );


  or
  g851
  (
    n540,
    n422,
    n230,
    n460,
    n497
  );


  and
  g852
  (
    n819,
    n171,
    n178,
    n219,
    n306
  );


  and
  g853
  (
    n778,
    n434,
    n281,
    n337,
    n388
  );


  or
  g854
  (
    n719,
    n460,
    n415,
    n482,
    n267
  );


  xnor
  g855
  (
    n610,
    n150,
    n238,
    n289,
    n340
  );


  nor
  g856
  (
    n737,
    n327,
    n144,
    n370,
    n147
  );


  and
  g857
  (
    n890,
    n534,
    n533
  );


  or
  g858
  (
    n891,
    n535,
    n537,
    n890,
    n536
  );


  and
  g859
  (
    n894,
    n545,
    n543,
    n548,
    n547
  );


  and
  g860
  (
    n895,
    n549,
    n891
  );


  and
  g861
  (
    n892,
    n538,
    n540,
    n891,
    n544
  );


  or
  g862
  (
    n893,
    n542,
    n539,
    n541,
    n546
  );


  not
  g863
  (
    n905,
    n892
  );


  not
  g864
  (
    n899,
    n893
  );


  not
  g865
  (
    n897,
    n894
  );


  not
  g866
  (
    n896,
    n895
  );


  buf
  g867
  (
    n901,
    n895
  );


  not
  g868
  (
    n898,
    n894
  );


  buf
  g869
  (
    n904,
    n893
  );


  buf
  g870
  (
    n902,
    n894
  );


  buf
  g871
  (
    n900,
    n892
  );


  xnor
  g872
  (
    n903,
    n895,
    n550
  );


  nor
  g873
  (
    n941,
    n584,
    n598,
    n611,
    n592
  );


  and
  g874
  (
    n930,
    n599,
    n897,
    n902,
    n898
  );


  xnor
  g875
  (
    n933,
    n585,
    n613,
    n596,
    n555
  );


  nand
  g876
  (
    n912,
    n582,
    n603,
    n598,
    n557
  );


  nor
  g877
  (
    n923,
    n903,
    n612,
    n567,
    n900
  );


  and
  g878
  (
    n931,
    n615,
    n903,
    n905,
    n588
  );


  nand
  g879
  (
    n932,
    n583,
    n591,
    n593,
    n610
  );


  nor
  g880
  (
    n920,
    n569,
    n901,
    n604,
    n898
  );


  xor
  g881
  (
    n906,
    n589,
    n583,
    n600,
    n610
  );


  or
  g882
  (
    n919,
    n595,
    n582,
    n586,
    n620
  );


  or
  g883
  (
    n915,
    n899,
    n587,
    n901,
    n565
  );


  or
  g884
  (
    n925,
    n601,
    n616,
    n580
  );


  or
  g885
  (
    n909,
    n618,
    n589,
    n896,
    n904
  );


  or
  g886
  (
    n935,
    n578,
    n572,
    n904,
    n599
  );


  xor
  g887
  (
    n910,
    n623,
    n898,
    n905,
    n619
  );


  and
  g888
  (
    n908,
    n562,
    n614,
    n896,
    n570
  );


  nand
  g889
  (
    n942,
    n553,
    n617,
    n560,
    n602
  );


  or
  g890
  (
    n924,
    n612,
    n593,
    n600,
    n579
  );


  or
  g891
  (
    KeyWire_0_55,
    n621,
    n897,
    n609,
    n575
  );


  xor
  g892
  (
    n926,
    n903,
    n605,
    n556,
    n601
  );


  xnor
  g893
  (
    n945,
    n618,
    n606,
    n622,
    n571
  );


  nand
  g894
  (
    n927,
    n591,
    n579,
    n590,
    n902
  );


  and
  g895
  (
    n914,
    n898,
    n606,
    n551,
    n559
  );


  or
  g896
  (
    n943,
    n620,
    n904,
    n619,
    n614
  );


  nor
  g897
  (
    n936,
    n896,
    n581,
    n613,
    n597
  );


  xnor
  g898
  (
    n939,
    n564,
    n576,
    n902,
    n585
  );


  or
  g899
  (
    n929,
    n901,
    n568,
    n899,
    n597
  );


  xor
  g900
  (
    n911,
    n615,
    n899,
    n578,
    n609
  );


  xnor
  g901
  (
    n928,
    n573,
    n577,
    n607,
    n900
  );


  nand
  g902
  (
    n917,
    n584,
    n901,
    n899,
    n897
  );


  nand
  g903
  (
    n913,
    n590,
    n587,
    n594,
    n611
  );


  and
  g904
  (
    n918,
    n602,
    n617,
    n904,
    n581
  );


  xor
  g905
  (
    n916,
    n577,
    n607,
    n905,
    n552
  );


  xnor
  g906
  (
    n938,
    n900,
    n902,
    n897,
    n586
  );


  xnor
  g907
  (
    n934,
    n596,
    n903,
    n621,
    n566
  );


  or
  g908
  (
    n907,
    n554,
    n900,
    n905,
    n605
  );


  or
  g909
  (
    n937,
    n603,
    n616,
    n558,
    n608
  );


  xnor
  g910
  (
    n944,
    n574,
    n604,
    n561,
    n896
  );


  nand
  g911
  (
    n921,
    n563,
    n594,
    n595,
    n592
  );


  nor
  g912
  (
    n940,
    n623,
    n622,
    n608,
    n588
  );


  and
  g913
  (
    n1078,
    n939,
    n725,
    n747,
    n788
  );


  and
  g914
  (
    n1063,
    n721,
    n934,
    n907,
    n738
  );


  or
  g915
  (
    n1091,
    n930,
    n913,
    n752,
    n918
  );


  xnor
  g916
  (
    n1104,
    n643,
    n781,
    n648,
    n924
  );


  or
  g917
  (
    n1014,
    n691,
    n673,
    n679,
    n632
  );


  nand
  g918
  (
    n1087,
    n708,
    n926,
    n653,
    n944
  );


  xor
  g919
  (
    n1101,
    n740,
    n762,
    n906,
    n774
  );


  nand
  g920
  (
    n1062,
    n777,
    n764,
    n756,
    n936
  );


  and
  g921
  (
    n1096,
    n705,
    n761,
    n684,
    n911
  );


  nand
  g922
  (
    n1054,
    n692,
    n693,
    n677,
    n758
  );


  or
  g923
  (
    n1073,
    n675,
    n663,
    n773,
    n654
  );


  nand
  g924
  (
    n983,
    n704,
    n659,
    n927,
    n733
  );


  nand
  g925
  (
    n1031,
    n774,
    n659,
    n760,
    n627
  );


  or
  g926
  (
    n1004,
    n728,
    n940,
    n944,
    n694
  );


  nor
  g927
  (
    n1035,
    n931,
    n752,
    n727
  );


  and
  g928
  (
    n965,
    n928,
    n639,
    n712,
    n933
  );


  and
  g929
  (
    n1055,
    n712,
    n733,
    n945,
    n748
  );


  xnor
  g930
  (
    n1013,
    n734,
    n655,
    n669,
    n664
  );


  xnor
  g931
  (
    n970,
    n923,
    n671,
    n702,
    n735
  );


  nand
  g932
  (
    n1043,
    n720,
    n678,
    n722,
    n641
  );


  xnor
  g933
  (
    n1030,
    n760,
    n627,
    n686,
    n937
  );


  xnor
  g934
  (
    n1081,
    n735,
    n763,
    n699,
    n939
  );


  xor
  g935
  (
    n1003,
    n686,
    n940,
    n647,
    n918
  );


  xor
  g936
  (
    n1069,
    n710,
    n715,
    n697,
    n911
  );


  nand
  g937
  (
    n975,
    n685,
    n731,
    n724,
    n790
  );


  xnor
  g938
  (
    n1077,
    n726,
    n650,
    n772,
    n679
  );


  or
  g939
  (
    n1008,
    n697,
    n649,
    n760,
    n775
  );


  and
  g940
  (
    n988,
    n681,
    n750,
    n722,
    n907
  );


  nand
  g941
  (
    n1097,
    n727,
    n756,
    n735,
    n694
  );


  and
  g942
  (
    n952,
    n921,
    n755,
    n753,
    n687
  );


  nor
  g943
  (
    n1079,
    n915,
    n941,
    n917,
    n762
  );


  nand
  g944
  (
    n1061,
    n689,
    n781,
    n652,
    n783
  );


  xor
  g945
  (
    n964,
    n684,
    n770,
    n701,
    n923
  );


  and
  g946
  (
    n977,
    n680,
    n914,
    n777,
    n909
  );


  or
  g947
  (
    n1011,
    n734,
    n674,
    n912,
    n636
  );


  or
  g948
  (
    n1056,
    n916,
    n938,
    n932,
    n778
  );


  nand
  g949
  (
    n1020,
    n787,
    n672,
    n709,
    n943
  );


  xnor
  g950
  (
    n1019,
    n782,
    n714,
    n934,
    n755
  );


  xnor
  g951
  (
    n1048,
    n633,
    n912,
    n911,
    n925
  );


  nand
  g952
  (
    n1095,
    n719,
    n755,
    n625,
    n713
  );


  xnor
  g953
  (
    n1088,
    n692,
    n786,
    n646,
    n728
  );


  nor
  g954
  (
    n1058,
    n932,
    n673,
    n703,
    n741
  );


  nand
  g955
  (
    n1037,
    n624,
    n912,
    n695,
    n908
  );


  or
  g956
  (
    n1100,
    n912,
    n917,
    n664,
    n688
  );


  nor
  g957
  (
    n966,
    n910,
    n729,
    n783,
    n745
  );


  and
  g958
  (
    n950,
    n939,
    n756,
    n906,
    n645
  );


  or
  g959
  (
    n1084,
    n906,
    n915,
    n665,
    n746
  );


  or
  g960
  (
    n1086,
    n697,
    n918,
    n683,
    n739
  );


  or
  g961
  (
    n987,
    n924,
    n753,
    n910,
    n649
  );


  nand
  g962
  (
    n999,
    n914,
    n685,
    n774,
    n687
  );


  xnor
  g963
  (
    n1082,
    n713,
    n925,
    n731,
    n921
  );


  or
  g964
  (
    n955,
    n738,
    n945,
    n757,
    n648
  );


  nand
  g965
  (
    n1049,
    n746,
    n754,
    n745,
    n769
  );


  xnor
  g966
  (
    n1015,
    n757,
    n909,
    n910,
    n941
  );


  or
  g967
  (
    n1006,
    n683,
    n908,
    n644,
    n767
  );


  xnor
  g968
  (
    n1093,
    n749,
    n710,
    n696,
    n701
  );


  and
  g969
  (
    n1072,
    n639,
    n681,
    n788,
    n624
  );


  xor
  g970
  (
    n1034,
    n692,
    n726,
    n917,
    n787
  );


  or
  g971
  (
    n974,
    n926,
    n768,
    n933,
    n784
  );


  nor
  g972
  (
    n1032,
    n687,
    n676,
    n938,
    n626
  );


  and
  g973
  (
    n1001,
    n754,
    n721,
    n695,
    n656
  );


  or
  g974
  (
    n1016,
    n928,
    n671,
    n738,
    n669
  );


  xnor
  g975
  (
    n1028,
    n933,
    n718,
    n906,
    n913
  );


  and
  g976
  (
    n1022,
    n675,
    n662,
    n945,
    n714
  );


  xor
  g977
  (
    n1017,
    n657,
    n922,
    n768,
    n700
  );


  nor
  g978
  (
    n1024,
    n772,
    n745,
    n942,
    n919
  );


  nand
  g979
  (
    n956,
    n695,
    n730,
    n723,
    n749
  );


  nand
  g980
  (
    n1036,
    n941,
    n748,
    n923,
    n712
  );


  and
  g981
  (
    n1105,
    n928,
    n935,
    n754,
    n936
  );


  and
  g982
  (
    n958,
    n909,
    n734,
    n927,
    n732
  );


  or
  g983
  (
    n1099,
    n653,
    n716,
    n920,
    n743
  );


  nor
  g984
  (
    n981,
    n629,
    n638,
    n625,
    n924
  );


  xor
  g985
  (
    n1044,
    n771,
    n646,
    n936,
    n707
  );


  and
  g986
  (
    n1040,
    n913,
    n776,
    n725,
    n682
  );


  nand
  g987
  (
    n978,
    n780,
    n929,
    n767,
    n751
  );


  xor
  g988
  (
    n1009,
    n634,
    n789,
    n742,
    n773
  );


  or
  g989
  (
    n954,
    n689,
    n678,
    n914,
    n702
  );


  nand
  g990
  (
    KeyWire_0_54,
    n660,
    n711,
    n666,
    n942
  );


  and
  g991
  (
    n1098,
    n661,
    n668,
    n706,
    n744
  );


  xor
  g992
  (
    n1065,
    n713,
    n664,
    n913,
    n704
  );


  nand
  g993
  (
    n962,
    n761,
    n667,
    n681,
    n643
  );


  nor
  g994
  (
    n1059,
    n743,
    n746,
    n909,
    n690
  );


  nor
  g995
  (
    n979,
    n736,
    n737,
    n654,
    n655
  );


  or
  g996
  (
    n1025,
    n660,
    n637,
    n940,
    n927
  );


  or
  g997
  (
    n1076,
    n652,
    n917,
    n709,
    n931
  );


  nor
  g998
  (
    n969,
    n736,
    n747,
    n705,
    n758
  );


  xor
  g999
  (
    n951,
    n672,
    n729,
    n717,
    n684
  );


  xor
  g1000
  (
    n1000,
    n698,
    n652,
    n709,
    n635
  );


  xor
  g1001
  (
    n957,
    n943,
    n934,
    n916,
    n724
  );


  xor
  g1002
  (
    n998,
    n677,
    n743,
    n922,
    n656
  );


  xor
  g1003
  (
    n1102,
    n931,
    n943,
    n789,
    n689
  );


  xnor
  g1004
  (
    n1057,
    n919,
    n908,
    n766,
    n626
  );


  and
  g1005
  (
    n1045,
    n766,
    n658,
    n929,
    n714
  );


  nor
  g1006
  (
    n973,
    n749,
    n628,
    n790,
    n915
  );


  and
  g1007
  (
    n1029,
    n767,
    n703,
    n634,
    n670
  );


  nor
  g1008
  (
    n1094,
    n744,
    n759,
    n727,
    n783
  );


  and
  g1009
  (
    n991,
    n726,
    n683,
    n662,
    n937
  );


  xnor
  g1010
  (
    n972,
    n724,
    n730,
    n665,
    n759
  );


  xor
  g1011
  (
    n990,
    n705,
    n706,
    n718,
    n742
  );


  nand
  g1012
  (
    n985,
    n744,
    n710,
    n930,
    n635
  );


  and
  g1013
  (
    n994,
    n930,
    n739,
    n700,
    n630
  );


  xor
  g1014
  (
    n1026,
    n700,
    n764,
    n944,
    n699
  );


  and
  g1015
  (
    n961,
    n721,
    n781,
    n764,
    n761
  );


  xnor
  g1016
  (
    n1046,
    n638,
    n670,
    n910,
    n711
  );


  nor
  g1017
  (
    n1005,
    n770,
    n720,
    n750,
    n628
  );


  nor
  g1018
  (
    n1027,
    n775,
    n667,
    n663,
    n650
  );


  xor
  g1019
  (
    n963,
    n790,
    n693,
    n660,
    n939
  );


  xor
  g1020
  (
    n1090,
    n785,
    n719,
    n716,
    n685
  );


  nand
  g1021
  (
    n984,
    n679,
    n779,
    n630
  );


  or
  g1022
  (
    n953,
    n702,
    n907,
    n908,
    n647
  );


  and
  g1023
  (
    n1042,
    n945,
    n658,
    n708,
    n911
  );


  or
  g1024
  (
    n949,
    n740,
    n640,
    n690,
    n686
  );


  nand
  g1025
  (
    n1068,
    n778,
    n923,
    n676,
    n747
  );


  xor
  g1026
  (
    n948,
    n935,
    n741,
    n920,
    n775
  );


  xor
  g1027
  (
    n1089,
    n650,
    n645,
    n642,
    n944
  );


  xnor
  g1028
  (
    KeyWire_0_52,
    n916,
    n631,
    n654,
    n732
  );


  xor
  g1029
  (
    n1085,
    n641,
    n653,
    n776,
    n920
  );


  nor
  g1030
  (
    n1067,
    n779,
    n707,
    n648,
    n914
  );


  nand
  g1031
  (
    n971,
    n927,
    n942,
    n729,
    n688
  );


  and
  g1032
  (
    n986,
    n930,
    n784,
    n682,
    n640
  );


  xnor
  g1033
  (
    n1018,
    n708,
    n926,
    n940,
    n675
  );


  or
  g1034
  (
    n989,
    n665,
    n785,
    n677,
    n730
  );


  and
  g1035
  (
    n967,
    n672,
    n765,
    n699,
    n733
  );


  nor
  g1036
  (
    n1041,
    n776,
    n651,
    n938,
    n723
  );


  or
  g1037
  (
    n980,
    n769,
    n657,
    n935,
    n780
  );


  or
  g1038
  (
    n946,
    n941,
    n937,
    n720,
    n715
  );


  xor
  g1039
  (
    n1047,
    n662,
    n762,
    n937,
    n676
  );


  nor
  g1040
  (
    n1023,
    n787,
    n765,
    n631,
    n763
  );


  xnor
  g1041
  (
    n1075,
    n784,
    n929,
    n771,
    n696
  );


  nor
  g1042
  (
    n1012,
    n732,
    n690,
    n786,
    n725
  );


  xnor
  g1043
  (
    n1071,
    n915,
    n632,
    n737,
    n668
  );


  or
  g1044
  (
    n1050,
    n691,
    n782,
    n919,
    n942
  );


  and
  g1045
  (
    n1066,
    n773,
    n678,
    n748,
    n651
  );


  or
  g1046
  (
    n959,
    n916,
    n642,
    n668,
    n661
  );


  or
  g1047
  (
    n1051,
    n636,
    n742,
    n707,
    n928
  );


  nand
  g1048
  (
    n1103,
    n682,
    n771,
    n661,
    n935
  );


  nand
  g1049
  (
    n1080,
    n737,
    n932,
    n651,
    n777
  );


  xnor
  g1050
  (
    n947,
    n751,
    n723,
    n759,
    n674
  );


  nor
  g1051
  (
    n1007,
    n785,
    n715,
    n696,
    n778
  );


  and
  g1052
  (
    n1033,
    n763,
    n659,
    n667,
    n655
  );


  and
  g1053
  (
    n1070,
    n657,
    n936,
    n698,
    n666
  );


  xnor
  g1054
  (
    n982,
    n931,
    n722,
    n921,
    n658
  );


  xor
  g1055
  (
    n976,
    n637,
    n929,
    n907,
    n768
  );


  nor
  g1056
  (
    n1053,
    n663,
    n644,
    n717,
    n680
  );


  nor
  g1057
  (
    n1092,
    n656,
    n758,
    n688,
    n766
  );


  xor
  g1058
  (
    n1038,
    n718,
    n691,
    n933,
    n788
  );


  nor
  g1059
  (
    n1002,
    n711,
    n934,
    n925,
    n701
  );


  or
  g1060
  (
    n968,
    n938,
    n671,
    n716,
    n694
  );


  or
  g1061
  (
    n996,
    n772,
    n731,
    n717,
    n924
  );


  and
  g1062
  (
    n1083,
    n925,
    n633,
    n920,
    n943
  );


  or
  g1063
  (
    n993,
    n757,
    n753,
    n669,
    n740
  );


  and
  g1064
  (
    n1060,
    n645,
    n789,
    n770,
    n693
  );


  xor
  g1065
  (
    n1039,
    n680,
    n706,
    n704,
    n674
  );


  or
  g1066
  (
    n960,
    n666,
    n919,
    n647,
    n786
  );


  xnor
  g1067
  (
    n997,
    n728,
    n703,
    n739,
    n922
  );


  or
  g1068
  (
    n1010,
    n649,
    n932,
    n741,
    n751
  );


  xnor
  g1069
  (
    n1021,
    n926,
    n670,
    n673,
    n782
  );


  and
  g1070
  (
    n995,
    n698,
    n780,
    n646,
    n719
  );


  xor
  g1071
  (
    n992,
    n750,
    n629,
    n922,
    n769
  );


  or
  g1072
  (
    n1074,
    n918,
    n765,
    n921,
    n736
  );


  nand
  g1073
  (
    n1106,
    n946,
    n791
  );


  or
  g1074
  (
    n1107,
    n1106,
    n792
  );


  not
  g1075
  (
    KeyWire_0_25,
    n1107
  );


  buf
  g1076
  (
    n1109,
    n1108
  );


  xnor
  g1077
  (
    n1113,
    n947,
    n1109,
    n950
  );


  and
  g1078
  (
    n1112,
    n949,
    n948,
    n950
  );


  nor
  g1079
  (
    n1111,
    n946,
    n947,
    n949,
    n1109
  );


  xor
  g1080
  (
    n1110,
    n951,
    n1109,
    n793
  );


  not
  g1081
  (
    n1115,
    n1106
  );


  nor
  g1082
  (
    n1114,
    n1112,
    n951,
    n1113
  );


  or
  g1083
  (
    n1117,
    n794,
    n796,
    n795,
    n1115
  );


  or
  g1084
  (
    n1116,
    n793,
    n795,
    n794
  );


  and
  g1085
  (
    n1118,
    n794,
    n1115,
    n1114,
    n796
  );


  and
  g1086
  (
    n1119,
    n952,
    n1117
  );


  and
  g1087
  (
    n1122,
    n1119,
    n796
  );


  xor
  g1088
  (
    n1120,
    n1118,
    n1119
  );


  and
  g1089
  (
    n1121,
    n1119,
    n1107
  );


  xor
  g1090
  (
    n1123,
    n1122,
    n798,
    n799
  );


  and
  g1091
  (
    n1126,
    n798,
    n1122,
    n800,
    n797
  );


  or
  g1092
  (
    n1125,
    n797,
    n798,
    n1121,
    n800
  );


  xor
  g1093
  (
    n1124,
    n799,
    n1120,
    n797,
    n800
  );


  buf
  g1094
  (
    n1130,
    n515
  );


  xor
  g1095
  (
    n1129,
    n1126,
    n506,
    n510,
    n1108
  );


  nand
  g1096
  (
    n1128,
    n507,
    n1108,
    n1125
  );


  nor
  g1097
  (
    n1140,
    n513,
    n508,
    n509,
    n1125
  );


  and
  g1098
  (
    n1134,
    n1124,
    n1119,
    n1125,
    n509
  );


  xnor
  g1099
  (
    n1127,
    n513,
    n507,
    n1113,
    n510
  );


  nor
  g1100
  (
    n1142,
    n507,
    n515,
    n1123
  );


  and
  g1101
  (
    n1132,
    n1126,
    n512,
    n513,
    n511
  );


  xnor
  g1102
  (
    n1138,
    n512,
    n513,
    n510,
    n511
  );


  nor
  g1103
  (
    n1135,
    n514,
    n511,
    n1126,
    n1123
  );


  xnor
  g1104
  (
    n1131,
    n506,
    n1124,
    n514,
    n511
  );


  and
  g1105
  (
    n1141,
    n505,
    n508,
    n1126,
    n1124
  );


  nand
  g1106
  (
    n1136,
    n512,
    n508,
    n1124,
    n1123
  );


  nand
  g1107
  (
    n1139,
    n506,
    n514,
    n507,
    n509
  );


  xor
  g1108
  (
    n1137,
    n506,
    n509,
    n515
  );


  xnor
  g1109
  (
    n1133,
    n510,
    n508,
    n514,
    n512
  );


  nand
  g1110
  (
    n1150,
    n855,
    n825,
    n837,
    n864
  );


  nor
  g1111
  (
    n1196,
    n812,
    n1132,
    n1133,
    n811
  );


  or
  g1112
  (
    n1191,
    n849,
    n803,
    n855,
    n1138
  );


  xor
  g1113
  (
    n1170,
    n824,
    n806,
    n1132
  );


  or
  g1114
  (
    n1153,
    n814,
    n823,
    n1139,
    n1140
  );


  xor
  g1115
  (
    n1200,
    n1129,
    n844,
    n1140
  );


  xnor
  g1116
  (
    n1201,
    n847,
    n1141,
    n830,
    n854
  );


  nor
  g1117
  (
    n1189,
    n802,
    n831,
    n824,
    n816
  );


  xnor
  g1118
  (
    n1194,
    n850,
    n860,
    n834,
    n839
  );


  and
  g1119
  (
    n1162,
    n858,
    n1137,
    n1133,
    n833
  );


  xnor
  g1120
  (
    n1169,
    n1141,
    n814,
    n838,
    n830
  );


  nand
  g1121
  (
    n1193,
    n844,
    n835,
    n852,
    n1137
  );


  xnor
  g1122
  (
    n1146,
    n856,
    n857,
    n1142,
    n1128
  );


  nor
  g1123
  (
    n1183,
    n856,
    n848,
    n1131,
    n809
  );


  xnor
  g1124
  (
    n1188,
    n857,
    n859,
    n1137,
    n841
  );


  xor
  g1125
  (
    n1178,
    n827,
    n823,
    n826,
    n803
  );


  nand
  g1126
  (
    n1159,
    n815,
    n847,
    n1136,
    n804
  );


  nand
  g1127
  (
    n1202,
    n821,
    n840,
    n839,
    n804
  );


  xor
  g1128
  (
    n1156,
    n838,
    n864,
    n807,
    n812
  );


  or
  g1129
  (
    n1144,
    n853,
    n843,
    n823,
    n1132
  );


  and
  g1130
  (
    n1147,
    n1131,
    n1133,
    n1135,
    n831
  );


  xor
  g1131
  (
    n1177,
    n818,
    n1135,
    n1142,
    n820
  );


  nor
  g1132
  (
    n1149,
    n1141,
    n811,
    n863
  );


  and
  g1133
  (
    n1204,
    n1135,
    n818,
    n832,
    n815
  );


  xor
  g1134
  (
    n1185,
    n808,
    n846,
    n814,
    n1132
  );


  nand
  g1135
  (
    n1143,
    n1134,
    n1130,
    n840,
    n862
  );


  nor
  g1136
  (
    KeyWire_0_58,
    n1136,
    n826,
    n861,
    n810
  );


  and
  g1137
  (
    n1158,
    n830,
    n802,
    n1134,
    n1139
  );


  xor
  g1138
  (
    n1151,
    n816,
    n1138,
    n819,
    n1130
  );


  xnor
  g1139
  (
    n1154,
    n850,
    n861,
    n838,
    n1135
  );


  nor
  g1140
  (
    n1190,
    n1127,
    n842,
    n807,
    n854
  );


  or
  g1141
  (
    n1205,
    n860,
    n837,
    n1129,
    n834
  );


  and
  g1142
  (
    KeyWire_0_32,
    n840,
    n845,
    n821,
    n835
  );


  or
  g1143
  (
    n1199,
    n825,
    n847,
    n801,
    n809
  );


  nand
  g1144
  (
    n1152,
    n842,
    n810,
    n864,
    n843
  );


  or
  g1145
  (
    n1180,
    n1131,
    n854,
    n1134,
    n817
  );


  xor
  g1146
  (
    n1187,
    n837,
    n825,
    n852,
    n805
  );


  or
  g1147
  (
    n1166,
    n829,
    n855,
    n806,
    n836
  );


  xnor
  g1148
  (
    n1167,
    n1128,
    n845,
    n853,
    n1129
  );


  xnor
  g1149
  (
    n1165,
    n842,
    n815,
    n819,
    n1137
  );


  xor
  g1150
  (
    n1175,
    n816,
    n841,
    n813,
    n826
  );


  or
  g1151
  (
    n1171,
    n824,
    n1142,
    n813,
    n843
  );


  or
  g1152
  (
    n1163,
    n805,
    n848,
    n844,
    n1127
  );


  and
  g1153
  (
    n1182,
    n849,
    n848,
    n860,
    n833
  );


  and
  g1154
  (
    n1206,
    n1128,
    n817,
    n850,
    n852
  );


  nand
  g1155
  (
    n1176,
    n853,
    n836,
    n808,
    n1141
  );


  nor
  g1156
  (
    n1186,
    n858,
    n1136,
    n821,
    n832
  );


  and
  g1157
  (
    n1179,
    n1133,
    n1142,
    n805,
    n858
  );


  and
  g1158
  (
    n1181,
    n863,
    n835,
    n828,
    n801
  );


  nand
  g1159
  (
    n1168,
    n859,
    n859,
    n846,
    n856
  );


  xor
  g1160
  (
    n1184,
    n1130,
    n828,
    n846,
    n809
  );


  and
  g1161
  (
    n1192,
    n1138,
    n1136,
    n862,
    n1134
  );


  and
  g1162
  (
    n1164,
    n863,
    n836,
    n834,
    n831
  );


  nand
  g1163
  (
    n1173,
    n822,
    n851,
    n839,
    n817
  );


  xor
  g1164
  (
    n1198,
    n820,
    n813,
    n1140,
    n833
  );


  xnor
  g1165
  (
    n1174,
    n1127,
    n803,
    n857,
    n822
  );


  xor
  g1166
  (
    n1155,
    n1139,
    n832,
    n819,
    n827
  );


  xor
  g1167
  (
    n1195,
    n808,
    n1127,
    n802,
    n851
  );


  nand
  g1168
  (
    KeyWire_0_35,
    n829,
    n1129,
    n827,
    n807
  );


  and
  g1169
  (
    n1161,
    n812,
    n861,
    n1128,
    n818
  );


  nand
  g1170
  (
    n1197,
    n801,
    n810,
    n1130,
    n1139
  );


  xnor
  g1171
  (
    n1145,
    n820,
    n822,
    n841,
    n804
  );


  or
  g1172
  (
    n1203,
    n851,
    n829,
    n1131,
    n862
  );


  nand
  g1173
  (
    n1157,
    n845,
    n1138,
    n828,
    n849
  );


  xnor
  g1174
  (
    n1236,
    n969,
    n1055,
    n1147,
    n1160
  );


  nor
  g1175
  (
    n1244,
    n1004,
    n985,
    n1189,
    n1050
  );


  and
  g1176
  (
    n1274,
    n1064,
    n969,
    n1183,
    n1071
  );


  nand
  g1177
  (
    n1273,
    n1199,
    n1070,
    n961,
    n1021
  );


  xor
  g1178
  (
    n1251,
    n1062,
    n1031,
    n1030,
    n1165
  );


  xnor
  g1179
  (
    n1264,
    n954,
    n1045,
    n1087,
    n1150
  );


  or
  g1180
  (
    n1309,
    n1175,
    n1166,
    n1199,
    n1000
  );


  and
  g1181
  (
    n1283,
    n871,
    n986,
    n1171,
    n1180
  );


  nor
  g1182
  (
    n1362,
    n1163,
    n1193,
    n995,
    n1204
  );


  and
  g1183
  (
    n1379,
    n964,
    n868,
    n1098,
    n1083
  );


  and
  g1184
  (
    n1226,
    n1069,
    n1192,
    n1015,
    n953
  );


  xor
  g1185
  (
    n1367,
    n1034,
    n1053,
    n1004,
    n1153
  );


  nand
  g1186
  (
    n1237,
    n1188,
    n1033,
    n1146,
    n981
  );


  and
  g1187
  (
    n1308,
    n1015,
    n1199,
    n1091,
    n1082
  );


  nand
  g1188
  (
    n1267,
    n1166,
    n1069,
    n1182,
    n867
  );


  xnor
  g1189
  (
    n1363,
    n1152,
    n1061,
    n1101,
    n1028
  );


  xnor
  g1190
  (
    n1254,
    n1148,
    n1077,
    n1094,
    n971
  );


  nor
  g1191
  (
    n1387,
    n967,
    n1159,
    n1089,
    n1072
  );


  xor
  g1192
  (
    n1381,
    n1064,
    n1043,
    n1073,
    n954
  );


  nor
  g1193
  (
    n1221,
    n1179,
    n1151,
    n1168,
    n998
  );


  nor
  g1194
  (
    n1338,
    n1166,
    n1153,
    n1077,
    n959
  );


  or
  g1195
  (
    n1208,
    n1000,
    n1066,
    n969,
    n1161
  );


  nor
  g1196
  (
    n1301,
    n1188,
    n1048,
    n978,
    n1097
  );


  nand
  g1197
  (
    n1317,
    n1175,
    n983,
    n1076,
    n1017
  );


  xnor
  g1198
  (
    n1365,
    n953,
    n1063,
    n1143,
    n1167
  );


  nor
  g1199
  (
    n1255,
    n1025,
    n970,
    n976,
    n1048
  );


  xnor
  g1200
  (
    n1329,
    n967,
    n1049,
    n1149,
    n1150
  );


  nand
  g1201
  (
    n1262,
    n1205,
    n1195,
    n982,
    n1054
  );


  or
  g1202
  (
    n1230,
    n1011,
    n1000,
    n1036,
    n1155
  );


  nor
  g1203
  (
    n1345,
    n1008,
    n1158,
    n1087,
    n961
  );


  xnor
  g1204
  (
    n1238,
    n1101,
    n1026,
    n1200,
    n984
  );


  xnor
  g1205
  (
    n1277,
    n1181,
    n1148,
    n1079,
    n1018
  );


  xnor
  g1206
  (
    n1311,
    n1025,
    n979,
    n1084,
    n988
  );


  nor
  g1207
  (
    n1354,
    n1177,
    n1035,
    n983,
    n1193
  );


  nand
  g1208
  (
    n1239,
    n1001,
    n1177,
    n1046,
    n867
  );


  xnor
  g1209
  (
    n1302,
    n1059,
    n1193,
    n1017,
    n1102
  );


  xnor
  g1210
  (
    n1253,
    n1154,
    n1148,
    n1160,
    n991
  );


  xnor
  g1211
  (
    n1326,
    n1154,
    n1197,
    n981,
    n1006
  );


  xnor
  g1212
  (
    n1209,
    n1194,
    n1074,
    n957,
    n1013
  );


  or
  g1213
  (
    n1335,
    n984,
    n1010,
    n1054,
    n1042
  );


  nor
  g1214
  (
    n1312,
    n1151,
    n1168,
    n1049,
    n1058
  );


  xor
  g1215
  (
    n1268,
    n960,
    n960,
    n865,
    n1052
  );


  nand
  g1216
  (
    n1313,
    n997,
    n1039,
    n870,
    n987
  );


  nor
  g1217
  (
    n1241,
    n1083,
    n1068,
    n988,
    n1074
  );


  xnor
  g1218
  (
    n1324,
    n994,
    n1047,
    n1065,
    n874
  );


  xnor
  g1219
  (
    n1216,
    n875,
    n1075,
    n1071
  );


  xnor
  g1220
  (
    n1242,
    n989,
    n1195,
    n1153,
    n1027
  );


  xnor
  g1221
  (
    n1280,
    n1005,
    n1080,
    n990,
    n997
  );


  nand
  g1222
  (
    n1278,
    n1088,
    n1058,
    n1196,
    n1160
  );


  xor
  g1223
  (
    n1359,
    n1191,
    n1040,
    n968,
    n1156
  );


  or
  g1224
  (
    n1248,
    n1149,
    n1015,
    n869,
    n1093
  );


  nor
  g1225
  (
    n1265,
    n1190,
    n1205,
    n1092,
    n978
  );


  and
  g1226
  (
    n1220,
    n1161,
    n993,
    n976,
    n1024
  );


  xnor
  g1227
  (
    n1364,
    n1075,
    n1147,
    n1143,
    n1192
  );


  xnor
  g1228
  (
    n1249,
    n1144,
    n866,
    n1073,
    n1008
  );


  nand
  g1229
  (
    KeyWire_0_30,
    n1016,
    n1148,
    n1185,
    n956
  );


  or
  g1230
  (
    n1351,
    n967,
    n1033,
    n1145,
    n1088
  );


  nand
  g1231
  (
    n1370,
    n1079,
    n1205,
    n982,
    n1047
  );


  nor
  g1232
  (
    n1256,
    n1003,
    n1185,
    n1011,
    n1191
  );


  xnor
  g1233
  (
    n1234,
    n1092,
    n1165,
    n1052,
    n1187
  );


  xnor
  g1234
  (
    n1247,
    n994,
    n974,
    n983,
    n1053
  );


  or
  g1235
  (
    n1232,
    n1035,
    n1095,
    n1160,
    n1100
  );


  xnor
  g1236
  (
    n1250,
    n1167,
    n974,
    n1188,
    n1001
  );


  nor
  g1237
  (
    n1371,
    n1031,
    n1182,
    n1009,
    n872
  );


  and
  g1238
  (
    n1288,
    n1098,
    n1023,
    n1030,
    n968
  );


  xor
  g1239
  (
    n1295,
    n1019,
    n1178,
    n1086,
    n1057
  );


  xor
  g1240
  (
    n1342,
    n1062,
    n1169,
    n1152,
    n1010
  );


  xor
  g1241
  (
    n1281,
    n1173,
    n1180,
    n1018,
    n1034
  );


  or
  g1242
  (
    n1304,
    n959,
    n1190,
    n963,
    n1184
  );


  xor
  g1243
  (
    n1382,
    n966,
    n998,
    n1167,
    n1170
  );


  and
  g1244
  (
    n1356,
    n1067,
    n1056,
    n1061,
    n957
  );


  or
  g1245
  (
    n1224,
    n1042,
    n1159,
    n1178,
    n1145
  );


  xnor
  g1246
  (
    n1388,
    n1078,
    n1029,
    n1065,
    n1197
  );


  nand
  g1247
  (
    n1337,
    n865,
    n1014,
    n1039
  );


  nor
  g1248
  (
    n1380,
    n1144,
    n1151,
    n984,
    n1145
  );


  and
  g1249
  (
    n1259,
    n1178,
    n1146,
    n1041,
    n1098
  );


  xnor
  g1250
  (
    n1210,
    n1201,
    n1147,
    n1169,
    n973
  );


  nor
  g1251
  (
    n1298,
    n873,
    n982,
    n1019,
    n1087
  );


  and
  g1252
  (
    n1266,
    n1016,
    n960,
    n1178,
    n994
  );


  or
  g1253
  (
    n1322,
    n1203,
    n1004,
    n1201,
    n1094
  );


  or
  g1254
  (
    n1252,
    n1187,
    n1159,
    n1018,
    n1155
  );


  nand
  g1255
  (
    n1214,
    n987,
    n1192,
    n1094,
    n992
  );


  xnor
  g1256
  (
    n1344,
    n1005,
    n1156,
    n1194,
    n1032
  );


  nand
  g1257
  (
    n1228,
    n1202,
    n871,
    n972,
    n999
  );


  xor
  g1258
  (
    n1331,
    n1155,
    n1023,
    n1189,
    n1201
  );


  nor
  g1259
  (
    n1330,
    n979,
    n1183,
    n1200,
    n1068
  );


  nand
  g1260
  (
    n1333,
    n1042,
    n1173,
    n1163,
    n1199
  );


  nand
  g1261
  (
    n1297,
    n1081,
    n1077,
    n1183,
    n1176
  );


  nand
  g1262
  (
    n1307,
    n1013,
    n1205,
    n1063,
    n996
  );


  or
  g1263
  (
    n1357,
    n1057,
    n1037,
    n1168,
    n958
  );


  nand
  g1264
  (
    n1325,
    n1186,
    n976,
    n995,
    n1006
  );


  xnor
  g1265
  (
    n1217,
    n970,
    n1184,
    n1177,
    n989
  );


  xor
  g1266
  (
    n1219,
    n1096,
    n1196,
    n1060,
    n1201
  );


  xor
  g1267
  (
    n1374,
    n1096,
    n1041,
    n977,
    n1091
  );


  or
  g1268
  (
    n1316,
    n1055,
    n1013,
    n1149,
    n1179
  );


  nand
  g1269
  (
    n1211,
    n1058,
    n1051,
    n1151,
    n1153
  );


  and
  g1270
  (
    n1373,
    n1086,
    n1069,
    n1066,
    n1193
  );


  xnor
  g1271
  (
    n1284,
    n1173,
    n1070,
    n987,
    n867
  );


  xor
  g1272
  (
    n1353,
    n1052,
    n1027,
    n1084,
    n977
  );


  xnor
  g1273
  (
    n1212,
    n1012,
    n1182,
    n1186,
    n1022
  );


  xor
  g1274
  (
    n1350,
    n1001,
    n1158,
    n997,
    n1177
  );


  nor
  g1275
  (
    n1332,
    n1046,
    n1157,
    n874,
    n1043
  );


  xnor
  g1276
  (
    n1290,
    n1165,
    n1186,
    n1204,
    n1061
  );


  xor
  g1277
  (
    n1240,
    n1017,
    n1002,
    n1196,
    n991
  );


  and
  g1278
  (
    n1361,
    n1090,
    n1051,
    n1063,
    n1174
  );


  or
  g1279
  (
    n1246,
    n1176,
    n1012,
    n1072,
    n1173
  );


  nand
  g1280
  (
    n1279,
    n1174,
    n1172,
    n1047,
    n1196
  );


  and
  g1281
  (
    n1276,
    n1179,
    n1200,
    n1020,
    n1038
  );


  or
  g1282
  (
    n1375,
    n1029,
    n1143,
    n1010,
    n1188
  );


  nor
  g1283
  (
    n1328,
    n1089,
    n1166,
    n871,
    n1078
  );


  nand
  g1284
  (
    n1355,
    n874,
    n1095,
    n1030,
    n1198
  );


  nand
  g1285
  (
    n1319,
    n1171,
    n875,
    n1203,
    n986
  );


  nor
  g1286
  (
    n1271,
    n1012,
    n973,
    n952,
    n1190
  );


  nor
  g1287
  (
    n1368,
    n1180,
    n962,
    n1068,
    n1161
  );


  xnor
  g1288
  (
    n1272,
    n1150,
    n1172,
    n1195,
    n1040
  );


  nor
  g1289
  (
    n1323,
    n989,
    n1051,
    n990,
    n1059
  );


  nand
  g1290
  (
    n1334,
    n1045,
    n1048,
    n1099,
    n1176
  );


  and
  g1291
  (
    n1285,
    n868,
    n1156,
    n1055,
    n1198
  );


  nor
  g1292
  (
    n1270,
    n986,
    n1163,
    n1146,
    n1158
  );


  or
  g1293
  (
    n1263,
    n963,
    n1060,
    n993
  );


  xor
  g1294
  (
    n1383,
    n1174,
    n866,
    n869,
    n1006
  );


  nand
  g1295
  (
    n1215,
    n961,
    n999,
    n985,
    n1065
  );


  nand
  g1296
  (
    n1366,
    n1081,
    n1189,
    n1032,
    n1074
  );


  and
  g1297
  (
    n1343,
    n1200,
    n972,
    n1197,
    n1049
  );


  xor
  g1298
  (
    n1321,
    n1147,
    n991,
    n964,
    n988
  );


  nor
  g1299
  (
    n1245,
    n962,
    n1076,
    n975,
    n966
  );


  nand
  g1300
  (
    n1289,
    n1025,
    n975,
    n965,
    n872
  );


  nor
  g1301
  (
    n1243,
    n1059,
    n1162,
    n1076,
    n965
  );


  xor
  g1302
  (
    KeyWire_0_12,
    n1169,
    n963,
    n980,
    n873
  );


  or
  g1303
  (
    n1231,
    n1089,
    n1162,
    n1100,
    n1066
  );


  nor
  g1304
  (
    n1358,
    n1097,
    n1204,
    n1062,
    n956
  );


  and
  g1305
  (
    n1218,
    n1060,
    n968,
    n977,
    n873
  );


  xnor
  g1306
  (
    n1261,
    n1203,
    n1090,
    n980,
    n1171
  );


  xor
  g1307
  (
    n1376,
    n1185,
    n975,
    n1167,
    n1146
  );


  xor
  g1308
  (
    n1336,
    n1164,
    n964,
    n1180,
    n1041
  );


  and
  g1309
  (
    n1360,
    n1157,
    n1007,
    n1172
  );


  or
  g1310
  (
    n1369,
    n1070,
    n1073,
    n1152,
    n1080
  );


  nor
  g1311
  (
    n1340,
    n1202,
    n999,
    n973,
    n866
  );


  nand
  g1312
  (
    n1385,
    n980,
    n1194,
    n1037,
    n1174
  );


  nor
  g1313
  (
    n1327,
    n992,
    n1085,
    n970,
    n1184
  );


  or
  g1314
  (
    n1282,
    n996,
    n1057,
    n1191,
    n1158
  );


  xor
  g1315
  (
    n1314,
    n1083,
    n1082,
    n996,
    n1186
  );


  and
  g1316
  (
    n1320,
    n1157,
    n870,
    n1091,
    n1092
  );


  nand
  g1317
  (
    n1299,
    n1169,
    n1171,
    n1035,
    n1026
  );


  xnor
  g1318
  (
    n1258,
    n1172,
    n1085,
    n1170,
    n1159
  );


  nand
  g1319
  (
    n1235,
    n1002,
    n1072,
    n1198,
    n1078
  );


  xnor
  g1320
  (
    n1303,
    n1192,
    n965,
    n1093,
    n1022
  );


  xnor
  g1321
  (
    n1300,
    n1050,
    n1040,
    n1183,
    n1194
  );


  nand
  g1322
  (
    n1257,
    n1190,
    n1014,
    n1085,
    n865
  );


  or
  g1323
  (
    n1222,
    n1154,
    n1007,
    n979,
    n870
  );


  nor
  g1324
  (
    n1386,
    n1028,
    n868,
    n1075,
    n955
  );


  nor
  g1325
  (
    n1318,
    n1143,
    n1189,
    n1090,
    n1144
  );


  and
  g1326
  (
    n1341,
    n1181,
    n971,
    n1162,
    n1021
  );


  nor
  g1327
  (
    n1310,
    n972,
    n1176,
    n1187,
    n1165
  );


  or
  g1328
  (
    n1225,
    n1197,
    n1029,
    n1203,
    n1099
  );


  xnor
  g1329
  (
    n1229,
    n1088,
    n1187,
    n1016,
    n1157
  );


  xnor
  g1330
  (
    n1349,
    n1023,
    n1164,
    n1038,
    n1020
  );


  xnor
  g1331
  (
    n1296,
    n1045,
    n1162,
    n1080,
    n1009
  );


  xnor
  g1332
  (
    n1223,
    n1033,
    n1026,
    n1079,
    n1182
  );


  nor
  g1333
  (
    n1305,
    n1164,
    n955,
    n869,
    n1054
  );


  xor
  g1334
  (
    n1260,
    n1096,
    n1050,
    n958,
    n1179
  );


  nand
  g1335
  (
    n1233,
    n1003,
    n1145,
    n1044,
    n1093
  );


  nor
  g1336
  (
    n1315,
    n966,
    n1043,
    n1027,
    n1144
  );


  and
  g1337
  (
    n1352,
    n998,
    n1020,
    n1086,
    n1164
  );


  xnor
  g1338
  (
    n1306,
    n974,
    n981,
    n1170,
    n1097
  );


  nand
  g1339
  (
    n1372,
    n1195,
    n978,
    n1155,
    n1181
  );


  xor
  g1340
  (
    n1378,
    n1021,
    n1154,
    n1082,
    n1067
  );


  xor
  g1341
  (
    n1339,
    n1036,
    n1031,
    n1101,
    n1161
  );


  nand
  g1342
  (
    n1275,
    n1056,
    n1037,
    n1168,
    n1084
  );


  nor
  g1343
  (
    n1287,
    n1008,
    n1022,
    n995,
    n1202
  );


  or
  g1344
  (
    n1293,
    n1175,
    n992,
    n1044,
    n1202
  );


  and
  g1345
  (
    n1213,
    n1185,
    n1170,
    n1064,
    n1024
  );


  and
  g1346
  (
    n1207,
    n1102,
    n1011,
    n1034,
    n1175
  );


  or
  g1347
  (
    n1227,
    n872,
    n1181,
    n971,
    n1163
  );


  xor
  g1348
  (
    n1294,
    n1002,
    n1081,
    n1152,
    n1095
  );


  nand
  g1349
  (
    n1292,
    n1184,
    n1019,
    n1150,
    n1005
  );


  nor
  g1350
  (
    n1347,
    n1009,
    n1191,
    n1032,
    n1156
  );


  nand
  g1351
  (
    n1291,
    n985,
    n1053,
    n1028,
    n1039
  );


  nor
  g1352
  (
    n1377,
    n1003,
    n1024,
    n1036,
    n1099
  );


  and
  g1353
  (
    n1384,
    n962,
    n1149,
    n1056,
    n1100
  );


  or
  g1354
  (
    n1346,
    n1204,
    n990,
    n1067,
    n1046
  );


  or
  g1355
  (
    n1348,
    n1198,
    n1044,
    n959,
    n1038
  );


  xnor
  g1356
  (
    n1551,
    n1210,
    n1352
  );


  and
  g1357
  (
    n1564,
    n1248,
    n1377
  );


  or
  g1358
  (
    n1473,
    n1262,
    n1252
  );


  and
  g1359
  (
    n1418,
    n1359,
    n1349
  );


  xnor
  g1360
  (
    n1395,
    n1301,
    n1253
  );


  and
  g1361
  (
    n1431,
    n1311,
    n1345
  );


  or
  g1362
  (
    n1584,
    n1228,
    n1300
  );


  xnor
  g1363
  (
    n1446,
    n1351,
    n1344
  );


  and
  g1364
  (
    n1548,
    n1256,
    n1354
  );


  xor
  g1365
  (
    n1403,
    n1307,
    n1383
  );


  or
  g1366
  (
    n1572,
    n1309,
    n1267
  );


  xor
  g1367
  (
    n1396,
    n1213,
    n1269
  );


  buf
  g1368
  (
    n1509,
    n1316
  );


  and
  g1369
  (
    n1390,
    n1248,
    n1227
  );


  xor
  g1370
  (
    n1500,
    n1261,
    n1319
  );


  xor
  g1371
  (
    n1480,
    n1237,
    n1306
  );


  xor
  g1372
  (
    n1592,
    n1264,
    n1233
  );


  xnor
  g1373
  (
    n1413,
    n1320,
    n1370
  );


  xnor
  g1374
  (
    n1408,
    n1369,
    n1349
  );


  nor
  g1375
  (
    n1513,
    n1247,
    n1303
  );


  xnor
  g1376
  (
    n1556,
    n1337,
    n1306
  );


  or
  g1377
  (
    n1432,
    n1238,
    n1218
  );


  xnor
  g1378
  (
    n1554,
    n1232,
    n1225
  );


  and
  g1379
  (
    n1412,
    n1278,
    n1263
  );


  or
  g1380
  (
    n1428,
    n1351,
    n1319
  );


  nand
  g1381
  (
    n1524,
    n1364,
    n1305
  );


  nand
  g1382
  (
    n1532,
    n1210,
    n1356
  );


  nand
  g1383
  (
    n1541,
    n1263,
    n1325
  );


  xnor
  g1384
  (
    n1424,
    n1277,
    n1343
  );


  xor
  g1385
  (
    KeyWire_0_63,
    n1221,
    n1372
  );


  nand
  g1386
  (
    n1489,
    n1276,
    n1343
  );


  xnor
  g1387
  (
    n1461,
    n1245,
    n1361
  );


  and
  g1388
  (
    n1518,
    n1358,
    n1331
  );


  or
  g1389
  (
    n1444,
    n1302,
    n1325
  );


  and
  g1390
  (
    n1561,
    n1209,
    n1327
  );


  or
  g1391
  (
    n1543,
    n1314,
    n1384
  );


  nand
  g1392
  (
    n1423,
    n1363,
    n1319
  );


  and
  g1393
  (
    n1420,
    n1378,
    n1277
  );


  xnor
  g1394
  (
    n1470,
    n1279,
    n1265
  );


  nor
  g1395
  (
    n1539,
    n1370,
    n1308
  );


  or
  g1396
  (
    n1492,
    n1333,
    n1307
  );


  xnor
  g1397
  (
    n1563,
    n1226,
    n1332
  );


  xnor
  g1398
  (
    n1544,
    n1223,
    n1333
  );


  or
  g1399
  (
    n1531,
    n1308,
    n1381
  );


  nor
  g1400
  (
    n1409,
    n1368,
    n1295
  );


  and
  g1401
  (
    n1579,
    n1214,
    n1263
  );


  nand
  g1402
  (
    n1406,
    n1228,
    n1282
  );


  and
  g1403
  (
    n1468,
    n1318,
    n1310
  );


  nand
  g1404
  (
    n1436,
    n1328,
    n1366
  );


  xnor
  g1405
  (
    n1471,
    n1317,
    n1383
  );


  and
  g1406
  (
    n1568,
    n1261,
    n1324
  );


  or
  g1407
  (
    n1586,
    n1322,
    n1239
  );


  nor
  g1408
  (
    n1570,
    n1297,
    n1362
  );


  and
  g1409
  (
    n1493,
    n1274,
    n1296
  );


  nand
  g1410
  (
    n1549,
    n1224,
    n1376
  );


  or
  g1411
  (
    n1407,
    n1231,
    n1338
  );


  nor
  g1412
  (
    n1434,
    n1256,
    n1311
  );


  nor
  g1413
  (
    n1402,
    n1374,
    n1266
  );


  xor
  g1414
  (
    n1397,
    n1245,
    n1340
  );


  nor
  g1415
  (
    n1478,
    n1338,
    n1219
  );


  xnor
  g1416
  (
    n1587,
    n1259,
    n1342
  );


  xnor
  g1417
  (
    n1523,
    n1287,
    n1227
  );


  xnor
  g1418
  (
    n1498,
    n1236,
    n1235
  );


  nand
  g1419
  (
    n1491,
    n1298,
    n1379
  );


  and
  g1420
  (
    n1445,
    n1226,
    n1262
  );


  nor
  g1421
  (
    n1569,
    n1251,
    n1277
  );


  xnor
  g1422
  (
    n1525,
    n1220,
    n1212
  );


  and
  g1423
  (
    n1439,
    n1340,
    n1245
  );


  nor
  g1424
  (
    n1466,
    n1341,
    n1334
  );


  and
  g1425
  (
    n1419,
    n1355,
    n1335
  );


  nor
  g1426
  (
    n1537,
    n1331,
    n1298
  );


  nor
  g1427
  (
    n1414,
    n1254,
    n1348
  );


  xor
  g1428
  (
    n1562,
    n1355,
    n1283
  );


  and
  g1429
  (
    n1574,
    n1314,
    n1256
  );


  and
  g1430
  (
    n1499,
    n1338,
    n1288
  );


  xor
  g1431
  (
    n1503,
    n1240,
    n1288
  );


  and
  g1432
  (
    n1451,
    n1346,
    n1233
  );


  xor
  g1433
  (
    n1526,
    n1216,
    n1345
  );


  xor
  g1434
  (
    n1501,
    n1242,
    n1358
  );


  and
  g1435
  (
    n1510,
    n1274,
    n1213
  );


  or
  g1436
  (
    n1512,
    n1211,
    n1288
  );


  xor
  g1437
  (
    n1448,
    n1242,
    n1329
  );


  nor
  g1438
  (
    n1467,
    n1241,
    n875
  );


  nand
  g1439
  (
    n1552,
    n1250,
    n1345
  );


  nand
  g1440
  (
    n1555,
    n1291,
    n1209
  );


  xor
  g1441
  (
    n1497,
    n1328,
    n1237
  );


  nand
  g1442
  (
    n1429,
    n1372,
    n1250
  );


  and
  g1443
  (
    n1494,
    n1291,
    n1292
  );


  nor
  g1444
  (
    n1573,
    n1384,
    n1218
  );


  xor
  g1445
  (
    n1426,
    n1220,
    n1279
  );


  nor
  g1446
  (
    n1496,
    n1381,
    n1223
  );


  and
  g1447
  (
    n1462,
    n1287,
    n1230
  );


  nor
  g1448
  (
    n1450,
    n1320,
    n1315
  );


  and
  g1449
  (
    n1575,
    n1216,
    n1267
  );


  and
  g1450
  (
    n1583,
    n1268,
    n1325
  );


  xnor
  g1451
  (
    n1458,
    n1330,
    n1234
  );


  and
  g1452
  (
    n1447,
    n1303,
    n1209
  );


  nor
  g1453
  (
    n1394,
    n1318,
    n1380
  );


  xor
  g1454
  (
    n1504,
    n1323,
    n1359
  );


  and
  g1455
  (
    n1442,
    n1230,
    n1262
  );


  xnor
  g1456
  (
    n1505,
    n1255,
    n1292
  );


  xnor
  g1457
  (
    n1533,
    n1240,
    n1312
  );


  nor
  g1458
  (
    n1438,
    n1258,
    n1283
  );


  and
  g1459
  (
    n1502,
    n1313,
    n1385
  );


  xor
  g1460
  (
    n1529,
    n1295,
    n1348
  );


  xnor
  g1461
  (
    n1515,
    n1364,
    n1280
  );


  xnor
  g1462
  (
    KeyWire_0_56,
    n1246,
    n1276
  );


  or
  g1463
  (
    n1460,
    n1221,
    n1321
  );


  nor
  g1464
  (
    n1511,
    n1265,
    n1290
  );


  nand
  g1465
  (
    n1536,
    n1235,
    n1329
  );


  nor
  g1466
  (
    n1484,
    n1323,
    n1367
  );


  and
  g1467
  (
    n1535,
    n1332,
    n1215
  );


  xor
  g1468
  (
    n1588,
    n1374,
    n1289
  );


  nor
  g1469
  (
    n1516,
    n1281,
    n1208
  );


  xnor
  g1470
  (
    n1559,
    n1247,
    n1270
  );


  or
  g1471
  (
    n1472,
    n1237,
    n1357
  );


  xnor
  g1472
  (
    n1459,
    n1255,
    n1265
  );


  nand
  g1473
  (
    n1411,
    n1295,
    n1217
  );


  or
  g1474
  (
    n1417,
    n1260,
    n1273
  );


  nand
  g1475
  (
    n1558,
    n1363,
    n1274
  );


  nand
  g1476
  (
    n1456,
    n1271,
    n1337
  );


  nor
  g1477
  (
    n1486,
    n1347,
    n1335
  );


  xor
  g1478
  (
    n1469,
    n1230,
    n1368
  );


  or
  g1479
  (
    n1405,
    n1292,
    n1331
  );


  or
  g1480
  (
    n1578,
    n1342,
    n1364
  );


  xor
  g1481
  (
    n1538,
    n1361,
    n1308
  );


  nor
  g1482
  (
    n1565,
    n1225,
    n1332
  );


  xnor
  g1483
  (
    n1528,
    n1297,
    n1366
  );


  and
  g1484
  (
    n1577,
    n1315,
    n1369
  );


  xnor
  g1485
  (
    n1443,
    n1322,
    n1249
  );


  nand
  g1486
  (
    n1589,
    n1271,
    n1207
  );


  xnor
  g1487
  (
    n1590,
    n1271,
    n1232
  );


  nor
  g1488
  (
    n1391,
    n1321,
    n1375
  );


  nor
  g1489
  (
    n1463,
    n1294,
    n1383
  );


  and
  g1490
  (
    n1410,
    n1229,
    n1299
  );


  nand
  g1491
  (
    n1440,
    n1270,
    n1259
  );


  nand
  g1492
  (
    n1520,
    n1290,
    n1309
  );


  and
  g1493
  (
    n1441,
    n1297,
    n1282
  );


  and
  g1494
  (
    n1557,
    n1323,
    n1339
  );


  nor
  g1495
  (
    n1454,
    n1215,
    n1348
  );


  and
  g1496
  (
    n1540,
    n1375,
    n1335,
    n1276,
    n1346
  );


  and
  g1497
  (
    n1465,
    n1311,
    n1212,
    n1275,
    n1296
  );


  nand
  g1498
  (
    n1479,
    n1300,
    n1309,
    n1318,
    n1235
  );


  nor
  g1499
  (
    n1449,
    n1217,
    n1315,
    n1324,
    n1243
  );


  xnor
  g1500
  (
    n1453,
    n1304,
    n1246,
    n1272,
    n1273
  );


  xor
  g1501
  (
    n1416,
    n1347,
    n1264,
    n1223,
    n1286
  );


  and
  g1502
  (
    n1425,
    n1341,
    n1234,
    n1349,
    n1252
  );


  nor
  g1503
  (
    n1401,
    n1302,
    n1222,
    n1229,
    n1371
  );


  nand
  g1504
  (
    n1427,
    n1289,
    n1268,
    n1270,
    n1334
  );


  and
  g1505
  (
    n1522,
    n1293,
    n1280,
    n1307,
    n1336
  );


  xor
  g1506
  (
    n1514,
    n1299,
    n1242,
    n1296,
    n1275
  );


  xor
  g1507
  (
    n1430,
    n1236,
    n1215,
    n1221,
    n1279
  );


  and
  g1508
  (
    n1415,
    n1358,
    n1353,
    n1232,
    n1228
  );


  nor
  g1509
  (
    n1389,
    n1246,
    n1312,
    n1233,
    n1310
  );


  and
  g1510
  (
    n1530,
    n1268,
    n1222,
    n1251,
    n1304
  );


  nand
  g1511
  (
    n1392,
    n1216,
    n1214,
    n1253,
    n1378
  );


  xnor
  g1512
  (
    n1567,
    n1231,
    n1381,
    n1224,
    n1244
  );


  nand
  g1513
  (
    n1400,
    n1301,
    n1384,
    n1272,
    n1356
  );


  and
  g1514
  (
    n1580,
    n1260,
    n1342,
    n1267,
    n1339
  );


  and
  g1515
  (
    KeyWire_0_27,
    n1346,
    n1257,
    n1376,
    n1343
  );


  nand
  g1516
  (
    n1545,
    n1214,
    n1236,
    n1347,
    n1374
  );


  xor
  g1517
  (
    n1482,
    n1258,
    n1378,
    n1252,
    n1293
  );


  xor
  g1518
  (
    n1546,
    n1333,
    n1282,
    n1357,
    n1285
  );


  and
  g1519
  (
    n1527,
    n1366,
    n1211,
    n1244,
    n1299
  );


  and
  g1520
  (
    n1553,
    n1377,
    n1361,
    n1284,
    n1324
  );


  and
  g1521
  (
    n1517,
    n1330,
    n1379,
    n1363,
    n1370
  );


  nor
  g1522
  (
    n1435,
    n1367,
    n1326,
    n1291,
    n1225
  );


  and
  g1523
  (
    n1542,
    n1257,
    n1334,
    n1326,
    n1344
  );


  xor
  g1524
  (
    n1519,
    n1377,
    n1368,
    n1219,
    n1313
  );


  xnor
  g1525
  (
    n1534,
    n1239,
    n1353,
    n1362,
    n1360
  );


  xnor
  g1526
  (
    n1455,
    n1251,
    n1365,
    n1327,
    n1322
  );


  nand
  g1527
  (
    n1477,
    n1301,
    n1317,
    n1211,
    n1320
  );


  xnor
  g1528
  (
    n1488,
    n1310,
    n1354,
    n1213,
    n1219
  );


  nand
  g1529
  (
    KeyWire_0_41,
    n1269,
    n1238,
    n1257,
    n1357
  );


  and
  g1530
  (
    n1521,
    n1208,
    n1359,
    n1249,
    n1373
  );


  xor
  g1531
  (
    n1437,
    n1360,
    n1241,
    n1336,
    n1275
  );


  xor
  g1532
  (
    n1481,
    n1327,
    n1224,
    n1293,
    n1336
  );


  xnor
  g1533
  (
    n1495,
    n1321,
    n1373,
    n1239,
    n1306
  );


  xor
  g1534
  (
    n1422,
    n1304,
    n1207,
    n1286,
    n1376
  );


  xor
  g1535
  (
    n1474,
    n1328,
    n1272,
    n1373,
    n1284
  );


  or
  g1536
  (
    n1571,
    n1380,
    n1305,
    n1302,
    n1371
  );


  xnor
  g1537
  (
    n1398,
    n1326,
    n1379,
    n1218,
    n1365
  );


  xnor
  g1538
  (
    n1475,
    n1266,
    n1356,
    n1300,
    n1289
  );


  xor
  g1539
  (
    n1591,
    n1340,
    n1240,
    n1290,
    n1316
  );


  and
  g1540
  (
    n1457,
    n1250,
    n1294,
    n1330,
    n1238
  );


  xnor
  g1541
  (
    n1566,
    n1360,
    n1369,
    n1350
  );


  nor
  g1542
  (
    n1485,
    n1258,
    n1249,
    n1222,
    n1229
  );


  or
  g1543
  (
    n1508,
    n1350,
    n1283,
    n1337,
    n1367
  );


  or
  g1544
  (
    n1404,
    n1254,
    n1382,
    n1220,
    n1227
  );


  xnor
  g1545
  (
    n1506,
    n1207,
    n1352,
    n1382,
    n1353
  );


  xor
  g1546
  (
    n1581,
    n1244,
    n1303,
    n1281,
    n1210
  );


  xor
  g1547
  (
    n1550,
    n1255,
    n1372,
    n1273,
    n1280
  );


  and
  g1548
  (
    n1399,
    n1281,
    n1351,
    n1329,
    n1344
  );


  and
  g1549
  (
    n1487,
    n1362,
    n1243,
    n1269,
    n1248
  );


  xnor
  g1550
  (
    n1507,
    n1339,
    n1285,
    n1294,
    n1243
  );


  nand
  g1551
  (
    n1490,
    n1354,
    n1266,
    n1226,
    n1355
  );


  and
  g1552
  (
    n1393,
    n1312,
    n1264,
    n1285,
    n1212
  );


  nor
  g1553
  (
    n1421,
    n1305,
    n1254,
    n1341,
    n1371
  );


  xor
  g1554
  (
    n1560,
    n1298,
    n1287,
    n1261,
    n1286
  );


  and
  g1555
  (
    n1582,
    n1317,
    n1278,
    n1260,
    n1382
  );


  and
  g1556
  (
    n1547,
    n1375,
    n1352,
    n1314,
    n1278
  );


  xnor
  g1557
  (
    n1483,
    n1259,
    n1217,
    n1313,
    n1208
  );


  nand
  g1558
  (
    n1452,
    n1231,
    n1234,
    n1241,
    n1365
  );


  or
  g1559
  (
    n1576,
    n1284,
    n1253,
    n1380,
    n1247
  );


  buf
  g1560
  (
    n1672,
    n1417
  );


  not
  g1561
  (
    n1708,
    n1422
  );


  not
  g1562
  (
    n1654,
    n1530
  );


  buf
  g1563
  (
    n1635,
    n1501
  );


  buf
  g1564
  (
    n1602,
    n1534
  );


  buf
  g1565
  (
    n1760,
    n1520
  );


  not
  g1566
  (
    n1818,
    n1445
  );


  buf
  g1567
  (
    n1814,
    n1514
  );


  buf
  g1568
  (
    n1712,
    n1540
  );


  buf
  g1569
  (
    n1711,
    n1464
  );


  buf
  g1570
  (
    n1605,
    n1562
  );


  not
  g1571
  (
    n1692,
    n1557
  );


  not
  g1572
  (
    n1757,
    n1541
  );


  not
  g1573
  (
    n1730,
    n1539
  );


  buf
  g1574
  (
    n1851,
    n1482
  );


  not
  g1575
  (
    n1669,
    n1466
  );


  not
  g1576
  (
    n1797,
    n1437
  );


  not
  g1577
  (
    n1778,
    n1503
  );


  not
  g1578
  (
    n1811,
    n1560
  );


  buf
  g1579
  (
    n1865,
    n1496
  );


  not
  g1580
  (
    n1850,
    n1540
  );


  buf
  g1581
  (
    n1603,
    n1419
  );


  not
  g1582
  (
    n1673,
    n1511
  );


  not
  g1583
  (
    n1598,
    n1427
  );


  not
  g1584
  (
    n1835,
    n1544
  );


  not
  g1585
  (
    n1699,
    n1415
  );


  buf
  g1586
  (
    n1724,
    n1429
  );


  buf
  g1587
  (
    n1836,
    n1497
  );


  buf
  g1588
  (
    n1819,
    n1553
  );


  buf
  g1589
  (
    n1722,
    n1500
  );


  not
  g1590
  (
    n1793,
    n1538
  );


  not
  g1591
  (
    n1655,
    n1520
  );


  not
  g1592
  (
    n1599,
    n1456
  );


  not
  g1593
  (
    n1728,
    n1474
  );


  not
  g1594
  (
    KeyWire_0_60,
    n1451
  );


  not
  g1595
  (
    n1769,
    n1426
  );


  buf
  g1596
  (
    n1600,
    n1490
  );


  buf
  g1597
  (
    n1718,
    n1400
  );


  not
  g1598
  (
    n1852,
    n1481
  );


  buf
  g1599
  (
    n1624,
    n1521
  );


  not
  g1600
  (
    n1806,
    n1507
  );


  not
  g1601
  (
    n1751,
    n1512
  );


  buf
  g1602
  (
    n1855,
    n1405
  );


  not
  g1603
  (
    n1798,
    n1425
  );


  buf
  g1604
  (
    n1616,
    n1444
  );


  buf
  g1605
  (
    n1857,
    n1505
  );


  not
  g1606
  (
    n1691,
    n1492
  );


  not
  g1607
  (
    n1842,
    n1552
  );


  buf
  g1608
  (
    n1813,
    n1533
  );


  not
  g1609
  (
    n1681,
    n1390
  );


  not
  g1610
  (
    n1833,
    n1551
  );


  buf
  g1611
  (
    n1713,
    n1510
  );


  buf
  g1612
  (
    n1860,
    n1467
  );


  not
  g1613
  (
    n1671,
    n1476
  );


  buf
  g1614
  (
    n1695,
    n1482
  );


  not
  g1615
  (
    n1731,
    n1465
  );


  not
  g1616
  (
    n1633,
    n1499
  );


  buf
  g1617
  (
    n1593,
    n1403
  );


  not
  g1618
  (
    n1758,
    n1517
  );


  buf
  g1619
  (
    n1763,
    n1446
  );


  buf
  g1620
  (
    n1774,
    n1396
  );


  not
  g1621
  (
    n1643,
    n1504
  );


  buf
  g1622
  (
    n1705,
    n1557
  );


  buf
  g1623
  (
    n1780,
    n1447
  );


  not
  g1624
  (
    n1662,
    n1415
  );


  buf
  g1625
  (
    n1843,
    n1433
  );


  not
  g1626
  (
    n1619,
    n1415
  );


  buf
  g1627
  (
    n1742,
    n1497
  );


  not
  g1628
  (
    n1826,
    n1404
  );


  not
  g1629
  (
    n1832,
    n1538
  );


  buf
  g1630
  (
    n1646,
    n1409
  );


  not
  g1631
  (
    n1638,
    n1523
  );


  not
  g1632
  (
    n1682,
    n1414
  );


  not
  g1633
  (
    n1644,
    n1494
  );


  not
  g1634
  (
    n1754,
    n1562
  );


  not
  g1635
  (
    n1773,
    n1542
  );


  buf
  g1636
  (
    n1837,
    n1500
  );


  not
  g1637
  (
    n1667,
    n1503
  );


  buf
  g1638
  (
    n1740,
    n1494
  );


  not
  g1639
  (
    n1815,
    n1520
  );


  buf
  g1640
  (
    n1665,
    n1515
  );


  not
  g1641
  (
    n1726,
    n1397
  );


  buf
  g1642
  (
    KeyWire_0_24,
    n1449
  );


  buf
  g1643
  (
    n1612,
    n1550
  );


  not
  g1644
  (
    n1765,
    n1438
  );


  buf
  g1645
  (
    n1653,
    n1473
  );


  buf
  g1646
  (
    n1663,
    n1509
  );


  buf
  g1647
  (
    KeyWire_0_1,
    n1490
  );


  not
  g1648
  (
    n1841,
    n1558
  );


  not
  g1649
  (
    n1861,
    n1464
  );


  not
  g1650
  (
    n1752,
    n1470
  );


  not
  g1651
  (
    n1767,
    n1476
  );


  buf
  g1652
  (
    n1783,
    n1523
  );


  not
  g1653
  (
    n1791,
    n1564
  );


  buf
  g1654
  (
    n1846,
    n1528
  );


  not
  g1655
  (
    n1739,
    n1453
  );


  buf
  g1656
  (
    n1684,
    n1416
  );


  not
  g1657
  (
    n1777,
    n1399
  );


  not
  g1658
  (
    n1776,
    n1493
  );


  not
  g1659
  (
    n1805,
    n1406
  );


  buf
  g1660
  (
    n1615,
    n1511
  );


  buf
  g1661
  (
    n1628,
    n1561
  );


  not
  g1662
  (
    n1702,
    n1430
  );


  buf
  g1663
  (
    n1735,
    n1462
  );


  not
  g1664
  (
    n1610,
    n1418
  );


  not
  g1665
  (
    n1634,
    n1565
  );


  not
  g1666
  (
    n1723,
    n1421
  );


  buf
  g1667
  (
    KeyWire_0_21,
    n1434
  );


  not
  g1668
  (
    n1747,
    n1428
  );


  buf
  g1669
  (
    n1642,
    n1516
  );


  not
  g1670
  (
    n1594,
    n1462
  );


  buf
  g1671
  (
    KeyWire_0_49,
    n1478
  );


  not
  g1672
  (
    n1622,
    n1539
  );


  buf
  g1673
  (
    n1750,
    n1533
  );


  buf
  g1674
  (
    n1649,
    n1543
  );


  not
  g1675
  (
    KeyWire_0_33,
    n1529
  );


  not
  g1676
  (
    n1845,
    n1442
  );


  not
  g1677
  (
    n1800,
    n1423
  );


  not
  g1678
  (
    n1741,
    n1502
  );


  not
  g1679
  (
    n1786,
    n1423
  );


  buf
  g1680
  (
    n1827,
    n1514
  );


  not
  g1681
  (
    n1686,
    n1446
  );


  not
  g1682
  (
    n1666,
    n1421
  );


  buf
  g1683
  (
    n1631,
    n1532
  );


  buf
  g1684
  (
    n1690,
    n1556
  );


  not
  g1685
  (
    n1796,
    n1531
  );


  not
  g1686
  (
    n1650,
    n1389
  );


  not
  g1687
  (
    n1744,
    n1443
  );


  not
  g1688
  (
    n1736,
    n1501
  );


  not
  g1689
  (
    n1737,
    n1489
  );


  not
  g1690
  (
    n1687,
    n1531
  );


  not
  g1691
  (
    n1660,
    n1470
  );


  not
  g1692
  (
    n1674,
    n1509
  );


  not
  g1693
  (
    n1721,
    n1552
  );


  not
  g1694
  (
    n1853,
    n1488
  );


  buf
  g1695
  (
    n1727,
    n1560
  );


  buf
  g1696
  (
    n1753,
    n1506
  );


  not
  g1697
  (
    n1659,
    n1566
  );


  buf
  g1698
  (
    n1606,
    n1529
  );


  buf
  g1699
  (
    n1762,
    n1412
  );


  not
  g1700
  (
    n1620,
    n1498
  );


  not
  g1701
  (
    n1738,
    n1431
  );


  not
  g1702
  (
    n1611,
    n1479
  );


  buf
  g1703
  (
    n1656,
    n1467
  );


  buf
  g1704
  (
    n1840,
    n1437
  );


  not
  g1705
  (
    n1632,
    n1432
  );


  not
  g1706
  (
    n1618,
    n1471
  );


  not
  g1707
  (
    n1657,
    n1414
  );


  not
  g1708
  (
    n1854,
    n1437
  );


  buf
  g1709
  (
    n1816,
    n1402
  );


  not
  g1710
  (
    n1733,
    n1479
  );


  buf
  g1711
  (
    n1658,
    n1546
  );


  buf
  g1712
  (
    n1637,
    n1473
  );


  not
  g1713
  (
    n1689,
    n1459
  );


  buf
  g1714
  (
    n1748,
    n1420
  );


  not
  g1715
  (
    n1802,
    n1528
  );


  not
  g1716
  (
    n1625,
    n1459
  );


  buf
  g1717
  (
    n1725,
    n1453
  );


  buf
  g1718
  (
    n1703,
    n1442
  );


  buf
  g1719
  (
    n1817,
    n1502
  );


  not
  g1720
  (
    n1788,
    n1409
  );


  buf
  g1721
  (
    n1867,
    n1391
  );


  buf
  g1722
  (
    n1781,
    n1496
  );


  not
  g1723
  (
    n1694,
    n1411
  );


  buf
  g1724
  (
    n1803,
    n1537
  );


  buf
  g1725
  (
    n1844,
    n1509
  );


  buf
  g1726
  (
    n1683,
    n1448
  );


  not
  g1727
  (
    KeyWire_0_53,
    n1450
  );


  not
  g1728
  (
    n1685,
    n1430
  );


  buf
  g1729
  (
    n1596,
    n1521
  );


  not
  g1730
  (
    n1848,
    n1516
  );


  buf
  g1731
  (
    n1809,
    n1547
  );


  not
  g1732
  (
    n1645,
    n1462
  );


  not
  g1733
  (
    n1864,
    n1543
  );


  not
  g1734
  (
    n1749,
    n1426
  );


  buf
  g1735
  (
    n1862,
    n1458
  );


  buf
  g1736
  (
    n1701,
    n1526
  );


  buf
  g1737
  (
    n1608,
    n1546
  );


  not
  g1738
  (
    n1785,
    n1510
  );


  buf
  g1739
  (
    n1678,
    n1407
  );


  buf
  g1740
  (
    n1661,
    n1525
  );


  not
  g1741
  (
    n1734,
    n1412
  );


  buf
  g1742
  (
    n1808,
    n1476
  );


  not
  g1743
  (
    n1828,
    n1528
  );


  buf
  g1744
  (
    n1787,
    n1477
  );


  buf
  g1745
  (
    n1770,
    n1439
  );


  buf
  g1746
  (
    n1648,
    n1406
  );


  not
  g1747
  (
    n1609,
    n1534
  );


  buf
  g1748
  (
    n1810,
    n1479
  );


  or
  g1749
  (
    n1697,
    n1485,
    n1506,
    n1465,
    n1555
  );


  xor
  g1750
  (
    n1676,
    n1484,
    n1552,
    n1478,
    n1424
  );


  and
  g1751
  (
    n1710,
    n1416,
    n1422,
    n1551,
    n1524
  );


  or
  g1752
  (
    n1772,
    n1503,
    n1452,
    n1486,
    n1457
  );


  xnor
  g1753
  (
    n1755,
    n1519,
    n1412,
    n1436,
    n1534
  );


  nand
  g1754
  (
    n1825,
    n1432,
    n1489,
    n1563,
    n1439
  );


  xnor
  g1755
  (
    n1714,
    n1428,
    n1425,
    n1430,
    n1407
  );


  xor
  g1756
  (
    n1823,
    n1495,
    n1549,
    n1405,
    n1441
  );


  nand
  g1757
  (
    n1720,
    n1544,
    n1541,
    n1475,
    n1429
  );


  xor
  g1758
  (
    n1789,
    n1452,
    n1474,
    n1513,
    n1435
  );


  nand
  g1759
  (
    n1807,
    n1463,
    n1494,
    n1487,
    n1466
  );


  nor
  g1760
  (
    n1623,
    n1469,
    n1558,
    n1391,
    n1481
  );


  and
  g1761
  (
    n1680,
    n1450,
    n1527,
    n1460,
    n1524
  );


  xnor
  g1762
  (
    n1626,
    n1389,
    n1404,
    n1393,
    n1390
  );


  xnor
  g1763
  (
    n1715,
    n1508,
    n1458,
    n1519,
    n1482
  );


  xor
  g1764
  (
    n1849,
    n1461,
    n1563,
    n1463,
    n1513
  );


  xor
  g1765
  (
    n1830,
    n1550,
    n1541,
    n1504,
    n1421
  );


  nor
  g1766
  (
    n1664,
    n1553,
    n1452,
    n1545,
    n1409
  );


  nand
  g1767
  (
    n1732,
    n1498,
    n1472,
    n1393,
    n1477
  );


  nand
  g1768
  (
    n1706,
    n1491,
    n1433,
    n1455,
    n1424
  );


  nor
  g1769
  (
    n1858,
    n1440,
    n1485,
    n1493,
    n1417
  );


  nor
  g1770
  (
    n1795,
    n1535,
    n1441,
    n1525,
    n1471
  );


  or
  g1771
  (
    n1696,
    n1440,
    n1488,
    n1553,
    n1471
  );


  nor
  g1772
  (
    n1759,
    n1527,
    n1426,
    n1450,
    n1521
  );


  or
  g1773
  (
    n1847,
    n1468,
    n1456,
    n1518,
    n1561
  );


  nor
  g1774
  (
    n1700,
    n1420,
    n1530,
    n1394,
    n1505
  );


  xnor
  g1775
  (
    n1829,
    n1456,
    n1473,
    n1545,
    n1424
  );


  and
  g1776
  (
    n1761,
    n1399,
    n1455,
    n1492,
    n1396
  );


  nor
  g1777
  (
    n1866,
    n1408,
    n1556,
    n1431,
    n1448
  );


  xor
  g1778
  (
    n1745,
    n1480,
    n1451,
    n1403,
    n1435
  );


  xor
  g1779
  (
    n1647,
    n1504,
    n1561,
    n1501,
    n1401
  );


  xnor
  g1780
  (
    n1804,
    n1522,
    n1545,
    n1533,
    n1414
  );


  xor
  g1781
  (
    n1693,
    n1453,
    n1438,
    n1394,
    n1562
  );


  xor
  g1782
  (
    n1709,
    n1543,
    n1530,
    n1532,
    n1536
  );


  or
  g1783
  (
    n1621,
    n1514,
    n1526,
    n1560,
    n1516
  );


  or
  g1784
  (
    n1613,
    n1392,
    n1563,
    n1519,
    n1554
  );


  nor
  g1785
  (
    n1636,
    n1550,
    n1487,
    n1432,
    n1434
  );


  and
  g1786
  (
    n1607,
    n1401,
    n1451,
    n1465,
    n1566
  );


  nand
  g1787
  (
    n1716,
    n1420,
    n1445,
    n1418,
    n1469
  );


  xnor
  g1788
  (
    n1668,
    n1495,
    n1441,
    n1413,
    n1508
  );


  and
  g1789
  (
    n1719,
    n1408,
    n1417,
    n1522,
    n1458
  );


  nand
  g1790
  (
    n1698,
    n1413,
    n1405,
    n1392,
    n1555
  );


  xor
  g1791
  (
    n1775,
    n1468,
    n1505,
    n1390,
    n1547
  );


  nand
  g1792
  (
    n1627,
    n1548,
    n1512,
    n1444,
    n1539
  );


  nand
  g1793
  (
    n1604,
    n1472,
    n1419,
    n1470,
    n1425
  );


  or
  g1794
  (
    n1756,
    n1435,
    n1461,
    n1510,
    n1422
  );


  nor
  g1795
  (
    n1717,
    n1478,
    n1525,
    n1439,
    n1445
  );


  or
  g1796
  (
    n1801,
    n1527,
    n1549,
    n1559,
    n1506
  );


  nor
  g1797
  (
    n1790,
    n1489,
    n1411,
    n1537,
    n1438
  );


  xor
  g1798
  (
    n1859,
    n1457,
    n1542,
    n1564,
    n1491
  );


  xnor
  g1799
  (
    n1704,
    n1472,
    n1536,
    n1443,
    n1499
  );


  xnor
  g1800
  (
    n1782,
    n1499,
    n1490,
    n1411,
    n1475
  );


  nor
  g1801
  (
    n1771,
    n1542,
    n1397,
    n1443,
    n1419
  );


  xnor
  g1802
  (
    n1595,
    n1449,
    n1410,
    n1507,
    n1531
  );


  nand
  g1803
  (
    n1768,
    n1475,
    n1400,
    n1555,
    n1559
  );


  xor
  g1804
  (
    n1784,
    n1565,
    n1401,
    n1398,
    n1544
  );


  xnor
  g1805
  (
    n1630,
    n1431,
    n1524,
    n1515,
    n1433
  );


  nand
  g1806
  (
    n1679,
    n1491,
    n1427,
    n1455,
    n1532
  );


  and
  g1807
  (
    n1764,
    n1446,
    n1444,
    n1495,
    n1485
  );


  and
  g1808
  (
    n1617,
    n1436,
    n1396,
    n1428,
    n1402
  );


  xor
  g1809
  (
    n1651,
    n1497,
    n1448,
    n1515,
    n1399
  );


  nand
  g1810
  (
    n1729,
    n1513,
    n1466,
    n1408,
    n1551
  );


  or
  g1811
  (
    n1834,
    n1486,
    n1535,
    n1410,
    n1454
  );


  nand
  g1812
  (
    n1707,
    n1449,
    n1467,
    n1461,
    n1538
  );


  nor
  g1813
  (
    n1820,
    n1454,
    n1398,
    n1395,
    n1564
  );


  and
  g1814
  (
    n1652,
    n1389,
    n1427,
    n1493,
    n1392
  );


  xnor
  g1815
  (
    n1792,
    n1537,
    n1395,
    n1463,
    n1464
  );


  xnor
  g1816
  (
    n1601,
    n1481,
    n1413,
    n1487,
    n1395
  );


  and
  g1817
  (
    n1766,
    n1529,
    n1502,
    n1517,
    n1404
  );


  xnor
  g1818
  (
    n1746,
    n1406,
    n1397,
    n1547,
    n1480
  );


  nor
  g1819
  (
    n1675,
    n1469,
    n1518,
    n1556,
    n1565
  );


  xor
  g1820
  (
    n1812,
    n1558,
    n1447,
    n1559,
    n1522
  );


  nand
  g1821
  (
    n1839,
    n1442,
    n1423,
    n1486,
    n1548
  );


  or
  g1822
  (
    n1677,
    n1410,
    n1500,
    n1418,
    n1483
  );


  xor
  g1823
  (
    n1821,
    n1511,
    n1554,
    n1557,
    n1483
  );


  nand
  g1824
  (
    KeyWire_0_51,
    n1429,
    n1468,
    n1457,
    n1540
  );


  and
  g1825
  (
    KeyWire_0_44,
    n1447,
    n1536,
    n1460,
    n1436
  );


  and
  g1826
  (
    n1629,
    n1554,
    n1488,
    n1496,
    n1407
  );


  xor
  g1827
  (
    n1688,
    n1548,
    n1400,
    n1480,
    n1523
  );


  xor
  g1828
  (
    n1641,
    n1507,
    n1526,
    n1394,
    n1474
  );


  nand
  g1829
  (
    n1838,
    n1460,
    n1512,
    n1393,
    n1403
  );


  xor
  g1830
  (
    KeyWire_0_2,
    n1484,
    n1517,
    n1535,
    n1454
  );


  or
  g1831
  (
    n1670,
    n1440,
    n1492,
    n1391,
    n1477
  );


  xnor
  g1832
  (
    n1856,
    n1498,
    n1549,
    n1546,
    n1434
  );


  nor
  g1833
  (
    n1743,
    n1416,
    n1402,
    n1483,
    n1518
  );


  nand
  g1834
  (
    n1614,
    n1484,
    n1459,
    n1508,
    n1398
  );


  or
  g1835
  (
    n2057,
    n1610,
    n1724,
    n1773
  );


  nor
  g1836
  (
    n1993,
    n1763,
    n1739,
    n1617,
    n1727
  );


  and
  g1837
  (
    n2054,
    n1750,
    n1764,
    n1767,
    n1778
  );


  xor
  g1838
  (
    n2095,
    n1615,
    n1651,
    n1810,
    n1769
  );


  xnor
  g1839
  (
    n1931,
    n1653,
    n1771,
    n1792,
    n1819
  );


  nand
  g1840
  (
    n1897,
    n1662,
    n1833,
    n1817,
    n1863
  );


  xnor
  g1841
  (
    n1919,
    n1785,
    n1831,
    n1847,
    n1651
  );


  nor
  g1842
  (
    n1962,
    n1751,
    n1802,
    n1786,
    n1853
  );


  nand
  g1843
  (
    n2096,
    n1640,
    n1699,
    n1655,
    n1826
  );


  nand
  g1844
  (
    n2004,
    n1638,
    n1867,
    n1809
  );


  or
  g1845
  (
    n2043,
    n1835,
    n1629,
    n1813,
    n1805
  );


  xor
  g1846
  (
    n2014,
    n1749,
    n1648,
    n1865,
    n1654
  );


  nand
  g1847
  (
    n1982,
    n1804,
    n1780,
    n1772,
    n1836
  );


  or
  g1848
  (
    n1901,
    n1689,
    n1851,
    n1726,
    n1724
  );


  xnor
  g1849
  (
    n2045,
    n1862,
    n1598,
    n1863,
    n1731
  );


  xnor
  g1850
  (
    n2023,
    n1738,
    n1647,
    n1794,
    n1743
  );


  and
  g1851
  (
    n2033,
    n1728,
    n1693,
    n1725,
    n1752
  );


  nand
  g1852
  (
    n1898,
    n1756,
    n1719,
    n1811,
    n1832
  );


  nand
  g1853
  (
    n1927,
    n1759,
    n1630,
    n1645,
    n1824
  );


  nor
  g1854
  (
    n2080,
    n1771,
    n1806,
    n1745,
    n1625
  );


  and
  g1855
  (
    n1921,
    n1771,
    n1670,
    n1793,
    n1617
  );


  nor
  g1856
  (
    n1913,
    n1818,
    n1852,
    n1694,
    n1771
  );


  or
  g1857
  (
    KeyWire_0_7,
    n1693,
    n1776,
    n1707,
    n1600
  );


  xnor
  g1858
  (
    n1974,
    n1594,
    n1717,
    n1643,
    n1618
  );


  or
  g1859
  (
    n2030,
    n1657,
    n1631,
    n1781,
    n1768
  );


  nand
  g1860
  (
    n1997,
    n1664,
    n1777,
    n1822,
    n1593
  );


  nand
  g1861
  (
    n1926,
    n1796,
    n1660,
    n1647,
    n1848
  );


  and
  g1862
  (
    n2021,
    n1821,
    n1814,
    n1692,
    n1798
  );


  and
  g1863
  (
    n1975,
    n1779,
    n1856,
    n1748,
    n1815
  );


  xnor
  g1864
  (
    n2031,
    n1838,
    n1832,
    n1763,
    n1825
  );


  xor
  g1865
  (
    KeyWire_0_47,
    n1851,
    n1646,
    n1601,
    n1742
  );


  or
  g1866
  (
    n2051,
    n1661,
    n1625,
    n1805,
    n1607
  );


  and
  g1867
  (
    n2044,
    n1678,
    n1717,
    n1750,
    n1744
  );


  xnor
  g1868
  (
    n1888,
    n1857,
    n1816,
    n1612,
    n1811
  );


  and
  g1869
  (
    n1960,
    n1746,
    n1837,
    n1666,
    n1735
  );


  xnor
  g1870
  (
    n2029,
    n1628,
    n1824,
    n1849,
    n1659
  );


  and
  g1871
  (
    n1949,
    n1806,
    n1847,
    n1732,
    n1858
  );


  xor
  g1872
  (
    n1992,
    n1702,
    n1711,
    n1622,
    n1817
  );


  xor
  g1873
  (
    n1900,
    n1821,
    n1732,
    n1709,
    n1635
  );


  nand
  g1874
  (
    n1968,
    n1773,
    n1866,
    n1598,
    n1698
  );


  nor
  g1875
  (
    n1877,
    n1663,
    n1741,
    n1840,
    n1666
  );


  xor
  g1876
  (
    n2099,
    n1866,
    n1620,
    n1692,
    n1769
  );


  nor
  g1877
  (
    n2022,
    n1815,
    n1604,
    n1643,
    n1647
  );


  xnor
  g1878
  (
    n2066,
    n1824,
    n1853,
    n1645,
    n1601
  );


  and
  g1879
  (
    n2105,
    n1858,
    n1787,
    n1661,
    n1750
  );


  nand
  g1880
  (
    n1943,
    n1614,
    n1758,
    n1768,
    n1836
  );


  nor
  g1881
  (
    n2053,
    n1792,
    n876,
    n1778,
    n1851
  );


  xor
  g1882
  (
    n2087,
    n1859,
    n1700,
    n1687,
    n1852
  );


  or
  g1883
  (
    n2058,
    n1616,
    n1766,
    n1836,
    n1644
  );


  nor
  g1884
  (
    n1893,
    n1854,
    n1854,
    n1638,
    n1773
  );


  xor
  g1885
  (
    n1933,
    n1688,
    n1807,
    n1637,
    n1772
  );


  or
  g1886
  (
    n2035,
    n1777,
    n1839,
    n1751,
    n1649
  );


  nand
  g1887
  (
    n1907,
    n1844,
    n1730,
    n1713,
    n1599
  );


  nand
  g1888
  (
    n2078,
    n1703,
    n1667,
    n1849,
    n1704
  );


  and
  g1889
  (
    n2089,
    n1672,
    n1678,
    n1755,
    n1744
  );


  xnor
  g1890
  (
    n1883,
    n1837,
    n1656,
    n1674,
    n1862
  );


  xor
  g1891
  (
    n1902,
    n1753,
    n1749,
    n1748,
    n1682
  );


  xor
  g1892
  (
    n1892,
    n1685,
    n1766,
    n1834,
    n1760
  );


  xor
  g1893
  (
    n1956,
    n1724,
    n1704,
    n1745,
    n1676
  );


  or
  g1894
  (
    n1872,
    n1846,
    n1719,
    n1842,
    n1693
  );


  nand
  g1895
  (
    n2050,
    n1780,
    n1708,
    n1727,
    n1624
  );


  and
  g1896
  (
    n1976,
    n1658,
    n1757,
    n1828,
    n1837
  );


  xor
  g1897
  (
    n2003,
    n1653,
    n1787,
    n1797,
    n1835
  );


  xor
  g1898
  (
    n1881,
    n1631,
    n1711,
    n1822,
    n1832
  );


  xnor
  g1899
  (
    n2040,
    n1689,
    n1810,
    n1619,
    n1625
  );


  xnor
  g1900
  (
    n2064,
    n1840,
    n1767,
    n1662,
    n1766
  );


  or
  g1901
  (
    n2032,
    n1859,
    n1609,
    n1646,
    n1780
  );


  nand
  g1902
  (
    n1991,
    n1609,
    n1861,
    n1845,
    n1732
  );


  xor
  g1903
  (
    n1894,
    n1644,
    n1850,
    n1715,
    n1646
  );


  or
  g1904
  (
    n1879,
    n1756,
    n1697,
    n1698,
    n1740
  );


  xnor
  g1905
  (
    n1905,
    n1708,
    n1736,
    n1810,
    n1638
  );


  and
  g1906
  (
    n1923,
    n1594,
    n1686,
    n1800,
    n1669
  );


  and
  g1907
  (
    n2083,
    n1619,
    n1700,
    n1841,
    n1636
  );


  nor
  g1908
  (
    n1918,
    n1839,
    n1769,
    n1793,
    n1829
  );


  xor
  g1909
  (
    n2055,
    n1857,
    n1630,
    n1850,
    n1602
  );


  nand
  g1910
  (
    n1970,
    n1783,
    n1765,
    n1800
  );


  and
  g1911
  (
    n1990,
    n1803,
    n1854,
    n1645,
    n1752
  );


  xor
  g1912
  (
    n2079,
    n1681,
    n1769,
    n1816,
    n1803
  );


  xor
  g1913
  (
    n2034,
    n1792,
    n1670,
    n1619,
    n1616
  );


  nand
  g1914
  (
    n1942,
    n1705,
    n1691,
    n1776,
    n1861
  );


  nand
  g1915
  (
    n1938,
    n1737,
    n1855,
    n1796,
    n1655
  );


  and
  g1916
  (
    n2093,
    n1667,
    n1791,
    n1668,
    n1752
  );


  nor
  g1917
  (
    n2009,
    n1606,
    n1595,
    n1776,
    n1781
  );


  nand
  g1918
  (
    n1920,
    n1828,
    n1798,
    n1637,
    n1751
  );


  nor
  g1919
  (
    n1891,
    n1622,
    n1815,
    n1747,
    n1783
  );


  nand
  g1920
  (
    n2097,
    n1790,
    n1652,
    n1856,
    n1678
  );


  nand
  g1921
  (
    n1939,
    n1627,
    n1617,
    n1768,
    n1754
  );


  nand
  g1922
  (
    n1945,
    n1721,
    n1705,
    n1758,
    n1599
  );


  nor
  g1923
  (
    n2102,
    n1747,
    n1728,
    n1839,
    n1827
  );


  nand
  g1924
  (
    n2075,
    n1740,
    n1614,
    n1597,
    n1630
  );


  xor
  g1925
  (
    n2008,
    n1746,
    n1675,
    n1687,
    n1629
  );


  or
  g1926
  (
    n2059,
    n1844,
    n1850,
    n1785,
    n1718
  );


  and
  g1927
  (
    n2047,
    n1616,
    n1844,
    n1773,
    n1671
  );


  or
  g1928
  (
    n1971,
    n1811,
    n1829,
    n1748,
    n1666
  );


  nor
  g1929
  (
    n2073,
    n1673,
    n1855,
    n1742,
    n1818
  );


  nand
  g1930
  (
    n1989,
    n1749,
    n1642,
    n1640,
    n1597
  );


  and
  g1931
  (
    n1870,
    n1731,
    n1593,
    n1814,
    n1603
  );


  or
  g1932
  (
    n2037,
    n876,
    n1790,
    n1757,
    n1793
  );


  or
  g1933
  (
    n1899,
    n1782,
    n1861,
    n1767,
    n1786
  );


  xor
  g1934
  (
    n2024,
    n1827,
    n1809,
    n1761,
    n1670
  );


  xor
  g1935
  (
    n2060,
    n1611,
    n1650,
    n1690,
    n1715
  );


  or
  g1936
  (
    n1996,
    n1794,
    n1777,
    n1774,
    n1845
  );


  xnor
  g1937
  (
    n1985,
    n1761,
    n1799,
    n1634,
    n1736
  );


  and
  g1938
  (
    n1908,
    n1661,
    n1809,
    n1755,
    n1720
  );


  xnor
  g1939
  (
    n2006,
    n1820,
    n1703,
    n1813,
    n1860
  );


  xor
  g1940
  (
    n2001,
    n1608,
    n1823,
    n1834,
    n1730
  );


  and
  g1941
  (
    n2109,
    n1741,
    n1747,
    n1701,
    n1743
  );


  and
  g1942
  (
    n1957,
    n1730,
    n1860,
    n1841,
    n1808
  );


  nor
  g1943
  (
    n1884,
    n1801,
    n1663,
    n1825,
    n1826
  );


  xnor
  g1944
  (
    n1961,
    n1743,
    n1802,
    n1715,
    n1753
  );


  nor
  g1945
  (
    n1986,
    n1750,
    n1679,
    n1827,
    n1798
  );


  and
  g1946
  (
    n2027,
    n1758,
    n1639,
    n1714,
    n1687
  );


  or
  g1947
  (
    n1914,
    n1796,
    n1861,
    n1823,
    n1784
  );


  xor
  g1948
  (
    n1965,
    n1680,
    n1831,
    n1760,
    n1801
  );


  xnor
  g1949
  (
    n1966,
    n1779,
    n1644,
    n1764,
    n1816
  );


  and
  g1950
  (
    n2063,
    n1694,
    n1657,
    n1611,
    n1814
  );


  nor
  g1951
  (
    n1922,
    n1680,
    n1867,
    n1658,
    n1846
  );


  and
  g1952
  (
    n1889,
    n1781,
    n1866,
    n1603,
    n1706
  );


  nand
  g1953
  (
    n1994,
    n1723,
    n1762,
    n1620,
    n1600
  );


  xor
  g1954
  (
    n1932,
    n1770,
    n1723,
    n1843,
    n1613
  );


  xor
  g1955
  (
    n2094,
    n1852,
    n1702,
    n1822,
    n1805
  );


  xor
  g1956
  (
    n2065,
    n1686,
    n1841,
    n1852,
    n1767
  );


  xor
  g1957
  (
    n1953,
    n1677,
    n1793,
    n1600,
    n1842
  );


  and
  g1958
  (
    n1959,
    n1720,
    n1780,
    n1669,
    n1795
  );


  nor
  g1959
  (
    n2077,
    n1800,
    n1681,
    n1599,
    n1736
  );


  or
  g1960
  (
    n1978,
    n1820,
    n1795,
    n1862,
    n1653
  );


  xor
  g1961
  (
    n1925,
    n1825,
    n1739,
    n1786,
    n1709
  );


  and
  g1962
  (
    n1885,
    n1754,
    n1620,
    n1855,
    n1709
  );


  nor
  g1963
  (
    n2015,
    n1833,
    n1598,
    n1795,
    n1839
  );


  and
  g1964
  (
    n1895,
    n1808,
    n1691,
    n1834,
    n1858
  );


  or
  g1965
  (
    n2071,
    n1792,
    n1702,
    n1740,
    n1765
  );


  nand
  g1966
  (
    n1874,
    n1830,
    n1819,
    n1854,
    n1853
  );


  nor
  g1967
  (
    n1930,
    n1662,
    n1648,
    n1602,
    n1712
  );


  xor
  g1968
  (
    n2026,
    n1779,
    n1731,
    n1716,
    n1787
  );


  nor
  g1969
  (
    n2005,
    n1706,
    n1744,
    n1805,
    n1681
  );


  nand
  g1970
  (
    n2098,
    n1679,
    n1615,
    n1783,
    n1634
  );


  xor
  g1971
  (
    n2061,
    n1635,
    n1742,
    n1609,
    n1778
  );


  nand
  g1972
  (
    n1929,
    n1833,
    n1757,
    n1789,
    n1716
  );


  xor
  g1973
  (
    n2062,
    n1745,
    n1824,
    n1831,
    n1711
  );


  xor
  g1974
  (
    n1904,
    n1853,
    n1735,
    n1733,
    n1808
  );


  xor
  g1975
  (
    n1967,
    n1679,
    n1747,
    n1838,
    n1845
  );


  or
  g1976
  (
    n2017,
    n1622,
    n1682,
    n1807,
    n1848
  );


  xor
  g1977
  (
    n2090,
    n1665,
    n1665,
    n1676,
    n1796
  );


  nand
  g1978
  (
    n1878,
    n1856,
    n1775,
    n1728,
    n1826
  );


  xor
  g1979
  (
    KeyWire_0_23,
    n1651,
    n1763,
    n1642,
    n1789
  );


  xor
  g1980
  (
    n2048,
    n1789,
    n1639,
    n1741,
    n1768
  );


  xor
  g1981
  (
    n1979,
    n1610,
    n1699,
    n1607,
    n1779
  );


  xor
  g1982
  (
    n2052,
    n1716,
    n1755,
    n1605
  );


  or
  g1983
  (
    n1999,
    n1718,
    n1688,
    n1772,
    n1728
  );


  nand
  g1984
  (
    n1868,
    n1836,
    n1722,
    n1596,
    n1672
  );


  xnor
  g1985
  (
    n2088,
    n1696,
    n1684,
    n1634,
    n1725
  );


  xnor
  g1986
  (
    n2081,
    n1683,
    n1812,
    n1766,
    n1735
  );


  xnor
  g1987
  (
    n2011,
    n1837,
    n1604,
    n1865,
    n1818
  );


  xnor
  g1988
  (
    n2108,
    n1631,
    n1636,
    n1683,
    n1727
  );


  xor
  g1989
  (
    n1935,
    n1737,
    n1738,
    n1729,
    n1843
  );


  xnor
  g1990
  (
    n1998,
    n1848,
    n1732,
    n1605,
    n1677
  );


  xnor
  g1991
  (
    n1951,
    n1821,
    n1632,
    n1849,
    n1734
  );


  or
  g1992
  (
    n1890,
    n1650,
    n1710,
    n1596,
    n1602
  );


  and
  g1993
  (
    n2039,
    n1621,
    n1759,
    n1751,
    n1774
  );


  or
  g1994
  (
    n2038,
    n1674,
    n1828,
    n1788
  );


  nand
  g1995
  (
    n1886,
    n1695,
    n1633,
    n1660,
    n1847
  );


  nand
  g1996
  (
    n2007,
    n1867,
    n1683,
    n1641,
    n1698
  );


  and
  g1997
  (
    n2085,
    n1731,
    n1640,
    n1812,
    n1794
  );


  xor
  g1998
  (
    n2068,
    n1659,
    n1833,
    n1627,
    n1611
  );


  nand
  g1999
  (
    n1928,
    n1803,
    n1695,
    n1774,
    n1760
  );


  xor
  g2000
  (
    n2049,
    n1733,
    n1739,
    n1626,
    n1760
  );


  xor
  g2001
  (
    n2104,
    n1817,
    n1648,
    n1772,
    n1729
  );


  nor
  g2002
  (
    n1948,
    n1825,
    n1729,
    n1593,
    n1813
  );


  or
  g2003
  (
    n2000,
    n1810,
    n1791,
    n1820,
    n1764
  );


  xor
  g2004
  (
    n1924,
    n1830,
    n1685,
    n1744,
    n1814
  );


  xnor
  g2005
  (
    n1980,
    n1596,
    n1633,
    n1710,
    n1729
  );


  nor
  g2006
  (
    n2074,
    n1850,
    n1864,
    n1673,
    n1804
  );


  nor
  g2007
  (
    n2018,
    n1691,
    n1739,
    n1684,
    n1781
  );


  xor
  g2008
  (
    n2067,
    n1746,
    n1735,
    n1822,
    n1668
  );


  xor
  g2009
  (
    n1969,
    n1841,
    n1775,
    n1860,
    n1655
  );


  xnor
  g2010
  (
    n2046,
    n1802,
    n1782,
    n1770,
    n1734
  );


  xnor
  g2011
  (
    n1950,
    n1753,
    n1675,
    n1829,
    n1797
  );


  nor
  g2012
  (
    n2082,
    n1690,
    n1806,
    n1712,
    n1743
  );


  xnor
  g2013
  (
    n2016,
    n1832,
    n1606,
    n1787,
    n1632
  );


  and
  g2014
  (
    n1958,
    n1817,
    n1788,
    n1756
  );


  nand
  g2015
  (
    n2106,
    n1774,
    n1749,
    n1838,
    n1758
  );


  or
  g2016
  (
    n1946,
    n1721,
    n1764,
    n1858,
    n1842
  );


  xor
  g2017
  (
    n2013,
    n1594,
    n1826,
    n1628,
    n1701
  );


  nand
  g2018
  (
    n2002,
    n1624,
    n1707,
    n1677,
    n1788
  );


  nor
  g2019
  (
    n1977,
    n1790,
    n1804,
    n1782,
    n1763
  );


  xor
  g2020
  (
    n1937,
    n1688,
    n1762,
    n1613,
    n1777
  );


  and
  g2021
  (
    n2107,
    n1829,
    n1656,
    n1799,
    n1652
  );


  or
  g2022
  (
    n1952,
    n1626,
    n1615,
    n1790,
    n1865
  );


  and
  g2023
  (
    n1995,
    n1862,
    n1671,
    n1664,
    n1714
  );


  nor
  g2024
  (
    n1873,
    n1799,
    n1765,
    n1797,
    n1848
  );


  or
  g2025
  (
    n2101,
    n1761,
    n1613,
    n1843,
    n1737
  );


  xor
  g2026
  (
    n2086,
    n1710,
    n1717,
    n1820,
    n1808
  );


  xnor
  g2027
  (
    n1912,
    n1775,
    n1610,
    n1612,
    n1601
  );


  and
  g2028
  (
    n2103,
    n1756,
    n1641,
    n1700,
    n1675
  );


  or
  g2029
  (
    n1876,
    n1784,
    n1633,
    n1778,
    n1801
  );


  xnor
  g2030
  (
    n1941,
    n1855,
    n1738,
    n1674,
    n1657
  );


  and
  g2031
  (
    n1903,
    n1618,
    n1673,
    n1621
  );


  and
  g2032
  (
    n1911,
    n1714,
    n1685,
    n1762,
    n1713
  );


  nand
  g2033
  (
    n2019,
    n1725,
    n1754,
    n1775,
    n1737
  );


  and
  g2034
  (
    n2041,
    n1863,
    n1618,
    n1605,
    n1761
  );


  xnor
  g2035
  (
    n2076,
    n1608,
    n1669,
    n1671,
    n1734
  );


  xor
  g2036
  (
    KeyWire_0_39,
    n1759,
    n1819,
    n1718,
    n1806
  );


  or
  g2037
  (
    n1906,
    n1804,
    n1838,
    n1746,
    n1639
  );


  xnor
  g2038
  (
    n1988,
    n1843,
    n1695,
    n1807,
    n1726
  );


  nor
  g2039
  (
    n2072,
    n1652,
    n1595,
    n1786,
    n1686
  );


  nand
  g2040
  (
    n2100,
    n1859,
    n1849,
    n1738,
    n1667
  );


  xnor
  g2041
  (
    n1940,
    n1704,
    n1864,
    n1623,
    n1707
  );


  and
  g2042
  (
    n2069,
    n1803,
    n1722,
    n1672,
    n1658
  );


  nor
  g2043
  (
    n2010,
    n1740,
    n1834,
    n1783,
    n1623
  );


  and
  g2044
  (
    n1983,
    n1723,
    n1851,
    n1641,
    n1847
  );


  nor
  g2045
  (
    n1936,
    n1776,
    n1665,
    n1608,
    n1595
  );


  nor
  g2046
  (
    n1947,
    n1840,
    n1656,
    n1720,
    n876
  );


  nor
  g2047
  (
    n1981,
    n1628,
    n1762,
    n1799,
    n1785
  );


  xor
  g2048
  (
    n2092,
    n1705,
    n1654,
    n1845,
    n1831
  );


  and
  g2049
  (
    n2028,
    n1835,
    n1818,
    n1789,
    n1629
  );


  xnor
  g2050
  (
    n2042,
    n1813,
    n1697,
    n1694,
    n1637
  );


  or
  g2051
  (
    n1910,
    n1752,
    n1701,
    n1866,
    n1753
  );


  nand
  g2052
  (
    n1916,
    n1741,
    n1604,
    n1736,
    n1807
  );


  xnor
  g2053
  (
    n1882,
    n1812,
    n1726,
    n1815,
    n1692
  );


  xnor
  g2054
  (
    n2070,
    n1865,
    n1830,
    n1734,
    n1800
  );


  nor
  g2055
  (
    n2036,
    n1597,
    n1795,
    n1770,
    n1797
  );


  or
  g2056
  (
    n1887,
    n1816,
    n1791,
    n1819,
    n1754
  );


  nand
  g2057
  (
    n1944,
    n1823,
    n1835,
    n1642,
    n1857
  );


  or
  g2058
  (
    n1973,
    n1730,
    n1636,
    n1770,
    n1624
  );


  or
  g2059
  (
    n2084,
    n1676,
    n1632,
    n1846,
    n1699
  );


  nand
  g2060
  (
    n2020,
    n1660,
    n1654,
    n1612,
    n1857
  );


  or
  g2061
  (
    n1963,
    n1842,
    n1650,
    n1856,
    n1860
  );


  nand
  g2062
  (
    n1869,
    n1643,
    n1680,
    n1614,
    n1757
  );


  nor
  g2063
  (
    n1917,
    n1649,
    n1844,
    n1719,
    n1713
  );


  nand
  g2064
  (
    n2091,
    n1682,
    n1712,
    n1823,
    n1802
  );


  xor
  g2065
  (
    n2012,
    n1703,
    n1627,
    n1708,
    n1785
  );


  nor
  g2066
  (
    n2056,
    n1784,
    n1668,
    n1859,
    n1684
  );


  and
  g2067
  (
    n1972,
    n1811,
    n1784,
    n1626,
    n1748
  );


  or
  g2068
  (
    n1955,
    n1663,
    n1690,
    n1697,
    n1649
  );


  xnor
  g2069
  (
    n1880,
    n1607,
    n1759,
    n1864,
    n1827
  );


  or
  g2070
  (
    n1984,
    n1798,
    n1840,
    n1864,
    n1689
  );


  nor
  g2071
  (
    n1954,
    n1794,
    n1782,
    n1812,
    n1733
  );


  xor
  g2072
  (
    n2025,
    n1863,
    n1623,
    n1659,
    n1742
  );


  xnor
  g2073
  (
    n1964,
    n1830,
    n1696,
    n1721,
    n1722
  );


  xnor
  g2074
  (
    n1896,
    n1821,
    n1846,
    n1696,
    n1791
  );


  xnor
  g2075
  (
    n1871,
    n1606,
    n1706,
    n1635,
    n1801
  );


  xnor
  g2076
  (
    n1934,
    n1664,
    n1603,
    n1745,
    n1733
  );


  not
  g2077
  (
    n2284,
    n1868
  );


  not
  g2078
  (
    n2346,
    n2077
  );


  buf
  g2079
  (
    n2214,
    n2107
  );


  buf
  g2080
  (
    n2369,
    n1928
  );


  buf
  g2081
  (
    n2210,
    n2029
  );


  buf
  g2082
  (
    n2187,
    n1874
  );


  buf
  g2083
  (
    n2192,
    n1947
  );


  buf
  g2084
  (
    n2287,
    n1940
  );


  not
  g2085
  (
    n2254,
    n1896
  );


  not
  g2086
  (
    n2349,
    n2083
  );


  buf
  g2087
  (
    n2286,
    n1936
  );


  not
  g2088
  (
    n2305,
    n2011
  );


  buf
  g2089
  (
    n2304,
    n2044
  );


  buf
  g2090
  (
    n2406,
    n2015
  );


  buf
  g2091
  (
    n2250,
    n1986
  );


  not
  g2092
  (
    n2405,
    n1984
  );


  not
  g2093
  (
    n2398,
    n1920
  );


  buf
  g2094
  (
    n2402,
    n1896
  );


  not
  g2095
  (
    n2249,
    n2039
  );


  not
  g2096
  (
    n2237,
    n1974
  );


  not
  g2097
  (
    n2124,
    n2073
  );


  buf
  g2098
  (
    n2117,
    n1995
  );


  buf
  g2099
  (
    n2309,
    n1990
  );


  not
  g2100
  (
    n2171,
    n2008
  );


  buf
  g2101
  (
    n2256,
    n1977
  );


  not
  g2102
  (
    n2179,
    n2057
  );


  buf
  g2103
  (
    KeyWire_0_18,
    n2019
  );


  not
  g2104
  (
    n2118,
    n2080
  );


  buf
  g2105
  (
    n2359,
    n2086
  );


  not
  g2106
  (
    n2191,
    n1905
  );


  not
  g2107
  (
    n2303,
    n2065
  );


  buf
  g2108
  (
    n2342,
    n2059
  );


  not
  g2109
  (
    n2135,
    n2011
  );


  not
  g2110
  (
    n2112,
    n2098
  );


  buf
  g2111
  (
    n2143,
    n1960
  );


  buf
  g2112
  (
    n2362,
    n2042
  );


  buf
  g2113
  (
    n2272,
    n2046
  );


  not
  g2114
  (
    n2340,
    n2104
  );


  buf
  g2115
  (
    n2306,
    n1873
  );


  not
  g2116
  (
    KeyWire_0_20,
    n2067
  );


  not
  g2117
  (
    n2266,
    n1993
  );


  buf
  g2118
  (
    n2157,
    n2062
  );


  not
  g2119
  (
    n2264,
    n1877
  );


  not
  g2120
  (
    n2328,
    n1991
  );


  buf
  g2121
  (
    n2391,
    n2103
  );


  buf
  g2122
  (
    n2227,
    n1917
  );


  not
  g2123
  (
    n2393,
    n2102
  );


  buf
  g2124
  (
    n2299,
    n1969
  );


  not
  g2125
  (
    n2113,
    n1998
  );


  not
  g2126
  (
    n2208,
    n2025
  );


  buf
  g2127
  (
    n2382,
    n1870
  );


  buf
  g2128
  (
    n2320,
    n2071
  );


  buf
  g2129
  (
    n2373,
    n2074
  );


  buf
  g2130
  (
    n2137,
    n1902
  );


  buf
  g2131
  (
    n2334,
    n1959
  );


  not
  g2132
  (
    n2324,
    n1912
  );


  not
  g2133
  (
    n2313,
    n1994
  );


  not
  g2134
  (
    n2374,
    n1970
  );


  buf
  g2135
  (
    n2132,
    n2101
  );


  not
  g2136
  (
    n2381,
    n1980
  );


  buf
  g2137
  (
    n2224,
    n1918
  );


  buf
  g2138
  (
    n2267,
    n2103
  );


  buf
  g2139
  (
    n2302,
    n2037
  );


  buf
  g2140
  (
    n2253,
    n2092
  );


  not
  g2141
  (
    n2273,
    n1926
  );


  not
  g2142
  (
    n2301,
    n2086
  );


  buf
  g2143
  (
    n2321,
    n1916
  );


  not
  g2144
  (
    n2408,
    n2076
  );


  buf
  g2145
  (
    n2206,
    n2106
  );


  buf
  g2146
  (
    n2262,
    n2079
  );


  buf
  g2147
  (
    n2240,
    n1927
  );


  buf
  g2148
  (
    n2186,
    n1964
  );


  not
  g2149
  (
    n2153,
    n2081
  );


  buf
  g2150
  (
    n2145,
    n1921
  );


  not
  g2151
  (
    KeyWire_0_11,
    n1929
  );


  not
  g2152
  (
    n2185,
    n1931
  );


  not
  g2153
  (
    n2258,
    n1906
  );


  buf
  g2154
  (
    n2167,
    n1963
  );


  not
  g2155
  (
    n2247,
    n1938
  );


  buf
  g2156
  (
    n2181,
    n2021
  );


  buf
  g2157
  (
    n2365,
    n1996
  );


  not
  g2158
  (
    n2239,
    n2093
  );


  buf
  g2159
  (
    n2177,
    n1952
  );


  buf
  g2160
  (
    n2379,
    n1999
  );


  buf
  g2161
  (
    n2163,
    n2095
  );


  not
  g2162
  (
    n2194,
    n2034
  );


  not
  g2163
  (
    n2372,
    n2103
  );


  buf
  g2164
  (
    n2139,
    n2024
  );


  buf
  g2165
  (
    n2400,
    n2098
  );


  buf
  g2166
  (
    n2169,
    n1982
  );


  buf
  g2167
  (
    n2188,
    n2026
  );


  not
  g2168
  (
    n2134,
    n1893
  );


  buf
  g2169
  (
    n2386,
    n1986
  );


  not
  g2170
  (
    n2230,
    n1909
  );


  not
  g2171
  (
    n2147,
    n2055
  );


  not
  g2172
  (
    n2389,
    n1957
  );


  not
  g2173
  (
    n2270,
    n2002
  );


  buf
  g2174
  (
    n2274,
    n2044
  );


  buf
  g2175
  (
    n2300,
    n1919
  );


  not
  g2176
  (
    n2407,
    n2076
  );


  not
  g2177
  (
    n2223,
    n2102
  );


  not
  g2178
  (
    n2367,
    n1981
  );


  buf
  g2179
  (
    n2291,
    n2038
  );


  not
  g2180
  (
    n2218,
    n1943
  );


  buf
  g2181
  (
    n2387,
    n1901
  );


  not
  g2182
  (
    n2268,
    n2003
  );


  buf
  g2183
  (
    n2245,
    n2012
  );


  buf
  g2184
  (
    n2330,
    n2061
  );


  buf
  g2185
  (
    n2332,
    n1991
  );


  not
  g2186
  (
    n2353,
    n2052
  );


  not
  g2187
  (
    n2385,
    n1984
  );


  not
  g2188
  (
    n2370,
    n1879
  );


  buf
  g2189
  (
    n2263,
    n2085
  );


  not
  g2190
  (
    n2115,
    n2006
  );


  buf
  g2191
  (
    n2326,
    n2073
  );


  not
  g2192
  (
    n2279,
    n2098
  );


  not
  g2193
  (
    n2165,
    n1923
  );


  buf
  g2194
  (
    n2388,
    n2027
  );


  not
  g2195
  (
    n2233,
    n2024
  );


  not
  g2196
  (
    n2255,
    n2010
  );


  buf
  g2197
  (
    n2246,
    n1988
  );


  buf
  g2198
  (
    n2390,
    n1932
  );


  not
  g2199
  (
    n2269,
    n1934
  );


  buf
  g2200
  (
    n2307,
    n1959
  );


  buf
  g2201
  (
    n2204,
    n1883
  );


  not
  g2202
  (
    n2184,
    n2107
  );


  nor
  g2203
  (
    n2198,
    n2042,
    n1899,
    n1894,
    n1998
  );


  xnor
  g2204
  (
    n2392,
    n2002,
    n1945,
    n2098,
    n1972
  );


  and
  g2205
  (
    n2211,
    n2051,
    n2007,
    n1966,
    n1954
  );


  nor
  g2206
  (
    n2325,
    n1903,
    n1997,
    n1895,
    n877
  );


  or
  g2207
  (
    n2238,
    n2094,
    n2085,
    n1918,
    n2000
  );


  and
  g2208
  (
    n2352,
    n2107,
    n2101,
    n1930,
    n1882
  );


  or
  g2209
  (
    n2114,
    n1972,
    n1921,
    n2042,
    n1891
  );


  nor
  g2210
  (
    n2158,
    n2031,
    n1988,
    n2104,
    n2106
  );


  xnor
  g2211
  (
    n2244,
    n1949,
    n2029,
    n1934,
    n1948
  );


  xnor
  g2212
  (
    n2354,
    n2082,
    n2094,
    n2030,
    n2054
  );


  or
  g2213
  (
    n2413,
    n1966,
    n2036,
    n1872,
    n1942
  );


  nand
  g2214
  (
    n2156,
    n2018,
    n1958,
    n2024,
    n2092
  );


  xnor
  g2215
  (
    n2275,
    n2009,
    n2003,
    n1994,
    n1933
  );


  xnor
  g2216
  (
    n2182,
    n1965,
    n2063,
    n2019,
    n2099
  );


  or
  g2217
  (
    n2345,
    n1891,
    n2009,
    n2078,
    n1975
  );


  xor
  g2218
  (
    n2251,
    n2004,
    n1880,
    n2093,
    n1995
  );


  xor
  g2219
  (
    n2271,
    n2091,
    n2019,
    n2030,
    n2087
  );


  nor
  g2220
  (
    n2358,
    n2056,
    n1884,
    n1881,
    n1927
  );


  xor
  g2221
  (
    n2197,
    n1936,
    n2038,
    n2075,
    n1946
  );


  nor
  g2222
  (
    n2375,
    n2104,
    n2088,
    n1971,
    n2020
  );


  xnor
  g2223
  (
    n2219,
    n2033,
    n2034,
    n2007,
    n2074
  );


  or
  g2224
  (
    n2243,
    n1958,
    n2031,
    n1987,
    n1922
  );


  xor
  g2225
  (
    n2162,
    n2034,
    n2013,
    n2020,
    n2007
  );


  nand
  g2226
  (
    n2414,
    n2016,
    n1932,
    n1968,
    n2018
  );


  nor
  g2227
  (
    n2344,
    n2026,
    n2008,
    n1973,
    n2083
  );


  or
  g2228
  (
    n2348,
    n1897,
    n2095,
    n2044,
    n2005
  );


  nand
  g2229
  (
    n2129,
    n1871,
    n1914,
    n1951,
    n1973
  );


  xor
  g2230
  (
    n2395,
    n2097,
    n2078,
    n2084,
    n1979
  );


  xnor
  g2231
  (
    n2292,
    n1874,
    n2043,
    n2002,
    n2030
  );


  xnor
  g2232
  (
    n2217,
    n2052,
    n2067,
    n1975,
    n2079
  );


  xor
  g2233
  (
    n2159,
    n1868,
    n2044,
    n1931,
    n1987
  );


  or
  g2234
  (
    n2199,
    n2033,
    n2008,
    n1877,
    n1953
  );


  nor
  g2235
  (
    n2277,
    n1878,
    n1955,
    n1893,
    n2054
  );


  and
  g2236
  (
    n2397,
    n2107,
    n1883,
    n2080,
    n1898
  );


  or
  g2237
  (
    n2282,
    n1890,
    n1887,
    n1953,
    n2091
  );


  or
  g2238
  (
    n2201,
    n1962,
    n1893,
    n1920,
    n2042
  );


  xnor
  g2239
  (
    n2294,
    n1913,
    n1983,
    n2006,
    n1924
  );


  xor
  g2240
  (
    n2280,
    n1935,
    n2033,
    n1905,
    n1922
  );


  xor
  g2241
  (
    n2415,
    n1908,
    n2035,
    n2001,
    n2052
  );


  nor
  g2242
  (
    n2203,
    n1948,
    n2068,
    n2055,
    n1900
  );


  and
  g2243
  (
    n2136,
    n2090,
    n1921,
    n2037,
    n1988
  );


  xnor
  g2244
  (
    n2371,
    n2078,
    n2028,
    n1895,
    n2069
  );


  xnor
  g2245
  (
    n2316,
    n1916,
    n1894,
    n1910,
    n2055
  );


  nor
  g2246
  (
    n2183,
    n1883,
    n2018,
    n2073,
    n2082
  );


  xor
  g2247
  (
    n2221,
    n1997,
    n2096,
    n2001,
    n2027
  );


  nor
  g2248
  (
    n2308,
    n2051,
    n2049,
    n1886,
    n2023
  );


  nand
  g2249
  (
    n2412,
    n1872,
    n2040,
    n1869,
    n2091
  );


  nand
  g2250
  (
    n2317,
    n2064,
    n1982,
    n2105,
    n2004
  );


  nand
  g2251
  (
    n2164,
    n1911,
    n1961,
    n1924,
    n2043
  );


  or
  g2252
  (
    n2399,
    n2000,
    n1981,
    n2083,
    n1938
  );


  nand
  g2253
  (
    n2131,
    n2101,
    n2057,
    n2010,
    n2015
  );


  xor
  g2254
  (
    n2232,
    n2052,
    n1869,
    n2000,
    n1906
  );


  nand
  g2255
  (
    n2138,
    n1917,
    n1873,
    n1897,
    n1903
  );


  and
  g2256
  (
    n2293,
    n1879,
    n1965,
    n2050,
    n1994
  );


  xnor
  g2257
  (
    n2285,
    n2022,
    n1994,
    n2017,
    n1967
  );


  and
  g2258
  (
    n2149,
    n2075,
    n1871,
    n1892,
    n2070
  );


  and
  g2259
  (
    KeyWire_0_62,
    n1943,
    n2049,
    n1983,
    n2105
  );


  nand
  g2260
  (
    n2207,
    n1897,
    n1925,
    n1991,
    n1944
  );


  and
  g2261
  (
    n2130,
    n2053,
    n1979,
    n1944,
    n2079
  );


  xnor
  g2262
  (
    n2228,
    n2047,
    n1928,
    n1907,
    n1920
  );


  nand
  g2263
  (
    n2261,
    n2027,
    n1933,
    n2077,
    n2072
  );


  nor
  g2264
  (
    n2189,
    n2037,
    n2071,
    n2012,
    n1938
  );


  xnor
  g2265
  (
    n2140,
    n2106,
    n1969,
    n2021
  );


  xnor
  g2266
  (
    n2222,
    n1945,
    n1875,
    n2007
  );


  nand
  g2267
  (
    KeyWire_0_3,
    n2053,
    n2066,
    n1992,
    n2022
  );


  nand
  g2268
  (
    n2120,
    n2001,
    n2018,
    n1892,
    n1978
  );


  xor
  g2269
  (
    n2172,
    n1986,
    n1971,
    n1901,
    n1929
  );


  and
  g2270
  (
    n2360,
    n2060,
    n1919,
    n2104,
    n2081
  );


  nand
  g2271
  (
    n2200,
    n1881,
    n1904,
    n1978,
    n2096
  );


  xor
  g2272
  (
    n2364,
    n2060,
    n1923,
    n1972,
    n1912
  );


  nor
  g2273
  (
    n2368,
    n2009,
    n2038,
    n2083,
    n2061
  );


  nand
  g2274
  (
    n2331,
    n1985,
    n1878,
    n1930,
    n1904
  );


  or
  g2275
  (
    n2110,
    n1892,
    n1936,
    n2050,
    n1980
  );


  and
  g2276
  (
    n2170,
    n2051,
    n1872,
    n1974,
    n1935
  );


  or
  g2277
  (
    n2376,
    n1993,
    n2068,
    n2026,
    n1917
  );


  xor
  g2278
  (
    n2155,
    n1992,
    n1965,
    n1997,
    n1990
  );


  and
  g2279
  (
    n2142,
    n1902,
    n1968,
    n2066,
    n2087
  );


  xnor
  g2280
  (
    n2377,
    n2011,
    n2092,
    n2093,
    n1954
  );


  nor
  g2281
  (
    n2336,
    n1899,
    n2090,
    n1999,
    n1934
  );


  nand
  g2282
  (
    n2161,
    n1970,
    n1989,
    n1990,
    n1941
  );


  xor
  g2283
  (
    n2409,
    n2005,
    n2087,
    n1873,
    n1944
  );


  or
  g2284
  (
    n2257,
    n2006,
    n1903,
    n2092,
    n2088
  );


  xnor
  g2285
  (
    n2178,
    n1879,
    n1959,
    n2040,
    n2036
  );


  and
  g2286
  (
    n2174,
    n2097,
    n2047,
    n1898,
    n1905
  );


  and
  g2287
  (
    n2416,
    n2047,
    n2037,
    n1925,
    n2059
  );


  or
  g2288
  (
    n2216,
    n2035,
    n2023,
    n1967,
    n1943
  );


  xor
  g2289
  (
    n2173,
    n2048,
    n1935,
    n1960,
    n1990
  );


  and
  g2290
  (
    n2241,
    n2054,
    n2033,
    n2079,
    n1949
  );


  nand
  g2291
  (
    n2327,
    n1998,
    n2059,
    n2045,
    n2100
  );


  nor
  g2292
  (
    n2314,
    n2022,
    n2045,
    n2090,
    n1962
  );


  and
  g2293
  (
    n2281,
    n1927,
    n1870,
    n1898,
    n1981
  );


  xnor
  g2294
  (
    n2160,
    n2053,
    n2028,
    n2066,
    n2058
  );


  xor
  g2295
  (
    n2151,
    n1977,
    n1885,
    n1924,
    n1884
  );


  nand
  g2296
  (
    n2252,
    n1891,
    n1962,
    n1933,
    n1889
  );


  xnor
  g2297
  (
    n2337,
    n2071,
    n2081,
    n2062,
    n1928
  );


  nand
  g2298
  (
    n2343,
    n1989,
    n1957,
    n2071,
    n2086
  );


  xor
  g2299
  (
    n2202,
    n1940,
    n2062,
    n2014,
    n2046
  );


  nand
  g2300
  (
    n2127,
    n2016,
    n1890,
    n1942,
    n2032
  );


  xnor
  g2301
  (
    n2290,
    n1996,
    n2072,
    n1956,
    n1888
  );


  nor
  g2302
  (
    n2394,
    n2016,
    n1922,
    n2063,
    n1887
  );


  nor
  g2303
  (
    n2351,
    n2070,
    n2019,
    n2047,
    n2058
  );


  xnor
  g2304
  (
    n2212,
    n1871,
    n1908,
    n2081,
    n1926
  );


  xor
  g2305
  (
    n2322,
    n1911,
    n2036,
    n1932,
    n2041
  );


  xnor
  g2306
  (
    n2209,
    n1947,
    n2075,
    n1915,
    n2093
  );


  nor
  g2307
  (
    n2288,
    n2028,
    n2014,
    n2001,
    n1961
  );


  xor
  g2308
  (
    n2361,
    n2040,
    n2077,
    n1929,
    n1937
  );


  or
  g2309
  (
    n2220,
    n2065,
    n2017,
    n2058,
    n2049
  );


  nand
  g2310
  (
    n2278,
    n1993,
    n1999,
    n2049,
    n1890
  );


  xnor
  g2311
  (
    n2411,
    n1945,
    n2059,
    n2105,
    n1888
  );


  xor
  g2312
  (
    n2338,
    n1992,
    n2065,
    n1884,
    n2009
  );


  nor
  g2313
  (
    n2311,
    n1952,
    n2089,
    n1907,
    n1971
  );


  or
  g2314
  (
    n2366,
    n1950,
    n2003,
    n1963,
    n1985
  );


  xnor
  g2315
  (
    n2154,
    n2102,
    n2065,
    n2023,
    n2046
  );


  nand
  g2316
  (
    n2180,
    n2057,
    n2036,
    n2090,
    n1916
  );


  and
  g2317
  (
    n2323,
    n2008,
    n2099,
    n1987
  );


  or
  g2318
  (
    n2190,
    n2074,
    n2105,
    n1910,
    n1997
  );


  xnor
  g2319
  (
    n2152,
    n2025,
    n1937,
    n1966,
    n2010
  );


  and
  g2320
  (
    n2410,
    n1878,
    n1910,
    n2050,
    n2082
  );


  xor
  g2321
  (
    KeyWire_0_57,
    n1951,
    n2004,
    n1961,
    n2063
  );


  and
  g2322
  (
    KeyWire_0_14,
    n2085,
    n2020,
    n1956,
    n1985
  );


  or
  g2323
  (
    n2235,
    n1876,
    n1925,
    n2055,
    n2099
  );


  nor
  g2324
  (
    n2333,
    n1942,
    n2102,
    n1900,
    n2056
  );


  xor
  g2325
  (
    n2403,
    n2015,
    n1967,
    n1912,
    n2014
  );


  nor
  g2326
  (
    n2248,
    n1913,
    n2000,
    n2108,
    n1911
  );


  nand
  g2327
  (
    n2123,
    n1882,
    n2069,
    n1956,
    n1996
  );


  or
  g2328
  (
    n2242,
    n1940,
    n1941,
    n2043,
    n2069
  );


  and
  g2329
  (
    n2296,
    n1876,
    n2029,
    n1902,
    n2074
  );


  xnor
  g2330
  (
    n2384,
    n1899,
    n1923,
    n1991,
    n2027
  );


  or
  g2331
  (
    n2350,
    n2076,
    n1987,
    n1979,
    n1889
  );


  and
  g2332
  (
    n2196,
    n2039,
    n2103,
    n2022,
    n2069
  );


  and
  g2333
  (
    n2205,
    n1869,
    n1947,
    n2031,
    n2097
  );


  or
  g2334
  (
    n2383,
    n2032,
    n2030,
    n2015,
    n1986
  );


  xnor
  g2335
  (
    n2318,
    n1887,
    n2005,
    n2072,
    n1983
  );


  and
  g2336
  (
    n2231,
    n1896,
    n1937,
    n1877,
    n1968
  );


  nand
  g2337
  (
    n2141,
    n1888,
    n1950,
    n2056,
    n1953
  );


  xnor
  g2338
  (
    KeyWire_0_4,
    n2011,
    n2032,
    n2064,
    n1985
  );


  nor
  g2339
  (
    n2312,
    n1875,
    n2048,
    n1973,
    n1868
  );


  and
  g2340
  (
    n2378,
    n1895,
    n2063,
    n1885,
    n2045
  );


  nor
  g2341
  (
    n2236,
    n2041,
    n1955,
    n1939,
    n1964
  );


  and
  g2342
  (
    n2335,
    n1867,
    n1984,
    n2035,
    n1992
  );


  nand
  g2343
  (
    n2289,
    n2076,
    n2041,
    n2051,
    n2046
  );


  and
  g2344
  (
    n2176,
    n2077,
    n1976,
    n2100,
    n1880
  );


  or
  g2345
  (
    n2144,
    n2091,
    n2005,
    n1998,
    n2057
  );


  nand
  g2346
  (
    n2276,
    n1995,
    n1900,
    n2080,
    n1915
  );


  or
  g2347
  (
    n2150,
    n2024,
    n2056,
    n2003,
    n1939
  );


  or
  g2348
  (
    n2116,
    n2041,
    n2073,
    n1960,
    n2070
  );


  nand
  g2349
  (
    n2111,
    n2017,
    n1984,
    n1976,
    n1948
  );


  xor
  g2350
  (
    n2166,
    n2043,
    n2014,
    n2089,
    n2013
  );


  nand
  g2351
  (
    n2341,
    n2082,
    n2061,
    n2048,
    n1885
  );


  xor
  g2352
  (
    n2283,
    n1914,
    n2064,
    n2072,
    n2020
  );


  nand
  g2353
  (
    n2265,
    n2032,
    n2038,
    n1988,
    n1880
  );


  xnor
  g2354
  (
    n2339,
    n1982,
    n2048,
    n1939,
    n1974
  );


  xor
  g2355
  (
    n2363,
    n2021,
    n1908,
    n1983,
    n1951
  );


  and
  g2356
  (
    n2401,
    n2086,
    n1886,
    n877,
    n2080
  );


  xnor
  g2357
  (
    n2126,
    n1913,
    n2028,
    n2067,
    n2021
  );


  and
  g2358
  (
    n2215,
    n1989,
    n1964,
    n1931,
    n1914
  );


  nor
  g2359
  (
    n2168,
    n2034,
    n2006,
    n2094
  );


  nor
  g2360
  (
    n2213,
    n2004,
    n1952,
    n1909,
    n1958
  );


  and
  g2361
  (
    n2357,
    n2012,
    n1881,
    n2016,
    n2064
  );


  xnor
  g2362
  (
    n2133,
    n2068,
    n1906,
    n2025,
    n2039
  );


  xnor
  g2363
  (
    n2122,
    n2023,
    n2088,
    n1889,
    n2066
  );


  or
  g2364
  (
    n2148,
    n1989,
    n2097,
    n2088,
    n2096
  );


  xor
  g2365
  (
    n2121,
    n1882,
    n1894,
    n1946,
    n2054
  );


  or
  g2366
  (
    n2310,
    n1930,
    n2031,
    n1999,
    n1955
  );


  xnor
  g2367
  (
    n2297,
    n2017,
    n1993,
    n2040,
    n1907
  );


  or
  g2368
  (
    n2315,
    n2002,
    n2106,
    n1963,
    n1918
  );


  nand
  g2369
  (
    n2195,
    n1946,
    n1909,
    n2078,
    n2084
  );


  xnor
  g2370
  (
    n2175,
    n2089,
    n2100,
    n1950,
    n2050
  );


  and
  g2371
  (
    n2319,
    n2039,
    n2084,
    n1904
  );


  or
  g2372
  (
    n2260,
    n2045,
    n2095,
    n1874,
    n2035
  );


  nand
  g2373
  (
    n2329,
    n1870,
    n2095,
    n2100,
    n1886
  );


  xor
  g2374
  (
    n2128,
    n1976,
    n1970,
    n1975,
    n2070
  );


  nand
  g2375
  (
    n2396,
    n2013,
    n2096,
    n2075,
    n2068
  );


  nand
  g2376
  (
    n2229,
    n1926,
    n1901,
    n2067,
    n2026
  );


  or
  g2377
  (
    n2347,
    n2101,
    n1941,
    n1954,
    n2060
  );


  or
  g2378
  (
    n2380,
    n2061,
    n2053,
    n1919,
    n2029
  );


  and
  g2379
  (
    n2146,
    n2085,
    n2058,
    n2087,
    n1977
  );


  and
  g2380
  (
    n2225,
    n1949,
    n2060,
    n2010,
    n2012
  );


  nand
  g2381
  (
    n2259,
    n1980,
    n1995,
    n2089,
    n1996
  );


  nor
  g2382
  (
    n2355,
    n2013,
    n2025,
    n2062,
    n1876
  );


  or
  g2383
  (
    n2356,
    n1978,
    n1915,
    n1957,
    n2108
  );


  xor
  g2384
  (
    n2611,
    n2154,
    n2290,
    n2210,
    n2216
  );


  xor
  g2385
  (
    n2585,
    n2126,
    n2344,
    n2132,
    n2284
  );


  xnor
  g2386
  (
    n2558,
    n2273,
    n2173,
    n2348,
    n2329
  );


  xor
  g2387
  (
    n2503,
    n2358,
    n2134,
    n2391,
    n1105
  );


  xnor
  g2388
  (
    n2653,
    n2155,
    n2240,
    n2254,
    n2413
  );


  and
  g2389
  (
    n2533,
    n2179,
    n2414,
    n2333,
    n2379
  );


  nor
  g2390
  (
    n2587,
    n2137,
    n2376,
    n2208,
    n2144
  );


  or
  g2391
  (
    n2651,
    n2298,
    n2411,
    n2128,
    n2402
  );


  xnor
  g2392
  (
    n2594,
    n2331,
    n2123,
    n2176,
    n2203
  );


  xnor
  g2393
  (
    n2449,
    n2127,
    n2394,
    n2322,
    n2403
  );


  or
  g2394
  (
    n2457,
    n2185,
    n2337,
    n2339,
    n2147
  );


  xnor
  g2395
  (
    n2561,
    n2225,
    n2175,
    n2113,
    n2223
  );


  and
  g2396
  (
    n2646,
    n2269,
    n2287,
    n2237,
    n2151
  );


  and
  g2397
  (
    n2513,
    n2316,
    n2264,
    n2374,
    n2158
  );


  xor
  g2398
  (
    n2479,
    n2252,
    n2253,
    n1386,
    n2371
  );


  xnor
  g2399
  (
    n2566,
    n2373,
    n2352,
    n2257,
    n2185
  );


  or
  g2400
  (
    n2429,
    n2382,
    n2148,
    n2120,
    n2256
  );


  or
  g2401
  (
    n2491,
    n2412,
    n2333,
    n2264,
    n2287
  );


  or
  g2402
  (
    n2575,
    n2343,
    n2304,
    n2138,
    n2158
  );


  and
  g2403
  (
    n2545,
    n2182,
    n2301,
    n2201,
    n2202
  );


  and
  g2404
  (
    n2649,
    n2128,
    n2158,
    n2127,
    n2320
  );


  nand
  g2405
  (
    n2450,
    n2117,
    n2136,
    n2238,
    n2389
  );


  nor
  g2406
  (
    n2514,
    n2186,
    n2266,
    n2349,
    n2408
  );


  nand
  g2407
  (
    n2422,
    n2171,
    n2244,
    n2250,
    n2309
  );


  or
  g2408
  (
    n2462,
    n2365,
    n2184,
    n2375,
    n2130
  );


  and
  g2409
  (
    n2528,
    n2320,
    n2332,
    n2347,
    n2266
  );


  or
  g2410
  (
    n2542,
    n2217,
    n2144,
    n2197,
    n2319
  );


  nand
  g2411
  (
    n2441,
    n2366,
    n2404,
    n2119,
    n2416
  );


  nor
  g2412
  (
    n2600,
    n2261,
    n2245,
    n2192,
    n2142
  );


  nor
  g2413
  (
    n2625,
    n2412,
    n2396,
    n2130,
    n2305
  );


  and
  g2414
  (
    n2492,
    n2312,
    n2160,
    n2192,
    n2336
  );


  or
  g2415
  (
    KeyWire_0_10,
    n2111,
    n2135,
    n2362,
    n2244
  );


  and
  g2416
  (
    n2568,
    n2399,
    n2368,
    n2365,
    n2194
  );


  nor
  g2417
  (
    n2552,
    n2380,
    n2156,
    n2357,
    n2214
  );


  and
  g2418
  (
    n2421,
    n2157,
    n2390,
    n2264,
    n2271
  );


  and
  g2419
  (
    n2632,
    n2290,
    n2349,
    n2191,
    n2122
  );


  nor
  g2420
  (
    n2650,
    n2411,
    n2315,
    n2366,
    n2140
  );


  nand
  g2421
  (
    n2475,
    n2327,
    n2202,
    n2218,
    n2392
  );


  xnor
  g2422
  (
    n2487,
    n2236,
    n2384,
    n2169,
    n2111
  );


  xnor
  g2423
  (
    n2430,
    n2387,
    n2347,
    n2413,
    n2126
  );


  xor
  g2424
  (
    n2631,
    n2390,
    n2379,
    n2397,
    n2255
  );


  xor
  g2425
  (
    n2486,
    n2268,
    n2274,
    n2284,
    n2350
  );


  xor
  g2426
  (
    n2620,
    n2329,
    n2278,
    n2201,
    n2272
  );


  xor
  g2427
  (
    KeyWire_0_42,
    n2112,
    n2230,
    n2267,
    n2332
  );


  nand
  g2428
  (
    n2589,
    n2407,
    n2281,
    n2141,
    n2412
  );


  xnor
  g2429
  (
    n2652,
    n2298,
    n2112,
    n2196,
    n2192
  );


  and
  g2430
  (
    n2613,
    n2321,
    n2115,
    n2223,
    n2409
  );


  xor
  g2431
  (
    n2621,
    n2213,
    n2223,
    n2169,
    n2398
  );


  or
  g2432
  (
    n2565,
    n2136,
    n2193,
    n2119,
    n2231
  );


  and
  g2433
  (
    n2628,
    n2196,
    n2165,
    n2255,
    n1104
  );


  and
  g2434
  (
    n2523,
    n2109,
    n2393,
    n2211,
    n2132
  );


  nand
  g2435
  (
    n2446,
    n2362,
    n2374,
    n2346,
    n2285
  );


  nand
  g2436
  (
    n2493,
    n2220,
    n2371,
    n2168,
    n2219
  );


  xor
  g2437
  (
    n2559,
    n2235,
    n2321,
    n2139,
    n2127
  );


  and
  g2438
  (
    n2629,
    n2163,
    n2355,
    n2178,
    n2133
  );


  nand
  g2439
  (
    n2444,
    n2287,
    n2265,
    n2299,
    n2391
  );


  nand
  g2440
  (
    n2543,
    n2351,
    n2241,
    n2313,
    n2328
  );


  or
  g2441
  (
    KeyWire_0_48,
    n2213,
    n2332,
    n2384,
    n2161
  );


  or
  g2442
  (
    n2435,
    n2164,
    n2386,
    n2278,
    n2275
  );


  xor
  g2443
  (
    n2602,
    n2126,
    n2212,
    n2367,
    n2228
  );


  and
  g2444
  (
    n2517,
    n2166,
    n2327,
    n2128,
    n2333
  );


  and
  g2445
  (
    n2541,
    n2258,
    n2338,
    n2115,
    n2260
  );


  nor
  g2446
  (
    n2531,
    n2293,
    n2359,
    n2306,
    n2340
  );


  and
  g2447
  (
    n2638,
    n2315,
    n2171,
    n2221,
    n2385
  );


  and
  g2448
  (
    KeyWire_0_16,
    n2400,
    n2131,
    n2293,
    n2309
  );


  and
  g2449
  (
    n2480,
    n2312,
    n2372,
    n2216,
    n2401
  );


  xnor
  g2450
  (
    n2630,
    n2240,
    n2328,
    n2199,
    n2265
  );


  nor
  g2451
  (
    n2560,
    n2222,
    n2315,
    n2250,
    n2259
  );


  or
  g2452
  (
    n2572,
    n2204,
    n2276,
    n2415,
    n2296
  );


  nand
  g2453
  (
    n2471,
    n2378,
    n2165,
    n2245,
    n2186
  );


  nand
  g2454
  (
    n2511,
    n2370,
    n2261,
    n2336,
    n2341
  );


  xor
  g2455
  (
    n2529,
    n2251,
    n2300,
    n2121,
    n2233
  );


  nand
  g2456
  (
    n2463,
    n2387,
    n2187,
    n2380,
    n2398
  );


  nor
  g2457
  (
    n2496,
    n2183,
    n2255,
    n2134,
    n2179
  );


  xor
  g2458
  (
    n2526,
    n2367,
    n2343,
    n2405,
    n2298
  );


  nor
  g2459
  (
    n2508,
    n2207,
    n2291,
    n2364,
    n2166
  );


  xnor
  g2460
  (
    n2488,
    n2180,
    n2289,
    n2195,
    n2279
  );


  and
  g2461
  (
    n2522,
    n2323,
    n2270,
    n2256,
    n2375
  );


  nand
  g2462
  (
    n2481,
    n2248,
    n2218,
    n2361,
    n2121
  );


  or
  g2463
  (
    n2527,
    n2278,
    n2206,
    n2221,
    n2294
  );


  and
  g2464
  (
    n2469,
    n2235,
    n2243,
    n2224,
    n2403
  );


  nor
  g2465
  (
    n2419,
    n2109,
    n2268,
    n2227,
    n2161
  );


  nor
  g2466
  (
    n2642,
    n2373,
    n2335,
    n2170,
    n2325
  );


  nor
  g2467
  (
    n2490,
    n2364,
    n2175,
    n2116,
    n2256
  );


  or
  g2468
  (
    n2442,
    n2351,
    n2124,
    n2247,
    n2386
  );


  xor
  g2469
  (
    n2618,
    n2227,
    n2182,
    n2409,
    n2391
  );


  nand
  g2470
  (
    n2549,
    n1386,
    n1385,
    n2311,
    n2370
  );


  or
  g2471
  (
    n2622,
    n2376,
    n2288,
    n2335,
    n2414
  );


  nand
  g2472
  (
    n2591,
    n2334,
    n2407,
    n2259,
    n2410
  );


  xor
  g2473
  (
    n2505,
    n2187,
    n2234,
    n2310,
    n2153
  );


  and
  g2474
  (
    n2612,
    n2195,
    n2242,
    n2198,
    n2217
  );


  xor
  g2475
  (
    n2518,
    n2152,
    n2361,
    n2177,
    n1386
  );


  or
  g2476
  (
    n2609,
    n2174,
    n2354,
    n2173,
    n2337
  );


  xnor
  g2477
  (
    n2601,
    n2379,
    n2197,
    n2388,
    n2303
  );


  xor
  g2478
  (
    n2473,
    n2129,
    n2188,
    n2143,
    n2364
  );


  xnor
  g2479
  (
    n2617,
    n2110,
    n2204,
    n2399,
    n2108
  );


  xnor
  g2480
  (
    n2521,
    n2236,
    n2363,
    n2157,
    n2208
  );


  xnor
  g2481
  (
    n2548,
    n2249,
    n2169,
    n2201,
    n2297
  );


  xor
  g2482
  (
    n2593,
    n2308,
    n2150,
    n2358,
    n2125
  );


  and
  g2483
  (
    n2453,
    n2398,
    n2316,
    n2221,
    n2143
  );


  and
  g2484
  (
    n2616,
    n2263,
    n2261,
    n2190,
    n2311
  );


  and
  g2485
  (
    n2418,
    n2330,
    n2150,
    n2402,
    n2342
  );


  or
  g2486
  (
    n2467,
    n2132,
    n2176,
    n2131,
    n2311
  );


  and
  g2487
  (
    n2468,
    n1104,
    n2205,
    n2178,
    n2356
  );


  or
  g2488
  (
    n2530,
    n2343,
    n2388,
    n2284,
    n2167
  );


  nor
  g2489
  (
    n2626,
    n2194,
    n2149,
    n2231,
    n2406
  );


  and
  g2490
  (
    n2489,
    n2281,
    n2151,
    n2129,
    n2395
  );


  xnor
  g2491
  (
    n2645,
    n2288,
    n2377,
    n2215,
    n2415
  );


  xor
  g2492
  (
    n2627,
    n2229,
    n2123,
    n1387,
    n2154
  );


  nand
  g2493
  (
    n2485,
    n2213,
    n2395,
    n2297,
    n2335
  );


  xnor
  g2494
  (
    n2569,
    n2205,
    n2153,
    n2330,
    n2408
  );


  or
  g2495
  (
    n2427,
    n2405,
    n2312,
    n2236,
    n1105
  );


  xnor
  g2496
  (
    n2448,
    n2325,
    n2167,
    n2302,
    n2331
  );


  or
  g2497
  (
    n2573,
    n2308,
    n2318,
    n2303,
    n2134
  );


  and
  g2498
  (
    n2581,
    n2345,
    n2152,
    n2283,
    n2207
  );


  and
  g2499
  (
    n2445,
    n2193,
    n2217,
    n2366,
    n2124
  );


  xor
  g2500
  (
    n2554,
    n2147,
    n2291,
    n2290,
    n2348
  );


  and
  g2501
  (
    n2556,
    n2322,
    n2340,
    n2145,
    n2176
  );


  nor
  g2502
  (
    n2464,
    n2237,
    n2414,
    n2356,
    n2232
  );


  nand
  g2503
  (
    n2562,
    n2413,
    n2214,
    n2262,
    n2318
  );


  xnor
  g2504
  (
    n2440,
    n2282,
    n2212,
    n2377,
    n2156
  );


  xor
  g2505
  (
    n2472,
    n2193,
    n2209,
    n2226,
    n2224
  );


  nand
  g2506
  (
    n2637,
    n2359,
    n2286,
    n2397,
    n2190
  );


  nor
  g2507
  (
    n2494,
    n2317,
    n2135,
    n1103,
    n2305
  );


  nand
  g2508
  (
    n2417,
    n2273,
    n2163,
    n2353,
    n2283
  );


  xor
  g2509
  (
    n2546,
    n2275,
    n2403,
    n2310,
    n2179
  );


  nor
  g2510
  (
    n2466,
    n2337,
    n2244,
    n2276,
    n2327
  );


  or
  g2511
  (
    n2534,
    n2381,
    n2344,
    n2365,
    n2165
  );


  or
  g2512
  (
    n2431,
    n2232,
    n2160,
    n2313,
    n2383
  );


  xnor
  g2513
  (
    n2470,
    n2401,
    n2295,
    n2307
  );


  nor
  g2514
  (
    n2595,
    n2410,
    n2189,
    n2339,
    n2280
  );


  or
  g2515
  (
    n2443,
    n2188,
    n2342,
    n2299,
    n2114
  );


  and
  g2516
  (
    n2578,
    n2378,
    n2168,
    n2184
  );


  xnor
  g2517
  (
    KeyWire_0_45,
    n2242,
    n2174,
    n2263,
    n2209
  );


  nor
  g2518
  (
    n2461,
    n2353,
    n2140,
    n1388,
    n2159
  );


  nand
  g2519
  (
    n2577,
    n2356,
    n2385,
    n2400,
    n2293
  );


  nand
  g2520
  (
    n2648,
    n2156,
    n2245,
    n2243,
    n2125
  );


  xnor
  g2521
  (
    n2557,
    n2381,
    n2357,
    n2250,
    n2406
  );


  xnor
  g2522
  (
    n2512,
    n2416,
    n2348,
    n2406,
    n2374
  );


  and
  g2523
  (
    n2623,
    n2140,
    n2282,
    n2136,
    n2279
  );


  nand
  g2524
  (
    n2465,
    n2392,
    n2225,
    n2265,
    n2108
  );


  xnor
  g2525
  (
    n2619,
    n2323,
    n2247,
    n2177,
    n2117
  );


  xnor
  g2526
  (
    n2586,
    n2144,
    n2411,
    n2294,
    n2277
  );


  nor
  g2527
  (
    n2570,
    n2342,
    n2252,
    n2302,
    n2188
  );


  nor
  g2528
  (
    n2606,
    n2393,
    n2355,
    n2345,
    n2206
  );


  nor
  g2529
  (
    n2439,
    n2248,
    n2190,
    n2229,
    n2404
  );


  nor
  g2530
  (
    n2598,
    n2185,
    n2164,
    n2272
  );


  nand
  g2531
  (
    n2634,
    n2191,
    n2141,
    n2274,
    n1102
  );


  nand
  g2532
  (
    n2588,
    n1104,
    n2334,
    n2155,
    n2353
  );


  xnor
  g2533
  (
    n2608,
    n2328,
    n2294,
    n2234,
    n2295
  );


  nand
  g2534
  (
    n2555,
    n2203,
    n2113,
    n2369,
    n2320
  );


  nor
  g2535
  (
    n2495,
    n2317,
    n2142,
    n2314,
    n2172
  );


  nand
  g2536
  (
    n2456,
    n2322,
    n2393,
    n2375,
    n2113
  );


  xor
  g2537
  (
    n2540,
    n2220,
    n2203,
    n2394,
    n2211
  );


  and
  g2538
  (
    n2455,
    n2181,
    n2277,
    n2180,
    n2253
  );


  nand
  g2539
  (
    n2624,
    n2402,
    n2280,
    n2116,
    n2198
  );


  and
  g2540
  (
    n2420,
    n2239,
    n2161,
    n2381,
    n2334
  );


  nand
  g2541
  (
    n2550,
    n2214,
    n2292,
    n1105,
    n2263
  );


  nand
  g2542
  (
    n2563,
    n2368,
    n2257,
    n2117,
    n2258
  );


  or
  g2543
  (
    n2576,
    n2230,
    n2267,
    n2272,
    n2247
  );


  and
  g2544
  (
    n2454,
    n2347,
    n2262,
    n2329,
    n2225
  );


  and
  g2545
  (
    n2516,
    n2219,
    n2210,
    n2246,
    n2331
  );


  nand
  g2546
  (
    n2483,
    n2326,
    n2149,
    n2345,
    n2385
  );


  xnor
  g2547
  (
    n2477,
    n2145,
    n2310,
    n2363,
    n2241
  );


  xor
  g2548
  (
    n2567,
    n2326,
    n2125,
    n2350,
    n2276
  );


  and
  g2549
  (
    n2423,
    n2195,
    n2330,
    n2415,
    n2196
  );


  xnor
  g2550
  (
    n2596,
    n2233,
    n2238,
    n2362,
    n2119
  );


  xnor
  g2551
  (
    n2520,
    n2355,
    n2110,
    n2338,
    n2215
  );


  or
  g2552
  (
    n2428,
    n2316,
    n2162,
    n2336,
    n2352
  );


  or
  g2553
  (
    KeyWire_0_5,
    n2409,
    n2118,
    n2183,
    n2154
  );


  nor
  g2554
  (
    n2532,
    n2218,
    n2383,
    n2254,
    n2153
  );


  or
  g2555
  (
    n2424,
    n2116,
    n2360,
    n1388,
    n2178
  );


  nand
  g2556
  (
    n2551,
    n2239,
    n2286,
    n2271,
    n2172
  );


  nand
  g2557
  (
    n2426,
    n2324,
    n2240,
    n2291,
    n2304
  );


  xnor
  g2558
  (
    n2547,
    n2254,
    n2155,
    n2200,
    n2368
  );


  xnor
  g2559
  (
    n2499,
    n2271,
    n2242,
    n2226,
    n2286
  );


  nand
  g2560
  (
    n2639,
    n2202,
    n2397,
    n2166,
    n2249
  );


  or
  g2561
  (
    n2509,
    n2267,
    n2159,
    n2118,
    n2371
  );


  and
  g2562
  (
    n2537,
    n2387,
    n2248,
    n2341,
    n2246
  );


  nor
  g2563
  (
    n2519,
    n2187,
    n2299,
    n2222,
    n2260
  );


  xnor
  g2564
  (
    n2610,
    n2243,
    n2401,
    n2360,
    n2131
  );


  xor
  g2565
  (
    n2647,
    n2354,
    n2112,
    n2139,
    n2177
  );


  xor
  g2566
  (
    n2536,
    n2377,
    n2210,
    n2157,
    n1385
  );


  nor
  g2567
  (
    n2535,
    n2160,
    n2122,
    n2110,
    n2251
  );


  and
  g2568
  (
    n2425,
    n2146,
    n2209,
    n2361,
    n2162
  );


  or
  g2569
  (
    n2476,
    n2258,
    n2124,
    n2349,
    n2259
  );


  nor
  g2570
  (
    n2438,
    n2138,
    n2319,
    n2307,
    n2249
  );


  nor
  g2571
  (
    n2460,
    n2172,
    n2212,
    n2369,
    n2289
  );


  or
  g2572
  (
    n2592,
    n2163,
    n2292,
    n2302,
    n2319
  );


  xnor
  g2573
  (
    n2564,
    n2118,
    n2251,
    n2301,
    n2123
  );


  xnor
  g2574
  (
    n2615,
    n2350,
    n2229,
    n2208,
    n1103
  );


  nand
  g2575
  (
    n2539,
    n2200,
    n2235,
    n2389,
    n2300
  );


  nor
  g2576
  (
    n2544,
    n2142,
    n2167,
    n2133,
    n2121
  );


  nand
  g2577
  (
    n2599,
    n2392,
    n2231,
    n2346,
    n2183
  );


  or
  g2578
  (
    n2590,
    n2238,
    n2180,
    n2308,
    n2386
  );


  nor
  g2579
  (
    n2583,
    n2115,
    n2273,
    n2400,
    n2146
  );


  nor
  g2580
  (
    n2641,
    n2309,
    n2388,
    n2219,
    n2120
  );


  nor
  g2581
  (
    n2644,
    n2344,
    n2300,
    n2162,
    n2232
  );


  or
  g2582
  (
    n2574,
    n2341,
    n2318,
    n2304,
    n2150
  );


  xor
  g2583
  (
    n2515,
    n2314,
    n2141,
    n2186,
    n2230
  );


  xnor
  g2584
  (
    n2607,
    n2369,
    n2148,
    n2285,
    n2292
  );


  nand
  g2585
  (
    n2497,
    n2222,
    n2111,
    n2227,
    n2171
  );


  or
  g2586
  (
    n2474,
    n2354,
    n2181,
    n2226,
    n1387
  );


  nor
  g2587
  (
    n2614,
    n2410,
    n2396,
    n2352,
    n2296
  );


  or
  g2588
  (
    n2571,
    n2280,
    n2376,
    n2270,
    n2224
  );


  nand
  g2589
  (
    n2507,
    n2296,
    n2306,
    n2130,
    n2338
  );


  nand
  g2590
  (
    n2525,
    n2253,
    n2404,
    n2269,
    n2326
  );


  nand
  g2591
  (
    n2604,
    n2215,
    n2216,
    n2198,
    n2137
  );


  and
  g2592
  (
    n2437,
    n2194,
    n2137,
    n2324,
    n2360
  );


  nand
  g2593
  (
    KeyWire_0_13,
    n2372,
    n2138,
    n2262,
    n2396
  );


  xnor
  g2594
  (
    n2579,
    n2149,
    n877,
    n2146,
    n2382
  );


  nand
  g2595
  (
    n2584,
    n2260,
    n2416,
    n2228,
    n2189
  );


  and
  g2596
  (
    n2451,
    n2173,
    n2357,
    n2241,
    n2289
  );


  and
  g2597
  (
    n2501,
    n2148,
    n2313,
    n2317,
    n2339
  );


  xor
  g2598
  (
    n2643,
    n1103,
    n2207,
    n2147,
    n2282
  );


  nor
  g2599
  (
    n2452,
    n2283,
    n2170,
    n2114,
    n2197
  );


  xnor
  g2600
  (
    n2603,
    n2122,
    n2191,
    n2200,
    n2129
  );


  and
  g2601
  (
    n2605,
    n2321,
    n2211,
    n2109,
    n2373
  );


  nor
  g2602
  (
    n2434,
    n2205,
    n2145,
    n2220,
    n2306
  );


  xnor
  g2603
  (
    n2482,
    n2152,
    n2380,
    n2384,
    n2407
  );


  xor
  g2604
  (
    n2484,
    n2257,
    n2297,
    n2275,
    n2204
  );


  nand
  g2605
  (
    n2580,
    n2303,
    n2378,
    n2159,
    n2358
  );


  or
  g2606
  (
    n2506,
    n2266,
    n2199,
    n2109,
    n2395
  );


  nand
  g2607
  (
    n2459,
    n2189,
    n2325,
    n2237,
    n2239
  );


  nand
  g2608
  (
    n2447,
    n2206,
    n2285,
    n2351,
    n2170
  );


  xnor
  g2609
  (
    n2538,
    n2175,
    n2405,
    n2305,
    n2363
  );


  xnor
  g2610
  (
    n2432,
    n2323,
    n2367,
    n2324,
    n2228
  );


  xnor
  g2611
  (
    n2524,
    n2399,
    n2382,
    n2408,
    n2370
  );


  nor
  g2612
  (
    n2478,
    n2279,
    n2277,
    n2135,
    n2174
  );


  xnor
  g2613
  (
    n2633,
    n2114,
    n2184,
    n2383,
    n2301
  );


  and
  g2614
  (
    n2436,
    n2139,
    n2233,
    n2346,
    n2181
  );


  or
  g2615
  (
    n2553,
    n2268,
    n2307,
    n2133,
    n2314
  );


  xor
  g2616
  (
    n2504,
    n2199,
    n2269,
    n2274,
    n2182
  );


  nor
  g2617
  (
    n2582,
    n2246,
    n1387,
    n2281,
    n2359
  );


  nand
  g2618
  (
    n2500,
    n2234,
    n2120,
    n2151,
    n2372
  );


  xor
  g2619
  (
    n2458,
    n2288,
    n2390,
    n2143,
    n2252
  );


  nor
  g2620
  (
    n2636,
    n2270,
    n2389,
    n2340,
    n2394
  );


  xnor
  g2621
  (
    n2676,
    n2484,
    n2599,
    n2649,
    n2623
  );


  or
  g2622
  (
    n2819,
    n2569,
    n879,
    n2494,
    n2602
  );


  nor
  g2623
  (
    n2666,
    n2533,
    n2593,
    n2496,
    n2541
  );


  nand
  g2624
  (
    n2793,
    n2472,
    n2569,
    n2435,
    n2521
  );


  xnor
  g2625
  (
    n2768,
    n2451,
    n2422,
    n2503,
    n2607
  );


  nand
  g2626
  (
    n2717,
    n2556,
    n2441,
    n2609,
    n2429
  );


  or
  g2627
  (
    n2688,
    n2600,
    n2422,
    n2602,
    n2529
  );


  nand
  g2628
  (
    n2689,
    n2622,
    n2423,
    n2638,
    n2630
  );


  xor
  g2629
  (
    n2674,
    n2609,
    n2571,
    n2469,
    n2642
  );


  or
  g2630
  (
    n2828,
    n2520,
    n2610,
    n2464,
    n2629
  );


  nand
  g2631
  (
    n2705,
    n2509,
    n2548,
    n2477,
    n2508
  );


  xor
  g2632
  (
    n2788,
    n2554,
    n2577,
    n2443,
    n2619
  );


  or
  g2633
  (
    n2687,
    n2595,
    n2563,
    n2591,
    n2597
  );


  nor
  g2634
  (
    n2701,
    n2501,
    n2569,
    n2455,
    n2459
  );


  nor
  g2635
  (
    n2781,
    n2466,
    n2417,
    n2496,
    n2575
  );


  xor
  g2636
  (
    n2778,
    n2504,
    n2510,
    n2612,
    n2464
  );


  or
  g2637
  (
    n2714,
    n2526,
    n2571,
    n2480,
    n2550
  );


  nand
  g2638
  (
    n2696,
    n2426,
    n2534,
    n2527,
    n2497
  );


  xor
  g2639
  (
    n2765,
    n2596,
    n2585,
    n2523,
    n2643
  );


  nor
  g2640
  (
    n2779,
    n2424,
    n2430,
    n2576,
    n2490
  );


  xnor
  g2641
  (
    n2709,
    n2458,
    n2448,
    n2534,
    n2419
  );


  xor
  g2642
  (
    n2809,
    n2538,
    n2450,
    n2582,
    n2572
  );


  nand
  g2643
  (
    n2817,
    n2537,
    n2611,
    n2455,
    n2540
  );


  or
  g2644
  (
    n2669,
    n2466,
    n2483,
    n2582,
    n2646
  );


  or
  g2645
  (
    n2762,
    n2531,
    n2500,
    n2424,
    n2623
  );


  nor
  g2646
  (
    n2690,
    n2454,
    n2433,
    n2496,
    n2513
  );


  nor
  g2647
  (
    n2823,
    n2518,
    n2634,
    n2546,
    n2433
  );


  nand
  g2648
  (
    n2710,
    n2425,
    n2613,
    n2488,
    n2560
  );


  nand
  g2649
  (
    n2731,
    n2440,
    n2501,
    n2616,
    n2527
  );


  nand
  g2650
  (
    n2825,
    n2565,
    n878,
    n2443,
    n2625
  );


  nand
  g2651
  (
    n2815,
    n2495,
    n2495,
    n2444,
    n2436
  );


  or
  g2652
  (
    n2749,
    n2429,
    n2593,
    n2468,
    n2618
  );


  nand
  g2653
  (
    n2826,
    n2451,
    n2536,
    n2492,
    n2465
  );


  nor
  g2654
  (
    n2816,
    n2454,
    n2422,
    n2584,
    n2554
  );


  xor
  g2655
  (
    n2777,
    n2603,
    n2461,
    n2449,
    n2428
  );


  nand
  g2656
  (
    n2744,
    n2439,
    n2458,
    n2608,
    n2651
  );


  xnor
  g2657
  (
    n2748,
    n2611,
    n2536,
    n2418,
    n2460
  );


  xor
  g2658
  (
    n2796,
    n2626,
    n2442,
    n2502,
    n2559
  );


  or
  g2659
  (
    n2831,
    n2594,
    n2434,
    n2574,
    n2626
  );


  xnor
  g2660
  (
    n2820,
    n2525,
    n2418,
    n2481,
    n2435
  );


  and
  g2661
  (
    n2798,
    n2651,
    n2545,
    n2549,
    n2625
  );


  xnor
  g2662
  (
    n2775,
    n2462,
    n2644,
    n2519,
    n2619
  );


  nor
  g2663
  (
    n2773,
    n2627,
    n2502,
    n2470,
    n2512
  );


  nand
  g2664
  (
    n2724,
    n2538,
    n2484,
    n2611,
    n2587
  );


  nor
  g2665
  (
    n2771,
    n2617,
    n2592,
    n2475,
    n2565
  );


  nand
  g2666
  (
    n2722,
    n2442,
    n2644,
    n2484,
    n2448
  );


  and
  g2667
  (
    n2716,
    n2438,
    n2648,
    n2554,
    n2612
  );


  xnor
  g2668
  (
    n2675,
    n2433,
    n2531,
    n2487,
    n2478
  );


  nand
  g2669
  (
    n2786,
    n2590,
    n2544,
    n2608,
    n2419
  );


  nor
  g2670
  (
    n2708,
    n2518,
    n2519,
    n2432,
    n2468
  );


  or
  g2671
  (
    n2660,
    n2498,
    n2588,
    n2508,
    n2601
  );


  xor
  g2672
  (
    n2830,
    n2602,
    n2558,
    n878,
    n2560
  );


  xor
  g2673
  (
    n2782,
    n2631,
    n2475,
    n2515,
    n2446
  );


  nand
  g2674
  (
    n2670,
    n2538,
    n2437,
    n2544,
    n2445
  );


  or
  g2675
  (
    n2769,
    n2636,
    n2633,
    n2592,
    n2453
  );


  nand
  g2676
  (
    n2734,
    n2516,
    n2483,
    n2617,
    n2437
  );


  and
  g2677
  (
    n2814,
    n2447,
    n2599,
    n2610,
    n2428
  );


  and
  g2678
  (
    n2752,
    n2530,
    n2638,
    n2583,
    n2462
  );


  nor
  g2679
  (
    n2730,
    n2500,
    n2622,
    n2518,
    n2524
  );


  xor
  g2680
  (
    n2702,
    n2457,
    n2629,
    n2461,
    n2580
  );


  xor
  g2681
  (
    n2797,
    n2417,
    n2628,
    n2506,
    n2607
  );


  and
  g2682
  (
    n2668,
    n2555,
    n2561,
    n2482,
    n2488
  );


  nor
  g2683
  (
    n2715,
    n2509,
    n2551,
    n2543,
    n2615
  );


  and
  g2684
  (
    n2792,
    n2520,
    n2588,
    n2478,
    n2603
  );


  xor
  g2685
  (
    n2754,
    n2568,
    n2577,
    n2623,
    n2512
  );


  and
  g2686
  (
    n2787,
    n2576,
    n2637,
    n2476
  );


  nand
  g2687
  (
    n2805,
    n2463,
    n2649,
    n2515,
    n2479
  );


  xor
  g2688
  (
    n2813,
    n2639,
    n2596,
    n2486,
    n2499
  );


  nor
  g2689
  (
    n2801,
    n2609,
    n2419,
    n2589,
    n1206
  );


  nor
  g2690
  (
    KeyWire_0_59,
    n2434,
    n2441,
    n2552,
    n2444
  );


  xor
  g2691
  (
    n2802,
    n2646,
    n2483,
    n2628,
    n2449
  );


  and
  g2692
  (
    n2758,
    n2452,
    n2566,
    n2501,
    n2469
  );


  nor
  g2693
  (
    n2753,
    n2586,
    n2594,
    n2524,
    n2606
  );


  or
  g2694
  (
    n2811,
    n2567,
    n2539,
    n2615,
    n2626
  );


  nand
  g2695
  (
    n2735,
    n2510,
    n2448,
    n2648,
    n2498
  );


  and
  g2696
  (
    n2683,
    n2578,
    n2504,
    n2426,
    n2487
  );


  or
  g2697
  (
    n2806,
    n2463,
    n2573,
    n2470,
    n2642
  );


  or
  g2698
  (
    n2803,
    n2642,
    n2539,
    n2562,
    n2621
  );


  or
  g2699
  (
    n2799,
    n2511,
    n2575,
    n2637,
    n2570
  );


  nand
  g2700
  (
    n2824,
    n2624,
    n2598,
    n2577,
    n2563
  );


  and
  g2701
  (
    n2742,
    n2514,
    n2456,
    n2428,
    n2507
  );


  or
  g2702
  (
    n2759,
    n2627,
    n2446,
    n2485,
    n2442
  );


  xnor
  g2703
  (
    n2700,
    n2631,
    n2652,
    n2482,
    n2561
  );


  xnor
  g2704
  (
    n2756,
    n2633,
    n2570,
    n2632,
    n2604
  );


  xnor
  g2705
  (
    n2719,
    n2561,
    n2479,
    n2425,
    n2616
  );


  and
  g2706
  (
    n2725,
    n2614,
    n2474,
    n2436,
    n2606
  );


  and
  g2707
  (
    n2659,
    n2651,
    n2530,
    n2539,
    n2421
  );


  or
  g2708
  (
    n2679,
    n2490,
    n2542,
    n2613,
    n2640
  );


  xnor
  g2709
  (
    n2692,
    n2636,
    n2600,
    n2421,
    n2650
  );


  or
  g2710
  (
    n2665,
    n2511,
    n2486,
    n2460,
    n2550
  );


  and
  g2711
  (
    n2750,
    n2455,
    n2439,
    n2508,
    n2517
  );


  or
  g2712
  (
    n2783,
    n2473,
    n2633,
    n2468,
    n2606
  );


  or
  g2713
  (
    n2755,
    n2528,
    n2427,
    n2634,
    n1206
  );


  and
  g2714
  (
    n2832,
    n2595,
    n2479,
    n2453,
    n2443
  );


  nor
  g2715
  (
    n2728,
    n2517,
    n2565,
    n2520,
    n2595
  );


  xor
  g2716
  (
    n2699,
    n2635,
    n2566,
    n2585,
    n2578
  );


  and
  g2717
  (
    n2808,
    n2535,
    n2489,
    n2641,
    n2526
  );


  or
  g2718
  (
    n2718,
    n1206,
    n2485,
    n2473,
    n2421
  );


  nand
  g2719
  (
    n2795,
    n2622,
    n2509,
    n2525,
    n2535
  );


  or
  g2720
  (
    n2655,
    n2570,
    n2562,
    n2584,
    n2432
  );


  xnor
  g2721
  (
    n2751,
    n2650,
    n2495,
    n2613,
    n2594
  );


  nand
  g2722
  (
    n2807,
    n2645,
    n2590,
    n2641
  );


  and
  g2723
  (
    n2761,
    n2457,
    n2477,
    n2619,
    n2548
  );


  or
  g2724
  (
    n2685,
    n2643,
    n2557,
    n2487
  );


  nand
  g2725
  (
    n2790,
    n2535,
    n2587,
    n2499,
    n2592
  );


  and
  g2726
  (
    n2721,
    n2548,
    n2431,
    n2469,
    n2584
  );


  xor
  g2727
  (
    n2703,
    n2578,
    n2627,
    n2436,
    n2446
  );


  or
  g2728
  (
    n2764,
    n2567,
    n2429,
    n2549,
    n2427
  );


  xnor
  g2729
  (
    n2791,
    n2572,
    n2536,
    n2473,
    n2506
  );


  nor
  g2730
  (
    n2760,
    n2599,
    n2634,
    n2492,
    n2647
  );


  nand
  g2731
  (
    n2827,
    n2470,
    n1566,
    n2639,
    n2630
  );


  nand
  g2732
  (
    n2726,
    n2519,
    n2425,
    n2581,
    n2653
  );


  xor
  g2733
  (
    n2767,
    n2562,
    n2471,
    n2608,
    n2420
  );


  nand
  g2734
  (
    n2681,
    n2457,
    n2516,
    n2643,
    n2494
  );


  or
  g2735
  (
    n2678,
    n2474,
    n2472,
    n2630,
    n2604
  );


  xor
  g2736
  (
    n2743,
    n2497,
    n1567,
    n2451,
    n2558
  );


  xnor
  g2737
  (
    n2664,
    n2452,
    n2645,
    n2581,
    n2540
  );


  xnor
  g2738
  (
    n2772,
    n2528,
    n2616,
    n2545,
    n2583
  );


  xor
  g2739
  (
    n2671,
    n2620,
    n2551,
    n2547,
    n2556
  );


  nor
  g2740
  (
    n2723,
    n2591,
    n2523,
    n2498,
    n2449
  );


  nand
  g2741
  (
    n2785,
    n2533,
    n2467,
    n2620,
    n2491
  );


  and
  g2742
  (
    n2804,
    n2420,
    n2568,
    n2640,
    n2522
  );


  nor
  g2743
  (
    n2695,
    n2574,
    n2447,
    n2459,
    n2553
  );


  nand
  g2744
  (
    n2784,
    n2441,
    n2579,
    n2632,
    n2499
  );


  xnor
  g2745
  (
    n2658,
    n2489,
    n2461,
    n2420,
    n2650
  );


  nand
  g2746
  (
    n2698,
    n2550,
    n2522,
    n2445,
    n2523
  );


  nand
  g2747
  (
    n2711,
    n2581,
    n2621,
    n2540,
    n2471
  );


  xor
  g2748
  (
    n2662,
    n2596,
    n2575,
    n2434,
    n2512
  );


  nand
  g2749
  (
    n2812,
    n2644,
    n2573,
    n2545,
    n2474
  );


  or
  g2750
  (
    n2720,
    n2423,
    n2532,
    n2649,
    n2537
  );


  and
  g2751
  (
    n2741,
    n2637,
    n2513,
    n2544,
    n2617
  );


  and
  g2752
  (
    n2686,
    n2490,
    n2628,
    n2583,
    n2563
  );


  and
  g2753
  (
    n2739,
    n2571,
    n2567,
    n2568,
    n2598
  );


  xor
  g2754
  (
    n2661,
    n2505,
    n2621,
    n2439,
    n2521
  );


  xnor
  g2755
  (
    n2677,
    n2580,
    n2471,
    n2638,
    n2527
  );


  xor
  g2756
  (
    n2737,
    n2505,
    n2603,
    n2480,
    n2465
  );


  and
  g2757
  (
    n2794,
    n2494,
    n2491,
    n2597,
    n2475
  );


  xor
  g2758
  (
    n2729,
    n2472,
    n2438,
    n2559
  );


  xor
  g2759
  (
    n2712,
    n2521,
    n2610,
    n2465,
    n2553
  );


  nor
  g2760
  (
    n2745,
    n2460,
    n2491,
    n2513,
    n2624
  );


  nand
  g2761
  (
    n2713,
    n2559,
    n2564,
    n2503,
    n2450
  );


  xor
  g2762
  (
    n2657,
    n2574,
    n2507,
    n2500,
    n2547
  );


  or
  g2763
  (
    n2763,
    n2546,
    n2418,
    n2614,
    n2493
  );


  nor
  g2764
  (
    n2707,
    n2601,
    n2588,
    n2564,
    n2566
  );


  nor
  g2765
  (
    n2746,
    n2510,
    n2576,
    n2564,
    n2615
  );


  nor
  g2766
  (
    n2780,
    n2542,
    n2462,
    n2528,
    n2556
  );


  nand
  g2767
  (
    n2704,
    n2459,
    n2607,
    n2593,
    n2552
  );


  nand
  g2768
  (
    n2822,
    n2551,
    n2456,
    n2517,
    n2645
  );


  xor
  g2769
  (
    n2776,
    n2618,
    n2605,
    n2629
  );


  xor
  g2770
  (
    n2684,
    n2552,
    n2456,
    n2424,
    n2514
  );


  xor
  g2771
  (
    n2738,
    n2532,
    n2529,
    n2635,
    n2453
  );


  and
  g2772
  (
    n2693,
    n2514,
    n2543,
    n2481,
    n2531
  );


  nand
  g2773
  (
    n2654,
    n2631,
    n2489,
    n2432,
    n2444
  );


  xnor
  g2774
  (
    n2757,
    n2541,
    n2426,
    n2493,
    n2635
  );


  nand
  g2775
  (
    n2833,
    n2591,
    n2431,
    n2601,
    n2605
  );


  nand
  g2776
  (
    n2732,
    n2620,
    n2586,
    n2437,
    n2476
  );


  nand
  g2777
  (
    n2727,
    n2625,
    n2597,
    n2486,
    n2612
  );


  xor
  g2778
  (
    n2747,
    n2485,
    n2640,
    n2585,
    n2572
  );


  or
  g2779
  (
    n2656,
    n2600,
    n2463,
    n2589,
    n2516
  );


  nor
  g2780
  (
    n2821,
    n2652,
    n2647,
    n2641,
    n878
  );


  xnor
  g2781
  (
    n2770,
    n2505,
    n2423,
    n2506,
    n2440
  );


  xor
  g2782
  (
    n2697,
    n2582,
    n2553,
    n2526,
    n2648
  );


  xnor
  g2783
  (
    n2733,
    n2653,
    n2507,
    n2492,
    n2546
  );


  nor
  g2784
  (
    n2691,
    n2558,
    n2580,
    n2547,
    n2555
  );


  or
  g2785
  (
    n2740,
    n2532,
    n2417,
    n2458,
    n2467
  );


  nor
  g2786
  (
    n2673,
    n2618,
    n2452,
    n2427,
    n2466
  );


  xnor
  g2787
  (
    n2694,
    n2431,
    n2632,
    n2515,
    n2598
  );


  xnor
  g2788
  (
    n2663,
    n2624,
    n2445,
    n2579,
    n2542
  );


  xor
  g2789
  (
    n2667,
    n2653,
    n2522,
    n2573,
    n2511
  );


  xor
  g2790
  (
    n2789,
    n2493,
    n2524,
    n2589,
    n2639
  );


  nor
  g2791
  (
    n2706,
    n2604,
    n2481,
    n2534,
    n2467
  );


  xnor
  g2792
  (
    n2818,
    n2435,
    n2477,
    n2478,
    n2430
  );


  or
  g2793
  (
    n2766,
    n2450,
    n2587,
    n2537,
    n2614
  );


  or
  g2794
  (
    n2810,
    n2503,
    n2646,
    n2529,
    n2560
  );


  xnor
  g2795
  (
    n2682,
    n2447,
    n2502,
    n2482,
    n2549
  );


  and
  g2796
  (
    n2736,
    n2557,
    n2636,
    n2430,
    n2504
  );


  xor
  g2797
  (
    n2800,
    n2530,
    n2533,
    n2497,
    n2652
  );


  nor
  g2798
  (
    n2672,
    n2543,
    n2586,
    n2454,
    n2579
  );


  xnor
  g2799
  (
    n2829,
    n2647,
    n2440,
    n2488,
    n2555
  );


  nand
  g2800
  (
    n2680,
    n2464,
    n2525,
    n2480,
    n2541
  );


  xnor
  g2801
  (
    n2897,
    n2679,
    n2792,
    n2657,
    n2795
  );


  xor
  g2802
  (
    n2899,
    n1588,
    n2708,
    n2742,
    n2684
  );


  nor
  g2803
  (
    n2925,
    n2775,
    n2663,
    n2796,
    n2818
  );


  or
  g2804
  (
    n2879,
    n2760,
    n2677,
    n2660,
    n2791
  );


  and
  g2805
  (
    n2910,
    n2790,
    n2736,
    n1587,
    n2793
  );


  nand
  g2806
  (
    n2916,
    n2832,
    n2823,
    n2786,
    n2746
  );


  xor
  g2807
  (
    n2924,
    n2812,
    n2706,
    n2687,
    n2757
  );


  or
  g2808
  (
    n2871,
    n2789,
    n2786,
    n2778,
    n2694
  );


  and
  g2809
  (
    n2956,
    n2719,
    n2667,
    n2790,
    n2754
  );


  and
  g2810
  (
    n2927,
    n1587,
    n1572,
    n2692,
    n2724
  );


  nand
  g2811
  (
    n2929,
    n1577,
    n1572,
    n2805,
    n2732
  );


  nand
  g2812
  (
    n2923,
    n2788,
    n1577,
    n2749,
    n2714
  );


  xor
  g2813
  (
    n2928,
    n2670,
    n2713,
    n2734,
    n2725
  );


  xnor
  g2814
  (
    n2937,
    n2712,
    n2776,
    n1592,
    n2819
  );


  nand
  g2815
  (
    n2900,
    n2809,
    n2692,
    n2743,
    n2693
  );


  xnor
  g2816
  (
    n2903,
    n2699,
    n2710,
    n2821,
    n2735
  );


  nor
  g2817
  (
    n2931,
    n2784,
    n2743,
    n2757,
    n2781
  );


  xor
  g2818
  (
    n2939,
    n2791,
    n1574,
    n2721,
    n2794
  );


  nor
  g2819
  (
    n2962,
    n1570,
    n2805,
    n2747,
    n2723
  );


  and
  g2820
  (
    n2907,
    n2676,
    n2806,
    n2815,
    n2747
  );


  xor
  g2821
  (
    n2866,
    n2792,
    n2763,
    n2807,
    n2683
  );


  xnor
  g2822
  (
    n2948,
    n2687,
    n2741,
    n2800,
    n2832
  );


  nor
  g2823
  (
    n2834,
    n1582,
    n2760,
    n2658,
    n2816
  );


  xor
  g2824
  (
    n2882,
    n2829,
    n2738,
    n2819,
    n1388
  );


  nor
  g2825
  (
    n2875,
    n2770,
    n2773,
    n2783,
    n1585
  );


  xnor
  g2826
  (
    n2947,
    n2750,
    n2772,
    n2667,
    n2739
  );


  and
  g2827
  (
    n2873,
    n2785,
    n2817,
    n2824,
    n1575
  );


  nand
  g2828
  (
    n2847,
    n2798,
    n2823,
    n2663,
    n2689
  );


  nor
  g2829
  (
    n2854,
    n2690,
    n1572,
    n2801,
    n2716
  );


  or
  g2830
  (
    n2932,
    n1568,
    n2808,
    n2765,
    n2712
  );


  xnor
  g2831
  (
    n2961,
    n2746,
    n1579,
    n2701,
    n2791
  );


  and
  g2832
  (
    n2853,
    n2654,
    n2808,
    n2779,
    n2767
  );


  or
  g2833
  (
    n2933,
    n2774,
    n2705,
    n2656,
    n2702
  );


  xor
  g2834
  (
    n2951,
    n1582,
    n2810,
    n1575,
    n2823
  );


  xor
  g2835
  (
    n2914,
    n2754,
    n2745,
    n1581,
    n2761
  );


  or
  g2836
  (
    n2902,
    n2731,
    n2660,
    n2798
  );


  xor
  g2837
  (
    n2930,
    n2696,
    n2802,
    n2707
  );


  nand
  g2838
  (
    n2890,
    n2714,
    n2655,
    n2778,
    n2674
  );


  and
  g2839
  (
    n2944,
    n1569,
    n1589,
    n2753,
    n2678
  );


  nand
  g2840
  (
    n2918,
    n2758,
    n2794,
    n2772
  );


  nor
  g2841
  (
    n2949,
    n2682,
    n2771,
    n2762,
    n2777
  );


  nand
  g2842
  (
    n2852,
    n2784,
    n2668,
    n2751,
    n2805
  );


  xnor
  g2843
  (
    n2936,
    n1388,
    n2768,
    n2674,
    n2779
  );


  and
  g2844
  (
    n2905,
    n2701,
    n2790,
    n2762,
    n2700
  );


  xor
  g2845
  (
    n2958,
    n2828,
    n2759,
    n2811,
    n2793
  );


  nor
  g2846
  (
    n2883,
    n2806,
    n2678,
    n2754,
    n2780
  );


  nand
  g2847
  (
    n2953,
    n2697,
    n2833,
    n2679,
    n2751
  );


  xnor
  g2848
  (
    n2880,
    n2811,
    n1590,
    n2812,
    n2722
  );


  and
  g2849
  (
    n2844,
    n2702,
    n2796,
    n2814,
    n2672
  );


  nand
  g2850
  (
    n2963,
    n2821,
    n2681,
    n2753,
    n2740
  );


  xnor
  g2851
  (
    n2955,
    n2806,
    n2688,
    n2820,
    n2744
  );


  nor
  g2852
  (
    n2915,
    n2703,
    n2819,
    n2682,
    n1588
  );


  xnor
  g2853
  (
    n2894,
    n2736,
    n2755,
    n2698,
    n2795
  );


  and
  g2854
  (
    n2940,
    n2771,
    n2704,
    n2768,
    n1580
  );


  xnor
  g2855
  (
    n2922,
    n2671,
    n2770,
    n2748,
    n1584
  );


  nand
  g2856
  (
    n2872,
    n2662,
    n1573,
    n2809,
    n2767
  );


  or
  g2857
  (
    n2887,
    n2815,
    n1586,
    n2796,
    n2831
  );


  and
  g2858
  (
    KeyWire_0_50,
    n2685,
    n1206,
    n1591,
    n2659
  );


  xnor
  g2859
  (
    n2843,
    n2770,
    n2799,
    n2737,
    n2673
  );


  nand
  g2860
  (
    n2850,
    n2721,
    n2720,
    n2697,
    n2758
  );


  or
  g2861
  (
    n2857,
    n1580,
    n2761,
    n2828,
    n2722
  );


  or
  g2862
  (
    n2891,
    n2740,
    n2813,
    n1586,
    n2737
  );


  xor
  g2863
  (
    n2935,
    n2696,
    n2807,
    n2832,
    n2759
  );


  or
  g2864
  (
    n2920,
    n2657,
    n2766,
    n2751,
    n2778
  );


  xnor
  g2865
  (
    n2898,
    n2753,
    n1590,
    n2658,
    n2720
  );


  nand
  g2866
  (
    n2950,
    n2730,
    n2707,
    n2782,
    n2795
  );


  or
  g2867
  (
    n2941,
    n2655,
    n2787,
    n2691,
    n2813
  );


  and
  g2868
  (
    n2846,
    n2808,
    n2757,
    n2748,
    n2680
  );


  nor
  g2869
  (
    n2919,
    n2724,
    n2734,
    n2777,
    n2773
  );


  or
  g2870
  (
    n2893,
    n1571,
    n2745,
    n2767,
    n2815
  );


  nand
  g2871
  (
    n2896,
    n2830,
    n2681,
    n2818,
    n2716
  );


  and
  g2872
  (
    n2865,
    n2695,
    n2729,
    n1583,
    n2727
  );


  xnor
  g2873
  (
    n2840,
    n2826,
    n2666,
    n2727,
    n2698
  );


  xnor
  g2874
  (
    n2888,
    n2675,
    n2706,
    n1585,
    n2726
  );


  xnor
  g2875
  (
    n2876,
    n1571,
    n2654,
    n2773,
    n1579
  );


  or
  g2876
  (
    n2851,
    n2659,
    n2782,
    n2809,
    n2764
  );


  nand
  g2877
  (
    n2926,
    n2662,
    n2781,
    n2826,
    n2717
  );


  or
  g2878
  (
    n2842,
    n2788,
    n2768,
    n2827,
    n2822
  );


  and
  g2879
  (
    n2895,
    n1591,
    n2684,
    n2829,
    n2675
  );


  and
  g2880
  (
    n2906,
    n2776,
    n2797,
    n2803,
    n2831
  );


  xnor
  g2881
  (
    n2889,
    n2829,
    n2792,
    n2816,
    n1582
  );


  xnor
  g2882
  (
    n2856,
    n2693,
    n2816,
    n2774,
    n2826
  );


  xnor
  g2883
  (
    n2943,
    n2766,
    n2784,
    n2756,
    n2813
  );


  and
  g2884
  (
    n2855,
    n2704,
    n2733,
    n2782,
    n2689
  );


  xor
  g2885
  (
    n2885,
    n1592,
    n1578,
    n2812,
    n2665
  );


  xor
  g2886
  (
    n2863,
    n2709,
    n2749,
    n2688,
    n2752
  );


  and
  g2887
  (
    n2909,
    n2787,
    n2825,
    n1586,
    n2800
  );


  and
  g2888
  (
    n2878,
    n2726,
    n2814,
    n2793,
    n2764
  );


  nor
  g2889
  (
    n2835,
    n2765,
    n1579,
    n2719,
    n2769
  );


  or
  g2890
  (
    n2959,
    n2804,
    n2775,
    n2661,
    n2690
  );


  and
  g2891
  (
    n2901,
    n2680,
    n2741,
    n2756,
    n2803
  );


  or
  g2892
  (
    n2862,
    n2774,
    n1576,
    n1578,
    n2668
  );


  xnor
  g2893
  (
    n2938,
    n2789,
    n2744,
    n2750,
    n1584
  );


  and
  g2894
  (
    n2861,
    n1574,
    n2723,
    n1576,
    n2801
  );


  nor
  g2895
  (
    n2841,
    n2708,
    n2691,
    n2824,
    n2811
  );


  nand
  g2896
  (
    n2908,
    n2728,
    n2664,
    n2755,
    n2665
  );


  nor
  g2897
  (
    n2837,
    n2822,
    n2831,
    n2787,
    n1581
  );


  xnor
  g2898
  (
    n2859,
    n1577,
    n2785,
    n2830,
    n1569
  );


  nor
  g2899
  (
    n2868,
    n2801,
    n2788,
    n2760,
    n2755
  );


  nor
  g2900
  (
    n2960,
    n2735,
    n2824,
    n1568,
    n2742
  );


  and
  g2901
  (
    n2877,
    n2725,
    n1583,
    n1573,
    n2717
  );


  xor
  g2902
  (
    n2934,
    n2817,
    n2686,
    n2699,
    n2827
  );


  nor
  g2903
  (
    n2869,
    n1589,
    n2676,
    n2762,
    n2803
  );


  and
  g2904
  (
    n2839,
    n2781,
    n2818,
    n2769,
    n2669
  );


  xor
  g2905
  (
    n2886,
    n2700,
    n1581,
    n2780,
    n2830
  );


  and
  g2906
  (
    n2946,
    n2810,
    n2661,
    n2817,
    n2711
  );


  and
  g2907
  (
    n2874,
    n2783,
    n2820,
    n2776,
    n2825
  );


  nand
  g2908
  (
    n2913,
    n2756,
    n2686,
    n2730,
    n2752
  );


  and
  g2909
  (
    n2858,
    n2814,
    n1578,
    n2821,
    n2670
  );


  xor
  g2910
  (
    n2848,
    n2677,
    n2695,
    n1585,
    n2763
  );


  nand
  g2911
  (
    n2945,
    n2799,
    n2833,
    n2669,
    n2777
  );


  nand
  g2912
  (
    n2870,
    n1570,
    n2807,
    n2783,
    n2656
  );


  nor
  g2913
  (
    n2921,
    n2710,
    n2664,
    n2750,
    n2765
  );


  and
  g2914
  (
    n2942,
    n2733,
    n1574,
    n2827,
    n2766
  );


  nand
  g2915
  (
    n2917,
    n1575,
    n2828,
    n2705,
    n1592
  );


  nor
  g2916
  (
    n2957,
    n1591,
    n2820,
    n2769,
    n2739
  );


  xnor
  g2917
  (
    n2954,
    n2825,
    n2713,
    n2694,
    n2731
  );


  nor
  g2918
  (
    n2867,
    n2759,
    n2715,
    n2804,
    n1589
  );


  xor
  g2919
  (
    n2912,
    n1580,
    n2800,
    n2683,
    n2685
  );


  xnor
  g2920
  (
    n2904,
    n2802,
    n2799,
    n1583,
    n2728
  );


  nand
  g2921
  (
    n2964,
    n2786,
    n1590,
    n1588,
    n2810
  );


  xnor
  g2922
  (
    n2881,
    n1584,
    n2732,
    n2711,
    n2772
  );


  xnor
  g2923
  (
    n2860,
    n2761,
    n2779,
    n2763,
    n1587
  );


  nor
  g2924
  (
    n2836,
    n2666,
    n1568,
    n2797
  );


  xnor
  g2925
  (
    n2849,
    n2789,
    n2833,
    n1573,
    n2752
  );


  nor
  g2926
  (
    n2892,
    n2804,
    n2715,
    n2672,
    n2738
  );


  xnor
  g2927
  (
    n2952,
    n2764,
    n2718,
    n1567,
    n2673
  );


  nand
  g2928
  (
    n2845,
    n2729,
    n2775,
    n2709,
    n1576
  );


  and
  g2929
  (
    n2884,
    n2718,
    n1571,
    n2771,
    n2780
  );


  nand
  g2930
  (
    n2864,
    n2671,
    n2703,
    n2785,
    n1567
  );


  nor
  g2931
  (
    n2838,
    n2758,
    n1570,
    n1569,
    n2822
  );


  or
  g2932
  (
    n2966,
    n2839,
    n2837,
    n2845,
    n2844
  );


  nand
  g2933
  (
    n2965,
    n2848,
    n2846,
    n2834,
    n2840
  );


  and
  g2934
  (
    n2968,
    n2849,
    n2836,
    n2842,
    n2838
  );


  xor
  g2935
  (
    n2967,
    n2843,
    n2841,
    n2835,
    n2847
  );


  xor
  g2936
  (
    n2971,
    n2850,
    n2966
  );


  buf
  g2937
  (
    n2969,
    n879
  );


  xor
  g2938
  (
    n2970,
    n2852,
    n2851,
    n2967,
    n2965
  );


  nor
  g2939
  (
    n2980,
    n2971,
    n2859,
    n2879,
    n2864
  );


  nand
  g2940
  (
    n2973,
    n2855,
    n2970,
    n2969,
    n2883
  );


  xor
  g2941
  (
    n2978,
    n2866,
    n2872,
    n2865,
    n2857
  );


  xor
  g2942
  (
    n2976,
    n2874,
    n2862,
    n2970,
    n2884
  );


  xnor
  g2943
  (
    n2982,
    n2971,
    n2880,
    n2853,
    n2869
  );


  nand
  g2944
  (
    n2972,
    n2871,
    n2971,
    n2969,
    n2876
  );


  xnor
  g2945
  (
    n2974,
    n2970,
    n2854,
    n2870,
    n2877
  );


  nor
  g2946
  (
    n2975,
    n2882,
    n2858,
    n2881,
    n2971
  );


  nor
  g2947
  (
    n2979,
    n2873,
    n2969,
    n2968,
    n2970
  );


  nand
  g2948
  (
    n2977,
    n2867,
    n2863,
    n2875,
    n2856
  );


  xor
  g2949
  (
    n2981,
    n2878,
    n2861,
    n2868,
    n2860
  );


  or
  g2950
  (
    n2983,
    n881,
    n880,
    n884,
    n883
  );


  nand
  g2951
  (
    n2985,
    n880,
    n882,
    n2975,
    n883
  );


  xor
  g2952
  (
    KeyWire_0_38,
    n880,
    n2972,
    n882
  );


  nor
  g2953
  (
    n2984,
    n2976,
    n881,
    n883,
    n2974
  );


  and
  g2954
  (
    n2986,
    n884,
    n884,
    n881,
    n2973
  );


  nand
  g2955
  (
    n2988,
    n2914,
    n2932,
    n2984,
    n2918
  );


  xor
  g2956
  (
    n2990,
    n2899,
    n2987,
    n2911,
    n885
  );


  xor
  g2957
  (
    n2997,
    n2923,
    n2906,
    n2908,
    n2886
  );


  xor
  g2958
  (
    n3006,
    n2981,
    n2980,
    n2983,
    n2888
  );


  nand
  g2959
  (
    n2999,
    n2987,
    n2902,
    n2910,
    n2983
  );


  or
  g2960
  (
    n3003,
    n2913,
    n2987,
    n2927,
    n2909
  );


  xor
  g2961
  (
    n3000,
    n2981,
    n2890,
    n2895,
    n2893
  );


  and
  g2962
  (
    n2998,
    n2903,
    n2920,
    n2985,
    n2924
  );


  xnor
  g2963
  (
    n2996,
    n2898,
    n2987,
    n2894,
    n2986
  );


  xor
  g2964
  (
    n3005,
    n2896,
    n2979,
    n2985,
    n2919
  );


  xnor
  g2965
  (
    n3002,
    n2912,
    n2929,
    n2986,
    n2926
  );


  nand
  g2966
  (
    n2995,
    n2930,
    n2983,
    n2986,
    n2907
  );


  xor
  g2967
  (
    n2993,
    n2915,
    n2933,
    n2887,
    n2984
  );


  xor
  g2968
  (
    n3001,
    n2982,
    n2901,
    n2921,
    n2885
  );


  and
  g2969
  (
    n2989,
    n2984,
    n2980,
    n2900,
    n2897
  );


  and
  g2970
  (
    n2992,
    n2892,
    n2985,
    n2889,
    n2980
  );


  xnor
  g2971
  (
    n3004,
    n2931,
    n2904,
    n2925,
    n2917
  );


  xnor
  g2972
  (
    n3007,
    n2981,
    n2977,
    n2984,
    n2985
  );


  xnor
  g2973
  (
    n2994,
    n2928,
    n2905,
    n2978,
    n2922
  );


  nor
  g2974
  (
    n2991,
    n2986,
    n2983,
    n2891,
    n2916
  );


  xor
  g2975
  (
    n3009,
    n2988,
    n2990,
    n2936,
    n2995
  );


  xor
  g2976
  (
    n3008,
    n2992,
    n2950,
    n3000,
    n2942
  );


  or
  g2977
  (
    n3012,
    n2935,
    n3001,
    n2941,
    n2989
  );


  nor
  g2978
  (
    n3014,
    n2939,
    n2934,
    n2945,
    n2948
  );


  xor
  g2979
  (
    n3010,
    n2946,
    n2993,
    n2943,
    n2940
  );


  nand
  g2980
  (
    n3011,
    n2991,
    n2949,
    n2997,
    n2944
  );


  nand
  g2981
  (
    n3015,
    n2994,
    n2951,
    n2937,
    n2998
  );


  nor
  g2982
  (
    n3013,
    n2938,
    n2947,
    n2999,
    n2996
  );


  or
  g2983
  (
    n3016,
    n2952,
    n2954,
    n3015,
    n2953
  );


  nand
  g2984
  (
    n3019,
    n2961,
    n2962,
    n2982
  );


  nand
  g2985
  (
    n3017,
    n3016,
    n3016,
    n2982,
    n2955
  );


  or
  g2986
  (
    n3018,
    n2959,
    n3016,
    n2960,
    n2958
  );


  nand
  g2987
  (
    n3020,
    n2963,
    n2956,
    n3016,
    n2957
  );


  and
  g2988
  (
    n3022,
    n887,
    n888,
    n886
  );


  nand
  g2989
  (
    n3023,
    n886,
    n887,
    n3019
  );


  or
  g2990
  (
    n3021,
    n3018,
    n885,
    n3017
  );


  buf
  g2991
  (
    n3024,
    n3022
  );


  not
  g2992
  (
    n3025,
    n3023
  );


  nor
  g2993
  (
    n3026,
    n889,
    n888,
    n3025
  );


  nor
  g2994
  (
    n3027,
    n3005,
    n3004,
    n3003,
    n3002
  );


  and
  g2995
  (
    n3028,
    n3006,
    n3007,
    n3026
  );


  buf
  g2996
  (
    n3030,
    n2964
  );


  buf
  g2997
  (
    n3029,
    n3028
  );


  xnor
  g2998
  (
    n3031,
    n3027,
    n3028
  );


  nand
  g2999
  (
    n3032,
    n3020,
    n889,
    n3031
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n527,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1831,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1640,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n2193,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n2298,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n2502,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n131,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1915,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n443,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n448,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n2597,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n2226,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1269,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n2510,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n2125,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n381,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n2433,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n517,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n2234,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n382,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n2404,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1863,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n92,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1909,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1799,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1108,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n651,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n1464,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n328,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n93,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n1286,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n257,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n1172,
    keyIn_0_32,
    KeyWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n1822,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n255,
    KeyNOTWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n1160,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n883,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n886,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n2987,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n1987,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n816,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n1585,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n2498,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n264,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n1824,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n2635,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n781,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n1875,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n2640,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n1597,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n2911,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n1794,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n1064,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n1639,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n1052,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n922,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n1433,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n2119,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n1148,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n2774,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n1779,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n809,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    n2295,
    keyIn_0_62,
    KeyWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n1476,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

