

module Stat_2000_205
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n889,
  n882,
  n883,
  n877,
  n890,
  n895,
  n881,
  n876,
  n892,
  n873,
  n891,
  n893,
  n874,
  n898,
  n886,
  n885,
  n875,
  n2020,
  n2025,
  n2021,
  n2029,
  n2030,
  n2024,
  n2031,
  n2028,
  n2019,
  n2022,
  n2026,
  n2027,
  n2018,
  n2032,
  n2023,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n889;
  output n882;
  output n883;
  output n877;
  output n890;
  output n895;
  output n881;
  output n876;
  output n892;
  output n873;
  output n891;
  output n893;
  output n874;
  output n898;
  output n886;
  output n885;
  output n875;
  output n2020;
  output n2025;
  output n2021;
  output n2029;
  output n2030;
  output n2024;
  output n2031;
  output n2028;
  output n2019;
  output n2022;
  output n2026;
  output n2027;
  output n2018;
  output n2032;
  output n2023;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n878;
  wire n879;
  wire n880;
  wire n884;
  wire n887;
  wire n888;
  wire n894;
  wire n896;
  wire n897;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    n43,
    n18
  );


  buf
  g1
  (
    n45,
    n16
  );


  buf
  g2
  (
    n120,
    n28
  );


  buf
  g3
  (
    n47,
    n22
  );


  buf
  g4
  (
    n104,
    n19
  );


  buf
  g5
  (
    n55,
    n10
  );


  buf
  g6
  (
    KeyWire_0_33,
    n14
  );


  not
  g7
  (
    n58,
    n24
  );


  not
  g8
  (
    n121,
    n28
  );


  buf
  g9
  (
    n95,
    n25
  );


  buf
  g10
  (
    n66,
    n3
  );


  buf
  g11
  (
    n89,
    n11
  );


  not
  g12
  (
    n141,
    n22
  );


  not
  g13
  (
    n35,
    n3
  );


  not
  g14
  (
    n144,
    n5
  );


  buf
  g15
  (
    n77,
    n28
  );


  buf
  g16
  (
    n96,
    n10
  );


  not
  g17
  (
    n112,
    n19
  );


  buf
  g18
  (
    n38,
    n13
  );


  not
  g19
  (
    n97,
    n8
  );


  not
  g20
  (
    n108,
    n6
  );


  buf
  g21
  (
    n114,
    n17
  );


  not
  g22
  (
    n102,
    n18
  );


  not
  g23
  (
    n75,
    n17
  );


  buf
  g24
  (
    n67,
    n1
  );


  buf
  g25
  (
    n80,
    n14
  );


  buf
  g26
  (
    n73,
    n10
  );


  buf
  g27
  (
    n125,
    n22
  );


  not
  g28
  (
    n113,
    n24
  );


  buf
  g29
  (
    n138,
    n6
  );


  not
  g30
  (
    n107,
    n21
  );


  buf
  g31
  (
    n123,
    n15
  );


  not
  g32
  (
    n131,
    n26
  );


  not
  g33
  (
    n64,
    n24
  );


  not
  g34
  (
    n70,
    n26
  );


  not
  g35
  (
    n86,
    n8
  );


  not
  g36
  (
    n44,
    n21
  );


  buf
  g37
  (
    n50,
    n4
  );


  buf
  g38
  (
    n33,
    n20
  );


  not
  g39
  (
    n100,
    n29
  );


  not
  g40
  (
    n118,
    n25
  );


  buf
  g41
  (
    n91,
    n8
  );


  buf
  g42
  (
    n93,
    n9
  );


  buf
  g43
  (
    n68,
    n23
  );


  buf
  g44
  (
    n111,
    n18
  );


  buf
  g45
  (
    n106,
    n7
  );


  not
  g46
  (
    n41,
    n16
  );


  buf
  g47
  (
    n99,
    n28
  );


  not
  g48
  (
    n39,
    n5
  );


  not
  g49
  (
    n132,
    n3
  );


  buf
  g50
  (
    n49,
    n2
  );


  not
  g51
  (
    n115,
    n15
  );


  buf
  g52
  (
    n94,
    n13
  );


  not
  g53
  (
    n81,
    n26
  );


  not
  g54
  (
    n88,
    n12
  );


  buf
  g55
  (
    n133,
    n16
  );


  buf
  g56
  (
    n61,
    n13
  );


  buf
  g57
  (
    n74,
    n17
  );


  buf
  g58
  (
    n142,
    n29
  );


  buf
  g59
  (
    n36,
    n6
  );


  not
  g60
  (
    n127,
    n20
  );


  buf
  g61
  (
    n136,
    n27
  );


  not
  g62
  (
    n69,
    n15
  );


  not
  g63
  (
    n116,
    n20
  );


  not
  g64
  (
    n40,
    n27
  );


  not
  g65
  (
    n130,
    n19
  );


  not
  g66
  (
    n124,
    n23
  );


  not
  g67
  (
    n76,
    n4
  );


  buf
  g68
  (
    n87,
    n11
  );


  not
  g69
  (
    n139,
    n15
  );


  not
  g70
  (
    n59,
    n12
  );


  buf
  g71
  (
    n72,
    n23
  );


  not
  g72
  (
    n82,
    n25
  );


  not
  g73
  (
    n42,
    n1
  );


  not
  g74
  (
    n140,
    n27
  );


  not
  g75
  (
    n54,
    n8
  );


  buf
  g76
  (
    n51,
    n20
  );


  not
  g77
  (
    n52,
    n1
  );


  buf
  g78
  (
    n145,
    n7
  );


  buf
  g79
  (
    n56,
    n12
  );


  buf
  g80
  (
    n105,
    n9
  );


  buf
  g81
  (
    n128,
    n24
  );


  not
  g82
  (
    n122,
    n9
  );


  not
  g83
  (
    n109,
    n2
  );


  not
  g84
  (
    n137,
    n10
  );


  buf
  g85
  (
    n143,
    n21
  );


  buf
  g86
  (
    n62,
    n17
  );


  not
  g87
  (
    n65,
    n21
  );


  not
  g88
  (
    n79,
    n1
  );


  buf
  g89
  (
    n117,
    n19
  );


  not
  g90
  (
    n71,
    n2
  );


  not
  g91
  (
    n46,
    n22
  );


  buf
  g92
  (
    n78,
    n13
  );


  buf
  g93
  (
    n90,
    n5
  );


  buf
  g94
  (
    n103,
    n7
  );


  buf
  g95
  (
    n135,
    n2
  );


  not
  g96
  (
    n134,
    n14
  );


  buf
  g97
  (
    n98,
    n12
  );


  buf
  g98
  (
    n60,
    n27
  );


  buf
  g99
  (
    n129,
    n5
  );


  buf
  g100
  (
    n37,
    n4
  );


  buf
  g101
  (
    n92,
    n25
  );


  buf
  g102
  (
    n146,
    n11
  );


  buf
  g103
  (
    n83,
    n6
  );


  buf
  g104
  (
    n63,
    n4
  );


  buf
  g105
  (
    n110,
    n9
  );


  buf
  g106
  (
    n119,
    n26
  );


  buf
  g107
  (
    n85,
    n16
  );


  not
  g108
  (
    n34,
    n11
  );


  not
  g109
  (
    n53,
    n14
  );


  buf
  g110
  (
    n57,
    n3
  );


  not
  g111
  (
    n48,
    n18
  );


  not
  g112
  (
    n126,
    n7
  );


  buf
  g113
  (
    n84,
    n23
  );


  buf
  g114
  (
    n567,
    n40
  );


  not
  g115
  (
    n493,
    n58
  );


  not
  g116
  (
    n511,
    n129
  );


  buf
  g117
  (
    n540,
    n110
  );


  buf
  g118
  (
    n422,
    n72
  );


  buf
  g119
  (
    n190,
    n124
  );


  buf
  g120
  (
    n296,
    n130
  );


  not
  g121
  (
    n242,
    n46
  );


  not
  g122
  (
    n485,
    n123
  );


  buf
  g123
  (
    n530,
    n136
  );


  not
  g124
  (
    n300,
    n44
  );


  not
  g125
  (
    n508,
    n111
  );


  buf
  g126
  (
    n550,
    n110
  );


  not
  g127
  (
    n239,
    n84
  );


  not
  g128
  (
    n324,
    n50
  );


  buf
  g129
  (
    n458,
    n89
  );


  not
  g130
  (
    n168,
    n92
  );


  buf
  g131
  (
    n435,
    n70
  );


  buf
  g132
  (
    n498,
    n107
  );


  buf
  g133
  (
    n566,
    n49
  );


  not
  g134
  (
    n198,
    n87
  );


  not
  g135
  (
    n288,
    n34
  );


  not
  g136
  (
    n526,
    n49
  );


  buf
  g137
  (
    n335,
    n142
  );


  not
  g138
  (
    n318,
    n133
  );


  buf
  g139
  (
    n248,
    n140
  );


  buf
  g140
  (
    n468,
    n104
  );


  not
  g141
  (
    n406,
    n42
  );


  buf
  g142
  (
    n419,
    n128
  );


  buf
  g143
  (
    n392,
    n57
  );


  buf
  g144
  (
    n174,
    n54
  );


  not
  g145
  (
    n428,
    n108
  );


  not
  g146
  (
    n203,
    n142
  );


  buf
  g147
  (
    n505,
    n87
  );


  not
  g148
  (
    n533,
    n143
  );


  not
  g149
  (
    n243,
    n37
  );


  not
  g150
  (
    n257,
    n46
  );


  buf
  g151
  (
    n373,
    n75
  );


  not
  g152
  (
    n399,
    n61
  );


  not
  g153
  (
    n184,
    n102
  );


  buf
  g154
  (
    n363,
    n143
  );


  not
  g155
  (
    n592,
    n35
  );


  buf
  g156
  (
    n453,
    n65
  );


  buf
  g157
  (
    n195,
    n142
  );


  not
  g158
  (
    n472,
    n70
  );


  buf
  g159
  (
    n587,
    n128
  );


  buf
  g160
  (
    n506,
    n67
  );


  buf
  g161
  (
    n438,
    n93
  );


  not
  g162
  (
    n416,
    n79
  );


  buf
  g163
  (
    n369,
    n71
  );


  not
  g164
  (
    n549,
    n42
  );


  not
  g165
  (
    n333,
    n126
  );


  not
  g166
  (
    n299,
    n104
  );


  not
  g167
  (
    n378,
    n64
  );


  not
  g168
  (
    n525,
    n130
  );


  buf
  g169
  (
    n451,
    n91
  );


  buf
  g170
  (
    n590,
    n137
  );


  not
  g171
  (
    KeyWire_0_35,
    n139
  );


  not
  g172
  (
    n444,
    n39
  );


  buf
  g173
  (
    n301,
    n122
  );


  not
  g174
  (
    n375,
    n40
  );


  not
  g175
  (
    n555,
    n121
  );


  buf
  g176
  (
    n338,
    n132
  );


  not
  g177
  (
    n230,
    n67
  );


  buf
  g178
  (
    n327,
    n83
  );


  not
  g179
  (
    n414,
    n39
  );


  not
  g180
  (
    n155,
    n109
  );


  not
  g181
  (
    n343,
    n46
  );


  not
  g182
  (
    n255,
    n66
  );


  not
  g183
  (
    n322,
    n131
  );


  not
  g184
  (
    n586,
    n36
  );


  not
  g185
  (
    n311,
    n112
  );


  not
  g186
  (
    n497,
    n65
  );


  not
  g187
  (
    n328,
    n88
  );


  not
  g188
  (
    n362,
    n102
  );


  buf
  g189
  (
    n261,
    n134
  );


  not
  g190
  (
    n353,
    n60
  );


  not
  g191
  (
    n377,
    n64
  );


  not
  g192
  (
    n185,
    n86
  );


  buf
  g193
  (
    n381,
    n85
  );


  not
  g194
  (
    n293,
    n133
  );


  buf
  g195
  (
    KeyWire_0_8,
    n36
  );


  buf
  g196
  (
    n359,
    n92
  );


  buf
  g197
  (
    n229,
    n113
  );


  not
  g198
  (
    n454,
    n85
  );


  buf
  g199
  (
    n517,
    n143
  );


  not
  g200
  (
    n187,
    n139
  );


  buf
  g201
  (
    n501,
    n121
  );


  buf
  g202
  (
    n361,
    n104
  );


  not
  g203
  (
    n431,
    n74
  );


  buf
  g204
  (
    n263,
    n62
  );


  buf
  g205
  (
    n319,
    n65
  );


  not
  g206
  (
    n394,
    n48
  );


  buf
  g207
  (
    n147,
    n34
  );


  not
  g208
  (
    KeyWire_0_11,
    n81
  );


  buf
  g209
  (
    n231,
    n89
  );


  not
  g210
  (
    n568,
    n78
  );


  not
  g211
  (
    n515,
    n137
  );


  buf
  g212
  (
    n595,
    n81
  );


  not
  g213
  (
    n447,
    n73
  );


  buf
  g214
  (
    n236,
    n81
  );


  buf
  g215
  (
    n320,
    n36
  );


  not
  g216
  (
    n214,
    n75
  );


  buf
  g217
  (
    n233,
    n128
  );


  buf
  g218
  (
    n286,
    n109
  );


  not
  g219
  (
    n461,
    n133
  );


  buf
  g220
  (
    n316,
    n120
  );


  not
  g221
  (
    n271,
    n67
  );


  buf
  g222
  (
    KeyWire_0_55,
    n96
  );


  not
  g223
  (
    n596,
    n42
  );


  not
  g224
  (
    n194,
    n33
  );


  not
  g225
  (
    n345,
    n66
  );


  buf
  g226
  (
    n516,
    n137
  );


  not
  g227
  (
    n332,
    n39
  );


  buf
  g228
  (
    n238,
    n138
  );


  buf
  g229
  (
    n507,
    n118
  );


  not
  g230
  (
    n417,
    n37
  );


  buf
  g231
  (
    n434,
    n141
  );


  not
  g232
  (
    n210,
    n56
  );


  buf
  g233
  (
    n425,
    n122
  );


  not
  g234
  (
    n509,
    n81
  );


  not
  g235
  (
    n561,
    n61
  );


  buf
  g236
  (
    n289,
    n62
  );


  not
  g237
  (
    n151,
    n91
  );


  buf
  g238
  (
    n235,
    n108
  );


  not
  g239
  (
    n499,
    n124
  );


  not
  g240
  (
    n348,
    n78
  );


  buf
  g241
  (
    n302,
    n113
  );


  not
  g242
  (
    n452,
    n143
  );


  buf
  g243
  (
    n269,
    n116
  );


  buf
  g244
  (
    n227,
    n103
  );


  not
  g245
  (
    n237,
    n145
  );


  not
  g246
  (
    n339,
    n131
  );


  not
  g247
  (
    n388,
    n43
  );


  buf
  g248
  (
    n266,
    n133
  );


  buf
  g249
  (
    n215,
    n136
  );


  not
  g250
  (
    n427,
    n95
  );


  not
  g251
  (
    n400,
    n107
  );


  not
  g252
  (
    n352,
    n84
  );


  buf
  g253
  (
    n351,
    n55
  );


  buf
  g254
  (
    n518,
    n119
  );


  not
  g255
  (
    n349,
    n73
  );


  not
  g256
  (
    n225,
    n116
  );


  buf
  g257
  (
    n284,
    n33
  );


  buf
  g258
  (
    n376,
    n125
  );


  not
  g259
  (
    n183,
    n40
  );


  not
  g260
  (
    n281,
    n145
  );


  buf
  g261
  (
    n481,
    n42
  );


  buf
  g262
  (
    n207,
    n59
  );


  buf
  g263
  (
    n186,
    n44
  );


  buf
  g264
  (
    n522,
    n117
  );


  buf
  g265
  (
    n455,
    n56
  );


  buf
  g266
  (
    n344,
    n34
  );


  not
  g267
  (
    n408,
    n76
  );


  buf
  g268
  (
    n330,
    n97
  );


  not
  g269
  (
    n448,
    n35
  );


  buf
  g270
  (
    n157,
    n83
  );


  not
  g271
  (
    n442,
    n87
  );


  not
  g272
  (
    n158,
    n139
  );


  not
  g273
  (
    n259,
    n137
  );


  not
  g274
  (
    n470,
    n74
  );


  not
  g275
  (
    n492,
    n43
  );


  buf
  g276
  (
    n169,
    n96
  );


  buf
  g277
  (
    n557,
    n124
  );


  not
  g278
  (
    KeyWire_0_62,
    n134
  );


  buf
  g279
  (
    n390,
    n94
  );


  not
  g280
  (
    n188,
    n58
  );


  buf
  g281
  (
    n209,
    n122
  );


  not
  g282
  (
    n382,
    n68
  );


  not
  g283
  (
    n254,
    n72
  );


  not
  g284
  (
    n486,
    n45
  );


  buf
  g285
  (
    n521,
    n127
  );


  not
  g286
  (
    n401,
    n57
  );


  buf
  g287
  (
    n383,
    n130
  );


  buf
  g288
  (
    n367,
    n92
  );


  not
  g289
  (
    n262,
    n118
  );


  not
  g290
  (
    n573,
    n115
  );


  not
  g291
  (
    n528,
    n95
  );


  buf
  g292
  (
    n380,
    n116
  );


  not
  g293
  (
    n212,
    n79
  );


  not
  g294
  (
    n432,
    n58
  );


  not
  g295
  (
    n273,
    n68
  );


  not
  g296
  (
    n563,
    n55
  );


  not
  g297
  (
    n467,
    n76
  );


  buf
  g298
  (
    n552,
    n48
  );


  buf
  g299
  (
    n163,
    n113
  );


  buf
  g300
  (
    n201,
    n118
  );


  buf
  g301
  (
    n177,
    n88
  );


  not
  g302
  (
    n405,
    n44
  );


  not
  g303
  (
    n576,
    n126
  );


  not
  g304
  (
    n487,
    n107
  );


  not
  g305
  (
    n479,
    n131
  );


  not
  g306
  (
    n265,
    n120
  );


  not
  g307
  (
    n436,
    n76
  );


  not
  g308
  (
    n379,
    n70
  );


  not
  g309
  (
    n170,
    n116
  );


  not
  g310
  (
    n189,
    n115
  );


  not
  g311
  (
    n433,
    n110
  );


  buf
  g312
  (
    n503,
    n41
  );


  buf
  g313
  (
    n274,
    n52
  );


  not
  g314
  (
    n173,
    n71
  );


  not
  g315
  (
    n409,
    n68
  );


  not
  g316
  (
    n331,
    n95
  );


  not
  g317
  (
    KeyWire_0_45,
    n79
  );


  buf
  g318
  (
    n290,
    n87
  );


  not
  g319
  (
    n558,
    n134
  );


  not
  g320
  (
    n370,
    n65
  );


  buf
  g321
  (
    n192,
    n140
  );


  not
  g322
  (
    n357,
    n97
  );


  buf
  g323
  (
    n253,
    n107
  );


  not
  g324
  (
    n553,
    n144
  );


  not
  g325
  (
    n488,
    n38
  );


  buf
  g326
  (
    n413,
    n125
  );


  not
  g327
  (
    n245,
    n38
  );


  buf
  g328
  (
    n366,
    n78
  );


  not
  g329
  (
    n474,
    n106
  );


  not
  g330
  (
    n536,
    n77
  );


  not
  g331
  (
    n329,
    n112
  );


  buf
  g332
  (
    n581,
    n43
  );


  not
  g333
  (
    n213,
    n129
  );


  not
  g334
  (
    n389,
    n77
  );


  buf
  g335
  (
    n222,
    n75
  );


  buf
  g336
  (
    n226,
    n130
  );


  buf
  g337
  (
    n205,
    n89
  );


  not
  g338
  (
    KeyWire_0_30,
    n83
  );


  buf
  g339
  (
    n456,
    n49
  );


  not
  g340
  (
    n386,
    n52
  );


  not
  g341
  (
    n597,
    n121
  );


  not
  g342
  (
    n465,
    n59
  );


  buf
  g343
  (
    n411,
    n41
  );


  buf
  g344
  (
    n478,
    n74
  );


  buf
  g345
  (
    n234,
    n123
  );


  not
  g346
  (
    n548,
    n68
  );


  buf
  g347
  (
    n494,
    n124
  );


  buf
  g348
  (
    n412,
    n135
  );


  buf
  g349
  (
    n384,
    n90
  );


  buf
  g350
  (
    n569,
    n66
  );


  buf
  g351
  (
    n572,
    n121
  );


  buf
  g352
  (
    n337,
    n129
  );


  buf
  g353
  (
    n580,
    n94
  );


  not
  g354
  (
    n420,
    n132
  );


  buf
  g355
  (
    n532,
    n45
  );


  not
  g356
  (
    n391,
    n99
  );


  buf
  g357
  (
    n223,
    n80
  );


  buf
  g358
  (
    n307,
    n123
  );


  buf
  g359
  (
    n276,
    n50
  );


  buf
  g360
  (
    n292,
    n140
  );


  buf
  g361
  (
    n407,
    n60
  );


  not
  g362
  (
    n202,
    n99
  );


  not
  g363
  (
    n310,
    n97
  );


  not
  g364
  (
    n559,
    n80
  );


  buf
  g365
  (
    n149,
    n47
  );


  not
  g366
  (
    n403,
    n37
  );


  not
  g367
  (
    n252,
    n46
  );


  buf
  g368
  (
    n181,
    n101
  );


  not
  g369
  (
    n208,
    n135
  );


  buf
  g370
  (
    KeyWire_0_29,
    n141
  );


  buf
  g371
  (
    n244,
    n91
  );


  not
  g372
  (
    n258,
    n59
  );


  buf
  g373
  (
    n342,
    n105
  );


  not
  g374
  (
    n277,
    n98
  );


  not
  g375
  (
    n534,
    n127
  );


  buf
  g376
  (
    n395,
    n106
  );


  buf
  g377
  (
    n228,
    n111
  );


  buf
  g378
  (
    n268,
    n86
  );


  buf
  g379
  (
    n176,
    n114
  );


  buf
  g380
  (
    KeyWire_0_24,
    n114
  );


  buf
  g381
  (
    n510,
    n48
  );


  not
  g382
  (
    n457,
    n63
  );


  buf
  g383
  (
    n500,
    n101
  );


  not
  g384
  (
    n421,
    n113
  );


  buf
  g385
  (
    n317,
    n82
  );


  buf
  g386
  (
    n314,
    n58
  );


  not
  g387
  (
    n398,
    n54
  );


  not
  g388
  (
    n476,
    n103
  );


  not
  g389
  (
    n346,
    n125
  );


  buf
  g390
  (
    n368,
    n88
  );


  buf
  g391
  (
    n221,
    n135
  );


  buf
  g392
  (
    KeyWire_0_52,
    n76
  );


  buf
  g393
  (
    n285,
    n86
  );


  not
  g394
  (
    n180,
    n71
  );


  not
  g395
  (
    KeyWire_0_53,
    n60
  );


  buf
  g396
  (
    n387,
    n82
  );


  not
  g397
  (
    n161,
    n62
  );


  not
  g398
  (
    n278,
    n108
  );


  not
  g399
  (
    n160,
    n108
  );


  buf
  g400
  (
    n484,
    n45
  );


  not
  g401
  (
    n179,
    n119
  );


  not
  g402
  (
    n547,
    n85
  );


  not
  g403
  (
    n374,
    n103
  );


  buf
  g404
  (
    n440,
    n99
  );


  buf
  g405
  (
    n150,
    n84
  );


  buf
  g406
  (
    n463,
    n105
  );


  not
  g407
  (
    n491,
    n102
  );


  buf
  g408
  (
    n464,
    n49
  );


  buf
  g409
  (
    n541,
    n71
  );


  buf
  g410
  (
    n460,
    n95
  );


  not
  g411
  (
    n445,
    n96
  );


  not
  g412
  (
    n588,
    n85
  );


  buf
  g413
  (
    n393,
    n74
  );


  buf
  g414
  (
    n410,
    n96
  );


  not
  g415
  (
    n582,
    n112
  );


  buf
  g416
  (
    n340,
    n132
  );


  not
  g417
  (
    n519,
    n61
  );


  buf
  g418
  (
    n371,
    n123
  );


  not
  g419
  (
    n341,
    n50
  );


  buf
  g420
  (
    n272,
    n41
  );


  buf
  g421
  (
    n154,
    n33
  );


  not
  g422
  (
    n219,
    n38
  );


  not
  g423
  (
    KeyWire_0_3,
    n53
  );


  not
  g424
  (
    n459,
    n144
  );


  buf
  g425
  (
    n305,
    n126
  );


  not
  g426
  (
    n217,
    n102
  );


  buf
  g427
  (
    n469,
    n55
  );


  buf
  g428
  (
    n294,
    n94
  );


  not
  g429
  (
    n267,
    n54
  );


  buf
  g430
  (
    KeyWire_0_27,
    n53
  );


  buf
  g431
  (
    n264,
    n69
  );


  buf
  g432
  (
    n424,
    n89
  );


  buf
  g433
  (
    n279,
    n119
  );


  buf
  g434
  (
    n336,
    n117
  );


  not
  g435
  (
    n247,
    n53
  );


  buf
  g436
  (
    n153,
    n126
  );


  buf
  g437
  (
    n167,
    n72
  );


  not
  g438
  (
    n315,
    n98
  );


  buf
  g439
  (
    n523,
    n106
  );


  buf
  g440
  (
    n483,
    n61
  );


  buf
  g441
  (
    n535,
    n82
  );


  buf
  g442
  (
    n313,
    n114
  );


  not
  g443
  (
    n449,
    n101
  );


  not
  g444
  (
    n397,
    n122
  );


  not
  g445
  (
    n303,
    n33
  );


  buf
  g446
  (
    n583,
    n145
  );


  buf
  g447
  (
    n175,
    n39
  );


  not
  g448
  (
    n275,
    n141
  );


  buf
  g449
  (
    n200,
    n34
  );


  buf
  g450
  (
    n439,
    n52
  );


  buf
  g451
  (
    n354,
    n47
  );


  buf
  g452
  (
    n490,
    n125
  );


  not
  g453
  (
    n495,
    n56
  );


  buf
  g454
  (
    n156,
    n111
  );


  not
  g455
  (
    n570,
    n138
  );


  buf
  g456
  (
    n556,
    n110
  );


  not
  g457
  (
    KeyWire_0_32,
    n111
  );


  not
  g458
  (
    n162,
    n135
  );


  not
  g459
  (
    n443,
    n104
  );


  not
  g460
  (
    n256,
    n141
  );


  buf
  g461
  (
    n304,
    n93
  );


  buf
  g462
  (
    n297,
    n138
  );


  buf
  g463
  (
    n415,
    n35
  );


  buf
  g464
  (
    n551,
    n118
  );


  buf
  g465
  (
    n197,
    n103
  );


  not
  g466
  (
    n446,
    n53
  );


  buf
  g467
  (
    n365,
    n75
  );


  not
  g468
  (
    n482,
    n101
  );


  not
  g469
  (
    n182,
    n51
  );


  not
  g470
  (
    n504,
    n105
  );


  not
  g471
  (
    n250,
    n35
  );


  not
  g472
  (
    n280,
    n64
  );


  buf
  g473
  (
    n591,
    n80
  );


  not
  g474
  (
    n441,
    n70
  );


  buf
  g475
  (
    n475,
    n79
  );


  buf
  g476
  (
    n172,
    n47
  );


  not
  g477
  (
    n246,
    n136
  );


  not
  g478
  (
    n196,
    n98
  );


  not
  g479
  (
    n358,
    n140
  );


  not
  g480
  (
    n512,
    n115
  );


  not
  g481
  (
    n270,
    n54
  );


  buf
  g482
  (
    n355,
    n91
  );


  not
  g483
  (
    n282,
    n45
  );


  buf
  g484
  (
    n199,
    n77
  );


  buf
  g485
  (
    n306,
    n59
  );


  buf
  g486
  (
    KeyWire_0_56,
    n90
  );


  buf
  g487
  (
    n321,
    n138
  );


  not
  g488
  (
    n159,
    n69
  );


  buf
  g489
  (
    n232,
    n47
  );


  not
  g490
  (
    n206,
    n105
  );


  buf
  g491
  (
    n423,
    n66
  );


  not
  g492
  (
    n562,
    n117
  );


  buf
  g493
  (
    n554,
    n78
  );


  not
  g494
  (
    n426,
    n134
  );


  not
  g495
  (
    n211,
    n119
  );


  buf
  g496
  (
    n249,
    n56
  );


  not
  g497
  (
    n496,
    n100
  );


  not
  g498
  (
    KeyWire_0_20,
    n82
  );


  buf
  g499
  (
    n334,
    n109
  );


  not
  g500
  (
    n527,
    n40
  );


  not
  g501
  (
    n579,
    n94
  );


  not
  g502
  (
    n347,
    n127
  );


  buf
  g503
  (
    n466,
    n136
  );


  not
  g504
  (
    n524,
    n144
  );


  buf
  g505
  (
    n513,
    n67
  );


  buf
  g506
  (
    n544,
    n99
  );


  buf
  g507
  (
    n204,
    n69
  );


  buf
  g508
  (
    n356,
    n90
  );


  buf
  g509
  (
    n295,
    n86
  );


  buf
  g510
  (
    n418,
    n57
  );


  buf
  g511
  (
    n193,
    n77
  );


  buf
  g512
  (
    n164,
    n57
  );


  not
  g513
  (
    n191,
    n63
  );


  not
  g514
  (
    n473,
    n83
  );


  buf
  g515
  (
    n538,
    n63
  );


  buf
  g516
  (
    n216,
    n73
  );


  not
  g517
  (
    n220,
    n63
  );


  not
  g518
  (
    n404,
    n62
  );


  not
  g519
  (
    n218,
    n97
  );


  buf
  g520
  (
    n241,
    n112
  );


  not
  g521
  (
    n260,
    n50
  );


  not
  g522
  (
    n539,
    n93
  );


  buf
  g523
  (
    n385,
    n48
  );


  not
  g524
  (
    n287,
    n93
  );


  not
  g525
  (
    n542,
    n109
  );


  not
  g526
  (
    n593,
    n69
  );


  buf
  g527
  (
    n543,
    n144
  );


  not
  g528
  (
    n574,
    n114
  );


  buf
  g529
  (
    n514,
    n64
  );


  not
  g530
  (
    n323,
    n120
  );


  not
  g531
  (
    n325,
    n117
  );


  buf
  g532
  (
    n471,
    n100
  );


  not
  g533
  (
    n565,
    n44
  );


  not
  g534
  (
    n450,
    n106
  );


  buf
  g535
  (
    n575,
    n84
  );


  not
  g536
  (
    n308,
    n51
  );


  not
  g537
  (
    n309,
    n43
  );


  not
  g538
  (
    n298,
    n115
  );


  buf
  g539
  (
    n350,
    n41
  );


  not
  g540
  (
    n531,
    n52
  );


  buf
  g541
  (
    KeyWire_0_31,
    n120
  );


  not
  g542
  (
    KeyWire_0_60,
    n92
  );


  buf
  g543
  (
    KeyWire_0_21,
    n36
  );


  buf
  g544
  (
    n594,
    n100
  );


  buf
  g545
  (
    n171,
    n131
  );


  not
  g546
  (
    n560,
    n80
  );


  buf
  g547
  (
    n152,
    n55
  );


  buf
  g548
  (
    n166,
    n128
  );


  not
  g549
  (
    n589,
    n127
  );


  not
  g550
  (
    n564,
    n139
  );


  buf
  g551
  (
    n489,
    n98
  );


  not
  g552
  (
    n251,
    n38
  );


  not
  g553
  (
    n312,
    n73
  );


  buf
  g554
  (
    n402,
    n60
  );


  not
  g555
  (
    n578,
    n51
  );


  not
  g556
  (
    n178,
    n129
  );


  buf
  g557
  (
    n480,
    n132
  );


  not
  g558
  (
    n372,
    n100
  );


  not
  g559
  (
    n283,
    n37
  );


  not
  g560
  (
    n584,
    n142
  );


  buf
  g561
  (
    n546,
    n72
  );


  not
  g562
  (
    n529,
    n51
  );


  not
  g563
  (
    n577,
    n88
  );


  not
  g564
  (
    n224,
    n90
  );


  buf
  g565
  (
    n848,
    n521
  );


  buf
  g566
  (
    n666,
    n448
  );


  not
  g567
  (
    n689,
    n481
  );


  buf
  g568
  (
    n767,
    n532
  );


  not
  g569
  (
    n851,
    n308
  );


  buf
  g570
  (
    n825,
    n518
  );


  not
  g571
  (
    n841,
    n247
  );


  not
  g572
  (
    n604,
    n325
  );


  buf
  g573
  (
    n749,
    n443
  );


  not
  g574
  (
    n631,
    n489
  );


  not
  g575
  (
    n691,
    n373
  );


  not
  g576
  (
    n834,
    n294
  );


  buf
  g577
  (
    n678,
    n402
  );


  not
  g578
  (
    n806,
    n451
  );


  buf
  g579
  (
    n667,
    n523
  );


  not
  g580
  (
    n725,
    n337
  );


  buf
  g581
  (
    n776,
    n454
  );


  buf
  g582
  (
    n758,
    n411
  );


  buf
  g583
  (
    n710,
    n248
  );


  buf
  g584
  (
    n813,
    n580
  );


  not
  g585
  (
    n673,
    n169
  );


  not
  g586
  (
    n619,
    n386
  );


  not
  g587
  (
    n621,
    n180
  );


  buf
  g588
  (
    n654,
    n535
  );


  buf
  g589
  (
    n800,
    n342
  );


  buf
  g590
  (
    n646,
    n491
  );


  buf
  g591
  (
    n865,
    n413
  );


  buf
  g592
  (
    n762,
    n539
  );


  buf
  g593
  (
    n761,
    n412
  );


  buf
  g594
  (
    n817,
    n378
  );


  buf
  g595
  (
    n795,
    n536
  );


  buf
  g596
  (
    n665,
    n485
  );


  not
  g597
  (
    n853,
    n447
  );


  not
  g598
  (
    n739,
    n254
  );


  buf
  g599
  (
    n637,
    n165
  );


  not
  g600
  (
    n692,
    n225
  );


  not
  g601
  (
    n858,
    n452
  );


  not
  g602
  (
    n752,
    n170
  );


  not
  g603
  (
    n849,
    n249
  );


  buf
  g604
  (
    n815,
    n334
  );


  not
  g605
  (
    n797,
    n503
  );


  not
  g606
  (
    n741,
    n548
  );


  not
  g607
  (
    n672,
    n502
  );


  not
  g608
  (
    n861,
    n359
  );


  not
  g609
  (
    n636,
    n561
  );


  not
  g610
  (
    n613,
    n528
  );


  buf
  g611
  (
    n660,
    n202
  );


  not
  g612
  (
    n799,
    n301
  );


  buf
  g613
  (
    n863,
    n398
  );


  and
  g614
  (
    n724,
    n446,
    n446,
    n363,
    n428
  );


  and
  g615
  (
    n757,
    n592,
    n524,
    n525,
    n538
  );


  and
  g616
  (
    n742,
    n376,
    n522,
    n534,
    n570
  );


  nor
  g617
  (
    n695,
    n392,
    n242,
    n517,
    n594
  );


  xor
  g618
  (
    n821,
    n526,
    n541,
    n567,
    n568
  );


  nor
  g619
  (
    n791,
    n534,
    n381,
    n516,
    n526
  );


  nand
  g620
  (
    n610,
    n538,
    n527,
    n236,
    n457
  );


  xnor
  g621
  (
    n789,
    n410,
    n589,
    n490,
    n314
  );


  or
  g622
  (
    n830,
    n563,
    n413,
    n213,
    n565
  );


  nand
  g623
  (
    n847,
    n372,
    n403,
    n283,
    n382
  );


  or
  g624
  (
    n671,
    n413,
    n505,
    n412,
    n550
  );


  and
  g625
  (
    n706,
    n548,
    n443,
    n449,
    n467
  );


  xnor
  g626
  (
    n779,
    n485,
    n229,
    n560,
    n431
  );


  and
  g627
  (
    n748,
    n450,
    n384,
    n333,
    n470
  );


  nand
  g628
  (
    n769,
    n424,
    n422,
    n582,
    n437
  );


  and
  g629
  (
    n811,
    n430,
    n411,
    n279,
    n380
  );


  xnor
  g630
  (
    n682,
    n302,
    n158,
    n391,
    n485
  );


  xor
  g631
  (
    n720,
    n597,
    n544,
    n431,
    n595
  );


  xnor
  g632
  (
    n778,
    n472,
    n420,
    n453,
    n538
  );


  xor
  g633
  (
    n722,
    n364,
    n273,
    n430,
    n418
  );


  or
  g634
  (
    n696,
    n583,
    n510,
    n512,
    n435
  );


  nand
  g635
  (
    n755,
    n584,
    n346,
    n403,
    n546
  );


  or
  g636
  (
    n838,
    n255,
    n477,
    n363,
    n434
  );


  xnor
  g637
  (
    n709,
    n292,
    n477,
    n524,
    n508
  );


  and
  g638
  (
    n788,
    n400,
    n423,
    n401,
    n516
  );


  xor
  g639
  (
    n738,
    n467,
    n235,
    n528,
    n265
  );


  nand
  g640
  (
    n836,
    n478,
    n354,
    n544,
    n398
  );


  nand
  g641
  (
    n822,
    n533,
    n351,
    n223,
    n191
  );


  or
  g642
  (
    n701,
    n311,
    n436,
    n495,
    n577
  );


  and
  g643
  (
    n625,
    n399,
    n488,
    n272,
    n552
  );


  nor
  g644
  (
    n772,
    n467,
    n581,
    n440,
    n408
  );


  or
  g645
  (
    n611,
    n375,
    n460,
    n281,
    n483
  );


  and
  g646
  (
    n831,
    n465,
    n562,
    n419,
    n585
  );


  or
  g647
  (
    n774,
    n568,
    n385,
    n591,
    n536
  );


  nand
  g648
  (
    n714,
    n231,
    n371,
    n457,
    n427
  );


  and
  g649
  (
    n649,
    n198,
    n388,
    n465,
    n470
  );


  xnor
  g650
  (
    n786,
    n529,
    n237,
    n564,
    n498
  );


  xor
  g651
  (
    n867,
    n483,
    n457,
    n446,
    n539
  );


  nor
  g652
  (
    n780,
    n527,
    n462,
    n415,
    n572
  );


  nand
  g653
  (
    n644,
    n358,
    n366,
    n452,
    n176
  );


  xor
  g654
  (
    n693,
    n556,
    n551,
    n428,
    n208
  );


  nand
  g655
  (
    n614,
    n511,
    n427,
    n487,
    n445
  );


  nor
  g656
  (
    n728,
    n296,
    n554,
    n375,
    n374
  );


  xnor
  g657
  (
    n603,
    n407,
    n271,
    n575,
    n186
  );


  nor
  g658
  (
    n763,
    n518,
    n305,
    n406,
    n567
  );


  xnor
  g659
  (
    n810,
    n432,
    n363,
    n257,
    n531
  );


  xor
  g660
  (
    KeyWire_0_26,
    n456,
    n396,
    n569,
    n575
  );


  xor
  g661
  (
    n743,
    n462,
    n268,
    n403,
    n570
  );


  xnor
  g662
  (
    KeyWire_0_63,
    n437,
    n444,
    n439,
    n420
  );


  xor
  g663
  (
    n681,
    n150,
    n415,
    n431,
    n356
  );


  and
  g664
  (
    n796,
    n417,
    n527,
    n164,
    n151
  );


  nor
  g665
  (
    n801,
    n264,
    n239,
    n352,
    n541
  );


  xor
  g666
  (
    n814,
    n537,
    n160,
    n435,
    n194
  );


  xnor
  g667
  (
    n664,
    n577,
    n559,
    n553,
    n387
  );


  or
  g668
  (
    n686,
    n477,
    n190,
    n393,
    n316
  );


  xnor
  g669
  (
    n860,
    n471,
    n541,
    n588,
    n286
  );


  and
  g670
  (
    n870,
    n453,
    n369,
    n379,
    n559
  );


  and
  g671
  (
    n775,
    n370,
    n378,
    n358,
    n591
  );


  nor
  g672
  (
    n804,
    n396,
    n569,
    n503,
    n590
  );


  xor
  g673
  (
    n617,
    n442,
    n354,
    n455,
    n581
  );


  or
  g674
  (
    n837,
    n429,
    n298,
    n529,
    n444
  );


  xnor
  g675
  (
    n598,
    n390,
    n368,
    n187,
    n497
  );


  xnor
  g676
  (
    n600,
    n495,
    n412,
    n270,
    n480
  );


  and
  g677
  (
    n717,
    n297,
    n377,
    n391,
    n367
  );


  xnor
  g678
  (
    n856,
    n590,
    n530,
    n499,
    n468
  );


  and
  g679
  (
    n805,
    n583,
    n354,
    n300,
    n593
  );


  nor
  g680
  (
    n684,
    n494,
    n310,
    n388,
    n461
  );


  and
  g681
  (
    n773,
    n212,
    n193,
    n352,
    n304
  );


  or
  g682
  (
    n793,
    n378,
    n253,
    n536,
    n433
  );


  xnor
  g683
  (
    n819,
    n463,
    n513,
    n260,
    n555
  );


  and
  g684
  (
    n826,
    n584,
    n371,
    n571,
    n537
  );


  xnor
  g685
  (
    n615,
    n449,
    n447,
    n383,
    n454
  );


  xor
  g686
  (
    n612,
    n479,
    n459,
    n390,
    n402
  );


  and
  g687
  (
    n705,
    n492,
    n463,
    n379,
    n423
  );


  nor
  g688
  (
    n658,
    n359,
    n321,
    n409,
    n175
  );


  and
  g689
  (
    n608,
    n507,
    n519,
    n544,
    n545
  );


  nor
  g690
  (
    n833,
    n441,
    n329,
    n153,
    n426
  );


  and
  g691
  (
    n662,
    n266,
    n240,
    n430,
    n578
  );


  or
  g692
  (
    n818,
    n357,
    n280,
    n543,
    n293
  );


  xnor
  g693
  (
    n781,
    n370,
    n375,
    n471,
    n540
  );


  nor
  g694
  (
    n629,
    n458,
    n489,
    n513,
    n576
  );


  nor
  g695
  (
    n694,
    n493,
    n514,
    n560,
    n422
  );


  xnor
  g696
  (
    n744,
    n207,
    n483,
    n174,
    n539
  );


  xnor
  g697
  (
    n816,
    n550,
    n552,
    n205,
    n400
  );


  xor
  g698
  (
    n711,
    n585,
    n418,
    n508,
    n480
  );


  xor
  g699
  (
    n634,
    n155,
    n557,
    n416,
    n425
  );


  nand
  g700
  (
    n783,
    n562,
    n197,
    n557,
    n409
  );


  nor
  g701
  (
    n768,
    n380,
    n443,
    n488,
    n276
  );


  xnor
  g702
  (
    n820,
    n473,
    n576,
    n475,
    n595
  );


  xor
  g703
  (
    n765,
    n499,
    n501,
    n303,
    n525
  );


  nand
  g704
  (
    n707,
    n177,
    n509,
    n404,
    n389
  );


  and
  g705
  (
    n845,
    n222,
    n515,
    n463,
    n360
  );


  nor
  g706
  (
    n754,
    n377,
    n407,
    n394,
    n379
  );


  xor
  g707
  (
    KeyWire_0_0,
    n401,
    n263,
    n374,
    n385
  );


  xor
  g708
  (
    n771,
    n184,
    n196,
    n238,
    n505
  );


  nand
  g709
  (
    n657,
    n432,
    n597,
    n458,
    n404
  );


  xnor
  g710
  (
    n623,
    n486,
    n494,
    n466,
    n358
  );


  and
  g711
  (
    n756,
    n396,
    n330,
    n596,
    n484
  );


  and
  g712
  (
    n843,
    n387,
    n448,
    n491,
    n521
  );


  nor
  g713
  (
    n835,
    n414,
    n324,
    n469,
    n384
  );


  xor
  g714
  (
    n651,
    n227,
    n547,
    n560,
    n555
  );


  nand
  g715
  (
    n683,
    n586,
    n434,
    n159,
    n183
  );


  nor
  g716
  (
    n713,
    n381,
    n335,
    n549,
    n554
  );


  xor
  g717
  (
    n659,
    n441,
    n464,
    n520,
    n148
  );


  nor
  g718
  (
    n864,
    n451,
    n573,
    n361,
    n582
  );


  nand
  g719
  (
    n626,
    n385,
    n390,
    n299,
    n362
  );


  or
  g720
  (
    n620,
    n199,
    n368,
    n408,
    n543
  );


  xnor
  g721
  (
    n868,
    n478,
    n377,
    n315,
    n251
  );


  xnor
  g722
  (
    n812,
    n429,
    n459,
    n274,
    n449
  );


  nor
  g723
  (
    n855,
    n345,
    n542,
    n350,
    n461
  );


  xor
  g724
  (
    n745,
    n547,
    n450,
    n585,
    n448
  );


  nand
  g725
  (
    n842,
    n306,
    n501,
    n285,
    n493
  );


  xnor
  g726
  (
    n854,
    n574,
    n168,
    n405,
    n482
  );


  xor
  g727
  (
    n648,
    n427,
    n566,
    n502,
    n512
  );


  nand
  g728
  (
    n829,
    n556,
    n474,
    n558,
    n521
  );


  and
  g729
  (
    n869,
    n152,
    n291,
    n267,
    n438
  );


  nand
  g730
  (
    n700,
    n484,
    n574,
    n421,
    n593
  );


  or
  g731
  (
    n787,
    n579,
    n171,
    n526,
    n204
  );


  or
  g732
  (
    n723,
    n423,
    n219,
    n371,
    n232
  );


  xnor
  g733
  (
    n712,
    n319,
    n275,
    n156,
    n466
  );


  nand
  g734
  (
    n699,
    n578,
    n497,
    n341,
    n573
  );


  or
  g735
  (
    n716,
    n438,
    n313,
    n386
  );


  xnor
  g736
  (
    n798,
    n250,
    n566,
    n252,
    n593
  );


  xnor
  g737
  (
    n753,
    n399,
    n484,
    n211,
    n410
  );


  xnor
  g738
  (
    n729,
    n440,
    n161,
    n520,
    n492
  );


  or
  g739
  (
    n703,
    n570,
    n209,
    n464,
    n417
  );


  xnor
  g740
  (
    n747,
    n571,
    n382,
    n393,
    n479
  );


  and
  g741
  (
    n827,
    n259,
    n589,
    n349,
    n534
  );


  xor
  g742
  (
    n764,
    n556,
    n424,
    n328,
    n157
  );


  nor
  g743
  (
    n866,
    n535,
    n586,
    n439,
    n517
  );


  and
  g744
  (
    n857,
    n374,
    n478,
    n332,
    n344
  );


  or
  g745
  (
    n688,
    n317,
    n203,
    n542,
    n234
  );


  and
  g746
  (
    n808,
    n482,
    n307,
    n498,
    n506
  );


  nand
  g747
  (
    n839,
    n529,
    n380,
    n465,
    n482
  );


  or
  g748
  (
    n677,
    n309,
    n530,
    n583,
    n426
  );


  nand
  g749
  (
    n785,
    n517,
    n533,
    n587,
    n258
  );


  and
  g750
  (
    n828,
    n395,
    n434,
    n528,
    n438
  );


  nor
  g751
  (
    n790,
    n473,
    n588,
    n246,
    n551
  );


  nor
  g752
  (
    n802,
    n553,
    n573,
    n486,
    n511
  );


  and
  g753
  (
    n645,
    n469,
    n577,
    n437,
    n474
  );


  or
  g754
  (
    n630,
    n489,
    n532,
    n419,
    n504
  );


  and
  g755
  (
    n731,
    n210,
    n361,
    n288,
    n578
  );


  xor
  g756
  (
    n633,
    n545,
    n564,
    n505,
    n163
  );


  xor
  g757
  (
    n674,
    n523,
    n405,
    n406,
    n565
  );


  xnor
  g758
  (
    n668,
    n394,
    n594,
    n456,
    n490
  );


  xor
  g759
  (
    n840,
    n497,
    n326,
    n581,
    n500
  );


  nand
  g760
  (
    n675,
    n422,
    n468,
    n353,
    n499
  );


  nand
  g761
  (
    n599,
    n269,
    n508,
    n359,
    n383
  );


  nand
  g762
  (
    n846,
    n318,
    n414,
    n531,
    n256
  );


  xnor
  g763
  (
    n832,
    n189,
    n574,
    n480,
    n503
  );


  xor
  g764
  (
    n809,
    n532,
    n473,
    n347,
    n546
  );


  xnor
  g765
  (
    n792,
    n504,
    n516,
    n243,
    n492
  );


  nor
  g766
  (
    n777,
    n429,
    n502,
    n185,
    n220
  );


  xnor
  g767
  (
    n607,
    n425,
    n356,
    n444,
    n388
  );


  xor
  g768
  (
    n702,
    n373,
    n436,
    n421,
    n355
  );


  or
  g769
  (
    n679,
    n481,
    n496,
    n525,
    n394
  );


  xor
  g770
  (
    n803,
    n450,
    n355,
    n523,
    n233
  );


  and
  g771
  (
    n751,
    n384,
    n506,
    n559,
    n230
  );


  nand
  g772
  (
    n844,
    n566,
    n472,
    n389,
    n590
  );


  nor
  g773
  (
    n642,
    n182,
    n571,
    n441,
    n244
  );


  and
  g774
  (
    n655,
    n367,
    n487,
    n558,
    n549
  );


  or
  g775
  (
    n737,
    n552,
    n512,
    n500,
    n216
  );


  and
  g776
  (
    n647,
    n224,
    n245,
    n365,
    n589
  );


  and
  g777
  (
    n632,
    n587,
    n392,
    n547,
    n462
  );


  nor
  g778
  (
    n734,
    n493,
    n511,
    n456,
    n166
  );


  or
  g779
  (
    n622,
    n540,
    n594,
    n537,
    n392
  );


  nand
  g780
  (
    n641,
    n565,
    n460,
    n351,
    n218
  );


  or
  g781
  (
    n643,
    n436,
    n543,
    n355,
    n356
  );


  xnor
  g782
  (
    n697,
    n509,
    n579,
    n339,
    n360
  );


  nand
  g783
  (
    n661,
    n553,
    n452,
    n432,
    n470
  );


  nor
  g784
  (
    n606,
    n535,
    n555,
    n393,
    n428
  );


  xnor
  g785
  (
    n746,
    n201,
    n458,
    n278,
    n439
  );


  and
  g786
  (
    n730,
    n391,
    n200,
    n596,
    n495
  );


  and
  g787
  (
    n605,
    n228,
    n322,
    n469,
    n466
  );


  nor
  g788
  (
    n823,
    n343,
    n383,
    n595,
    n221
  );


  or
  g789
  (
    n676,
    n416,
    n445,
    n460,
    n282
  );


  nand
  g790
  (
    n627,
    n592,
    n364,
    n348,
    n564
  );


  xor
  g791
  (
    n718,
    n472,
    n395,
    n414,
    n411
  );


  or
  g792
  (
    n794,
    n471,
    n580,
    n389,
    n241
  );


  nand
  g793
  (
    n624,
    n447,
    n408,
    n365,
    n284
  );


  and
  g794
  (
    n638,
    n365,
    n362,
    n476,
    n442
  );


  nand
  g795
  (
    n687,
    n353,
    n475,
    n504,
    n481
  );


  nor
  g796
  (
    n708,
    n376,
    n453,
    n588,
    n531
  );


  nand
  g797
  (
    n721,
    n507,
    n597,
    n217,
    n382
  );


  or
  g798
  (
    n807,
    n558,
    n178,
    n400,
    n188
  );


  and
  g799
  (
    n736,
    n206,
    n367,
    n533,
    n515
  );


  nand
  g800
  (
    n704,
    n518,
    n490,
    n474,
    n501
  );


  nor
  g801
  (
    n656,
    n522,
    n510,
    n407,
    n459
  );


  and
  g802
  (
    n685,
    n561,
    n401,
    n320,
    n586
  );


  nand
  g803
  (
    n727,
    n398,
    n154,
    n451,
    n486
  );


  and
  g804
  (
    n733,
    n506,
    n562,
    n419,
    n417
  );


  nor
  g805
  (
    n635,
    n338,
    n500,
    n361,
    n399
  );


  nand
  g806
  (
    n715,
    n397,
    n406,
    n426,
    n277
  );


  xnor
  g807
  (
    n750,
    n476,
    n494,
    n563,
    n510
  );


  xor
  g808
  (
    n670,
    n487,
    n353,
    n519,
    n425
  );


  or
  g809
  (
    n618,
    n545,
    n455,
    n352,
    n395
  );


  xnor
  g810
  (
    n652,
    n587,
    n418,
    n520,
    n369
  );


  xnor
  g811
  (
    n719,
    n387,
    n323,
    n496,
    n287
  );


  and
  g812
  (
    n663,
    n445,
    n563,
    n397,
    n366
  );


  or
  g813
  (
    n669,
    n491,
    n515,
    n579,
    n226
  );


  xor
  g814
  (
    n824,
    n468,
    n568,
    n475,
    n179
  );


  nor
  g815
  (
    n784,
    n327,
    n554,
    n369,
    n340
  );


  xor
  g816
  (
    n770,
    n397,
    n370,
    n368,
    n488
  );


  nor
  g817
  (
    n735,
    n421,
    n567,
    n455,
    n214
  );


  or
  g818
  (
    n859,
    n433,
    n454,
    n295,
    n357
  );


  or
  g819
  (
    n852,
    n336,
    n498,
    n167,
    n351
  );


  xnor
  g820
  (
    n698,
    n173,
    n181,
    n591,
    n360
  );


  xor
  g821
  (
    n850,
    n435,
    n376,
    n366,
    n542
  );


  nand
  g822
  (
    n650,
    n215,
    n550,
    n557,
    n514
  );


  nor
  g823
  (
    n653,
    n476,
    n548,
    n192,
    n172
  );


  or
  g824
  (
    n740,
    n596,
    n572,
    n540,
    n561
  );


  and
  g825
  (
    n759,
    n364,
    n546,
    n530,
    n402
  );


  or
  g826
  (
    n862,
    n575,
    n357,
    n551,
    n461
  );


  xor
  g827
  (
    n726,
    n513,
    n312,
    n147,
    n524
  );


  xnor
  g828
  (
    n760,
    n442,
    n372,
    n405,
    n424
  );


  xor
  g829
  (
    n732,
    n592,
    n464,
    n373,
    n409
  );


  xor
  g830
  (
    n766,
    n522,
    n519,
    n149,
    n381
  );


  xnor
  g831
  (
    n628,
    n507,
    n290,
    n582,
    n162
  );


  and
  g832
  (
    n602,
    n195,
    n514,
    n549,
    n479
  );


  xor
  g833
  (
    n640,
    n569,
    n496,
    n576,
    n509
  );


  or
  g834
  (
    n609,
    n372,
    n261,
    n415,
    n331
  );


  nand
  g835
  (
    n616,
    n262,
    n433,
    n362,
    n420
  );


  nand
  g836
  (
    n601,
    n404,
    n572,
    n580,
    n410
  );


  xor
  g837
  (
    n680,
    n440,
    n584,
    n289,
    n416
  );


  buf
  g838
  (
    n871,
    n614
  );


  not
  g839
  (
    n897,
    n604
  );


  buf
  g840
  (
    n872,
    n598
  );


  buf
  g841
  (
    n898,
    n610
  );


  buf
  g842
  (
    n883,
    n603
  );


  buf
  g843
  (
    n879,
    n621
  );


  buf
  g844
  (
    n878,
    n609
  );


  not
  g845
  (
    n887,
    n624
  );


  not
  g846
  (
    n873,
    n613
  );


  buf
  g847
  (
    n874,
    n601
  );


  not
  g848
  (
    n888,
    n619
  );


  buf
  g849
  (
    n886,
    n616
  );


  buf
  g850
  (
    n884,
    n615
  );


  not
  g851
  (
    n877,
    n625
  );


  not
  g852
  (
    n894,
    n620
  );


  not
  g853
  (
    n882,
    n599
  );


  buf
  g854
  (
    n893,
    n605
  );


  not
  g855
  (
    n889,
    n611
  );


  buf
  g856
  (
    n892,
    n606
  );


  not
  g857
  (
    n875,
    n600
  );


  not
  g858
  (
    n895,
    n612
  );


  buf
  g859
  (
    n881,
    n617
  );


  buf
  g860
  (
    n890,
    n618
  );


  not
  g861
  (
    n885,
    n623
  );


  not
  g862
  (
    n880,
    n608
  );


  not
  g863
  (
    n876,
    n607
  );


  not
  g864
  (
    KeyWire_0_38,
    n602
  );


  buf
  g865
  (
    n891,
    n622
  );


  not
  g866
  (
    n919,
    n890
  );


  not
  g867
  (
    n900,
    n887
  );


  not
  g868
  (
    n936,
    n889
  );


  not
  g869
  (
    n908,
    n884
  );


  not
  g870
  (
    n921,
    n888
  );


  buf
  g871
  (
    n934,
    n871
  );


  not
  g872
  (
    n915,
    n880
  );


  not
  g873
  (
    n918,
    n883
  );


  buf
  g874
  (
    n925,
    n877
  );


  not
  g875
  (
    n903,
    n881
  );


  not
  g876
  (
    n937,
    n874
  );


  not
  g877
  (
    n923,
    n888
  );


  not
  g878
  (
    n902,
    n897
  );


  not
  g879
  (
    n924,
    n882
  );


  buf
  g880
  (
    n939,
    n891
  );


  buf
  g881
  (
    n938,
    n885
  );


  buf
  g882
  (
    n935,
    n881
  );


  buf
  g883
  (
    n901,
    n872
  );


  buf
  g884
  (
    n912,
    n890
  );


  buf
  g885
  (
    n917,
    n884
  );


  buf
  g886
  (
    n945,
    n895
  );


  buf
  g887
  (
    n929,
    n889
  );


  buf
  g888
  (
    n920,
    n896
  );


  not
  g889
  (
    n932,
    n883
  );


  buf
  g890
  (
    n944,
    n893
  );


  buf
  g891
  (
    n941,
    n887
  );


  not
  g892
  (
    n904,
    n895
  );


  not
  g893
  (
    n899,
    n875
  );


  not
  g894
  (
    n913,
    n879
  );


  buf
  g895
  (
    n907,
    n894
  );


  not
  g896
  (
    n922,
    n878
  );


  not
  g897
  (
    n926,
    n878
  );


  buf
  g898
  (
    n909,
    n882
  );


  buf
  g899
  (
    n930,
    n885
  );


  buf
  g900
  (
    n946,
    n894
  );


  buf
  g901
  (
    n931,
    n879
  );


  not
  g902
  (
    n940,
    n877
  );


  buf
  g903
  (
    n910,
    n891
  );


  buf
  g904
  (
    n943,
    n880
  );


  buf
  g905
  (
    n933,
    n876
  );


  not
  g906
  (
    n942,
    n896
  );


  buf
  g907
  (
    n916,
    n886
  );


  buf
  g908
  (
    n906,
    n873
  );


  not
  g909
  (
    n927,
    n886
  );


  not
  g910
  (
    n928,
    n892
  );


  buf
  g911
  (
    n905,
    n897
  );


  buf
  g912
  (
    n911,
    n893
  );


  not
  g913
  (
    n914,
    n892
  );


  not
  g914
  (
    n1020,
    n934
  );


  not
  g915
  (
    n960,
    n932
  );


  not
  g916
  (
    n1002,
    n925
  );


  buf
  g917
  (
    n1041,
    n932
  );


  buf
  g918
  (
    n1004,
    n910
  );


  not
  g919
  (
    n1050,
    n935
  );


  not
  g920
  (
    n989,
    n934
  );


  not
  g921
  (
    n953,
    n918
  );


  not
  g922
  (
    n1027,
    n925
  );


  buf
  g923
  (
    n976,
    n916
  );


  not
  g924
  (
    n972,
    n899
  );


  not
  g925
  (
    n1084,
    n905
  );


  buf
  g926
  (
    n1066,
    n920
  );


  not
  g927
  (
    n949,
    n911
  );


  buf
  g928
  (
    n1063,
    n908
  );


  not
  g929
  (
    n969,
    n912
  );


  not
  g930
  (
    n967,
    n928
  );


  not
  g931
  (
    n964,
    n904
  );


  buf
  g932
  (
    n965,
    n933
  );


  not
  g933
  (
    n958,
    n908
  );


  not
  g934
  (
    n1012,
    n925
  );


  not
  g935
  (
    n1053,
    n927
  );


  buf
  g936
  (
    n1057,
    n909
  );


  not
  g937
  (
    n1052,
    n937
  );


  buf
  g938
  (
    n1061,
    n921
  );


  buf
  g939
  (
    n1043,
    n928
  );


  not
  g940
  (
    n1013,
    n901
  );


  not
  g941
  (
    n978,
    n933
  );


  buf
  g942
  (
    n1074,
    n906
  );


  not
  g943
  (
    n1068,
    n900
  );


  buf
  g944
  (
    n1036,
    n937
  );


  not
  g945
  (
    n1062,
    n921
  );


  not
  g946
  (
    n1016,
    n918
  );


  buf
  g947
  (
    n1009,
    n913
  );


  buf
  g948
  (
    KeyWire_0_36,
    n922
  );


  buf
  g949
  (
    n981,
    n923
  );


  buf
  g950
  (
    n1045,
    n915
  );


  buf
  g951
  (
    n1003,
    n920
  );


  buf
  g952
  (
    n1007,
    n920
  );


  buf
  g953
  (
    KeyWire_0_4,
    n902
  );


  buf
  g954
  (
    n957,
    n901
  );


  buf
  g955
  (
    n948,
    n936
  );


  not
  g956
  (
    n1011,
    n918
  );


  not
  g957
  (
    n1025,
    n926
  );


  not
  g958
  (
    n970,
    n901
  );


  buf
  g959
  (
    n988,
    n932
  );


  buf
  g960
  (
    n959,
    n930
  );


  buf
  g961
  (
    n1046,
    n931
  );


  buf
  g962
  (
    KeyWire_0_57,
    n907
  );


  buf
  g963
  (
    n985,
    n931
  );


  buf
  g964
  (
    n1081,
    n919
  );


  not
  g965
  (
    n1021,
    n914
  );


  buf
  g966
  (
    n950,
    n922
  );


  buf
  g967
  (
    n1071,
    n923
  );


  buf
  g968
  (
    n1024,
    n936
  );


  not
  g969
  (
    n1047,
    n929
  );


  not
  g970
  (
    n995,
    n916
  );


  not
  g971
  (
    n974,
    n918
  );


  buf
  g972
  (
    n986,
    n921
  );


  not
  g973
  (
    n968,
    n902
  );


  not
  g974
  (
    n1055,
    n917
  );


  not
  g975
  (
    n954,
    n927
  );


  not
  g976
  (
    n1006,
    n915
  );


  buf
  g977
  (
    n1001,
    n936
  );


  buf
  g978
  (
    n1070,
    n935
  );


  buf
  g979
  (
    n987,
    n914
  );


  buf
  g980
  (
    n1019,
    n926
  );


  buf
  g981
  (
    n1073,
    n903
  );


  not
  g982
  (
    n952,
    n911
  );


  not
  g983
  (
    n980,
    n928
  );


  not
  g984
  (
    n997,
    n902
  );


  not
  g985
  (
    n1014,
    n914
  );


  buf
  g986
  (
    n966,
    n904
  );


  buf
  g987
  (
    n975,
    n907
  );


  buf
  g988
  (
    KeyWire_0_13,
    n930
  );


  buf
  g989
  (
    n1075,
    n929
  );


  buf
  g990
  (
    n971,
    n915
  );


  buf
  g991
  (
    n977,
    n930
  );


  buf
  g992
  (
    n1072,
    n909
  );


  not
  g993
  (
    n1065,
    n905
  );


  not
  g994
  (
    n1067,
    n912
  );


  not
  g995
  (
    n1026,
    n916
  );


  not
  g996
  (
    n983,
    n919
  );


  not
  g997
  (
    n1040,
    n930
  );


  buf
  g998
  (
    KeyWire_0_49,
    n924
  );


  not
  g999
  (
    n1082,
    n929
  );


  not
  g1000
  (
    n994,
    n905
  );


  buf
  g1001
  (
    n951,
    n903
  );


  not
  g1002
  (
    n992,
    n926
  );


  not
  g1003
  (
    n973,
    n934
  );


  not
  g1004
  (
    KeyWire_0_43,
    n913
  );


  not
  g1005
  (
    n956,
    n924
  );


  buf
  g1006
  (
    n991,
    n923
  );


  buf
  g1007
  (
    n1058,
    n923
  );


  buf
  g1008
  (
    n1015,
    n903
  );


  buf
  g1009
  (
    n1042,
    n907
  );


  not
  g1010
  (
    n955,
    n929
  );


  not
  g1011
  (
    n1083,
    n922
  );


  buf
  g1012
  (
    KeyWire_0_23,
    n933
  );


  not
  g1013
  (
    n1054,
    n931
  );


  not
  g1014
  (
    KeyWire_0_41,
    n900
  );


  buf
  g1015
  (
    n979,
    n916
  );


  buf
  g1016
  (
    n982,
    n900
  );


  buf
  g1017
  (
    n1010,
    n919
  );


  not
  g1018
  (
    n1038,
    n935
  );


  not
  g1019
  (
    n1037,
    n908
  );


  buf
  g1020
  (
    KeyWire_0_15,
    n931
  );


  buf
  g1021
  (
    n1017,
    n924
  );


  not
  g1022
  (
    n1044,
    n932
  );


  buf
  g1023
  (
    n1008,
    n899
  );


  not
  g1024
  (
    n1033,
    n910
  );


  not
  g1025
  (
    n996,
    n910
  );


  buf
  g1026
  (
    n1018,
    n925
  );


  buf
  g1027
  (
    n1000,
    n904
  );


  buf
  g1028
  (
    n963,
    n937
  );


  not
  g1029
  (
    n1030,
    n936
  );


  buf
  g1030
  (
    n984,
    n917
  );


  buf
  g1031
  (
    n1080,
    n917
  );


  not
  g1032
  (
    n1049,
    n935
  );


  not
  g1033
  (
    n1076,
    n927
  );


  buf
  g1034
  (
    n1060,
    n926
  );


  not
  g1035
  (
    n962,
    n906
  );


  buf
  g1036
  (
    n1032,
    n909
  );


  buf
  g1037
  (
    n1028,
    n906
  );


  not
  g1038
  (
    n1077,
    n921
  );


  buf
  g1039
  (
    n1022,
    n911
  );


  not
  g1040
  (
    n993,
    n924
  );


  buf
  g1041
  (
    n1056,
    n912
  );


  not
  g1042
  (
    n1048,
    n913
  );


  buf
  g1043
  (
    n961,
    n920
  );


  not
  g1044
  (
    n1029,
    n919
  );


  not
  g1045
  (
    n1034,
    n927
  );


  not
  g1046
  (
    n1039,
    n933
  );


  buf
  g1047
  (
    n1051,
    n917
  );


  buf
  g1048
  (
    n947,
    n922
  );


  not
  g1049
  (
    n1023,
    n934
  );


  not
  g1050
  (
    n1064,
    n928
  );


  not
  g1051
  (
    n1005,
    n899
  );


  xor
  g1052
  (
    n1086,
    n635,
    n699,
    n956,
    n701
  );


  and
  g1053
  (
    n1089,
    n709,
    n637,
    n688,
    n650
  );


  or
  g1054
  (
    n1122,
    n713,
    n989,
    n655,
    n693
  );


  xor
  g1055
  (
    n1102,
    n669,
    n715,
    n653,
    n960
  );


  and
  g1056
  (
    n1098,
    n950,
    n986,
    n741,
    n983
  );


  xor
  g1057
  (
    n1085,
    n979,
    n672,
    n959,
    n726
  );


  xor
  g1058
  (
    n1104,
    n628,
    n740,
    n642,
    n717
  );


  nor
  g1059
  (
    n1108,
    n953,
    n649,
    n657,
    n630
  );


  nor
  g1060
  (
    n1105,
    n640,
    n962,
    n984,
    n739
  );


  or
  g1061
  (
    n1118,
    n690,
    n676,
    n694,
    n711
  );


  or
  g1062
  (
    n1096,
    n728,
    n719,
    n948,
    n660
  );


  nor
  g1063
  (
    n1097,
    n667,
    n712,
    n662,
    n966
  );


  nor
  g1064
  (
    n1099,
    n663,
    n968,
    n696,
    n648
  );


  and
  g1065
  (
    n1116,
    n703,
    n702,
    n656,
    n951
  );


  xor
  g1066
  (
    n1124,
    n666,
    n691,
    n737,
    n722
  );


  nor
  g1067
  (
    n1088,
    n949,
    n671,
    n714,
    n980
  );


  or
  g1068
  (
    n1101,
    n705,
    n684,
    n708,
    n718
  );


  xor
  g1069
  (
    n1109,
    n632,
    n668,
    n686,
    n981
  );


  nor
  g1070
  (
    n1120,
    n678,
    n674,
    n698,
    n689
  );


  xnor
  g1071
  (
    n1113,
    n629,
    n990,
    n679,
    n700
  );


  xnor
  g1072
  (
    n1107,
    n704,
    n736,
    n735,
    n724
  );


  xnor
  g1073
  (
    n1119,
    n692,
    n720,
    n947,
    n634
  );


  or
  g1074
  (
    n1103,
    n627,
    n727,
    n961,
    n658
  );


  xor
  g1075
  (
    n1093,
    n977,
    n978,
    n639,
    n738
  );


  and
  g1076
  (
    n1111,
    n647,
    n644,
    n665,
    n652
  );


  xnor
  g1077
  (
    n1090,
    n971,
    n988,
    n670,
    n682
  );


  nand
  g1078
  (
    n1106,
    n641,
    n952,
    n731,
    n976
  );


  and
  g1079
  (
    n1114,
    n973,
    n673,
    n710,
    n957
  );


  xor
  g1080
  (
    n1094,
    n683,
    n729,
    n958,
    n967
  );


  nand
  g1081
  (
    n1121,
    n645,
    n636,
    n685,
    n733
  );


  and
  g1082
  (
    n1092,
    n638,
    n730,
    n964,
    n646
  );


  nand
  g1083
  (
    n1112,
    n985,
    n721,
    n955,
    n677
  );


  and
  g1084
  (
    n1095,
    n633,
    n969,
    n659,
    n631
  );


  xor
  g1085
  (
    n1087,
    n695,
    n725,
    n716,
    n626
  );


  xnor
  g1086
  (
    n1110,
    n664,
    n706,
    n643,
    n972
  );


  xor
  g1087
  (
    n1100,
    n675,
    n661,
    n723,
    n697
  );


  or
  g1088
  (
    n1123,
    n680,
    n687,
    n654,
    n651
  );


  xor
  g1089
  (
    n1117,
    n963,
    n954,
    n681,
    n975
  );


  or
  g1090
  (
    n1091,
    n732,
    n734,
    n974,
    n707
  );


  xnor
  g1091
  (
    n1115,
    n970,
    n982,
    n965,
    n987
  );


  buf
  g1092
  (
    n1131,
    n1091
  );


  buf
  g1093
  (
    n1125,
    n1088
  );


  not
  g1094
  (
    n1133,
    n1090
  );


  buf
  g1095
  (
    n1127,
    n1087
  );


  buf
  g1096
  (
    n1130,
    n1089
  );


  not
  g1097
  (
    n1129,
    n1094
  );


  not
  g1098
  (
    n1128,
    n1092
  );


  not
  g1099
  (
    n1134,
    n1093
  );


  buf
  g1100
  (
    n1126,
    n1085
  );


  buf
  g1101
  (
    n1132,
    n1086
  );


  buf
  g1102
  (
    n1150,
    n1125
  );


  not
  g1103
  (
    n1140,
    n938
  );


  buf
  g1104
  (
    n1146,
    n1129
  );


  not
  g1105
  (
    n1136,
    n1125
  );


  not
  g1106
  (
    n1145,
    n1127
  );


  buf
  g1107
  (
    n1147,
    n1128
  );


  not
  g1108
  (
    n1148,
    n1129
  );


  not
  g1109
  (
    n1144,
    n1126
  );


  not
  g1110
  (
    n1135,
    n938
  );


  not
  g1111
  (
    n1152,
    n1125
  );


  buf
  g1112
  (
    n1138,
    n1127
  );


  buf
  g1113
  (
    n1142,
    n1126
  );


  not
  g1114
  (
    n1143,
    n938
  );


  buf
  g1115
  (
    n1149,
    n1125
  );


  buf
  g1116
  (
    n1137,
    n1128
  );


  buf
  g1117
  (
    n1153,
    n1128
  );


  buf
  g1118
  (
    n1139,
    n1126
  );


  nor
  g1119
  (
    n1151,
    n938,
    n1127,
    n1129
  );


  nor
  g1120
  (
    n1141,
    n1127,
    n1126,
    n937,
    n1128
  );


  nor
  g1121
  (
    n1159,
    n993,
    n1048,
    n1054,
    n1042
  );


  or
  g1122
  (
    n1155,
    n1136,
    n1057,
    n1054,
    n1016
  );


  nand
  g1123
  (
    n1163,
    n1138,
    n1004,
    n1139,
    n997
  );


  nor
  g1124
  (
    n1170,
    n1138,
    n1137,
    n1043,
    n998
  );


  nand
  g1125
  (
    n1165,
    n1055,
    n1139,
    n1012,
    n1030
  );


  and
  g1126
  (
    n1171,
    n1000,
    n996,
    n1053,
    n1024
  );


  and
  g1127
  (
    KeyWire_0_7,
    n1015,
    n1058,
    n1140,
    n1007
  );


  xnor
  g1128
  (
    n1173,
    n1029,
    n1139,
    n1141,
    n1020
  );


  or
  g1129
  (
    n1161,
    n1002,
    n1140,
    n1135,
    n1059
  );


  or
  g1130
  (
    n1179,
    n1035,
    n1013,
    n1038,
    n1045
  );


  or
  g1131
  (
    n1160,
    n1058,
    n1017,
    n1008,
    n1055
  );


  and
  g1132
  (
    n1164,
    n1142,
    n1010,
    n1141,
    n999
  );


  or
  g1133
  (
    n1169,
    n1019,
    n1136,
    n1039,
    n1009
  );


  nand
  g1134
  (
    n1154,
    n1057,
    n1011,
    n1050,
    n1036
  );


  xor
  g1135
  (
    n1174,
    n1056,
    n1028,
    n1141,
    n1034
  );


  nor
  g1136
  (
    n1166,
    n1049,
    n1058,
    n1051,
    n1135
  );


  xnor
  g1137
  (
    n1176,
    n1140,
    n1052,
    n1056,
    n1023
  );


  xor
  g1138
  (
    n1167,
    n1046,
    n995,
    n1021,
    n1001
  );


  xor
  g1139
  (
    n1178,
    n1053,
    n1137,
    n1003,
    n1014
  );


  xor
  g1140
  (
    n1162,
    n1059,
    n994,
    n1140,
    n1044
  );


  nand
  g1141
  (
    n1168,
    n1033,
    n1138,
    n1037
  );


  xnor
  g1142
  (
    n1172,
    n1041,
    n1040,
    n991,
    n1006
  );


  xnor
  g1143
  (
    n1177,
    n1022,
    n1135,
    n1005,
    n1027
  );


  xor
  g1144
  (
    n1157,
    n1032,
    n1026,
    n1047,
    n1136
  );


  or
  g1145
  (
    n1156,
    n992,
    n1031,
    n1139,
    n1018
  );


  and
  g1146
  (
    n1158,
    n1025,
    n1141,
    n1059,
    n1137
  );


  buf
  g1147
  (
    n1216,
    n1142
  );


  buf
  g1148
  (
    n1213,
    n1163
  );


  not
  g1149
  (
    n1219,
    n1105
  );


  not
  g1150
  (
    n1198,
    n1160
  );


  buf
  g1151
  (
    n1191,
    n1075
  );


  buf
  g1152
  (
    n1184,
    n1065
  );


  nor
  g1153
  (
    n1199,
    n1165,
    n1103,
    n1111,
    n1076
  );


  xor
  g1154
  (
    n1222,
    n1164,
    n1073,
    n1166,
    n1104
  );


  or
  g1155
  (
    n1211,
    n1079,
    n1070,
    n1122,
    n1067
  );


  nor
  g1156
  (
    n1208,
    n1072,
    n939,
    n1068,
    n1166
  );


  xor
  g1157
  (
    n1194,
    n1065,
    n940,
    n1061,
    n939
  );


  and
  g1158
  (
    n1215,
    n1069,
    n1108,
    n1067,
    n1068
  );


  xor
  g1159
  (
    n1203,
    n1121,
    n1159,
    n1063,
    n1164
  );


  or
  g1160
  (
    n1204,
    n940,
    n1063,
    n1144,
    n1116
  );


  nor
  g1161
  (
    n1201,
    n1072,
    n1112,
    n1073,
    n1164
  );


  and
  g1162
  (
    n1221,
    n1161,
    n1117,
    n1095,
    n1110
  );


  xnor
  g1163
  (
    n1217,
    n1159,
    n1071,
    n1145,
    n1078
  );


  and
  g1164
  (
    n1209,
    n1060,
    n1163,
    n1167,
    n1162
  );


  and
  g1165
  (
    n1196,
    n1163,
    n1065,
    n1115,
    n1096
  );


  or
  g1166
  (
    n1186,
    n1076,
    n1076,
    n1170,
    n939
  );


  nor
  g1167
  (
    n1185,
    n1160,
    n1161,
    n1060,
    n1143
  );


  nand
  g1168
  (
    n1187,
    n1062,
    n1077,
    n1145,
    n1168
  );


  nor
  g1169
  (
    n1200,
    n1156,
    n1162,
    n1168,
    n1169
  );


  xor
  g1170
  (
    KeyWire_0_50,
    n1079,
    n1124,
    n1167,
    n1120
  );


  xnor
  g1171
  (
    n1205,
    n1142,
    n1071,
    n940,
    n1107
  );


  or
  g1172
  (
    n1192,
    n1066,
    n1156,
    n1060,
    n1166
  );


  nor
  g1173
  (
    n1206,
    n1158,
    n1100,
    n1077
  );


  nor
  g1174
  (
    n1202,
    n1170,
    n1066,
    n1075,
    n1157
  );


  nand
  g1175
  (
    n1180,
    n1068,
    n1075,
    n940,
    n1144
  );


  and
  g1176
  (
    n1188,
    n1145,
    n742,
    n1070,
    n1119
  );


  and
  g1177
  (
    n1190,
    n1067,
    n939,
    n1101,
    n1106
  );


  and
  g1178
  (
    n1195,
    n1063,
    n1162,
    n1097,
    n1167
  );


  nand
  g1179
  (
    n1197,
    n1155,
    n1158,
    n1144,
    n1073
  );


  nand
  g1180
  (
    n1207,
    n1143,
    n1069,
    n1161,
    n1062
  );


  nor
  g1181
  (
    n1220,
    n1113,
    n1155,
    n1114,
    n1169
  );


  xnor
  g1182
  (
    n1223,
    n1145,
    n1169,
    n1061,
    n1168
  );


  and
  g1183
  (
    n1183,
    n1071,
    n1154,
    n1069,
    n1078
  );


  xor
  g1184
  (
    n1214,
    n1109,
    n1123,
    n1118,
    n1154
  );


  or
  g1185
  (
    n1210,
    n1078,
    n1143,
    n1074
  );


  or
  g1186
  (
    n1218,
    n1064,
    n1142,
    n1074,
    n1066
  );


  xor
  g1187
  (
    n1189,
    n743,
    n1157,
    n1099,
    n1062
  );


  xor
  g1188
  (
    n1212,
    n1061,
    n1144,
    n1064,
    n1070
  );


  nor
  g1189
  (
    n1181,
    n1074,
    n1102,
    n1064,
    n1165
  );


  xnor
  g1190
  (
    n1193,
    n1072,
    n1098,
    n1160,
    n1165
  );


  buf
  g1191
  (
    KeyWire_0_5,
    n944
  );


  not
  g1192
  (
    n1225,
    n1187
  );


  buf
  g1193
  (
    n1239,
    n1130
  );


  not
  g1194
  (
    n1238,
    n1214
  );


  buf
  g1195
  (
    n1246,
    n1152
  );


  buf
  g1196
  (
    n1244,
    n1150
  );


  or
  g1197
  (
    n1261,
    n1150,
    n1134,
    n898
  );


  or
  g1198
  (
    n1258,
    n1149,
    n1133,
    n1219
  );


  xnor
  g1199
  (
    KeyWire_0_46,
    n1196,
    n1222,
    n1131
  );


  nor
  g1200
  (
    n1234,
    n1210,
    n1080,
    n1146
  );


  xnor
  g1201
  (
    n1249,
    n1133,
    n898,
    n1148
  );


  or
  g1202
  (
    n1251,
    n1202,
    n1152,
    n1131
  );


  nand
  g1203
  (
    n1263,
    n1180,
    n944,
    n1148
  );


  xnor
  g1204
  (
    n1262,
    n1189,
    n1205,
    n944
  );


  and
  g1205
  (
    KeyWire_0_48,
    n1129,
    n1081,
    n1134
  );


  and
  g1206
  (
    n1228,
    n1215,
    n1134,
    n1206
  );


  and
  g1207
  (
    n1240,
    n941,
    n1216,
    n1081
  );


  or
  g1208
  (
    n1226,
    n942,
    n1130,
    n1211
  );


  or
  g1209
  (
    n1259,
    n1151,
    n1195,
    n1185
  );


  xnor
  g1210
  (
    n1253,
    n1079,
    n1132,
    n1082
  );


  and
  g1211
  (
    KeyWire_0_12,
    n1149,
    n1192,
    n1146
  );


  or
  g1212
  (
    n1227,
    n1081,
    n1220,
    n1151
  );


  and
  g1213
  (
    n1245,
    n1183,
    n1221,
    n1150
  );


  xnor
  g1214
  (
    n1229,
    n1147,
    n1193,
    n1149
  );


  xnor
  g1215
  (
    n1265,
    n1200,
    n1147,
    n1149
  );


  nand
  g1216
  (
    n1233,
    n1181,
    n941,
    n943
  );


  or
  g1217
  (
    n1252,
    n1190,
    n1130,
    n1223
  );


  and
  g1218
  (
    n1241,
    n1146,
    n1213,
    n1188
  );


  or
  g1219
  (
    n1224,
    n1207,
    n1131,
    n1209
  );


  xnor
  g1220
  (
    KeyWire_0_58,
    n1134,
    n1182,
    n943
  );


  or
  g1221
  (
    n1231,
    n1212,
    n1197,
    n944
  );


  xnor
  g1222
  (
    n1237,
    n1208,
    n1132
  );


  nand
  g1223
  (
    n1243,
    n1150,
    n1133,
    n943
  );


  and
  g1224
  (
    n1257,
    n1204,
    n1147,
    n1151
  );


  xnor
  g1225
  (
    KeyWire_0_17,
    n1201,
    n1133,
    n943
  );


  and
  g1226
  (
    n1242,
    n1151,
    n942,
    n1146
  );


  nor
  g1227
  (
    n1248,
    n942,
    n1186,
    n1203
  );


  nand
  g1228
  (
    n1236,
    n1148,
    n1080,
    n1199
  );


  nand
  g1229
  (
    n1266,
    n1218,
    n941,
    n1194
  );


  and
  g1230
  (
    n1232,
    n1147,
    n1131,
    n1148
  );


  or
  g1231
  (
    n1230,
    n941,
    n942,
    n1132
  );


  and
  g1232
  (
    n1254,
    n1184,
    n1198,
    n1217
  );


  xnor
  g1233
  (
    n1235,
    n1130,
    n1080,
    n1191
  );


  buf
  g1234
  (
    n1367,
    n1260
  );


  buf
  g1235
  (
    n1270,
    n1153
  );


  not
  g1236
  (
    n1330,
    n1236
  );


  not
  g1237
  (
    n1353,
    n1239
  );


  not
  g1238
  (
    n1340,
    n1243
  );


  buf
  g1239
  (
    n1377,
    n1232
  );


  buf
  g1240
  (
    n1351,
    n1236
  );


  buf
  g1241
  (
    n1293,
    n1247
  );


  not
  g1242
  (
    n1281,
    n1255
  );


  not
  g1243
  (
    n1357,
    n1230
  );


  not
  g1244
  (
    n1335,
    n1237
  );


  not
  g1245
  (
    n1333,
    n1249
  );


  buf
  g1246
  (
    n1374,
    n1153
  );


  buf
  g1247
  (
    n1317,
    n1255
  );


  not
  g1248
  (
    n1364,
    n1228
  );


  buf
  g1249
  (
    n1301,
    n1225
  );


  buf
  g1250
  (
    n1288,
    n1249
  );


  buf
  g1251
  (
    n1310,
    n1234
  );


  not
  g1252
  (
    n1300,
    n1234
  );


  buf
  g1253
  (
    n1343,
    n1260
  );


  buf
  g1254
  (
    n1360,
    n1246
  );


  not
  g1255
  (
    n1295,
    n1226
  );


  buf
  g1256
  (
    n1287,
    n1235
  );


  not
  g1257
  (
    n1312,
    n1259
  );


  not
  g1258
  (
    n1277,
    n1245
  );


  buf
  g1259
  (
    n1365,
    n1250
  );


  not
  g1260
  (
    n1323,
    n1238
  );


  buf
  g1261
  (
    n1373,
    n1241
  );


  not
  g1262
  (
    n1303,
    n1244
  );


  buf
  g1263
  (
    n1363,
    n1248
  );


  buf
  g1264
  (
    n1368,
    n1251
  );


  not
  g1265
  (
    n1361,
    n1239
  );


  not
  g1266
  (
    n1337,
    n1247
  );


  not
  g1267
  (
    n1372,
    n1229
  );


  buf
  g1268
  (
    n1332,
    n1226
  );


  not
  g1269
  (
    n1328,
    n1258
  );


  not
  g1270
  (
    n1354,
    n1226
  );


  buf
  g1271
  (
    n1267,
    n1252
  );


  buf
  g1272
  (
    n1345,
    n1231
  );


  not
  g1273
  (
    n1316,
    n1227
  );


  buf
  g1274
  (
    n1307,
    n1244
  );


  buf
  g1275
  (
    n1304,
    n1242
  );


  not
  g1276
  (
    n1355,
    n1230
  );


  buf
  g1277
  (
    n1331,
    n1227
  );


  not
  g1278
  (
    n1291,
    n1256
  );


  not
  g1279
  (
    n1375,
    n1231
  );


  not
  g1280
  (
    n1336,
    n1233
  );


  buf
  g1281
  (
    n1376,
    n1258
  );


  buf
  g1282
  (
    n1362,
    n1152
  );


  buf
  g1283
  (
    n1338,
    n1260
  );


  buf
  g1284
  (
    n1369,
    n1228
  );


  buf
  g1285
  (
    n1348,
    n1235
  );


  buf
  g1286
  (
    n1314,
    n1243
  );


  not
  g1287
  (
    n1326,
    n1225
  );


  not
  g1288
  (
    n1329,
    n1252
  );


  buf
  g1289
  (
    n1276,
    n1238
  );


  not
  g1290
  (
    n1346,
    n1259
  );


  buf
  g1291
  (
    n1290,
    n1233
  );


  not
  g1292
  (
    n1278,
    n1152
  );


  not
  g1293
  (
    KeyWire_0_16,
    n1253
  );


  buf
  g1294
  (
    n1286,
    n1237
  );


  buf
  g1295
  (
    n1269,
    n1229
  );


  not
  g1296
  (
    n1275,
    n1237
  );


  not
  g1297
  (
    n1358,
    n1242
  );


  buf
  g1298
  (
    n1320,
    n1259
  );


  not
  g1299
  (
    n1321,
    n1233
  );


  buf
  g1300
  (
    n1319,
    n1229
  );


  not
  g1301
  (
    n1297,
    n1232
  );


  not
  g1302
  (
    n1313,
    n1252
  );


  not
  g1303
  (
    n1282,
    n1241
  );


  buf
  g1304
  (
    n1324,
    n1236
  );


  not
  g1305
  (
    n1318,
    n1242
  );


  buf
  g1306
  (
    KeyWire_0_22,
    n1227
  );


  buf
  g1307
  (
    n1366,
    n1256
  );


  buf
  g1308
  (
    n1272,
    n1254
  );


  buf
  g1309
  (
    n1280,
    n1248
  );


  buf
  g1310
  (
    n1344,
    n1248
  );


  buf
  g1311
  (
    n1311,
    n1247
  );


  buf
  g1312
  (
    n1315,
    n1257
  );


  not
  g1313
  (
    n1325,
    n1239
  );


  not
  g1314
  (
    n1302,
    n1224
  );


  not
  g1315
  (
    n1294,
    n1225
  );


  buf
  g1316
  (
    n1378,
    n1255
  );


  buf
  g1317
  (
    n1284,
    n1250
  );


  not
  g1318
  (
    n1322,
    n1243
  );


  buf
  g1319
  (
    n1334,
    n1258
  );


  not
  g1320
  (
    n1341,
    n1240
  );


  buf
  g1321
  (
    n1289,
    n1240
  );


  not
  g1322
  (
    n1371,
    n1238
  );


  not
  g1323
  (
    KeyWire_0_39,
    n1257
  );


  buf
  g1324
  (
    n1352,
    n1228
  );


  not
  g1325
  (
    n1308,
    n1253
  );


  buf
  g1326
  (
    n1370,
    n1230
  );


  buf
  g1327
  (
    n1283,
    n1254
  );


  buf
  g1328
  (
    n1285,
    n1232
  );


  buf
  g1329
  (
    n1309,
    n1257
  );


  buf
  g1330
  (
    n1327,
    n1257
  );


  buf
  g1331
  (
    n1356,
    n1259
  );


  buf
  g1332
  (
    n1342,
    n1251
  );


  buf
  g1333
  (
    n1299,
    n1254
  );


  not
  g1334
  (
    n1349,
    n1250
  );


  not
  g1335
  (
    n1350,
    n1258
  );


  not
  g1336
  (
    n1273,
    n1231
  );


  not
  g1337
  (
    n1268,
    n1241
  );


  buf
  g1338
  (
    n1306,
    n1153
  );


  not
  g1339
  (
    n1305,
    n1245
  );


  buf
  g1340
  (
    n1296,
    n1246
  );


  not
  g1341
  (
    n1271,
    n1246
  );


  not
  g1342
  (
    n1279,
    n1249
  );


  not
  g1343
  (
    n1292,
    n1253
  );


  xor
  g1344
  (
    n1347,
    n1251,
    n1245,
    n1240,
    n1153
  );


  xnor
  g1345
  (
    n1274,
    n1234,
    n1244,
    n1235,
    n1256
  );


  buf
  g1346
  (
    n1675,
    n1317
  );


  buf
  g1347
  (
    n1523,
    n1179
  );


  buf
  g1348
  (
    n1445,
    n1338
  );


  not
  g1349
  (
    n1387,
    n1277
  );


  buf
  g1350
  (
    n1742,
    n1328
  );


  not
  g1351
  (
    n1729,
    n1316
  );


  buf
  g1352
  (
    n1667,
    n1311
  );


  not
  g1353
  (
    KeyWire_0_14,
    n1326
  );


  not
  g1354
  (
    n1391,
    n1342
  );


  buf
  g1355
  (
    n1733,
    n1354
  );


  buf
  g1356
  (
    n1715,
    n1351
  );


  not
  g1357
  (
    n1638,
    n1284
  );


  buf
  g1358
  (
    n1741,
    n1267
  );


  buf
  g1359
  (
    n1662,
    n1314
  );


  not
  g1360
  (
    n1753,
    n1305
  );


  not
  g1361
  (
    n1583,
    n1311
  );


  not
  g1362
  (
    n1587,
    n1350
  );


  buf
  g1363
  (
    n1637,
    n1294
  );


  not
  g1364
  (
    n1511,
    n1348
  );


  not
  g1365
  (
    n1656,
    n1287
  );


  not
  g1366
  (
    n1562,
    n1344
  );


  buf
  g1367
  (
    n1503,
    n1313
  );


  buf
  g1368
  (
    n1427,
    n1324
  );


  not
  g1369
  (
    n1507,
    n1331
  );


  not
  g1370
  (
    n1575,
    n1320
  );


  buf
  g1371
  (
    n1747,
    n1355
  );


  not
  g1372
  (
    n1695,
    n1332
  );


  buf
  g1373
  (
    n1532,
    n1323
  );


  not
  g1374
  (
    n1451,
    n1275
  );


  not
  g1375
  (
    n1605,
    n1297
  );


  buf
  g1376
  (
    n1526,
    n1349
  );


  buf
  g1377
  (
    n1564,
    n1307
  );


  buf
  g1378
  (
    n1443,
    n1173
  );


  buf
  g1379
  (
    n1740,
    n1299
  );


  buf
  g1380
  (
    n1702,
    n1291
  );


  buf
  g1381
  (
    n1433,
    n1294
  );


  buf
  g1382
  (
    n1654,
    n1283
  );


  not
  g1383
  (
    n1636,
    n1338
  );


  not
  g1384
  (
    n1652,
    n1175
  );


  not
  g1385
  (
    n1446,
    n1325
  );


  buf
  g1386
  (
    n1722,
    n1347
  );


  not
  g1387
  (
    n1726,
    n1348
  );


  not
  g1388
  (
    n1506,
    n1270
  );


  not
  g1389
  (
    n1645,
    n1336
  );


  buf
  g1390
  (
    n1593,
    n1276
  );


  not
  g1391
  (
    n1477,
    n1293
  );


  buf
  g1392
  (
    n1743,
    n1281
  );


  not
  g1393
  (
    n1669,
    n1282
  );


  not
  g1394
  (
    n1533,
    n1340
  );


  buf
  g1395
  (
    KeyWire_0_28,
    n1334
  );


  buf
  g1396
  (
    n1501,
    n1178
  );


  not
  g1397
  (
    n1724,
    n1334
  );


  not
  g1398
  (
    n1746,
    n1285
  );


  buf
  g1399
  (
    n1582,
    n1321
  );


  buf
  g1400
  (
    n1534,
    n1274
  );


  buf
  g1401
  (
    n1671,
    n1344
  );


  not
  g1402
  (
    n1509,
    n1269
  );


  not
  g1403
  (
    n1705,
    n1340
  );


  buf
  g1404
  (
    n1479,
    n1293
  );


  not
  g1405
  (
    n1467,
    n1301
  );


  not
  g1406
  (
    n1612,
    n1357
  );


  not
  g1407
  (
    n1437,
    n1289
  );


  buf
  g1408
  (
    n1685,
    n1357
  );


  not
  g1409
  (
    n1417,
    n1275
  );


  buf
  g1410
  (
    n1469,
    n1290
  );


  not
  g1411
  (
    n1674,
    n1303
  );


  buf
  g1412
  (
    n1418,
    n1287
  );


  buf
  g1413
  (
    n1725,
    n1361
  );


  buf
  g1414
  (
    n1383,
    n1306
  );


  not
  g1415
  (
    n1500,
    n1270
  );


  buf
  g1416
  (
    n1466,
    n1288
  );


  buf
  g1417
  (
    n1713,
    n1283
  );


  buf
  g1418
  (
    n1599,
    n1323
  );


  not
  g1419
  (
    n1397,
    n1305
  );


  not
  g1420
  (
    n1390,
    n1278
  );


  buf
  g1421
  (
    n1557,
    n1292
  );


  buf
  g1422
  (
    n1472,
    n1349
  );


  buf
  g1423
  (
    n1623,
    n1329
  );


  not
  g1424
  (
    n1580,
    n1319
  );


  buf
  g1425
  (
    n1571,
    n1284
  );


  not
  g1426
  (
    n1629,
    n1343
  );


  not
  g1427
  (
    n1749,
    n1316
  );


  not
  g1428
  (
    n1520,
    n1322
  );


  buf
  g1429
  (
    n1738,
    n1359
  );


  not
  g1430
  (
    n1595,
    n1315
  );


  buf
  g1431
  (
    n1596,
    n1347
  );


  buf
  g1432
  (
    n1584,
    n1298
  );


  buf
  g1433
  (
    n1395,
    n1279
  );


  not
  g1434
  (
    n1690,
    n1319
  );


  buf
  g1435
  (
    n1586,
    n1282
  );


  buf
  g1436
  (
    n1428,
    n1174
  );


  not
  g1437
  (
    n1402,
    n1083
  );


  buf
  g1438
  (
    n1478,
    n1301
  );


  not
  g1439
  (
    n1542,
    n1338
  );


  buf
  g1440
  (
    n1706,
    n1331
  );


  not
  g1441
  (
    n1535,
    n1296
  );


  buf
  g1442
  (
    n1613,
    n1309
  );


  buf
  g1443
  (
    n1615,
    n1273
  );


  not
  g1444
  (
    n1622,
    n1342
  );


  not
  g1445
  (
    n1463,
    n1176
  );


  buf
  g1446
  (
    n1727,
    n1276
  );


  not
  g1447
  (
    n1687,
    n1352
  );


  not
  g1448
  (
    n1496,
    n1346
  );


  not
  g1449
  (
    n1611,
    n1311
  );


  buf
  g1450
  (
    n1589,
    n1296
  );


  buf
  g1451
  (
    n1739,
    n1290
  );


  not
  g1452
  (
    n1540,
    n1342
  );


  not
  g1453
  (
    n1384,
    n1310
  );


  buf
  g1454
  (
    n1488,
    n1337
  );


  not
  g1455
  (
    n1409,
    n1325
  );


  not
  g1456
  (
    n1604,
    n1278
  );


  not
  g1457
  (
    n1399,
    n1306
  );


  not
  g1458
  (
    n1415,
    n1271
  );


  not
  g1459
  (
    n1686,
    n1279
  );


  buf
  g1460
  (
    n1392,
    n1333
  );


  buf
  g1461
  (
    n1386,
    n1312
  );


  not
  g1462
  (
    n1620,
    n1301
  );


  buf
  g1463
  (
    n1730,
    n1347
  );


  not
  g1464
  (
    n1655,
    n1271
  );


  buf
  g1465
  (
    n1452,
    n1327
  );


  not
  g1466
  (
    n1665,
    n1275
  );


  buf
  g1467
  (
    n1525,
    n1309
  );


  buf
  g1468
  (
    n1572,
    n1172
  );


  buf
  g1469
  (
    n1538,
    n1339
  );


  not
  g1470
  (
    n1708,
    n1289
  );


  buf
  g1471
  (
    n1563,
    n1325
  );


  buf
  g1472
  (
    n1630,
    n1325
  );


  not
  g1473
  (
    n1720,
    n1318
  );


  buf
  g1474
  (
    n1592,
    n1267
  );


  not
  g1475
  (
    n1432,
    n1320
  );


  buf
  g1476
  (
    n1748,
    n1269
  );


  not
  g1477
  (
    n1545,
    n1357
  );


  buf
  g1478
  (
    n1541,
    n1326
  );


  buf
  g1479
  (
    n1552,
    n1179
  );


  buf
  g1480
  (
    n1554,
    n1312
  );


  buf
  g1481
  (
    n1628,
    n1298
  );


  not
  g1482
  (
    n1579,
    n1309
  );


  buf
  g1483
  (
    n1698,
    n1285
  );


  buf
  g1484
  (
    n1524,
    n1274
  );


  not
  g1485
  (
    n1414,
    n1174
  );


  not
  g1486
  (
    n1585,
    n1288
  );


  buf
  g1487
  (
    n1718,
    n1272
  );


  not
  g1488
  (
    n1588,
    n1296
  );


  buf
  g1489
  (
    n1388,
    n1279
  );


  buf
  g1490
  (
    n1699,
    n1173
  );


  not
  g1491
  (
    n1617,
    n1311
  );


  not
  g1492
  (
    n1703,
    n1340
  );


  not
  g1493
  (
    n1490,
    n1353
  );


  not
  g1494
  (
    n1517,
    n1278
  );


  not
  g1495
  (
    n1473,
    n1307
  );


  not
  g1496
  (
    n1664,
    n1273
  );


  not
  g1497
  (
    n1597,
    n1328
  );


  not
  g1498
  (
    n1416,
    n1312
  );


  not
  g1499
  (
    n1561,
    n1339
  );


  not
  g1500
  (
    n1701,
    n1314
  );


  not
  g1501
  (
    n1430,
    n1358
  );


  buf
  g1502
  (
    n1491,
    n1286
  );


  not
  g1503
  (
    n1606,
    n1282
  );


  buf
  g1504
  (
    n1553,
    n1319
  );


  buf
  g1505
  (
    n1465,
    n1289
  );


  buf
  g1506
  (
    n1462,
    n1319
  );


  not
  g1507
  (
    n1653,
    n1082
  );


  not
  g1508
  (
    n1470,
    n1276
  );


  buf
  g1509
  (
    n1398,
    n1323
  );


  buf
  g1510
  (
    n1548,
    n1312
  );


  not
  g1511
  (
    n1751,
    n1295
  );


  not
  g1512
  (
    n1505,
    n1360
  );


  buf
  g1513
  (
    n1646,
    n1324
  );


  buf
  g1514
  (
    n1547,
    n1335
  );


  not
  g1515
  (
    n1419,
    n1317
  );


  buf
  g1516
  (
    KeyWire_0_37,
    n1178
  );


  not
  g1517
  (
    n1504,
    n1349
  );


  buf
  g1518
  (
    n1471,
    n1316
  );


  not
  g1519
  (
    n1661,
    n1280
  );


  not
  g1520
  (
    n1448,
    n1330
  );


  not
  g1521
  (
    n1567,
    n1343
  );


  buf
  g1522
  (
    n1401,
    n1310
  );


  buf
  g1523
  (
    n1408,
    n1353
  );


  buf
  g1524
  (
    n1435,
    n1296
  );


  not
  g1525
  (
    n1457,
    n1295
  );


  not
  g1526
  (
    n1735,
    n1329
  );


  buf
  g1527
  (
    n1558,
    n1343
  );


  not
  g1528
  (
    n1403,
    n1286
  );


  buf
  g1529
  (
    n1420,
    n1307
  );


  buf
  g1530
  (
    n1529,
    n1084
  );


  buf
  g1531
  (
    n1484,
    n1304
  );


  not
  g1532
  (
    n1453,
    n1344
  );


  not
  g1533
  (
    n1438,
    n1273
  );


  not
  g1534
  (
    n1481,
    n1346
  );


  buf
  g1535
  (
    n1644,
    n1326
  );


  buf
  g1536
  (
    n1696,
    n1356
  );


  buf
  g1537
  (
    n1590,
    n1327
  );


  buf
  g1538
  (
    n1521,
    n1334
  );


  not
  g1539
  (
    n1732,
    n1356
  );


  not
  g1540
  (
    n1624,
    n1360
  );


  buf
  g1541
  (
    n1700,
    n1315
  );


  not
  g1542
  (
    n1512,
    n1333
  );


  not
  g1543
  (
    n1704,
    n1320
  );


  buf
  g1544
  (
    KeyWire_0_18,
    n1171
  );


  buf
  g1545
  (
    n1568,
    n1340
  );


  buf
  g1546
  (
    n1577,
    n1301
  );


  buf
  g1547
  (
    n1413,
    n1276
  );


  not
  g1548
  (
    n1618,
    n1295
  );


  not
  g1549
  (
    n1736,
    n1344
  );


  not
  g1550
  (
    n1489,
    n1291
  );


  not
  g1551
  (
    n1677,
    n1306
  );


  not
  g1552
  (
    n1627,
    n1302
  );


  buf
  g1553
  (
    n1440,
    n1298
  );


  not
  g1554
  (
    n1607,
    n1297
  );


  not
  g1555
  (
    n1518,
    n1274
  );


  buf
  g1556
  (
    KeyWire_0_1,
    n1308
  );


  buf
  g1557
  (
    n1380,
    n1346
  );


  not
  g1558
  (
    n1406,
    n1082
  );


  buf
  g1559
  (
    n1404,
    n1318
  );


  buf
  g1560
  (
    n1639,
    n1291
  );


  buf
  g1561
  (
    n1632,
    n1171
  );


  not
  g1562
  (
    n1626,
    n1273
  );


  not
  g1563
  (
    n1694,
    n1268
  );


  not
  g1564
  (
    n1673,
    n1329
  );


  not
  g1565
  (
    n1672,
    n1083
  );


  not
  g1566
  (
    n1716,
    n1083
  );


  not
  g1567
  (
    n1487,
    n1175
  );


  not
  g1568
  (
    n1728,
    n1279
  );


  not
  g1569
  (
    n1423,
    n1334
  );


  buf
  g1570
  (
    n1556,
    n1271
  );


  not
  g1571
  (
    n1519,
    n1341
  );


  buf
  g1572
  (
    KeyWire_0_61,
    n1299
  );


  buf
  g1573
  (
    n1546,
    n1355
  );


  not
  g1574
  (
    n1449,
    n1175
  );


  not
  g1575
  (
    n1711,
    n1326
  );


  buf
  g1576
  (
    n1551,
    n1303
  );


  buf
  g1577
  (
    n1689,
    n1305
  );


  buf
  g1578
  (
    n1570,
    n1350
  );


  not
  g1579
  (
    n1666,
    n1318
  );


  not
  g1580
  (
    n1441,
    n1293
  );


  buf
  g1581
  (
    n1485,
    n1281
  );


  buf
  g1582
  (
    n1543,
    n1278
  );


  not
  g1583
  (
    n1731,
    n1298
  );


  not
  g1584
  (
    n1609,
    n1345
  );


  not
  g1585
  (
    n1410,
    n1269
  );


  not
  g1586
  (
    n1560,
    n1322
  );


  buf
  g1587
  (
    n1684,
    n1286
  );


  not
  g1588
  (
    n1566,
    n1302
  );


  not
  g1589
  (
    n1522,
    n1342
  );


  buf
  g1590
  (
    n1555,
    n1333
  );


  buf
  g1591
  (
    KeyWire_0_44,
    n1308
  );


  buf
  g1592
  (
    n1389,
    n1176
  );


  buf
  g1593
  (
    n1536,
    n1350
  );


  not
  g1594
  (
    n1679,
    n1336
  );


  buf
  g1595
  (
    n1752,
    n1290
  );


  not
  g1596
  (
    n1544,
    n1337
  );


  not
  g1597
  (
    n1411,
    n1170
  );


  not
  g1598
  (
    n1381,
    n1284
  );


  buf
  g1599
  (
    n1625,
    n1281
  );


  buf
  g1600
  (
    n1591,
    n1267
  );


  buf
  g1601
  (
    n1527,
    n1346
  );


  buf
  g1602
  (
    n1480,
    n1356
  );


  buf
  g1603
  (
    n1447,
    n1332
  );


  buf
  g1604
  (
    n1614,
    n1297
  );


  buf
  g1605
  (
    n1693,
    n1280
  );


  buf
  g1606
  (
    n1635,
    n1172
  );


  not
  g1607
  (
    n1603,
    n1347
  );


  buf
  g1608
  (
    n1464,
    n1327
  );


  buf
  g1609
  (
    n1429,
    n1299
  );


  not
  g1610
  (
    n1723,
    n1310
  );


  buf
  g1611
  (
    n1755,
    n1314
  );


  not
  g1612
  (
    n1621,
    n1314
  );


  buf
  g1613
  (
    KeyWire_0_51,
    n1335
  );


  not
  g1614
  (
    n1594,
    n1358
  );


  buf
  g1615
  (
    n1610,
    n1355
  );


  not
  g1616
  (
    n1565,
    n1316
  );


  not
  g1617
  (
    n1717,
    n1271
  );


  not
  g1618
  (
    n1598,
    n1359
  );


  not
  g1619
  (
    n1709,
    n1308
  );


  buf
  g1620
  (
    n1549,
    n1179
  );


  buf
  g1621
  (
    n1657,
    n1280
  );


  not
  g1622
  (
    n1712,
    n1281
  );


  buf
  g1623
  (
    n1474,
    n1321
  );


  buf
  g1624
  (
    n1659,
    n1351
  );


  not
  g1625
  (
    n1649,
    n1269
  );


  not
  g1626
  (
    n1710,
    n1345
  );


  buf
  g1627
  (
    n1502,
    n1272
  );


  not
  g1628
  (
    n1576,
    n1353
  );


  not
  g1629
  (
    n1642,
    n1324
  );


  buf
  g1630
  (
    n1660,
    n1270
  );


  buf
  g1631
  (
    n1510,
    n1299
  );


  buf
  g1632
  (
    n1707,
    n1297
  );


  buf
  g1633
  (
    n1734,
    n1324
  );


  not
  g1634
  (
    n1385,
    n1308
  );


  not
  g1635
  (
    n1499,
    n1327
  );


  buf
  g1636
  (
    n1631,
    n1359
  );


  buf
  g1637
  (
    n1407,
    n1352
  );


  not
  g1638
  (
    n1460,
    n1345
  );


  buf
  g1639
  (
    n1573,
    n1172
  );


  buf
  g1640
  (
    n1434,
    n1320
  );


  buf
  g1641
  (
    n1396,
    n1349
  );


  not
  g1642
  (
    n1678,
    n1358
  );


  buf
  g1643
  (
    n1550,
    n1306
  );


  not
  g1644
  (
    n1458,
    n1272
  );


  buf
  g1645
  (
    n1486,
    n1176
  );


  not
  g1646
  (
    n1497,
    n1318
  );


  buf
  g1647
  (
    n1682,
    n1272
  );


  buf
  g1648
  (
    n1658,
    n1292
  );


  buf
  g1649
  (
    n1559,
    n1294
  );


  not
  g1650
  (
    n1691,
    n1330
  );


  not
  g1651
  (
    n1382,
    n1285
  );


  not
  g1652
  (
    n1539,
    n1333
  );


  buf
  g1653
  (
    n1641,
    n1289
  );


  buf
  g1654
  (
    n1608,
    n1356
  );


  not
  g1655
  (
    n1668,
    n1177
  );


  buf
  g1656
  (
    n1600,
    n1084
  );


  buf
  g1657
  (
    n1643,
    n1277
  );


  buf
  g1658
  (
    n1714,
    n1359
  );


  not
  g1659
  (
    n1681,
    n1322
  );


  not
  g1660
  (
    n1495,
    n1315
  );


  buf
  g1661
  (
    n1601,
    n1268
  );


  not
  g1662
  (
    n1650,
    n1328
  );


  not
  g1663
  (
    n1578,
    n1084
  );


  not
  g1664
  (
    n1744,
    n1341
  );


  buf
  g1665
  (
    n1648,
    n1337
  );


  buf
  g1666
  (
    n1459,
    n1354
  );


  not
  g1667
  (
    n1721,
    n1302
  );


  not
  g1668
  (
    n1676,
    n1361
  );


  buf
  g1669
  (
    n1442,
    n1305
  );


  buf
  g1670
  (
    n1476,
    n1274
  );


  not
  g1671
  (
    n1697,
    n1357
  );


  not
  g1672
  (
    n1450,
    n1300
  );


  not
  g1673
  (
    n1412,
    n1277
  );


  buf
  g1674
  (
    n1516,
    n1355
  );


  not
  g1675
  (
    n1683,
    n1304
  );


  not
  g1676
  (
    n1574,
    n1335
  );


  not
  g1677
  (
    n1455,
    n1332
  );


  buf
  g1678
  (
    n1513,
    n1288
  );


  buf
  g1679
  (
    n1680,
    n1294
  );


  not
  g1680
  (
    n1537,
    n1350
  );


  buf
  g1681
  (
    n1634,
    n1337
  );


  not
  g1682
  (
    n1602,
    n1317
  );


  buf
  g1683
  (
    n1498,
    n1304
  );


  buf
  g1684
  (
    n1647,
    n1341
  );


  not
  g1685
  (
    n1400,
    n1315
  );


  not
  g1686
  (
    n1405,
    n1285
  );


  not
  g1687
  (
    n1515,
    n1288
  );


  not
  g1688
  (
    KeyWire_0_19,
    n1300
  );


  buf
  g1689
  (
    n1581,
    n1354
  );


  not
  g1690
  (
    n1493,
    n1177
  );


  not
  g1691
  (
    n1456,
    n1348
  );


  not
  g1692
  (
    n1393,
    n1280
  );


  not
  g1693
  (
    n1670,
    n1332
  );


  not
  g1694
  (
    KeyWire_0_47,
    n1313
  );


  not
  g1695
  (
    n1745,
    n1307
  );


  not
  g1696
  (
    n1421,
    n1277
  );


  not
  g1697
  (
    n1394,
    n1352
  );


  buf
  g1698
  (
    n1640,
    n1317
  );


  buf
  g1699
  (
    n1379,
    n1323
  );


  not
  g1700
  (
    n1530,
    n1292
  );


  not
  g1701
  (
    n1492,
    n1330
  );


  not
  g1702
  (
    n1483,
    n1353
  );


  not
  g1703
  (
    n1475,
    n1268
  );


  not
  g1704
  (
    n1444,
    n1300
  );


  buf
  g1705
  (
    n1425,
    n1295
  );


  not
  g1706
  (
    n1439,
    n1360
  );


  not
  g1707
  (
    n1692,
    n1173
  );


  not
  g1708
  (
    n1531,
    n1341
  );


  not
  g1709
  (
    n1461,
    n1339
  );


  nand
  g1710
  (
    n1422,
    n1171,
    n1303,
    n1293,
    n1270
  );


  and
  g1711
  (
    n1619,
    n1360,
    n1275,
    n1304,
    n1352
  );


  nand
  g1712
  (
    n1426,
    n1361,
    n1291,
    n1268,
    n1338
  );


  xnor
  g1713
  (
    n1754,
    n1343,
    n1336,
    n1358,
    n1329
  );


  nor
  g1714
  (
    n1651,
    n1330,
    n1300,
    n1322,
    n1351
  );


  nor
  g1715
  (
    n1424,
    n1290,
    n1284,
    n1174,
    n1345
  );


  nor
  g1716
  (
    n1719,
    n1282,
    n1328,
    n1339,
    n1313
  );


  nand
  g1717
  (
    n1468,
    n1336,
    n1351,
    n1331,
    n1302
  );


  and
  g1718
  (
    n1436,
    n1292,
    n1331,
    n1321,
    n1309
  );


  nand
  g1719
  (
    n1616,
    n1283,
    n1313,
    n1267,
    n1348
  );


  xor
  g1720
  (
    n1663,
    n1310,
    n1303,
    n1178,
    n1283
  );


  nand
  g1721
  (
    n1528,
    n1287,
    n1177,
    n1321,
    n1286
  );


  and
  g1722
  (
    n1633,
    n1354,
    n1361,
    n1287,
    n1335
  );


  not
  g1723
  (
    KeyWire_0_59,
    n1382
  );


  buf
  g1724
  (
    n1756,
    n1381
  );


  buf
  g1725
  (
    n1757,
    n1380
  );


  not
  g1726
  (
    n1759,
    n1379
  );


  xnor
  g1727
  (
    n1764,
    n1262,
    n1265,
    n751,
    n1757
  );


  xnor
  g1728
  (
    n1760,
    n747,
    n1758,
    n756,
    n1264
  );


  and
  g1729
  (
    n1762,
    n1758,
    n1263,
    n1757,
    n1264
  );


  or
  g1730
  (
    n1766,
    n1756,
    n755,
    n945,
    n1266
  );


  and
  g1731
  (
    n1768,
    n1265,
    n1759,
    n745,
    n750
  );


  and
  g1732
  (
    n1761,
    n1756,
    n1262,
    n752
  );


  or
  g1733
  (
    n1769,
    n1261,
    n1266,
    n1758,
    n1264
  );


  xor
  g1734
  (
    n1767,
    n1758,
    n748,
    n1266,
    n1263
  );


  xnor
  g1735
  (
    n1772,
    n753,
    n1261,
    n945
  );


  and
  g1736
  (
    n1773,
    n754,
    n1263,
    n1757
  );


  xor
  g1737
  (
    n1770,
    n945,
    n1264,
    n1262,
    n1263
  );


  or
  g1738
  (
    n1763,
    n1261,
    n746,
    n1759,
    n1260
  );


  nor
  g1739
  (
    n1771,
    n1266,
    n1265,
    n1759
  );


  nand
  g1740
  (
    n1765,
    n945,
    n744,
    n1759,
    n749
  );


  buf
  g1741
  (
    n1791,
    n1767
  );


  not
  g1742
  (
    n1810,
    n1362
  );


  buf
  g1743
  (
    n1792,
    n1765
  );


  not
  g1744
  (
    n1785,
    n1369
  );


  buf
  g1745
  (
    n1799,
    n1762
  );


  not
  g1746
  (
    n1795,
    n30
  );


  buf
  g1747
  (
    n1826,
    n1768
  );


  buf
  g1748
  (
    n1780,
    n1365
  );


  buf
  g1749
  (
    n1782,
    n1769
  );


  buf
  g1750
  (
    n1796,
    n1768
  );


  not
  g1751
  (
    n1823,
    n1366
  );


  not
  g1752
  (
    n1822,
    n1762
  );


  not
  g1753
  (
    n1794,
    n1769
  );


  not
  g1754
  (
    n1778,
    n1770
  );


  not
  g1755
  (
    n1818,
    n1374
  );


  buf
  g1756
  (
    n1788,
    n1365
  );


  not
  g1757
  (
    n1827,
    n1762
  );


  not
  g1758
  (
    n1802,
    n1369
  );


  buf
  g1759
  (
    n1787,
    n1767
  );


  buf
  g1760
  (
    n1783,
    n1378
  );


  not
  g1761
  (
    n1775,
    n31
  );


  buf
  g1762
  (
    n1784,
    n1368
  );


  not
  g1763
  (
    n1828,
    n1363
  );


  not
  g1764
  (
    n1801,
    n1364
  );


  not
  g1765
  (
    KeyWire_0_42,
    n1768
  );


  buf
  g1766
  (
    n1779,
    n1378
  );


  not
  g1767
  (
    n1808,
    n1377
  );


  buf
  g1768
  (
    n1805,
    n1764
  );


  and
  g1769
  (
    n1829,
    n29,
    n1760
  );


  nor
  g1770
  (
    n1812,
    n1770,
    n31,
    n1368,
    n1764
  );


  or
  g1771
  (
    n1798,
    n1373,
    n1761,
    n1366,
    n1763
  );


  xnor
  g1772
  (
    n1811,
    n1772,
    n1765,
    n31,
    n1768
  );


  xnor
  g1773
  (
    KeyWire_0_9,
    n1760,
    n1366,
    n1767,
    n1368
  );


  or
  g1774
  (
    n1797,
    n1373,
    n1377,
    n1773,
    n1376
  );


  xnor
  g1775
  (
    n1776,
    n1764,
    n1362,
    n1376,
    n31
  );


  nand
  g1776
  (
    n1817,
    n32,
    n1370,
    n1363,
    n1371
  );


  xor
  g1777
  (
    n1786,
    n1772,
    n1763,
    n1760,
    n1376
  );


  or
  g1778
  (
    n1816,
    n1767,
    n1771,
    n30,
    n1766
  );


  xnor
  g1779
  (
    n1821,
    n1378,
    n1770,
    n1367,
    n1370
  );


  xor
  g1780
  (
    n1804,
    n1375,
    n1375,
    n1377,
    n1373
  );


  xnor
  g1781
  (
    n1825,
    n1371,
    n1375,
    n1374,
    n1761
  );


  or
  g1782
  (
    n1774,
    n1760,
    n1764,
    n1771,
    n32
  );


  or
  g1783
  (
    n1815,
    n1761,
    n1365,
    n1367,
    n1769
  );


  xnor
  g1784
  (
    n1803,
    n1374,
    n1370,
    n1369
  );


  xnor
  g1785
  (
    n1789,
    n1366,
    n1376,
    n1773,
    n1364
  );


  nand
  g1786
  (
    n1781,
    n1363,
    n1772,
    n1372
  );


  nor
  g1787
  (
    n1777,
    n1773,
    n1377,
    n1365,
    n1769
  );


  or
  g1788
  (
    n1790,
    n1761,
    n1368,
    n1375,
    n1364
  );


  xor
  g1789
  (
    n1800,
    n1362,
    n1371,
    n1367,
    n1363
  );


  nand
  g1790
  (
    KeyWire_0_40,
    n1362,
    n1367,
    n1763,
    n1762
  );


  nand
  g1791
  (
    n1809,
    n29,
    n32,
    n1372
  );


  xor
  g1792
  (
    n1824,
    n1364,
    n1372,
    n30,
    n1378
  );


  and
  g1793
  (
    n1814,
    n1771,
    n1766,
    n1765,
    n1773
  );


  or
  g1794
  (
    n1820,
    n1372,
    n1766,
    n1771,
    n1371
  );


  and
  g1795
  (
    n1807,
    n1770,
    n1373,
    n30,
    n1763
  );


  nor
  g1796
  (
    n1813,
    n1765,
    n1369,
    n1766,
    n1374
  );


  xor
  g1797
  (
    n1877,
    n1575,
    n1406,
    n1818,
    n1780
  );


  and
  g1798
  (
    n1933,
    n1778,
    n1721,
    n1658,
    n1803
  );


  xor
  g1799
  (
    n1832,
    n1808,
    n1812,
    n1793,
    n1822
  );


  or
  g1800
  (
    n1884,
    n1713,
    n1533,
    n1742,
    n1418
  );


  xor
  g1801
  (
    n1915,
    n1618,
    n1781,
    n1403,
    n1537
  );


  nand
  g1802
  (
    n1927,
    n1801,
    n1489,
    n1683,
    n1396
  );


  nand
  g1803
  (
    n1955,
    n1498,
    n1682,
    n1800,
    n1745
  );


  or
  g1804
  (
    n1848,
    n1414,
    n1790,
    n1434,
    n1677
  );


  nor
  g1805
  (
    n1913,
    n1755,
    n1469,
    n1827,
    n1467
  );


  nand
  g1806
  (
    n1830,
    n1566,
    n1426,
    n1799,
    n1724
  );


  and
  g1807
  (
    n1842,
    n1648,
    n1780,
    n1811,
    n1613
  );


  nor
  g1808
  (
    n1947,
    n1420,
    n1829,
    n1716,
    n1826
  );


  or
  g1809
  (
    n1882,
    n1488,
    n1617,
    n1573,
    n1718
  );


  nor
  g1810
  (
    n1909,
    n1774,
    n1816,
    n1546,
    n1725
  );


  xor
  g1811
  (
    n1843,
    n1383,
    n1398,
    n1819,
    n1800
  );


  nand
  g1812
  (
    n1836,
    n1815,
    n1561,
    n1644,
    n1726
  );


  and
  g1813
  (
    n1856,
    n1503,
    n1810,
    n1435,
    n1776
  );


  xor
  g1814
  (
    n1914,
    n1652,
    n1661,
    n1564,
    n1740
  );


  xor
  g1815
  (
    n1865,
    n1823,
    n1438,
    n1822,
    n1656
  );


  and
  g1816
  (
    n1932,
    n1696,
    n1730,
    n1782,
    n1394
  );


  nor
  g1817
  (
    n1860,
    n1814,
    n1534,
    n1508,
    n1574
  );


  or
  g1818
  (
    n1931,
    n1810,
    n1585,
    n1712,
    n1802
  );


  nor
  g1819
  (
    n1907,
    n1807,
    n1442,
    n1423,
    n1568
  );


  xor
  g1820
  (
    n1926,
    n1807,
    n1697,
    n1794,
    n1808
  );


  nor
  g1821
  (
    n1916,
    n1684,
    n1825,
    n1622,
    n1640
  );


  nor
  g1822
  (
    n1896,
    n1823,
    n1501,
    n1527,
    n1389
  );


  xor
  g1823
  (
    n1859,
    n1616,
    n1693,
    n1480,
    n1560
  );


  xnor
  g1824
  (
    n1840,
    n1675,
    n1731,
    n1593,
    n1487
  );


  xnor
  g1825
  (
    n1944,
    n1607,
    n1719,
    n1750,
    n1789
  );


  nor
  g1826
  (
    n1930,
    n1540,
    n1462,
    n1803,
    n1387
  );


  and
  g1827
  (
    n1831,
    n1634,
    n1710,
    n1809,
    n1649
  );


  and
  g1828
  (
    n1904,
    n1802,
    n1526,
    n1650,
    n1624
  );


  xor
  g1829
  (
    n1910,
    n1541,
    n1500,
    n1587,
    n1544
  );


  xor
  g1830
  (
    n1873,
    n1797,
    n1805,
    n1465,
    n1586
  );


  or
  g1831
  (
    n1920,
    n1601,
    n1795,
    n1687,
    n1804
  );


  xnor
  g1832
  (
    n1869,
    n1729,
    n1497,
    n1553,
    n1657
  );


  or
  g1833
  (
    n1887,
    n1819,
    n1623,
    n1817,
    n1645
  );


  xor
  g1834
  (
    n1900,
    n1579,
    n1548,
    n1749,
    n1393
  );


  or
  g1835
  (
    KeyWire_0_6,
    n1779,
    n1820,
    n1476,
    n1612
  );


  or
  g1836
  (
    n1841,
    n1673,
    n1776,
    n1827,
    n1576
  );


  or
  g1837
  (
    n1919,
    n1754,
    n1775,
    n1805,
    n1654
  );


  xor
  g1838
  (
    n1908,
    n1631,
    n1452,
    n1698,
    n1603
  );


  and
  g1839
  (
    n1936,
    n1399,
    n1391,
    n1814,
    n1605
  );


  xor
  g1840
  (
    n1953,
    n1592,
    n1744,
    n1786,
    n1664
  );


  xor
  g1841
  (
    n1885,
    n1787,
    n1388,
    n1449,
    n1801
  );


  xor
  g1842
  (
    n1847,
    n1798,
    n1691,
    n1514,
    n1679
  );


  xnor
  g1843
  (
    n1892,
    n1415,
    n1709,
    n1825,
    n1826
  );


  xnor
  g1844
  (
    n1923,
    n1819,
    n1545,
    n1717,
    n1690
  );


  nor
  g1845
  (
    n1911,
    n1680,
    n1791,
    n1582,
    n1600
  );


  xor
  g1846
  (
    n1867,
    n1453,
    n1795,
    n1565,
    n1419
  );


  nor
  g1847
  (
    n1861,
    n1507,
    n1407,
    n1461,
    n1794
  );


  and
  g1848
  (
    n1934,
    n1412,
    n1470,
    n1815,
    n1425
  );


  xor
  g1849
  (
    n1862,
    n1620,
    n1824,
    n1828,
    n1424
  );


  xor
  g1850
  (
    n1852,
    n1522,
    n1525,
    n1813,
    n1792
  );


  xor
  g1851
  (
    n1928,
    n1633,
    n1793,
    n1451,
    n1610
  );


  xnor
  g1852
  (
    n1834,
    n1433,
    n1641,
    n1584,
    n1796
  );


  nand
  g1853
  (
    n1952,
    n1450,
    n1824,
    n1655,
    n1444
  );


  or
  g1854
  (
    n1835,
    n1737,
    n1543,
    n1598,
    n1695
  );


  nor
  g1855
  (
    n1851,
    n1663,
    n1395,
    n1783,
    n1520
  );


  or
  g1856
  (
    n1837,
    n1483,
    n1400,
    n1723,
    n1630
  );


  xor
  g1857
  (
    n1949,
    n1384,
    n1386,
    n946,
    n1531
  );


  and
  g1858
  (
    n1922,
    n1676,
    n1828,
    n1557,
    n1827
  );


  xnor
  g1859
  (
    n1954,
    n146,
    n1689,
    n1428,
    n1806
  );


  nor
  g1860
  (
    n1871,
    n1704,
    n1529,
    n1536,
    n146
  );


  or
  g1861
  (
    n1864,
    n1702,
    n1608,
    n1551,
    n1632
  );


  or
  g1862
  (
    n1925,
    n1468,
    n1647,
    n1809,
    n145
  );


  xor
  g1863
  (
    n1945,
    n1778,
    n1441,
    n1705,
    n1817
  );


  nand
  g1864
  (
    n1897,
    n1552,
    n1429,
    n1542,
    n1826
  );


  nor
  g1865
  (
    n1921,
    n1475,
    n1604,
    n946,
    n1459
  );


  nor
  g1866
  (
    n1950,
    n1707,
    n1523,
    n1596,
    n1401
  );


  xor
  g1867
  (
    n1937,
    n1473,
    n1660,
    n1495,
    n1578
  );


  and
  g1868
  (
    n1838,
    n1621,
    n1590,
    n1829,
    n1782
  );


  xor
  g1869
  (
    n1938,
    n1738,
    n1588,
    n1797,
    n1785
  );


  nor
  g1870
  (
    n1941,
    n1591,
    n1477,
    n758,
    n1739
  );


  nand
  g1871
  (
    n1888,
    n1443,
    n1491,
    n1637,
    n1678
  );


  nor
  g1872
  (
    n1850,
    n1518,
    n1615,
    n1589,
    n1486
  );


  xor
  g1873
  (
    n1854,
    n1812,
    n1741,
    n1736,
    n1818
  );


  xor
  g1874
  (
    n1948,
    n1625,
    n1580,
    n1509,
    n1667
  );


  or
  g1875
  (
    n1898,
    n1516,
    n1505,
    n1550,
    n1668
  );


  xor
  g1876
  (
    n1878,
    n1517,
    n1484,
    n1478,
    n946
  );


  xor
  g1877
  (
    n1857,
    n1774,
    n1562,
    n1427,
    n1671
  );


  and
  g1878
  (
    KeyWire_0_25,
    n1790,
    n1385,
    n1510,
    n1494
  );


  and
  g1879
  (
    n1833,
    n1639,
    n1437,
    n1781,
    n1492
  );


  or
  g1880
  (
    n1893,
    n1570,
    n1555,
    n1688,
    n1554
  );


  nand
  g1881
  (
    n1844,
    n1569,
    n1445,
    n1563,
    n1446
  );


  xor
  g1882
  (
    n1935,
    n1822,
    n1829,
    n1458,
    n1669
  );


  xor
  g1883
  (
    n1924,
    n1519,
    n1735,
    n1804,
    n757
  );


  nor
  g1884
  (
    n1883,
    n1703,
    n1397,
    n1493,
    n1422
  );


  nor
  g1885
  (
    n1903,
    n1583,
    n1408,
    n1811,
    n1820
  );


  nor
  g1886
  (
    n1855,
    n1699,
    n1471,
    n1672,
    n1777
  );


  xnor
  g1887
  (
    n1905,
    n1485,
    n1466,
    n1413,
    n1464
  );


  and
  g1888
  (
    n1866,
    n1558,
    n1722,
    n1390,
    n1472
  );


  xor
  g1889
  (
    n1863,
    n1504,
    n1751,
    n1559,
    n1594
  );


  or
  g1890
  (
    n1917,
    n1789,
    n1816,
    n1474,
    n1692
  );


  xor
  g1891
  (
    n1891,
    n1430,
    n1662,
    n1417,
    n1506
  );


  or
  g1892
  (
    n1858,
    n1643,
    n1821,
    n1595,
    n1436
  );


  xor
  g1893
  (
    n1846,
    n1511,
    n1567,
    n1635,
    n1431
  );


  xor
  g1894
  (
    n1951,
    n1447,
    n1496,
    n1481,
    n1490
  );


  or
  g1895
  (
    n1902,
    n1609,
    n1747,
    n1817,
    n1611
  );


  or
  g1896
  (
    n1839,
    n1685,
    n1440,
    n1681,
    n1798
  );


  or
  g1897
  (
    n1957,
    n1666,
    n1821,
    n1820,
    n1670
  );


  or
  g1898
  (
    n1874,
    n1785,
    n1602,
    n1629,
    n1828
  );


  and
  g1899
  (
    n1889,
    n1777,
    n1614,
    n1411,
    n1825
  );


  xnor
  g1900
  (
    n1956,
    n1792,
    n1402,
    n1784,
    n1665
  );


  or
  g1901
  (
    n1895,
    n1788,
    n146,
    n1775,
    n1708
  );


  and
  g1902
  (
    n1849,
    n1524,
    n1727,
    n1535,
    n1732
  );


  or
  g1903
  (
    n1879,
    n1528,
    n1457,
    n1455,
    n1513
  );


  and
  g1904
  (
    n1929,
    n1571,
    n946,
    n1448,
    n1636
  );


  and
  g1905
  (
    n1870,
    n1720,
    n1743,
    n1824,
    n1786
  );


  or
  g1906
  (
    n1880,
    n1502,
    n1463,
    n1572,
    n1556
  );


  xnor
  g1907
  (
    n1946,
    n1538,
    n1752,
    n1549,
    n1815
  );


  and
  g1908
  (
    n1886,
    n1456,
    n1432,
    n1482,
    n1714
  );


  xnor
  g1909
  (
    n1940,
    n1821,
    n1753,
    n1628,
    n1734
  );


  and
  g1910
  (
    n1939,
    n1701,
    n1597,
    n1405,
    n1748
  );


  or
  g1911
  (
    n1875,
    n1653,
    n1577,
    n1746,
    n1694
  );


  nand
  g1912
  (
    n1853,
    n1409,
    n1659,
    n1799,
    n1796
  );


  xnor
  g1913
  (
    n1901,
    n1686,
    n1521,
    n1651,
    n1706
  );


  nand
  g1914
  (
    n1881,
    n1784,
    n1606,
    n1813,
    n146
  );


  xor
  g1915
  (
    KeyWire_0_2,
    n1512,
    n1532,
    n1814,
    n1806
  );


  xnor
  g1916
  (
    n1912,
    n1392,
    n1779,
    n1816,
    n1479
  );


  or
  g1917
  (
    n1894,
    n1410,
    n1646,
    n1787,
    n1547
  );


  xor
  g1918
  (
    n1918,
    n1421,
    n1823,
    n1619,
    n1728
  );


  or
  g1919
  (
    n1942,
    n1715,
    n1788,
    n1581,
    n1642
  );


  nor
  g1920
  (
    KeyWire_0_54,
    n1416,
    n1404,
    n1539,
    n1626
  );


  or
  g1921
  (
    n1872,
    n1439,
    n1454,
    n1638,
    n1460
  );


  and
  g1922
  (
    n1943,
    n1515,
    n1733,
    n1627,
    n1711
  );


  nand
  g1923
  (
    KeyWire_0_10,
    n1674,
    n1530,
    n1818,
    n1499
  );


  nor
  g1924
  (
    n1868,
    n1791,
    n1783,
    n1599,
    n1700
  );


  xor
  g1925
  (
    n1995,
    n1834,
    n775,
    n1893,
    n817
  );


  and
  g1926
  (
    n2010,
    n1830,
    n762,
    n820,
    n786
  );


  and
  g1927
  (
    n2013,
    n805,
    n1896,
    n763,
    n1868
  );


  xor
  g1928
  (
    n1994,
    n822,
    n797,
    n1882,
    n1895
  );


  and
  g1929
  (
    n1958,
    n862,
    n1954,
    n1929,
    n773
  );


  and
  g1930
  (
    n1999,
    n1885,
    n1859,
    n1948,
    n1837
  );


  xor
  g1931
  (
    n1983,
    n836,
    n841,
    n864,
    n850
  );


  xor
  g1932
  (
    n2006,
    n837,
    n1899,
    n1866,
    n1857
  );


  xor
  g1933
  (
    n1963,
    n764,
    n829,
    n809,
    n1840
  );


  nand
  g1934
  (
    n1997,
    n828,
    n1924,
    n1922,
    n802
  );


  xnor
  g1935
  (
    n1991,
    n1841,
    n1853,
    n1928,
    n1874
  );


  and
  g1936
  (
    n1986,
    n814,
    n1887,
    n839,
    n1911
  );


  xnor
  g1937
  (
    n2016,
    n819,
    n1955,
    n1873,
    n799
  );


  xnor
  g1938
  (
    n2008,
    n1867,
    n846,
    n816,
    n791
  );


  and
  g1939
  (
    n2009,
    n1860,
    n1943,
    n794,
    n778
  );


  xnor
  g1940
  (
    n2015,
    n1903,
    n1915,
    n770,
    n857
  );


  nand
  g1941
  (
    n2014,
    n813,
    n821,
    n1862,
    n1890
  );


  xnor
  g1942
  (
    n1976,
    n1869,
    n868,
    n790,
    n1888
  );


  and
  g1943
  (
    n1969,
    n843,
    n803,
    n1855,
    n826
  );


  and
  g1944
  (
    n1984,
    n1880,
    n1925,
    n870,
    n845
  );


  xor
  g1945
  (
    n1988,
    n801,
    n842,
    n1864,
    n781
  );


  nor
  g1946
  (
    n1978,
    n1849,
    n1956,
    n1953,
    n761
  );


  xnor
  g1947
  (
    n1967,
    n1920,
    n1898,
    n1883,
    n1884
  );


  nand
  g1948
  (
    n2017,
    n1901,
    n830,
    n1886,
    n766
  );


  nor
  g1949
  (
    n1965,
    n804,
    n1905,
    n1847,
    n1832
  );


  xor
  g1950
  (
    n2001,
    n1909,
    n834,
    n1831,
    n772
  );


  nand
  g1951
  (
    n2003,
    n1846,
    n1845,
    n865,
    n1892
  );


  nand
  g1952
  (
    n1979,
    n760,
    n838,
    n840,
    n815
  );


  nand
  g1953
  (
    n1968,
    n1937,
    n811,
    n1930,
    n796
  );


  xor
  g1954
  (
    n1989,
    n1900,
    n860,
    n769,
    n784
  );


  and
  g1955
  (
    n2005,
    n1833,
    n1916,
    n1839,
    n861
  );


  or
  g1956
  (
    n2004,
    n1945,
    n1940,
    n1904,
    n780
  );


  xnor
  g1957
  (
    n1970,
    n1854,
    n1894,
    n793,
    n852
  );


  xnor
  g1958
  (
    n1993,
    n1856,
    n806,
    n1835,
    n1912
  );


  xnor
  g1959
  (
    n2002,
    n1889,
    n800,
    n808,
    n825
  );


  and
  g1960
  (
    n1973,
    n1913,
    n1861,
    n1842,
    n789
  );


  or
  g1961
  (
    n1998,
    n818,
    n810,
    n782,
    n774
  );


  and
  g1962
  (
    n1980,
    n1897,
    n1951,
    n1875,
    n1942
  );


  and
  g1963
  (
    n1962,
    n831,
    n787,
    n776,
    n863
  );


  and
  g1964
  (
    n1974,
    n1848,
    n824,
    n854,
    n1933
  );


  and
  g1965
  (
    n1981,
    n1947,
    n777,
    n823,
    n783
  );


  nor
  g1966
  (
    n1977,
    n1844,
    n771,
    n1952,
    n1957
  );


  nor
  g1967
  (
    n2012,
    n1935,
    n1858,
    n768,
    n851
  );


  xnor
  g1968
  (
    n2000,
    n1836,
    n1950,
    n1938,
    n1871
  );


  xor
  g1969
  (
    n1996,
    n812,
    n858,
    n853,
    n827
  );


  xnor
  g1970
  (
    n1964,
    n807,
    n1914,
    n1941,
    n1852
  );


  xor
  g1971
  (
    n1985,
    n848,
    n759,
    n1870,
    n1879
  );


  nor
  g1972
  (
    n1975,
    n1863,
    n1902,
    n844,
    n1891
  );


  and
  g1973
  (
    n1961,
    n855,
    n869,
    n856,
    n1936
  );


  xor
  g1974
  (
    KeyWire_0_34,
    n1908,
    n1881,
    n1932,
    n832
  );


  nand
  g1975
  (
    n1982,
    n1927,
    n1851,
    n767,
    n1926
  );


  nor
  g1976
  (
    n2007,
    n1838,
    n859,
    n1907,
    n1878
  );


  or
  g1977
  (
    n1992,
    n1843,
    n765,
    n1949,
    n1931
  );


  xor
  g1978
  (
    n1971,
    n867,
    n1850,
    n833,
    n1921
  );


  xor
  g1979
  (
    n1990,
    n1865,
    n1910,
    n849,
    n847
  );


  or
  g1980
  (
    n1987,
    n1906,
    n1917,
    n1939,
    n788
  );


  nor
  g1981
  (
    n1959,
    n1919,
    n1934,
    n1946,
    n795
  );


  xor
  g1982
  (
    n1960,
    n1872,
    n1918,
    n785,
    n798
  );


  xnor
  g1983
  (
    n1966,
    n1876,
    n792,
    n1923,
    n1877
  );


  or
  g1984
  (
    n2011,
    n1944,
    n779,
    n835,
    n866
  );


  and
  g1985
  (
    n2025,
    n1973,
    n1996,
    n2001,
    n2016
  );


  and
  g1986
  (
    n2019,
    n1984,
    n1976,
    n1962,
    n2002
  );


  nor
  g1987
  (
    n2027,
    n1981,
    n1988,
    n1975,
    n1989
  );


  or
  g1988
  (
    n2032,
    n1985,
    n2012,
    n1969,
    n1958
  );


  xor
  g1989
  (
    n2031,
    n1963,
    n1967,
    n2011,
    n1972
  );


  and
  g1990
  (
    n2023,
    n1978,
    n1987,
    n1961,
    n1983
  );


  xnor
  g1991
  (
    n2030,
    n2010,
    n2003,
    n1980,
    n2004
  );


  nand
  g1992
  (
    n2028,
    n2013,
    n1982,
    n1999,
    n1970
  );


  or
  g1993
  (
    n2020,
    n1971,
    n2014,
    n1960,
    n2009
  );


  xnor
  g1994
  (
    n2026,
    n1990,
    n1965,
    n2017,
    n2000
  );


  nor
  g1995
  (
    n2021,
    n1994,
    n2006,
    n1993,
    n1977
  );


  and
  g1996
  (
    n2018,
    n1964,
    n2007,
    n1997,
    n1974
  );


  xor
  g1997
  (
    n2024,
    n1992,
    n1966,
    n1968,
    n1991
  );


  or
  g1998
  (
    n2022,
    n1979,
    n2008,
    n2005,
    n1995
  );


  nand
  g1999
  (
    n2029,
    n1986,
    n1959,
    n2015,
    n1998
  );


  xor
  KeyGate_0_0
  (
    n690,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1482,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n1906,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n165,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1079,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1264,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n1845,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1175,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n240,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n1793,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1876,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n360,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1255,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n998,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1431,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n1035,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n1339,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n1260,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1688,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1737,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n571,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n396,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n1298,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n999,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n430,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1890,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n782,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n437,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1750,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n502,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n545,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n291,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n462,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n101,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n1972,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n585,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n990,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    n1494,
    keyIn_0_37,
    KeyWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    n896,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n1359,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n1806,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n1069,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n1819,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n1031,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n1569,
    keyIn_0_44,
    KeyWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n148,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n1247,
    KeyNOTWire_0_46
  );


  xor
  KeyGate_0_47
  (
    n1514,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n1250,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n1078,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n1182,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n1454,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n520,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n364,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n1899,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n477,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n326,
    KeyNOTWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n1059,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n1256,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n1758,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n537,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n1508,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n429,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n639,
    KeyNOTWire_0_63
  );


endmodule

