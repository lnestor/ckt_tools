

module Stat_100_49
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n96,
  n107,
  n118,
  n110,
  n98,
  n106,
  n113,
  n121,
  n99,
  n111,
  n109,
  n97,
  n114,
  n93,
  n88,
  n119,
  n116,
  n101,
  n120,
  n103,
  n87,
  n108,
  n104,
  n115,
  n123,
  n128,
  n127,
  n129,
  n126,
  n124,
  n132,
  n131,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n96;
  output n107;
  output n118;
  output n110;
  output n98;
  output n106;
  output n113;
  output n121;
  output n99;
  output n111;
  output n109;
  output n97;
  output n114;
  output n93;
  output n88;
  output n119;
  output n116;
  output n101;
  output n120;
  output n103;
  output n87;
  output n108;
  output n104;
  output n115;
  output n123;
  output n128;
  output n127;
  output n129;
  output n126;
  output n124;
  output n132;
  output n131;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n94;
  wire n95;
  wire n100;
  wire n102;
  wire n105;
  wire n112;
  wire n117;
  wire n122;
  wire n125;
  wire n130;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  buf
  g0
  (
    n39,
    n19
  );


  not
  g1
  (
    KeyWire_0_53,
    n27
  );


  buf
  g2
  (
    KeyWire_0_45,
    n5
  );


  buf
  g3
  (
    KeyWire_0_9,
    n32
  );


  buf
  g4
  (
    KeyWire_0_42,
    n28
  );


  buf
  g5
  (
    KeyWire_0_34,
    n31
  );


  not
  g6
  (
    KeyWire_0_40,
    n21
  );


  not
  g7
  (
    n33,
    n10
  );


  not
  g8
  (
    KeyWire_0_26,
    n15
  );


  buf
  g9
  (
    KeyWire_0_6,
    n2
  );


  buf
  g10
  (
    KeyWire_0_31,
    n3
  );


  buf
  g11
  (
    KeyWire_0_11,
    n26
  );


  buf
  g12
  (
    KeyWire_0_39,
    n29
  );


  buf
  g13
  (
    n35,
    n20
  );


  not
  g14
  (
    KeyWire_0_57,
    n26
  );


  buf
  g15
  (
    n45,
    n16
  );


  buf
  g16
  (
    KeyWire_0_4,
    n26
  );


  buf
  g17
  (
    KeyWire_0_24,
    n24
  );


  not
  g18
  (
    n70,
    n13
  );


  buf
  g19
  (
    n78,
    n8
  );


  not
  g20
  (
    KeyWire_0_54,
    n25
  );


  buf
  g21
  (
    n73,
    n17
  );


  not
  g22
  (
    KeyWire_0_59,
    n24
  );


  buf
  g23
  (
    n72,
    n18
  );


  not
  g24
  (
    n68,
    n28
  );


  not
  g25
  (
    KeyWire_0_55,
    n29
  );


  buf
  g26
  (
    n66,
    n27
  );


  not
  g27
  (
    KeyWire_0_27,
    n11
  );


  buf
  g28
  (
    n67,
    n14
  );


  not
  g29
  (
    n62,
    n12
  );


  buf
  g30
  (
    KeyWire_0_49,
    n25
  );


  buf
  g31
  (
    KeyWire_0_56,
    n4
  );


  buf
  g32
  (
    n65,
    n31
  );


  not
  g33
  (
    KeyWire_0_62,
    n23
  );


  buf
  g34
  (
    n64,
    n30
  );


  buf
  g35
  (
    KeyWire_0_18,
    n27
  );


  buf
  g36
  (
    n82,
    n30
  );


  not
  g37
  (
    KeyWire_0_60,
    n25
  );


  not
  g38
  (
    KeyWire_0_50,
    n22
  );


  not
  g39
  (
    n41,
    n32
  );


  buf
  g40
  (
    n48,
    n29
  );


  buf
  g41
  (
    n71,
    n32
  );


  not
  g42
  (
    KeyWire_0_32,
    n28
  );


  buf
  g43
  (
    KeyWire_0_19,
    n1
  );


  buf
  g44
  (
    n44,
    n6
  );


  not
  g45
  (
    n40,
    n7
  );


  buf
  g46
  (
    KeyWire_0_8,
    n31
  );


  not
  g47
  (
    n50,
    n24
  );


  not
  g48
  (
    KeyWire_0_28,
    n9
  );


  not
  g49
  (
    KeyWire_0_51,
    n30
  );


  or
  g50
  (
    KeyWire_0_41,
    n61,
    n47,
    n36,
    n37
  );


  nand
  g51
  (
    KeyWire_0_38,
    n53,
    n55,
    n78,
    n75
  );


  or
  g52
  (
    n86,
    n73,
    n50,
    n65,
    n51
  );


  nand
  g53
  (
    KeyWire_0_33,
    n39,
    n56,
    n51,
    n37
  );


  xnor
  g54
  (
    KeyWire_0_25,
    n79,
    n50,
    n70,
    n39
  );


  nand
  g55
  (
    KeyWire_0_12,
    n35,
    n63,
    n33,
    n68
  );


  or
  g56
  (
    KeyWire_0_1,
    n40,
    n80,
    n72,
    n39
  );


  nor
  g57
  (
    KeyWire_0_7,
    n73,
    n74,
    n77,
    n38
  );


  nand
  g58
  (
    KeyWire_0_63,
    n44,
    n67,
    n66
  );


  nor
  g59
  (
    KeyWire_0_58,
    n65,
    n45,
    n79,
    n35
  );


  xnor
  g60
  (
    KeyWire_0_14,
    n42,
    n59,
    n60,
    n77
  );


  and
  g61
  (
    n117,
    n55,
    n33,
    n67,
    n58
  );


  or
  g62
  (
    KeyWire_0_5,
    n72,
    n58,
    n56,
    n79
  );


  or
  g63
  (
    KeyWire_0_10,
    n75,
    n66,
    n37,
    n47
  );


  or
  g64
  (
    n97,
    n62,
    n78,
    n48,
    n41
  );


  nor
  g65
  (
    n119,
    n67,
    n52,
    n78
  );


  nand
  g66
  (
    n94,
    n65,
    n70,
    n71
  );


  xor
  g67
  (
    n105,
    n57,
    n59,
    n68,
    n62
  );


  xnor
  g68
  (
    KeyWire_0_23,
    n53,
    n74,
    n63,
    n35
  );


  and
  g69
  (
    n107,
    n61,
    n50,
    n75,
    n76
  );


  and
  g70
  (
    KeyWire_0_17,
    n68,
    n44,
    n71,
    n69
  );


  or
  g71
  (
    KeyWire_0_48,
    n46,
    n68,
    n67,
    n36
  );


  nand
  g72
  (
    n109,
    n64,
    n76,
    n34
  );


  nor
  g73
  (
    KeyWire_0_21,
    n57,
    n44,
    n46,
    n41
  );


  or
  g74
  (
    n118,
    n54,
    n45,
    n41,
    n74
  );


  xor
  g75
  (
    KeyWire_0_30,
    n49,
    n71,
    n46,
    n43
  );


  nand
  g76
  (
    KeyWire_0_22,
    n78,
    n45,
    n40,
    n65
  );


  xnor
  g77
  (
    KeyWire_0_20,
    n76,
    n42,
    n74
  );


  xor
  g78
  (
    KeyWire_0_2,
    n54,
    n49,
    n64,
    n53
  );


  nor
  g79
  (
    n122,
    n66,
    n48,
    n56,
    n70
  );


  nand
  g80
  (
    n96,
    n60,
    n69,
    n77,
    n52
  );


  or
  g81
  (
    KeyWire_0_36,
    n73,
    n38,
    n75,
    n69
  );


  xnor
  g82
  (
    n87,
    n69,
    n71,
    n60,
    n64
  );


  xnor
  g83
  (
    KeyWire_0_52,
    n72,
    n58,
    n64,
    n54
  );


  or
  g84
  (
    KeyWire_0_44,
    n34,
    n36,
    n63,
    n55
  );


  nor
  g85
  (
    KeyWire_0_16,
    n61,
    n73,
    n51,
    n38
  );


  xnor
  g86
  (
    KeyWire_0_46,
    n48,
    n72,
    n77,
    n43
  );


  xnor
  g87
  (
    KeyWire_0_35,
    n63,
    n43,
    n79,
    n40
  );


  xor
  g88
  (
    KeyWire_0_15,
    n62,
    n57,
    n49,
    n47
  );


  xnor
  g89
  (
    KeyWire_0_13,
    n59,
    n34,
    n80,
    n33
  );


  or
  g90
  (
    KeyWire_0_47,
    n81,
    n115,
    n82
  );


  xnor
  g91
  (
    KeyWire_0_37,
    n82,
    n110,
    n117
  );


  xor
  g92
  (
    KeyWire_0_43,
    n120,
    n119,
    n121
  );


  nand
  g93
  (
    n126,
    n81,
    n122,
    n116
  );


  nor
  g94
  (
    KeyWire_0_0,
    n113,
    n80,
    n82
  );


  xor
  g95
  (
    KeyWire_0_29,
    n81,
    n114,
    n109
  );


  xor
  g96
  (
    n130,
    n81,
    n82,
    n80,
    n108
  );


  or
  g97
  (
    n129,
    n112,
    n118,
    n107,
    n111
  );


  buf
  g98
  (
    KeyWire_0_61,
    n130
  );


  buf
  g99
  (
    KeyWire_0_3,
    n129
  );


  xor
  KeyGate_0_0
  (
    n128,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n101,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n110,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n131,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n75,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n120,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n76,
    KeyNOTWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n106,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n63,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n55,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n91,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n81,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n104,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n99,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n121,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n92,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n108,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n89,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n56,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n74,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n90,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n95,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n88,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n113,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n61,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n84,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n46,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n60,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n37,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n124,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n85,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n53,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n57,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n93,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n34,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n111,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n115,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n127,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n114,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    n69,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n51,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n100,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n42,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n123,
    keyIn_0_43,
    KeyWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n83,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n59,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n112,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n125,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n98,
    KeyNOTWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n54,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n77,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n38,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n103,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n49,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n52,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n43,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n47,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n36,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n102,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n58,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n79,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n132,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n80,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n116,
    KeyNOTWire_0_63
  );


endmodule

