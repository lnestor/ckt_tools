// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_105 written by SynthGen on 2021/04/05 11:08:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_105 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n518, n382, n542, n459, n399, n425, n435, n390,
 n407, n445, n383, n362, n487, n553, n426, n403,
 n917, n915, n1022, n1019, n1023, n1030, n1024, n1028,
 n1032, n1025, n1020, n1031, n1021, n1027, n1026, n1029);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n518, n382, n542, n459, n399, n425, n435, n390,
 n407, n445, n383, n362, n487, n553, n426, n403,
 n917, n915, n1022, n1019, n1023, n1030, n1024, n1028,
 n1032, n1025, n1020, n1031, n1021, n1027, n1026, n1029;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n384, n385, n386, n387,
 n388, n389, n391, n392, n393, n394, n395, n396,
 n397, n398, n400, n401, n402, n404, n405, n406,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n427, n428, n429, n430, n431, n432, n433,
 n434, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n460,
 n461, n462, n463, n464, n465, n466, n467, n468,
 n469, n470, n471, n472, n473, n474, n475, n476,
 n477, n478, n479, n480, n481, n482, n483, n484,
 n485, n486, n488, n489, n490, n491, n492, n493,
 n494, n495, n496, n497, n498, n499, n500, n501,
 n502, n503, n504, n505, n506, n507, n508, n509,
 n510, n511, n512, n513, n514, n515, n516, n517,
 n519, n520, n521, n522, n523, n524, n525, n526,
 n527, n528, n529, n530, n531, n532, n533, n534,
 n535, n536, n537, n538, n539, n540, n541, n543,
 n544, n545, n546, n547, n548, n549, n550, n551,
 n552, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n916, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018;

buf  g0 (n63, n1);
buf  g1 (n50, n11);
buf  g2 (n43, n10);
buf  g3 (n105, n20);
not  g4 (n70, n18);
not  g5 (n110, n10);
not  g6 (n44, n19);
not  g7 (n109, n7);
not  g8 (n112, n15);
buf  g9 (n71, n8);
buf  g10 (n79, n13);
buf  g11 (n60, n19);
not  g12 (n95, n13);
buf  g13 (n83, n3);
not  g14 (n34, n5);
not  g15 (n65, n12);
buf  g16 (n38, n18);
buf  g17 (n67, n14);
not  g18 (n107, n15);
not  g19 (n81, n15);
not  g20 (n47, n16);
not  g21 (n96, n19);
not  g22 (n94, n6);
not  g23 (n80, n18);
buf  g24 (n39, n4);
not  g25 (n84, n5);
buf  g26 (n59, n5);
not  g27 (n89, n8);
buf  g28 (n88, n5);
buf  g29 (n75, n6);
buf  g30 (n46, n21);
not  g31 (n49, n11);
not  g32 (n35, n4);
buf  g33 (n92, n6);
not  g34 (n113, n7);
buf  g35 (n48, n9);
not  g36 (n85, n15);
buf  g37 (n55, n13);
not  g38 (n104, n10);
buf  g39 (n86, n17);
not  g40 (n52, n17);
not  g41 (n82, n14);
not  g42 (n114, n10);
buf  g43 (n53, n14);
buf  g44 (n97, n16);
not  g45 (n57, n8);
not  g46 (n111, n17);
not  g47 (n91, n9);
buf  g48 (n77, n20);
buf  g49 (n69, n11);
buf  g50 (n68, n7);
not  g51 (n99, n9);
buf  g52 (n90, n11);
not  g53 (n73, n21);
not  g54 (n33, n12);
not  g55 (n36, n3);
buf  g56 (n72, n3);
not  g57 (n101, n2);
not  g58 (n45, n14);
buf  g59 (n40, n16);
not  g60 (n58, n19);
not  g61 (n51, n6);
buf  g62 (n42, n12);
buf  g63 (n108, n4);
not  g64 (n41, n1);
not  g65 (n54, n7);
buf  g66 (n78, n2);
not  g67 (n100, n13);
buf  g68 (n102, n9);
not  g69 (n103, n8);
not  g70 (n66, n18);
not  g71 (n93, n17);
buf  g72 (n76, n20);
not  g73 (n37, n2);
not  g74 (n56, n3);
buf  g75 (n87, n16);
buf  g76 (n61, n20);
not  g77 (n64, n1);
not  g78 (n106, n1);
not  g79 (n74, n12);
buf  g80 (n98, n4);
buf  g81 (n62, n2);
not  g82 (n296, n62);
not  g83 (n312, n90);
not  g84 (n245, n83);
not  g85 (n220, n48);
buf  g86 (n134, n88);
not  g87 (n284, n45);
not  g88 (n208, n40);
not  g89 (n353, n58);
buf  g90 (n299, n72);
not  g91 (n189, n51);
not  g92 (n146, n60);
buf  g93 (n230, n92);
not  g94 (n244, n44);
not  g95 (n117, n37);
not  g96 (n168, n61);
buf  g97 (n211, n50);
not  g98 (n276, n36);
not  g99 (n138, n40);
not  g100 (n232, n37);
not  g101 (n300, n49);
not  g102 (n221, n39);
buf  g103 (n132, n38);
not  g104 (n185, n75);
buf  g105 (n354, n93);
not  g106 (n147, n66);
buf  g107 (n273, n44);
not  g108 (n202, n53);
buf  g109 (n278, n45);
buf  g110 (n125, n62);
not  g111 (n324, n68);
buf  g112 (n256, n68);
buf  g113 (n348, n76);
not  g114 (n148, n49);
not  g115 (n281, n47);
buf  g116 (n274, n35);
buf  g117 (n163, n82);
buf  g118 (n293, n45);
not  g119 (n340, n83);
not  g120 (n235, n66);
buf  g121 (n266, n37);
buf  g122 (n155, n56);
buf  g123 (n135, n90);
buf  g124 (n257, n72);
not  g125 (n305, n53);
buf  g126 (n292, n85);
buf  g127 (n227, n49);
not  g128 (n175, n60);
not  g129 (n171, n66);
buf  g130 (n314, n86);
not  g131 (n250, n42);
buf  g132 (n166, n86);
not  g133 (n344, n75);
not  g134 (n150, n55);
not  g135 (n294, n94);
not  g136 (n204, n88);
not  g137 (n201, n65);
not  g138 (n288, n93);
not  g139 (n167, n52);
buf  g140 (n270, n77);
buf  g141 (n228, n67);
not  g142 (n269, n61);
not  g143 (n341, n82);
buf  g144 (n213, n79);
buf  g145 (n283, n63);
buf  g146 (n309, n89);
buf  g147 (n291, n52);
buf  g148 (n161, n69);
not  g149 (n355, n93);
not  g150 (n264, n41);
buf  g151 (n303, n34);
not  g152 (n311, n68);
not  g153 (n209, n60);
buf  g154 (n219, n59);
not  g155 (n304, n86);
buf  g156 (n237, n88);
not  g157 (n131, n36);
not  g158 (n316, n72);
buf  g159 (n308, n41);
not  g160 (n216, n47);
buf  g161 (n328, n89);
buf  g162 (n258, n84);
not  g163 (n319, n42);
not  g164 (n289, n67);
buf  g165 (n122, n74);
not  g166 (n149, n39);
not  g167 (n129, n63);
buf  g168 (n287, n44);
not  g169 (n279, n74);
not  g170 (n121, n51);
not  g171 (n246, n43);
not  g172 (n141, n54);
not  g173 (n295, n38);
not  g174 (n140, n94);
not  g175 (n158, n74);
buf  g176 (n322, n34);
not  g177 (n180, n56);
buf  g178 (n210, n85);
not  g179 (n315, n63);
not  g180 (n212, n90);
not  g181 (n162, n56);
not  g182 (n137, n48);
not  g183 (n261, n73);
buf  g184 (n152, n78);
not  g185 (n238, n39);
buf  g186 (n127, n91);
not  g187 (n133, n47);
buf  g188 (n164, n77);
not  g189 (n192, n65);
buf  g190 (n351, n77);
buf  g191 (n318, n70);
buf  g192 (n115, n61);
not  g193 (n145, n79);
buf  g194 (n203, n75);
not  g195 (n259, n81);
not  g196 (n242, n90);
not  g197 (n290, n86);
not  g198 (n345, n70);
not  g199 (n241, n36);
not  g200 (n251, n53);
buf  g201 (n225, n59);
buf  g202 (n275, n54);
buf  g203 (n332, n76);
buf  g204 (n126, n48);
buf  g205 (n352, n58);
buf  g206 (n123, n91);
not  g207 (n174, n50);
not  g208 (n195, n63);
not  g209 (n179, n80);
not  g210 (n249, n69);
not  g211 (n338, n71);
buf  g212 (n160, n42);
not  g213 (n306, n38);
buf  g214 (n247, n60);
buf  g215 (n262, n64);
buf  g216 (n196, n48);
not  g217 (n254, n67);
buf  g218 (n159, n33);
not  g219 (n265, n84);
buf  g220 (n243, n46);
not  g221 (n165, n55);
not  g222 (n329, n91);
buf  g223 (n142, n53);
buf  g224 (n178, n64);
buf  g225 (n120, n62);
buf  g226 (n337, n92);
not  g227 (n226, n35);
buf  g228 (n184, n73);
not  g229 (n233, n37);
buf  g230 (n151, n85);
not  g231 (n218, n43);
not  g232 (n214, n66);
buf  g233 (n325, n83);
not  g234 (n177, n92);
not  g235 (n143, n87);
not  g236 (n130, n57);
not  g237 (n224, n43);
buf  g238 (n191, n80);
not  g239 (n154, n58);
buf  g240 (n116, n80);
not  g241 (n286, n71);
not  g242 (n231, n87);
buf  g243 (n200, n35);
buf  g244 (n326, n73);
not  g245 (n268, n57);
buf  g246 (n118, n41);
buf  g247 (n124, n59);
not  g248 (n298, n42);
buf  g249 (n334, n65);
not  g250 (n183, n88);
not  g251 (n190, n81);
buf  g252 (n248, n71);
buf  g253 (n206, n46);
buf  g254 (n207, n71);
not  g255 (n347, n39);
buf  g256 (n217, n50);
buf  g257 (n157, n33);
not  g258 (n277, n73);
not  g259 (n313, n81);
buf  g260 (n169, n52);
not  g261 (n272, n55);
not  g262 (n139, n79);
buf  g263 (n346, n34);
not  g264 (n282, n94);
not  g265 (n188, n82);
not  g266 (n172, n46);
not  g267 (n343, n78);
buf  g268 (n310, n70);
buf  g269 (n222, n61);
buf  g270 (n255, n82);
not  g271 (n331, n35);
buf  g272 (n156, n94);
not  g273 (n285, n87);
buf  g274 (n170, n89);
buf  g275 (n327, n38);
not  g276 (n128, n75);
buf  g277 (n223, n62);
not  g278 (n229, n77);
not  g279 (n119, n43);
buf  g280 (n215, n50);
buf  g281 (n333, n49);
buf  g282 (n187, n74);
not  g283 (n350, n34);
not  g284 (n271, n84);
not  g285 (n240, n46);
buf  g286 (n323, n76);
not  g287 (n253, n93);
buf  g288 (n349, n64);
buf  g289 (n176, n36);
not  g290 (n181, n41);
not  g291 (n301, n68);
not  g292 (n205, n64);
not  g293 (n267, n52);
not  g294 (n321, n33);
not  g295 (n280, n54);
not  g296 (n297, n56);
not  g297 (n186, n69);
buf  g298 (n336, n80);
buf  g299 (n136, n92);
not  g300 (n335, n51);
buf  g301 (n194, n65);
not  g302 (n197, n47);
buf  g303 (n198, n70);
buf  g304 (n173, n76);
not  g305 (n302, n55);
not  g306 (n193, n78);
not  g307 (n144, n58);
not  g308 (n234, n44);
buf  g309 (n252, n40);
buf  g310 (n317, n51);
buf  g311 (n330, n69);
buf  g312 (n199, n91);
not  g313 (n182, n78);
buf  g314 (n260, n40);
buf  g315 (n356, n67);
buf  g316 (n320, n87);
buf  g317 (n342, n84);
buf  g318 (n153, n54);
not  g319 (n339, n72);
not  g320 (n239, n95);
nand g321 (n263, n81, n79);
and  g322 (n236, n57, n83, n45, n85);
xnor g323 (n307, n33, n89, n59, n57);
or   g324 (n397, n213, n137, n305, n248);
and  g325 (n360, n272, n231, n227, n151);
nor  g326 (n419, n133, n165, n317, n163);
nand g327 (n505, n147, n301, n180, n313);
or   g328 (n441, n212, n163, n215, n198);
and  g329 (n506, n196, n237, n174, n173);
nor  g330 (n547, n224, n232, n193, n168);
nand g331 (n539, n195, n219, n137, n259);
xnor g332 (n518, n220, n264, n139, n224);
or   g333 (n434, n190, n284, n289, n279);
and  g334 (n359, n194, n237, n135, n244);
xnor g335 (n552, n313, n202, n198, n226);
nand g336 (n494, n138, n139, n301, n160);
and  g337 (n430, n282, n164, n188, n211);
or   g338 (n414, n209, n208, n293, n229);
nand g339 (n386, n208, n300, n232, n296);
xnor g340 (n501, n201, n268, n159, n175);
nand g341 (n527, n217, n125, n199, n184);
xor  g342 (n504, n274, n305, n284, n291);
nand g343 (n377, n241, n292, n255, n141);
xor  g344 (n517, n287, n157, n145, n308);
and  g345 (n471, n320, n264, n207, n314);
or   g346 (n451, n237, n249, n159, n162);
nand g347 (n442, n303, n199, n157, n178);
xnor g348 (n523, n228, n214, n136, n300);
xor  g349 (n492, n183, n154, n287, n115);
nand g350 (n387, n131, n251, n268, n219);
xnor g351 (n555, n168, n133, n259, n295);
and  g352 (n376, n158, n191, n314, n186);
xor  g353 (n393, n179, n141, n310, n166);
or   g354 (n440, n149, n215, n218, n221);
nand g355 (n454, n191, n162, n278, n159);
xnor g356 (n367, n195, n148, n228, n185);
xnor g357 (n533, n265, n263, n233, n246);
nand g358 (n467, n204, n309, n130, n301);
xnor g359 (n540, n221, n254, n175, n281);
nand g360 (n511, n283, n171, n162, n252);
and  g361 (n398, n253, n186, n286, n257);
nor  g362 (n390, n284, n188, n219, n250);
or   g363 (n401, n127, n304, n143, n243);
xor  g364 (n381, n149, n160, n144, n261);
nor  g365 (n427, n194, n223, n163, n191);
or   g366 (n514, n296, n258, n138, n247);
nand g367 (n509, n272, n258, n318, n224);
nand g368 (n510, n178, n307, n214, n204);
and  g369 (n546, n156, n203, n245, n239);
xnor g370 (n415, n274, n178, n194, n279);
xor  g371 (n469, n149, n312, n217, n235);
xor  g372 (n529, n253, n316, n269, n281);
nor  g373 (n416, n221, n147, n297, n293);
or   g374 (n364, n262, n130, n267, n192);
nand g375 (n538, n183, n260, n294, n118);
xor  g376 (n537, n267, n176, n315, n233);
xor  g377 (n425, n261, n212, n216, n161);
and  g378 (n490, n311, n249, n209, n164);
xor  g379 (n443, n292, n250, n147, n311);
and  g380 (n524, n256, n140, n224, n226);
or   g381 (n502, n128, n320, n206, n171);
and  g382 (n435, n117, n275, n201, n161);
nor  g383 (n431, n315, n304, n167, n264);
xor  g384 (n358, n300, n185, n126, n306);
nand g385 (n519, n226, n289, n190, n189);
and  g386 (n531, n251, n273, n218, n208);
or   g387 (n495, n173, n127, n144, n235);
nand g388 (n521, n275, n299, n242, n123);
or   g389 (n460, n261, n264, n212, n294);
xor  g390 (n410, n197, n195, n296, n265);
xor  g391 (n497, n145, n305, n126, n221);
and  g392 (n468, n129, n267, n225, n287);
xor  g393 (n421, n306, n182, n127, n277);
xnor g394 (n449, n293, n161, n309, n240);
xnor g395 (n473, n176, n172, n120, n255);
xnor g396 (n369, n171, n183, n204, n124);
and  g397 (n459, n306, n148, n193, n200);
or   g398 (n428, n177, n174, n181, n286);
nand g399 (n450, n239, n266, n136, n257);
xnor g400 (n404, n231, n164, n292, n163);
nand g401 (n389, n236, n230, n176, n273);
xor  g402 (n462, n123, n271, n243, n155);
xor  g403 (n516, n238, n188, n260, n120);
nand g404 (n361, n253, n148, n230, n220);
or   g405 (n500, n190, n172, n151, n316);
nand g406 (n370, n146, n238, n244, n302);
xor  g407 (n423, n251, n254, n185, n261);
nand g408 (n508, n227, n231, n137, n271);
or   g409 (n545, n247, n263, n206, n205);
nand g410 (n422, n281, n270, n218, n257);
nor  g411 (n452, n246, n270, n303, n248);
nand g412 (n405, n288, n284, n238, n234);
xor  g413 (n528, n279, n216, n241, n135);
xnor g414 (n493, n202, n310, n134, n203);
nand g415 (n382, n289, n267, n247, n311);
xnor g416 (n526, n280, n256, n207, n158);
xnor g417 (n420, n303, n211, n229, n225);
and  g418 (n472, n242, n190, n157, n238);
and  g419 (n543, n318, n150, n302, n256);
and  g420 (n515, n154, n281, n260, n191);
xor  g421 (n470, n150, n129, n298, n179);
xnor g422 (n384, n246, n239, n198, n236);
or   g423 (n498, n148, n288, n184, n205);
and  g424 (n365, n182, n226, n280, n275);
xor  g425 (n550, n188, n175, n210, n259);
nand g426 (n433, n130, n162, n248, n202);
xor  g427 (n484, n176, n174, n132, n156);
xnor g428 (n513, n259, n244, n166, n199);
xnor g429 (n407, n311, n151, n132, n203);
xnor g430 (n392, n201, n192, n256, n207);
nor  g431 (n503, n193, n297, n302, n116);
xor  g432 (n388, n195, n287, n266, n225);
and  g433 (n378, n179, n199, n169, n309);
nor  g434 (n463, n159, n143, n152, n296);
xor  g435 (n432, n135, n160, n133, n245);
xor  g436 (n489, n167, n140, n293, n228);
nand g437 (n487, n134, n128, n197, n304);
xor  g438 (n525, n157, n155, n222, n170);
xnor g439 (n448, n165, n169, n290, n317);
xor  g440 (n399, n234, n185, n166, n319);
nor  g441 (n379, n142, n265, n282, n290);
nand g442 (n554, n135, n285, n160, n312);
xor  g443 (n458, n131, n297, n254, n242);
xor  g444 (n411, n290, n230, n181, n215);
xnor g445 (n391, n172, n275, n165, n164);
xnor g446 (n486, n121, n314, n235, n260);
xor  g447 (n402, n245, n262, n292, n145);
or   g448 (n542, n187, n181, n299, n205);
nor  g449 (n474, n270, n258, n288, n172);
xnor g450 (n453, n282, n298, n269, n247);
and  g451 (n373, n317, n147, n268, n228);
nor  g452 (n362, n215, n126, n273, n282);
xor  g453 (n444, n126, n149, n173, n153);
and  g454 (n483, n143, n181, n271, n312);
xnor g455 (n374, n183, n277, n189, n216);
xnor g456 (n412, n309, n182, n294, n202);
nor  g457 (n400, n318, n258, n180, n156);
nor  g458 (n541, n187, n280, n205, n312);
xnor g459 (n480, n206, n142, n121, n129);
nand g460 (n465, n294, n276, n307, n150);
nor  g461 (n408, n189, n252, n239, n169);
xor  g462 (n520, n142, n140, n222, n223);
and  g463 (n475, n132, n317, n129, n196);
nand g464 (n551, n319, n158, n115, n127);
or   g465 (n534, n268, n223, n308, n177);
xnor g466 (n488, n222, n209, n186, n136);
xnor g467 (n438, n213, n285, n130, n194);
nor  g468 (n417, n243, n316, n234, n170);
nor  g469 (n548, n290, n316, n236, n279);
or   g470 (n366, n241, n236, n174, n122);
nand g471 (n395, n263, n295, n125, n198);
or   g472 (n544, n214, n201, n237, n273);
and  g473 (n485, n168, n146, n301, n308);
nand g474 (n530, n278, n276, n227, n308);
nor  g475 (n357, n182, n184, n298, n150);
or   g476 (n457, n153, n289, n213, n138);
or   g477 (n536, n178, n167, n291, n165);
nor  g478 (n549, n142, n229, n200, n197);
nor  g479 (n437, n118, n153, n291, n251);
or   g480 (n396, n179, n153, n154, n197);
xnor g481 (n418, n233, n231, n319, n134);
nand g482 (n522, n192, n288, n180, n286);
nand g483 (n380, n119, n146, n240, n277);
nand g484 (n385, n152, n269, n141, n136);
nor  g485 (n464, n246, n196, n277, n243);
nand g486 (n371, n204, n128, n313, n170);
xnor g487 (n447, n116, n143, n156, n171);
xor  g488 (n507, n210, n214, n310, n207);
or   g489 (n439, n274, n257, n139, n161);
nor  g490 (n496, n240, n170, n193, n285);
xnor g491 (n461, n232, n291, n285, n300);
or   g492 (n479, n152, n184, n269, n212);
xnor g493 (n409, n280, n304, n154, n177);
nor  g494 (n406, n245, n283, n265, n252);
xor  g495 (n477, n145, n196, n255, n319);
xnor g496 (n512, n248, n298, n235, n295);
xnor g497 (n535, n305, n180, n225, n217);
or   g498 (n499, n169, n262, n263, n166);
xor  g499 (n426, n250, n167, n271, n315);
xor  g500 (n375, n187, n152, n217, n318);
xor  g501 (n436, n302, n177, n299, n283);
xor  g502 (n372, n262, n131, n144, n133);
nor  g503 (n363, n232, n266, n134, n155);
or   g504 (n456, n227, n229, n295, n315);
and  g505 (n455, n233, n140, n203, n230);
nor  g506 (n413, n208, n216, n146, n234);
nor  g507 (n394, n187, n220, n117, n306);
or   g508 (n478, n283, n137, n173, n254);
or   g509 (n403, n250, n192, n278, n122);
and  g510 (n466, n297, n314, n244, n249);
xor  g511 (n446, n223, n252, n274, n151);
xor  g512 (n481, n313, n286, n303, n200);
and  g513 (n445, n128, n200, n242, n276);
nand g514 (n476, n131, n144, n218, n138);
xor  g515 (n424, n158, n272, n307, n141);
and  g516 (n429, n220, n175, n206, n189);
and  g517 (n368, n278, n210, n186, n240);
xnor g518 (n553, n209, n213, n310, n249);
xnor g519 (n383, n119, n241, n139, n211);
nand g520 (n491, n255, n270, n210, n299);
xor  g521 (n532, n124, n132, n222, n272);
and  g522 (n482, n168, n211, n219, n155);
nand g523 (n556, n307, n276, n266, n253);
or   g524 (n620, n457, n547, n371, n29);
nand g525 (n648, n520, n540, n449, n337);
xnor g526 (n756, n443, n348, n415, n416);
xor  g527 (n608, n326, n438, n423, n502);
xor  g528 (n565, n497, n488, n462, n518);
nor  g529 (n715, n334, n468, n439, n329);
xnor g530 (n662, n367, n517, n321, n432);
and  g531 (n577, n329, n498, n371, n433);
and  g532 (n622, n400, n364, n22, n424);
or   g533 (n694, n387, n449, n473, n339);
and  g534 (n769, n543, n434, n437, n499);
and  g535 (n579, n472, n369, n389, n476);
or   g536 (n619, n26, n385, n544, n333);
nand g537 (n617, n553, n471, n425, n331);
xnor g538 (n661, n328, n467, n505);
xnor g539 (n765, n459, n456, n523, n439);
nor  g540 (n712, n546, n548, n516, n531);
nand g541 (n602, n531, n334, n365, n28);
or   g542 (n768, n450, n468, n401, n540);
nor  g543 (n777, n343, n403, n395, n459);
and  g544 (n735, n482, n403, n343, n523);
and  g545 (n586, n542, n427, n446, n526);
or   g546 (n611, n101, n473, n407, n511);
nor  g547 (n754, n410, n479, n495, n430);
xor  g548 (n666, n447, n552, n99, n453);
and  g549 (n567, n346, n472, n426, n386);
nand g550 (n750, n437, n491, n492, n400);
nand g551 (n651, n471, n530, n439);
xnor g552 (n612, n370, n544, n502, n500);
and  g553 (n560, n407, n330, n446, n99);
nor  g554 (n582, n536, n419, n511, n490);
and  g555 (n701, n541, n521, n24, n554);
xor  g556 (n587, n497, n493, n400, n31);
and  g557 (n600, n518, n407, n503, n533);
nand g558 (n594, n411, n490, n369, n541);
xor  g559 (n685, n469, n320, n100, n444);
xor  g560 (n734, n445, n397, n327, n496);
xnor g561 (n656, n358, n367, n525, n451);
xnor g562 (n650, n553, n510, n343, n397);
and  g563 (n705, n419, n378, n362, n390);
or   g564 (n764, n97, n535, n100, n329);
or   g565 (n590, n330, n329, n442, n545);
nand g566 (n606, n515, n489, n498, n516);
xor  g567 (n732, n453, n403, n537, n493);
nor  g568 (n779, n411, n528, n448, n434);
and  g569 (n647, n494, n396, n394, n552);
xor  g570 (n737, n440, n537, n346, n349);
xor  g571 (n585, n489, n405, n402, n521);
xor  g572 (n566, n323, n30, n455, n373);
or   g573 (n706, n31, n401, n548, n449);
and  g574 (n702, n372, n400, n551, n408);
xnor g575 (n760, n410, n450, n527);
and  g576 (n634, n420, n461, n440, n30);
nand g577 (n595, n96, n430, n435, n462);
nand g578 (n716, n342, n494, n395, n382);
nand g579 (n564, n414, n24, n337, n442);
nor  g580 (n778, n491, n523, n381, n412);
nand g581 (n676, n339, n388, n359, n428);
nor  g582 (n641, n413, n463, n535, n29);
or   g583 (n758, n27, n478, n96, n336);
and  g584 (n708, n527, n465, n22, n393);
or   g585 (n767, n494, n528, n423, n475);
nor  g586 (n751, n339, n417, n404, n493);
nor  g587 (n629, n433, n429, n21, n381);
nor  g588 (n729, n546, n406, n460);
xor  g589 (n783, n375, n399, n471, n514);
and  g590 (n605, n408, n447, n415, n409);
xnor g591 (n589, n404, n483, n418, n332);
and  g592 (n730, n459, n549, n357, n534);
nor  g593 (n621, n422, n506, n366, n398);
nor  g594 (n637, n446, n425, n344, n380);
and  g595 (n693, n463, n501, n505, n525);
nand g596 (n578, n328, n451, n396, n462);
or   g597 (n686, n374, n435, n527, n455);
or   g598 (n563, n516, n473, n320, n423);
xnor g599 (n644, n331, n538, n532, n443);
xor  g600 (n725, n488, n514, n444, n501);
or   g601 (n678, n348, n495, n508, n532);
xnor g602 (n721, n403, n518, n321, n501);
xnor g603 (n742, n422, n513, n424, n551);
or   g604 (n616, n443, n483, n467, n493);
nand g605 (n575, n409, n456, n455, n542);
xor  g606 (n752, n321, n521, n445, n330);
xnor g607 (n630, n486, n518, n443, n497);
nor  g608 (n749, n504, n411, n341, n398);
xnor g609 (n649, n431, n479, n532, n23);
nand g610 (n741, n337, n498, n531, n417);
and  g611 (n573, n470, n340, n458, n539);
or   g612 (n763, n368, n31, n524, n464);
or   g613 (n659, n499, n473, n505, n446);
nand g614 (n664, n445, n543, n453, n402);
or   g615 (n574, n484, n455, n447, n338);
and  g616 (n653, n531, n543, n469, n472);
xnor g617 (n632, n441, n448, n454, n341);
or   g618 (n633, n537, n99, n440, n429);
or   g619 (n562, n492, n466, n512, n442);
xnor g620 (n727, n418, n533, n492, n396);
or   g621 (n696, n429, n401, n344, n477);
and  g622 (n736, n536, n525, n30, n503);
nand g623 (n603, n441, n523, n549, n345);
nand g624 (n726, n333, n515, n343, n451);
xor  g625 (n709, n342, n519, n347, n529);
nand g626 (n739, n325, n421, n513);
nor  g627 (n609, n376, n477, n480, n461);
xor  g628 (n628, n437, n422, n485, n508);
xor  g629 (n703, n97, n338, n495, n472);
xnor g630 (n627, n522, n420, n524, n431);
nand g631 (n746, n508, n468, n529, n341);
nand g632 (n688, n417, n96, n509, n422);
xnor g633 (n680, n342, n509, n437, n541);
or   g634 (n770, n504, n530, n525);
xor  g635 (n669, n25, n402, n483);
nor  g636 (n720, n474, n504, n360, n480);
nand g637 (n635, n499, n486, n325, n517);
nand g638 (n642, n477, n427, n332, n374);
xnor g639 (n675, n331, n390, n496, n398);
and  g640 (n668, n373, n512, n460, n524);
and  g641 (n569, n344, n101, n413, n428);
xor  g642 (n583, n545, n550, n542, n485);
xnor g643 (n673, n25, n475, n532, n330);
or   g644 (n724, n509, n378, n438, n368);
xor  g645 (n719, n24, n551, n510, n102);
xnor g646 (n618, n456, n95, n444, n397);
nor  g647 (n599, n384, n482, n545, n503);
or   g648 (n631, n470, n511, n29, n456);
or   g649 (n753, n361, n526, n500, n372);
xor  g650 (n652, n364, n539, n322, n418);
and  g651 (n643, n384, n419, n334, n548);
nor  g652 (n707, n462, n370, n460, n435);
nor  g653 (n657, n98, n332, n336, n491);
nand g654 (n782, n481, n380, n467, n375);
xor  g655 (n744, n348, n552, n410, n506);
or   g656 (n593, n510, n449, n102, n508);
or   g657 (n740, n331, n22, n539, n24);
and  g658 (n674, n538, n528, n444, n428);
xor  g659 (n568, n513, n522, n427, n486);
or   g660 (n762, n545, n358, n416, n487);
nor  g661 (n723, n346, n481, n338, n552);
or   g662 (n759, n347, n460, n327, n506);
or   g663 (n717, n379, n438, n491, n359);
nor  g664 (n683, n471, n475, n534, n28);
xnor g665 (n679, n101, n98, n326, n379);
xnor g666 (n646, n447, n549, n543, n345);
xor  g667 (n580, n515, n463, n334, n404);
and  g668 (n667, n414, n429, n326, n457);
nand g669 (n581, n31, n32, n464, n554);
xor  g670 (n601, n490, n335, n533, n463);
and  g671 (n695, n480, n405, n487, n396);
xor  g672 (n614, n324, n499, n551, n410);
and  g673 (n772, n27, n496, n520, n454);
nor  g674 (n626, n436, n328, n489, n496);
and  g675 (n692, n480, n100, n433, n534);
and  g676 (n761, n482, n442, n340, n452);
or   g677 (n636, n519, n327, n476, n424);
xor  g678 (n638, n478, n507, n502, n30);
xnor g679 (n691, n479, n448, n324, n452);
xor  g680 (n597, n519, n399, n393, n395);
nand g681 (n766, n417, n528, n486, n101);
nand g682 (n745, n324, n539, n546, n412);
or   g683 (n698, n494, n340, n500, n428);
nand g684 (n584, n519, n535, n498, n28);
xnor g685 (n610, n363, n484, n406, n21);
xor  g686 (n728, n506, n507, n500, n404);
nand g687 (n558, n341, n464, n323, n465);
xor  g688 (n660, n322, n509, n420, n522);
nor  g689 (n684, n524, n415, n438, n454);
xor  g690 (n592, n432, n481, n469, n391);
nor  g691 (n714, n398, n515, n477, n490);
and  g692 (n718, n399, n448, n345, n349);
nor  g693 (n780, n492, n392, n323, n324);
xor  g694 (n771, n347, n344, n389, n466);
xor  g695 (n604, n526, n336, n432, n408);
xnor g696 (n591, n414, n95, n452, n100);
or   g697 (n623, n453, n411, n335, n365);
nand g698 (n561, n474, n25, n517, n497);
nand g699 (n654, n26, n395, n550, n388);
xnor g700 (n687, n335, n409, n439, n445);
xnor g701 (n624, n452, n360, n327, n383);
and  g702 (n570, n461, n458, n541, n337);
or   g703 (n640, n99, n435, n514, n454);
or   g704 (n748, n501, n421, n431, n28);
nor  g705 (n755, n464, n465, n336, n357);
or   g706 (n690, n507, n489, n502, n366);
nand g707 (n598, n413, n458, n436, n511);
nor  g708 (n559, n32, n419, n26, n425);
nand g709 (n697, n512, n325, n468, n363);
nor  g710 (n775, n459, n426, n96, n485);
nand g711 (n738, n25, n97, n430, n326);
xor  g712 (n639, n516, n478, n26, n482);
and  g713 (n615, n550, n430, n547, n554);
nand g714 (n713, n32, n322, n547, n361);
nand g715 (n663, n377, n391, n457, n538);
nand g716 (n743, n348, n394, n333, n23);
and  g717 (n572, n451, n323, n409, n520);
or   g718 (n710, n434, n421, n414, n426);
xor  g719 (n747, n423, n416, n550, n476);
xnor g720 (n576, n475, n529, n335, n440);
nor  g721 (n670, n549, n32, n362, n397);
nor  g722 (n571, n547, n97, n377, n420);
nor  g723 (n700, n481, n479, n544, n469);
xor  g724 (n699, n465, n553, n421, n349);
xor  g725 (n681, n533, n376, n347, n536);
nand g726 (n757, n441, n425, n540, n488);
nand g727 (n613, n383, n333, n548, n520);
xnor g728 (n645, n441, n487, n98, n434);
nor  g729 (n731, n495, n424, n466, n488);
nand g730 (n596, n457, n485, n514, n385);
and  g731 (n711, n427, n436, n484, n503);
or   g732 (n722, n433, n392, n415, n535);
nand g733 (n625, n458, n412, n401, n483);
xnor g734 (n776, n470, n461, n538, n431);
and  g735 (n655, n405, n27, n321, n349);
and  g736 (n672, n487, n529, n544, n416);
and  g737 (n774, n325, n406, n328, n474);
nor  g738 (n689, n436, n399, n27, n405);
or   g739 (n665, n432, n426, n484, n534);
nand g740 (n682, n470, n474, n408, n540);
nand g741 (n671, n412, n342, n478, n23);
nand g742 (n557, n450, n23, n322, n339);
nor  g743 (n658, n387, n467, n29, n382);
and  g744 (n588, n95, n526, n476, n332);
nand g745 (n773, n527, n407, n536, n542);
nor  g746 (n704, n386, n546, n504, n340);
xor  g747 (n607, n98, n512, n510, n466);
xor  g748 (n781, n346, n522, n413, n418);
nor  g749 (n677, n345, n507, n553, n537);
and  g750 (n733, n338, n22, n517, n521);
or   g751 (n793, n686, n629, n617, n626);
and  g752 (n822, n668, n580, n619, n620);
or   g753 (n808, n670, n678, n567, n689);
xnor g754 (n827, n651, n594, n624, n593);
or   g755 (n812, n608, n105, n690, n637);
and  g756 (n825, n667, n577, n589, n106);
or   g757 (n785, n672, n102, n639, n566);
xor  g758 (n818, n681, n633, n606, n604);
nand g759 (n819, n602, n103, n582, n568);
xor  g760 (n799, n659, n572, n614, n350);
or   g761 (n817, n352, n682, n103, n585);
and  g762 (n811, n104, n597, n351, n592);
xnor g763 (n829, n687, n674, n352, n575);
xor  g764 (n788, n685, n646, n605, n350);
or   g765 (n790, n611, n105, n662, n688);
xnor g766 (n797, n654, n105, n621, n600);
xor  g767 (n820, n644, n652, n667, n627);
and  g768 (n798, n607, n658, n691, n622);
and  g769 (n828, n107, n676, n673);
xor  g770 (n815, n636, n351, n686, n649);
xnor g771 (n802, n102, n685, n578, n642);
nand g772 (n804, n671, n591, n681, n647);
nor  g773 (n807, n668, n106, n351, n666);
nor  g774 (n794, n571, n352, n623, n596);
xor  g775 (n830, n573, n692, n590, n584);
nor  g776 (n787, n616, n350, n680, n625);
xnor g777 (n806, n628, n613, n678, n107);
nor  g778 (n809, n640, n565, n105, n103);
and  g779 (n800, n660, n672, n609, n691);
nor  g780 (n805, n650, n618, n684, n631);
or   g781 (n816, n630, n574, n106, n599);
nor  g782 (n796, n103, n583, n641, n653);
nand g783 (n823, n648, n104, n576, n684);
nor  g784 (n814, n569, n595, n673, n682);
xor  g785 (n813, n689, n645, n670, n665);
or   g786 (n784, n104, n677, n692, n581);
xor  g787 (n824, n107, n352, n615, n688);
and  g788 (n821, n351, n675, n669, n601);
or   g789 (n826, n598, n683, n579, n632);
nor  g790 (n789, n104, n107, n664, n612);
xnor g791 (n786, n661, n106, n663, n677);
nor  g792 (n803, n669, n655, n603, n680);
xor  g793 (n792, n657, n638, n635, n679);
nor  g794 (n810, n690, n634, n610, n675);
nand g795 (n795, n656, n588, n587, n683);
xnor g796 (n791, n687, n674, n586, n643);
xnor g797 (n801, n570, n350, n671, n679);
buf  g798 (n875, n798);
not  g799 (n864, n794);
buf  g800 (n840, n109);
buf  g801 (n847, n805);
buf  g802 (n859, n804);
buf  g803 (n862, n793);
buf  g804 (n865, n114);
buf  g805 (n869, n112);
not  g806 (n844, n113);
buf  g807 (n831, n787);
not  g808 (n832, n108);
not  g809 (n866, n113);
buf  g810 (n836, n111);
buf  g811 (n860, n113);
buf  g812 (n876, n806);
buf  g813 (n849, n787);
buf  g814 (n845, n795);
buf  g815 (n872, n791);
not  g816 (n871, n801);
buf  g817 (n868, n803);
not  g818 (n834, n790);
buf  g819 (n878, n808);
not  g820 (n873, n785);
not  g821 (n877, n795);
not  g822 (n880, n802);
buf  g823 (n870, n109);
buf  g824 (n838, n112);
not  g825 (n848, n803);
buf  g826 (n846, n801);
not  g827 (n835, n788);
buf  g828 (n857, n797);
not  g829 (n861, n793);
buf  g830 (n867, n788);
not  g831 (n841, n112);
not  g832 (n837, n108);
not  g833 (n858, n110);
not  g834 (n853, n792);
not  g835 (n874, n792);
buf  g836 (n850, n807);
buf  g837 (n843, n791);
xnor g838 (n839, n796, n789);
nor  g839 (n856, n112, n808, n790, n108);
nand g840 (n852, n802, n809, n786, n789);
nand g841 (n851, n109, n806, n108, n796);
and  g842 (n863, n109, n799, n804, n785);
nor  g843 (n879, n797, n114, n786, n111);
nor  g844 (n842, n807, n110, n111);
xor  g845 (n855, n784, n110, n805, n798);
nand g846 (n854, n113, n800, n794);
xnor g847 (n833, n799, n111, n114);
nor  g848 (n915, n856, n864, n847, n870);
xnor g849 (n884, n849, n854, n846, n862);
xnor g850 (n886, n851, n853, n849, n836);
and  g851 (n885, n872, n859, n869, n842);
nor  g852 (n900, n849, n861, n854, n871);
nor  g853 (n911, n832, n831, n833, n843);
nand g854 (n904, n850, n856, n852, n869);
or   g855 (n903, n835, n852, n844, n865);
xnor g856 (n896, n864, n833, n834);
nand g857 (n914, n864, n834, n866, n863);
xnor g858 (n891, n845, n861, n841, n865);
nor  g859 (n916, n848, n859, n845, n870);
xnor g860 (n890, n860, n849, n832, n855);
xor  g861 (n881, n862, n855, n837, n840);
or   g862 (n919, n863, n848, n861, n868);
nor  g863 (n920, n854, n845, n855, n862);
xor  g864 (n905, n838, n852, n864, n843);
nand g865 (n902, n857, n843, n842, n868);
nand g866 (n899, n867, n865, n844, n850);
nand g867 (n922, n850, n869, n834, n836);
xor  g868 (n913, n867, n871, n851, n866);
or   g869 (n907, n839, n861, n853, n847);
or   g870 (n906, n841, n857, n858);
and  g871 (n888, n863, n859, n832, n836);
or   g872 (n912, n870, n860, n835, n837);
xor  g873 (n882, n848, n846, n868, n872);
nor  g874 (n889, n866, n837, n853, n839);
nand g875 (n883, n840, n835, n859, n872);
or   g876 (n887, n843, n841, n872, n858);
xnor g877 (n894, n871, n839, n850, n848);
xor  g878 (n909, n835, n836, n860, n866);
xnor g879 (n895, n871, n851, n831, n870);
xnor g880 (n892, n833, n838, n869, n840);
nand g881 (n898, n842, n854, n834, n857);
nand g882 (n921, n867, n852, n858, n841);
and  g883 (n901, n846, n855, n844);
or   g884 (n893, n867, n858, n860, n863);
nand g885 (n917, n847, n862, n840, n873);
or   g886 (n897, n865, n851, n837, n838);
xor  g887 (n918, n868, n845, n839, n856);
or   g888 (n908, n853, n832, n873, n842);
xnor g889 (n910, n847, n846, n838, n856);
xnor g890 (n936, n885, n353, n878, n715);
nand g891 (n925, n877, n874, n719, n704);
xnor g892 (n931, n880, n915, n917, n721);
xnor g893 (n932, n725, n353, n900, n724);
xor  g894 (n955, n896, n724, n708, n701);
nand g895 (n949, n877, n722, n721, n711);
nand g896 (n937, n909, n875, n700, n879);
or   g897 (n959, n695, n356, n702, n694);
and  g898 (n961, n874, n918, n702, n876);
nand g899 (n951, n879, n895, n723, n556);
or   g900 (n926, n355, n875, n697, n889);
nor  g901 (n950, n884, n904, n696, n717);
xor  g902 (n956, n877, n353, n693, n901);
xor  g903 (n940, n880, n712, n911);
or   g904 (n927, n880, n707, n716, n710);
xor  g905 (n948, n354, n709, n718, n903);
nand g906 (n953, n908, n899, n878, n913);
and  g907 (n933, n879, n716, n887, n556);
xor  g908 (n943, n696, n705, n888, n706);
nor  g909 (n928, n704, n922, n700, n698);
or   g910 (n935, n897, n722, n919, n723);
nand g911 (n962, n891, n906, n709, n698);
nor  g912 (n934, n910, n555, n705, n898);
xnor g913 (n923, n878, n878, n355, n894);
nand g914 (n947, n720, n354, n876);
nor  g915 (n960, n905, n556, n880, n356);
nand g916 (n954, n875, n916, n694, n902);
xnor g917 (n924, n714, n355, n877, n875);
or   g918 (n939, n717, n713, n555);
nand g919 (n929, n719, n879, n695, n715);
xnor g920 (n942, n714, n876, n873, n893);
nor  g921 (n941, n554, n883, n706, n707);
xnor g922 (n944, n720, n701, n555, n699);
xor  g923 (n938, n699, n873, n555, n556);
xor  g924 (n958, n708, n718, n892, n356);
nand g925 (n952, n874, n693, n354, n912);
and  g926 (n930, n354, n921, n703, n356);
or   g927 (n957, n886, n874, n355, n907);
nand g928 (n946, n914, n890, n920, n697);
and  g929 (n945, n710, n711, n353, n703);
nor  g930 (n1010, n941, n930, n827, n748);
and  g931 (n987, n732, n764, n932, n774);
nor  g932 (n976, n933, n761, n951, n952);
nand g933 (n1016, n955, n753, n778, n777);
xnor g934 (n977, n742, n823, n819, n945);
or   g935 (n998, n953, n735, n947, n959);
xnor g936 (n969, n775, n812, n954, n952);
or   g937 (n979, n811, n778, n751, n735);
xor  g938 (n972, n934, n779, n936, n738);
xor  g939 (n964, n926, n768, n781, n772);
or   g940 (n986, n809, n738, n938, n759);
xor  g941 (n1001, n825, n943, n762, n814);
or   g942 (n993, n755, n754, n816, n744);
xor  g943 (n1003, n780, n743, n820, n948);
nor  g944 (n980, n741, n771, n824, n773);
xor  g945 (n971, n731, n820, n828, n783);
xor  g946 (n1015, n960, n810, n734, n782);
and  g947 (n997, n955, n775, n821, n928);
and  g948 (n1012, n727, n773, n761, n956);
nor  g949 (n978, n756, n827, n829, n822);
xnor g950 (n983, n729, n925, n733, n817);
nor  g951 (n1000, n733, n757, n931, n772);
xnor g952 (n1018, n740, n754, n760, n826);
xnor g953 (n985, n755, n927, n781, n828);
xor  g954 (n996, n748, n825, n935, n951);
xnor g955 (n1009, n745, n741, n771, n830);
xnor g956 (n992, n962, n818, n817, n739);
and  g957 (n1013, n929, n760, n937, n737);
and  g958 (n994, n746, n756, n774, n757);
or   g959 (n1006, n822, n734, n946, n777);
or   g960 (n968, n942, n766, n725, n826);
or   g961 (n963, n766, n769, n758, n816);
xnor g962 (n1007, n954, n780, n749, n763);
xnor g963 (n990, n949, n783, n744, n823);
and  g964 (n975, n812, n811, n818, n739);
nor  g965 (n1008, n813, n737, n939, n751);
xor  g966 (n974, n728, n747, n829, n957);
and  g967 (n988, n815, n829, n923, n727);
and  g968 (n1017, n736, n828, n731, n776);
nor  g969 (n981, n747, n813, n764, n752);
xor  g970 (n984, n762, n940, n948, n827);
nor  g971 (n1005, n749, n829, n726);
and  g972 (n995, n830, n770, n736, n776);
xnor g973 (n965, n759, n830, n959, n769);
xor  g974 (n966, n824, n746, n830, n752);
xor  g975 (n989, n949, n740, n770, n958);
nand g976 (n1004, n767, n810, n730, n815);
xnor g977 (n982, n729, n758, n742, n950);
nor  g978 (n970, n768, n950, n765, n728);
xnor g979 (n999, n814, n767, n753, n782);
nor  g980 (n1011, n956, n962, n961);
xor  g981 (n1014, n750, n953, n819, n924);
and  g982 (n973, n827, n730, n957, n743);
and  g983 (n1002, n944, n763, n821, n960);
and  g984 (n991, n958, n750, n745, n765);
nand g985 (n967, n828, n947, n779, n732);
or   g986 (n1026, n967, n1008, n977, n1006);
nand g987 (n1027, n985, n1011, n997, n1004);
nor  g988 (n1031, n995, n1002, n1000, n966);
xor  g989 (n1029, n980, n989, n1003, n964);
xor  g990 (n1024, n994, n1005, n1007, n1012);
and  g991 (n1032, n976, n1013, n983, n998);
xor  g992 (n1022, n992, n990, n969, n968);
and  g993 (n1030, n1018, n986, n970, n1015);
and  g994 (n1025, n1014, n988, n1001, n978);
and  g995 (n1020, n972, n982, n971, n987);
xor  g996 (n1023, n984, n981, n991, n999);
xnor g997 (n1019, n1010, n1017, n974, n965);
xor  g998 (n1021, n979, n1009, n973, n1016);
xnor g999 (n1028, n963, n996, n993, n975);
endmodule
