// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_821_382 written by SynthGen on 2021/05/24 19:48:30
module Stat_821_382( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19,
 n571, n767, n766, n764, n760, n765, n770, n762,
 n768, n771, n759, n758, n796, n798, n803, n802,
 n811, n815, n828, n832, n833, n839, n840);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19;

output n571, n767, n766, n764, n760, n765, n770, n762,
 n768, n771, n759, n758, n796, n798, n803, n802,
 n811, n815, n828, n832, n833, n839, n840;

wire n20, n21, n22, n23, n24, n25, n26, n27,
 n28, n29, n30, n31, n32, n33, n34, n35,
 n36, n37, n38, n39, n40, n41, n42, n43,
 n44, n45, n46, n47, n48, n49, n50, n51,
 n52, n53, n54, n55, n56, n57, n58, n59,
 n60, n61, n62, n63, n64, n65, n66, n67,
 n68, n69, n70, n71, n72, n73, n74, n75,
 n76, n77, n78, n79, n80, n81, n82, n83,
 n84, n85, n86, n87, n88, n89, n90, n91,
 n92, n93, n94, n95, n96, n97, n98, n99,
 n100, n101, n102, n103, n104, n105, n106, n107,
 n108, n109, n110, n111, n112, n113, n114, n115,
 n116, n117, n118, n119, n120, n121, n122, n123,
 n124, n125, n126, n127, n128, n129, n130, n131,
 n132, n133, n134, n135, n136, n137, n138, n139,
 n140, n141, n142, n143, n144, n145, n146, n147,
 n148, n149, n150, n151, n152, n153, n154, n155,
 n156, n157, n158, n159, n160, n161, n162, n163,
 n164, n165, n166, n167, n168, n169, n170, n171,
 n172, n173, n174, n175, n176, n177, n178, n179,
 n180, n181, n182, n183, n184, n185, n186, n187,
 n188, n189, n190, n191, n192, n193, n194, n195,
 n196, n197, n198, n199, n200, n201, n202, n203,
 n204, n205, n206, n207, n208, n209, n210, n211,
 n212, n213, n214, n215, n216, n217, n218, n219,
 n220, n221, n222, n223, n224, n225, n226, n227,
 n228, n229, n230, n231, n232, n233, n234, n235,
 n236, n237, n238, n239, n240, n241, n242, n243,
 n244, n245, n246, n247, n248, n249, n250, n251,
 n252, n253, n254, n255, n256, n257, n258, n259,
 n260, n261, n262, n263, n264, n265, n266, n267,
 n268, n269, n270, n271, n272, n273, n274, n275,
 n276, n277, n278, n279, n280, n281, n282, n283,
 n284, n285, n286, n287, n288, n289, n290, n291,
 n292, n293, n294, n295, n296, n297, n298, n299,
 n300, n301, n302, n303, n304, n305, n306, n307,
 n308, n309, n310, n311, n312, n313, n314, n315,
 n316, n317, n318, n319, n320, n321, n322, n323,
 n324, n325, n326, n327, n328, n329, n330, n331,
 n332, n333, n334, n335, n336, n337, n338, n339,
 n340, n341, n342, n343, n344, n345, n346, n347,
 n348, n349, n350, n351, n352, n353, n354, n355,
 n356, n357, n358, n359, n360, n361, n362, n363,
 n364, n365, n366, n367, n368, n369, n370, n371,
 n372, n373, n374, n375, n376, n377, n378, n379,
 n380, n381, n382, n383, n384, n385, n386, n387,
 n388, n389, n390, n391, n392, n393, n394, n395,
 n396, n397, n398, n399, n400, n401, n402, n403,
 n404, n405, n406, n407, n408, n409, n410, n411,
 n412, n413, n414, n415, n416, n417, n418, n419,
 n420, n421, n422, n423, n424, n425, n426, n427,
 n428, n429, n430, n431, n432, n433, n434, n435,
 n436, n437, n438, n439, n440, n441, n442, n443,
 n444, n445, n446, n447, n448, n449, n450, n451,
 n452, n453, n454, n455, n456, n457, n458, n459,
 n460, n461, n462, n463, n464, n465, n466, n467,
 n468, n469, n470, n471, n472, n473, n474, n475,
 n476, n477, n478, n479, n480, n481, n482, n483,
 n484, n485, n486, n487, n488, n489, n490, n491,
 n492, n493, n494, n495, n496, n497, n498, n499,
 n500, n501, n502, n503, n504, n505, n506, n507,
 n508, n509, n510, n511, n512, n513, n514, n515,
 n516, n517, n518, n519, n520, n521, n522, n523,
 n524, n525, n526, n527, n528, n529, n530, n531,
 n532, n533, n534, n535, n536, n537, n538, n539,
 n540, n541, n542, n543, n544, n545, n546, n547,
 n548, n549, n550, n551, n552, n553, n554, n555,
 n556, n557, n558, n559, n560, n561, n562, n563,
 n564, n565, n566, n567, n568, n569, n570, n572,
 n573, n574, n575, n576, n577, n578, n579, n580,
 n581, n582, n583, n584, n585, n586, n587, n588,
 n589, n590, n591, n592, n593, n594, n595, n596,
 n597, n598, n599, n600, n601, n602, n603, n604,
 n605, n606, n607, n608, n609, n610, n611, n612,
 n613, n614, n615, n616, n617, n618, n619, n620,
 n621, n622, n623, n624, n625, n626, n627, n628,
 n629, n630, n631, n632, n633, n634, n635, n636,
 n637, n638, n639, n640, n641, n642, n643, n644,
 n645, n646, n647, n648, n649, n650, n651, n652,
 n653, n654, n655, n656, n657, n658, n659, n660,
 n661, n662, n663, n664, n665, n666, n667, n668,
 n669, n670, n671, n672, n673, n674, n675, n676,
 n677, n678, n679, n680, n681, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n701, n702, n703, n704, n705, n706, n707, n708,
 n709, n710, n711, n712, n713, n714, n715, n716,
 n717, n718, n719, n720, n721, n722, n723, n724,
 n725, n726, n727, n728, n729, n730, n731, n732,
 n733, n734, n735, n736, n737, n738, n739, n740,
 n741, n742, n743, n744, n745, n746, n747, n748,
 n749, n750, n751, n752, n753, n754, n755, n756,
 n757, n761, n763, n769, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n794, n795, n797, n799, n800, n801,
 n804, n805, n806, n807, n808, n809, n810, n812,
 n813, n814, n816, n817, n818, n819, n820, n821,
 n822, n823, n824, n825, n826, n827, n829, n830,
 n831, n834, n835, n836, n837, n838;

buf  g0 (n32, n7);
buf  g1 (n89, n9);
buf  g2 (n64, n18);
buf  g3 (n42, n6);
not  g4 (n54, n6);
buf  g5 (n90, n15);
buf  g6 (n22, n19);
buf  g7 (n67, n19);
buf  g8 (n36, n17);
not  g9 (n71, n3);
buf  g10 (n33, n12);
not  g11 (n52, n2);
buf  g12 (n44, n10);
buf  g13 (n28, n19);
buf  g14 (n20, n16);
buf  g15 (n46, n18);
not  g16 (n94, n8);
buf  g17 (n25, n17);
not  g18 (n24, n8);
buf  g19 (n91, n13);
buf  g20 (n70, n6);
not  g21 (n57, n16);
not  g22 (n84, n12);
not  g23 (n85, n10);
buf  g24 (n48, n1);
buf  g25 (n88, n14);
buf  g26 (n50, n2);
buf  g27 (n75, n13);
buf  g28 (n30, n7);
not  g29 (n79, n2);
not  g30 (n56, n18);
buf  g31 (n77, n14);
not  g32 (n87, n4);
not  g33 (n51, n5);
not  g34 (n39, n14);
not  g35 (n45, n8);
not  g36 (n23, n9);
buf  g37 (n72, n18);
not  g38 (n93, n6);
buf  g39 (n73, n14);
not  g40 (n78, n12);
buf  g41 (n60, n15);
buf  g42 (n41, n4);
not  g43 (n61, n8);
not  g44 (n63, n17);
buf  g45 (n95, n2);
not  g46 (n81, n4);
not  g47 (n34, n11);
buf  g48 (n38, n5);
not  g49 (n40, n3);
not  g50 (n59, n13);
buf  g51 (n69, n16);
buf  g52 (n35, n9);
buf  g53 (n27, n3);
not  g54 (n68, n5);
not  g55 (n76, n4);
not  g56 (n49, n17);
not  g57 (n47, n11);
buf  g58 (n58, n15);
not  g59 (n37, n7);
not  g60 (n83, n11);
buf  g61 (n82, n15);
not  g62 (n21, n7);
not  g63 (n86, n10);
buf  g64 (n74, n1);
not  g65 (n65, n12);
not  g66 (n29, n1);
buf  g67 (n43, n13);
buf  g68 (n55, n3);
not  g69 (n66, n11);
not  g70 (n53, n10);
not  g71 (n31, n19);
buf  g72 (n80, n1);
not  g73 (n62, n9);
buf  g74 (n26, n16);
not  g75 (n92, n5);
buf  g76 (n339, n73);
buf  g77 (n137, n23);
not  g78 (n219, n26);
buf  g79 (n112, n20);
buf  g80 (n125, n53);
buf  g81 (n244, n70);
not  g82 (n308, n69);
not  g83 (n202, n24);
not  g84 (n126, n70);
buf  g85 (n325, n59);
buf  g86 (n225, n37);
not  g87 (n314, n71);
not  g88 (n114, n81);
not  g89 (n343, n59);
buf  g90 (n212, n85);
not  g91 (n352, n71);
buf  g92 (n159, n22);
buf  g93 (n139, n21);
buf  g94 (n122, n41);
buf  g95 (n100, n23);
buf  g96 (n330, n42);
buf  g97 (n111, n21);
buf  g98 (n163, n58);
buf  g99 (n151, n28);
not  g100 (n260, n90);
not  g101 (n318, n47);
buf  g102 (n108, n88);
not  g103 (n104, n82);
buf  g104 (n121, n48);
buf  g105 (n147, n84);
not  g106 (n350, n89);
not  g107 (n313, n25);
not  g108 (n205, n22);
buf  g109 (n256, n37);
buf  g110 (n110, n88);
buf  g111 (n236, n46);
not  g112 (n182, n48);
buf  g113 (n134, n49);
buf  g114 (n243, n67);
not  g115 (n266, n67);
not  g116 (n380, n68);
not  g117 (n262, n55);
buf  g118 (n378, n61);
buf  g119 (n310, n38);
buf  g120 (n162, n77);
buf  g121 (n117, n36);
buf  g122 (n297, n87);
not  g123 (n257, n43);
not  g124 (n322, n31);
not  g125 (n274, n60);
buf  g126 (n319, n55);
buf  g127 (n148, n54);
buf  g128 (n311, n76);
buf  g129 (n307, n74);
buf  g130 (n127, n45);
not  g131 (n279, n34);
not  g132 (n269, n58);
buf  g133 (n255, n39);
not  g134 (n119, n36);
buf  g135 (n200, n24);
not  g136 (n348, n43);
not  g137 (n193, n69);
buf  g138 (n99, n67);
buf  g139 (n216, n41);
buf  g140 (n240, n36);
not  g141 (n101, n38);
not  g142 (n364, n30);
not  g143 (n359, n47);
buf  g144 (n340, n25);
not  g145 (n323, n42);
buf  g146 (n238, n39);
buf  g147 (n250, n50);
not  g148 (n172, n33);
buf  g149 (n227, n22);
buf  g150 (n189, n29);
not  g151 (n371, n87);
not  g152 (n267, n70);
buf  g153 (n366, n76);
buf  g154 (n261, n31);
not  g155 (n303, n70);
not  g156 (n105, n64);
not  g157 (n334, n66);
buf  g158 (n210, n51);
not  g159 (n248, n80);
buf  g160 (n146, n40);
not  g161 (n342, n74);
buf  g162 (n284, n34);
not  g163 (n177, n56);
not  g164 (n170, n80);
buf  g165 (n191, n45);
not  g166 (n158, n68);
not  g167 (n188, n46);
not  g168 (n229, n82);
buf  g169 (n135, n82);
not  g170 (n226, n24);
buf  g171 (n301, n86);
buf  g172 (n192, n34);
buf  g173 (n120, n49);
buf  g174 (n207, n30);
buf  g175 (n259, n60);
buf  g176 (n183, n66);
not  g177 (n263, n60);
buf  g178 (n252, n40);
buf  g179 (n335, n22);
buf  g180 (n357, n50);
buf  g181 (n295, n43);
buf  g182 (n345, n35);
not  g183 (n132, n85);
buf  g184 (n312, n51);
buf  g185 (n361, n40);
buf  g186 (n228, n55);
not  g187 (n247, n52);
buf  g188 (n285, n85);
not  g189 (n201, n31);
buf  g190 (n116, n49);
buf  g191 (n195, n75);
buf  g192 (n281, n59);
not  g193 (n254, n86);
not  g194 (n271, n24);
buf  g195 (n234, n32);
not  g196 (n346, n63);
buf  g197 (n175, n75);
not  g198 (n242, n35);
buf  g199 (n180, n46);
not  g200 (n272, n44);
buf  g201 (n290, n84);
buf  g202 (n324, n30);
not  g203 (n153, n45);
not  g204 (n160, n54);
not  g205 (n249, n88);
buf  g206 (n245, n35);
buf  g207 (n214, n63);
not  g208 (n265, n50);
buf  g209 (n376, n28);
not  g210 (n333, n74);
not  g211 (n296, n32);
not  g212 (n231, n77);
buf  g213 (n369, n56);
not  g214 (n109, n46);
not  g215 (n161, n62);
not  g216 (n143, n52);
not  g217 (n288, n89);
not  g218 (n302, n53);
not  g219 (n351, n28);
buf  g220 (n298, n45);
not  g221 (n115, n79);
not  g222 (n239, n66);
not  g223 (n128, n90);
not  g224 (n203, n47);
buf  g225 (n331, n91);
buf  g226 (n184, n81);
not  g227 (n332, n78);
buf  g228 (n190, n86);
buf  g229 (n368, n61);
buf  g230 (n118, n65);
buf  g231 (n168, n57);
buf  g232 (n291, n82);
not  g233 (n321, n71);
not  g234 (n251, n65);
buf  g235 (n338, n21);
buf  g236 (n198, n47);
not  g237 (n140, n39);
not  g238 (n370, n44);
buf  g239 (n286, n77);
not  g240 (n181, n87);
not  g241 (n154, n31);
buf  g242 (n336, n56);
buf  g243 (n379, n57);
buf  g244 (n164, n77);
not  g245 (n123, n43);
buf  g246 (n316, n20);
not  g247 (n133, n40);
buf  g248 (n169, n33);
not  g249 (n152, n72);
buf  g250 (n98, n54);
buf  g251 (n355, n71);
buf  g252 (n241, n74);
not  g253 (n328, n61);
not  g254 (n171, n62);
not  g255 (n194, n37);
buf  g256 (n309, n80);
buf  g257 (n124, n38);
buf  g258 (n329, n64);
not  g259 (n280, n84);
not  g260 (n317, n67);
not  g261 (n287, n61);
buf  g262 (n213, n59);
not  g263 (n220, n73);
not  g264 (n344, n20);
not  g265 (n306, n51);
not  g266 (n327, n83);
not  g267 (n206, n23);
not  g268 (n320, n76);
not  g269 (n142, n87);
not  g270 (n246, n27);
not  g271 (n103, n69);
buf  g272 (n315, n33);
not  g273 (n136, n34);
not  g274 (n326, n73);
buf  g275 (n337, n79);
buf  g276 (n106, n91);
buf  g277 (n282, n42);
buf  g278 (n157, n29);
buf  g279 (n372, n80);
buf  g280 (n176, n26);
not  g281 (n173, n29);
buf  g282 (n349, n83);
not  g283 (n197, n32);
not  g284 (n299, n66);
not  g285 (n382, n78);
buf  g286 (n276, n72);
not  g287 (n373, n36);
buf  g288 (n365, n64);
not  g289 (n300, n72);
buf  g290 (n293, n65);
not  g291 (n253, n78);
not  g292 (n199, n42);
buf  g293 (n196, n25);
not  g294 (n289, n54);
not  g295 (n150, n32);
buf  g296 (n341, n75);
not  g297 (n165, n53);
not  g298 (n167, n64);
buf  g299 (n264, n89);
not  g300 (n149, n78);
not  g301 (n278, n23);
buf  g302 (n97, n65);
not  g303 (n374, n53);
buf  g304 (n347, n63);
buf  g305 (n131, n84);
not  g306 (n353, n85);
buf  g307 (n178, n56);
buf  g308 (n96, n30);
buf  g309 (n179, n72);
not  g310 (n218, n29);
not  g311 (n215, n27);
buf  g312 (n367, n86);
not  g313 (n208, n39);
buf  g314 (n305, n91);
not  g315 (n277, n81);
buf  g316 (n155, n58);
buf  g317 (n356, n41);
not  g318 (n230, n52);
buf  g319 (n360, n35);
not  g320 (n221, n62);
buf  g321 (n224, n27);
not  g322 (n283, n89);
not  g323 (n145, n58);
buf  g324 (n294, n37);
not  g325 (n102, n26);
not  g326 (n363, n73);
not  g327 (n268, n48);
not  g328 (n237, n68);
buf  g329 (n107, n21);
not  g330 (n113, n51);
buf  g331 (n375, n88);
buf  g332 (n235, n79);
buf  g333 (n304, n26);
not  g334 (n174, n83);
not  g335 (n129, n68);
buf  g336 (n233, n33);
buf  g337 (n258, n38);
not  g338 (n377, n62);
buf  g339 (n187, n57);
buf  g340 (n186, n57);
not  g341 (n144, n63);
buf  g342 (n381, n79);
buf  g343 (n138, n69);
buf  g344 (n292, n90);
buf  g345 (n275, n44);
not  g346 (n362, n60);
buf  g347 (n217, n81);
not  g348 (n141, n76);
buf  g349 (n211, n25);
not  g350 (n166, n55);
not  g351 (n354, n50);
buf  g352 (n222, n20);
buf  g353 (n358, n83);
not  g354 (n130, n41);
not  g355 (n204, n28);
not  g356 (n273, n52);
not  g357 (n232, n27);
not  g358 (n209, n90);
buf  g359 (n223, n75);
buf  g360 (n185, n48);
buf  g361 (n270, n49);
buf  g362 (n156, n44);
buf  g363 (n493, n134);
buf  g364 (n496, n101);
buf  g365 (n428, n107);
not  g366 (n384, n208);
buf  g367 (n441, n129);
not  g368 (n474, n123);
not  g369 (n407, n138);
buf  g370 (n383, n111);
not  g371 (n410, n113);
buf  g372 (n417, n136);
not  g373 (n397, n195);
not  g374 (n477, n178);
buf  g375 (n473, n110);
not  g376 (n448, n96);
not  g377 (n423, n179);
buf  g378 (n475, n186);
not  g379 (n454, n166);
buf  g380 (n486, n102);
buf  g381 (n433, n106);
not  g382 (n459, n148);
buf  g383 (n395, n172);
not  g384 (n430, n205);
not  g385 (n385, n156);
buf  g386 (n472, n190);
not  g387 (n398, n127);
not  g388 (n427, n118);
not  g389 (n403, n109);
buf  g390 (n438, n206);
not  g391 (n451, n202);
not  g392 (n396, n177);
not  g393 (n445, n146);
buf  g394 (n484, n188);
buf  g395 (n447, n126);
buf  g396 (n411, n97);
buf  g397 (n388, n122);
not  g398 (n401, n204);
buf  g399 (n429, n100);
buf  g400 (n476, n198);
not  g401 (n482, n183);
buf  g402 (n439, n163);
not  g403 (n400, n170);
buf  g404 (n444, n191);
buf  g405 (n487, n207);
buf  g406 (n413, n193);
buf  g407 (n479, n135);
not  g408 (n471, n174);
not  g409 (n489, n209);
buf  g410 (n440, n168);
not  g411 (n488, n104);
buf  g412 (n421, n200);
buf  g413 (n463, n171);
buf  g414 (n446, n120);
not  g415 (n394, n133);
buf  g416 (n412, n162);
not  g417 (n453, n128);
buf  g418 (n452, n151);
not  g419 (n460, n119);
buf  g420 (n478, n192);
not  g421 (n455, n203);
not  g422 (n422, n189);
not  g423 (n409, n181);
not  g424 (n464, n141);
buf  g425 (n490, n167);
not  g426 (n443, n132);
buf  g427 (n420, n196);
buf  g428 (n461, n152);
not  g429 (n434, n153);
not  g430 (n470, n98);
not  g431 (n457, n160);
not  g432 (n492, n155);
buf  g433 (n469, n164);
buf  g434 (n418, n149);
buf  g435 (n467, n161);
not  g436 (n416, n142);
not  g437 (n495, n115);
buf  g438 (n392, n103);
buf  g439 (n432, n150);
buf  g440 (n419, n199);
buf  g441 (n481, n185);
not  g442 (n437, n180);
not  g443 (n480, n112);
not  g444 (n415, n182);
buf  g445 (n431, n157);
buf  g446 (n390, n154);
not  g447 (n386, n173);
buf  g448 (n425, n99);
not  g449 (n414, n158);
buf  g450 (n435, n175);
not  g451 (n442, n130);
not  g452 (n402, n184);
buf  g453 (n462, n147);
buf  g454 (n391, n131);
buf  g455 (n456, n187);
buf  g456 (n408, n121);
buf  g457 (n436, n159);
buf  g458 (n491, n108);
not  g459 (n387, n124);
not  g460 (n494, n145);
not  g461 (n449, n117);
buf  g462 (n458, n143);
buf  g463 (n405, n144);
not  g464 (n404, n125);
not  g465 (n483, n169);
buf  g466 (n468, n197);
buf  g467 (n465, n137);
buf  g468 (n399, n114);
buf  g469 (n424, n140);
buf  g470 (n393, n116);
buf  g471 (n450, n201);
buf  g472 (n426, n105);
not  g473 (n466, n194);
buf  g474 (n406, n165);
not  g475 (n485, n176);
buf  g476 (n389, n139);
or   g477 (n501, n423, n417, n386, n416);
nand g478 (n518, n413, n387, n391, n403);
xor  g479 (n508, n420, n385, n425, n394);
and  g480 (n510, n422, n397, n393, n390);
nand g481 (n511, n408, n419, n389, n406);
nand g482 (n507, n399, n415, n422, n384);
xnor g483 (n500, n412, n397, n387, n392);
xor  g484 (n515, n386, n405, n425, n407);
nand g485 (n505, n409, n409, n408, n388);
nand g486 (n498, n418, n398, n399, n407);
nor  g487 (n509, n394, n412, n393, n402);
and  g488 (n506, n417, n426, n398, n411);
or   g489 (n503, n388, n413, n400);
xnor g490 (n497, n384, n396, n427, n410);
or   g491 (n517, n396, n406, n418, n421);
xnor g492 (n513, n395, n421, n416, n426);
or   g493 (n499, n404, n385, n420, n403);
xnor g494 (n502, n390, n424, n404, n401);
or   g495 (n516, n391, n419, n415, n423);
nor  g496 (n512, n410, n401, n383, n392);
nand g497 (n504, n389, n402, n414, n405);
nand g498 (n514, n395, n411, n414, n424);
buf  g499 (n522, n499);
buf  g500 (n528, n504);
not  g501 (n523, n502);
not  g502 (n521, n507);
buf  g503 (n520, n500);
not  g504 (n519, n498);
not  g505 (n527, n501);
not  g506 (n525, n506);
buf  g507 (n524, n503);
xor  g508 (n526, n505, n497);
not  g509 (n537, n524);
buf  g510 (n531, n520);
buf  g511 (n533, n521);
buf  g512 (n536, n523);
not  g513 (n532, n525);
not  g514 (n529, n522);
buf  g515 (n535, n519);
buf  g516 (n534, n527);
not  g517 (n530, n526);
not  g518 (n542, n214);
buf  g519 (n546, n533);
xnor g520 (n539, n229, n530, n213, n242);
xnor g521 (n550, n235, n210, n530, n220);
and  g522 (n548, n225, n238, n221, n533);
xor  g523 (n544, n234, n532, n228);
xnor g524 (n540, n240, n239, n534, n212);
xnor g525 (n547, n223, n232, n237, n533);
nand g526 (n538, n211, n224, n215, n533);
or   g527 (n545, n230, n529, n218, n227);
or   g528 (n549, n241, n219, n531, n217);
or   g529 (n541, n236, n216, n226, n531);
nor  g530 (n543, n222, n534, n233, n231);
nand g531 (n562, n445, n538, n543, n430);
nand g532 (n554, n244, n445, n539, n439);
nand g533 (n560, n541, n443, n540, n428);
xor  g534 (n557, n544, n443, n542, n245);
or   g535 (n558, n444, n541, n441, n538);
nor  g536 (n552, n543, n431, n247, n539);
nor  g537 (n551, n429, n540, n440, n434);
xor  g538 (n559, n435, n436, n440, n446);
or   g539 (n555, n433, n442, n432, n542);
or   g540 (n561, n544, n437, n246, n248);
and  g541 (n564, n434, n442, n545, n437);
xor  g542 (n563, n441, n430, n428, n433);
and  g543 (n565, n439, n429, n243, n427);
nor  g544 (n553, n436, n431, n432, n435);
nand g545 (n556, n446, n438, n444);
xnor g546 (n569, n563, n565, n553, n253);
nand g547 (n581, n551, n272, n258, n289);
xor  g548 (n577, n264, n259, n260, n292);
nor  g549 (n566, n254, n564, n558, n559);
xor  g550 (n575, n556, n280, n285, n279);
nor  g551 (n576, n283, n273, n261, n278);
xor  g552 (n580, n267, n266, n296, n557);
xor  g553 (n579, n269, n562, n277, n560);
nor  g554 (n578, n270, n286, n565, n555);
nand g555 (n567, n295, n282, n256, n255);
or   g556 (n574, n291, n249, n271, n288);
and  g557 (n570, n268, n275, n265, n294);
xor  g558 (n572, n257, n561, n284, n274);
xor  g559 (n571, n552, n251, n262, n293);
nor  g560 (n573, n554, n290, n281, n250);
or   g561 (n568, n252, n263, n276, n287);
buf  g562 (n613, n450);
buf  g563 (n619, n476);
buf  g564 (n607, n473);
not  g565 (n597, n570);
not  g566 (n609, n573);
not  g567 (n594, n453);
buf  g568 (n588, n465);
buf  g569 (n623, n576);
buf  g570 (n617, n458);
not  g571 (n601, n460);
not  g572 (n583, n567);
not  g573 (n602, n465);
buf  g574 (n608, n572);
not  g575 (n626, n468);
not  g576 (n598, n451);
not  g577 (n604, n458);
xor  g578 (n621, n471, n468);
nand g579 (n620, n469, n572, n452, n463);
xor  g580 (n618, n478, n472, n484, n464);
nor  g581 (n589, n460, n575, n482, n566);
or   g582 (n593, n489, n568, n455, n478);
xnor g583 (n603, n487, n570, n566, n568);
xor  g584 (n610, n575, n574, n450, n571);
xor  g585 (n615, n453, n566, n492, n569);
nor  g586 (n611, n576, n467, n569);
nand g587 (n595, n470, n577, n483, n459);
nand g588 (n587, n577, n571, n463, n459);
or   g589 (n614, n487, n448, n477, n485);
nand g590 (n605, n488, n572, n452, n569);
nor  g591 (n627, n451, n569, n457, n567);
xor  g592 (n592, n568, n573, n570, n477);
nand g593 (n628, n577, n462, n574, n479);
or   g594 (n599, n456, n490, n447, n480);
or   g595 (n586, n568, n474, n567, n489);
xor  g596 (n591, n574, n461, n466, n475);
nor  g597 (n590, n469, n449, n472, n576);
or   g598 (n585, n479, n571, n481);
xnor g599 (n596, n490, n572, n475, n575);
or   g600 (n582, n456, n576, n574, n491);
xnor g601 (n584, n470, n571, n454, n573);
xor  g602 (n600, n567, n471, n491, n575);
or   g603 (n616, n447, n455, n573, n486);
nor  g604 (n612, n464, n474, n473, n482);
and  g605 (n606, n485, n454, n476, n577);
xnor g606 (n622, n483, n449, n484, n570);
nor  g607 (n624, n488, n462, n457, n486);
or   g608 (n625, n448, n466, n461, n480);
not  g609 (n630, n591);
buf  g610 (n635, n584);
not  g611 (n633, n597);
not  g612 (n638, n583);
not  g613 (n629, n598);
buf  g614 (n637, n593);
nor  g615 (n631, n589, n590);
and  g616 (n636, n587, n596, n595, n598);
xnor g617 (n634, n596, n586, n592, n594);
or   g618 (n632, n595, n588, n597, n585);
buf  g619 (n642, n606);
buf  g620 (n647, n606);
nor  g621 (n641, n637, n610);
nand g622 (n640, n631, n630, n607, n632);
xnor g623 (n648, n638, n603, n599, n602);
nor  g624 (n649, n492, n638, n602, n600);
nand g625 (n646, n604, n599, n600, n608);
or   g626 (n639, n607, n601, n610);
nor  g627 (n643, n603, n605, n608, n635);
xor  g628 (n644, n604, n609, n605);
and  g629 (n645, n633, n629, n634, n636);
not  g630 (n666, n643);
not  g631 (n670, n308);
buf  g632 (n657, n322);
not  g633 (n678, n508);
not  g634 (n689, n642);
buf  g635 (n668, n309);
not  g636 (n677, n611);
buf  g637 (n671, n648);
not  g638 (n655, n647);
not  g639 (n676, n641);
not  g640 (n669, n649);
not  g641 (n674, n648);
buf  g642 (n662, n644);
not  g643 (n651, n319);
buf  g644 (n686, n327);
not  g645 (n681, n645);
buf  g646 (n656, n303);
not  g647 (n688, n649);
buf  g648 (n690, n640);
not  g649 (n665, n644);
not  g650 (n658, n611);
buf  g651 (n683, n647);
buf  g652 (n679, n616);
buf  g653 (n692, n645);
not  g654 (n652, n648);
not  g655 (n663, n318);
nor  g656 (n673, n644, n639);
nor  g657 (n672, n617, n613, n534, n301);
xnor g658 (n661, n512, n614, n314, n642);
xnor g659 (n687, n649, n614, n640, n325);
xnor g660 (n653, n513, n643, n645, n305);
nand g661 (n680, n640, n641, n509, n647);
and  g662 (n650, n615, n320, n317, n311);
nand g663 (n660, n315, n612, n298);
nor  g664 (n691, n639, n645, n646, n321);
or   g665 (n675, n534, n299, n313, n312);
and  g666 (n684, n642, n646, n511, n310);
xnor g667 (n667, n640, n326, n641, n324);
and  g668 (n664, n510, n297, n646, n316);
nand g669 (n685, n647, n306, n646, n323);
or   g670 (n693, n307, n649, n643, n304);
and  g671 (n654, n644, n615, n616, n639);
nor  g672 (n659, n643, n642, n613, n641);
xnor g673 (n682, n300, n639, n648, n302);
buf  g674 (n710, n336);
buf  g675 (n728, n674);
buf  g676 (n734, n680);
buf  g677 (n711, n535);
not  g678 (n736, n496);
buf  g679 (n703, n659);
buf  g680 (n696, n665);
not  g681 (n733, n689);
buf  g682 (n708, n670);
not  g683 (n724, n494);
buf  g684 (n741, n618);
buf  g685 (n718, n536);
not  g686 (n705, n536);
not  g687 (n697, n658);
not  g688 (n720, n693);
not  g689 (n706, n681);
xnor g690 (n699, n656, n683);
xnor g691 (n716, n679, n686, n682, n662);
nand g692 (n702, n673, n545, n680, n332);
nand g693 (n719, n536, n518, n687, n671);
and  g694 (n713, n339, n328, n653, n514);
nor  g695 (n709, n537, n689, n676, n549);
nand g696 (n739, n684, n692, n579, n650);
nor  g697 (n725, n677, n495, n651, n493);
xnor g698 (n715, n618, n338, n688, n546);
xor  g699 (n722, n342, n550, n330, n678);
xnor g700 (n695, n578, n684, n516, n580);
xnor g701 (n737, n537, n621, n691);
xnor g702 (n738, n578, n334, n495, n654);
xnor g703 (n700, n675, n580, n617, n579);
nand g704 (n723, n691, n682, n528, n331);
xor  g705 (n714, n579, n547, n535, n620);
nor  g706 (n727, n676, n536, n664, n672);
nor  g707 (n704, n335, n620, n578, n344);
nand g708 (n698, n579, n546, n687, n535);
nand g709 (n701, n580, n690, n581, n679);
xnor g710 (n726, n681, n581, n693, n91);
xnor g711 (n735, n580, n669, n667, n494);
xnor g712 (n717, n690, n550, n581, n677);
nand g713 (n730, n652, n329, n663, n678);
nor  g714 (n740, n537, n581, n333, n340);
xnor g715 (n732, n661, n578, n493, n548);
or   g716 (n712, n657, n692, n337, n686);
xnor g717 (n729, n619, n549, n683, n537);
and  g718 (n694, n548, n341, n666, n517);
nor  g719 (n731, n660, n515, n619, n535);
or   g720 (n721, n343, n668, n688, n685);
nor  g721 (n707, n685, n496, n547, n655);
not  g722 (n744, n694);
buf  g723 (n742, n696);
xor  g724 (n743, n695, n697);
or   g725 (n745, n744, n742, n743);
not  g726 (n746, n745);
not  g727 (n747, n745);
not  g728 (n755, n746);
not  g729 (n749, n746);
not  g730 (n753, n747);
not  g731 (n751, n746);
buf  g732 (n748, n746);
not  g733 (n750, n747);
buf  g734 (n752, n747);
not  g735 (n754, n747);
nor  g736 (n770, n626, n703, n748, n713);
or   g737 (n760, n729, n705, n626, n727);
and  g738 (n764, n754, n721, n753, n752);
xnor g739 (n758, n750, n708, n719, n753);
or   g740 (n762, n720, n710, n716, n699);
nand g741 (n768, n623, n711, n751, n715);
and  g742 (n771, n755, n702, n725, n751);
or   g743 (n763, n622, n714, n754, n700);
nand g744 (n766, n712, n717, n730, n698);
and  g745 (n767, n624, n709, n752, n724);
nor  g746 (n756, n728, n750, n726, n731);
nand g747 (n761, n749, n701, n754, n723);
and  g748 (n769, n749, n748, n718, n707);
or   g749 (n757, n755, n623, n624, n704);
xor  g750 (n759, n722, n625, n755, n706);
nor  g751 (n765, n755, n622, n625, n732);
not  g752 (n773, n767);
buf  g753 (n775, n770);
not  g754 (n776, n771);
buf  g755 (n772, n345);
nand g756 (n774, n768, n769);
buf  g757 (n789, n346);
buf  g758 (n777, n776);
not  g759 (n787, n93);
not  g760 (n792, n92);
buf  g761 (n793, n351);
not  g762 (n778, n774);
not  g763 (n784, n354);
buf  g764 (n791, n93);
xnor g765 (n794, n773, n353);
or   g766 (n783, n94, n734, n735, n347);
or   g767 (n779, n348, n352, n95, n772);
xor  g768 (n790, n93, n94, n92, n776);
xor  g769 (n786, n94, n776, n349, n92);
or   g770 (n788, n774, n775, n773);
nand g771 (n781, n773, n94, n772, n775);
xor  g772 (n785, n93, n95, n774);
nand g773 (n782, n773, n774, n95, n775);
nor  g774 (n780, n733, n350, n776, n92);
not  g775 (n795, n778);
not  g776 (n798, n779);
buf  g777 (n797, n780);
not  g778 (n796, n777);
nand g779 (n799, n781, n797, n798, n780);
buf  g780 (n800, n799);
buf  g781 (n801, n799);
not  g782 (n803, n801);
and  g783 (n802, n801, n800, n355);
and  g784 (n804, n801, n357, n800, n356);
nand g785 (n805, n804, n782, n781);
buf  g786 (n807, n805);
not  g787 (n809, n784);
nand g788 (n808, n783, n358, n805, n785);
nand g789 (n806, n784, n783, n805);
buf  g790 (n810, n806);
not  g791 (n811, n806);
or   g792 (n812, n811, n359);
buf  g793 (n814, n812);
buf  g794 (n813, n812);
and  g795 (n815, n785, n786, n812);
and  g796 (n816, n814, n787, n788, n815);
nor  g797 (n817, n788, n627, n787, n786);
nand g798 (n819, n807, n807, n816, n366);
and  g799 (n825, n361, n365, n808, n809);
xnor g800 (n820, n360, n809, n817);
xor  g801 (n821, n370, n816, n807);
xnor g802 (n818, n364, n817, n368, n816);
xnor g803 (n823, n369, n808, n362, n809);
xor  g804 (n822, n808, n808, n627, n817);
xnor g805 (n824, n807, n367, n363, n817);
or   g806 (n827, n823, n825, n824);
nand g807 (n826, n822, n821, n824, n820);
xnor g808 (n828, n819, n371, n372, n818);
xor  g809 (n830, n790, n789, n828);
nor  g810 (n829, n827, n790, n791);
or   g811 (n832, n793, n830, n738, n792);
or   g812 (n831, n829, n793, n736, n830);
nor  g813 (n833, n830, n830, n737, n792);
and  g814 (n834, n374, n373, n628, n833);
or   g815 (n837, n376, n375, n380, n382);
nand g816 (n836, n381, n834, n379, n377);
nor  g817 (n838, n739, n740, n834, n628);
xor  g818 (n835, n794, n378, n834);
nand g819 (n839, n837, n837, n838, n836);
and  g820 (n840, n741, n835, n838, n794);
endmodule
