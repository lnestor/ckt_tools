

module Stat_923_296
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n75,
  n35,
  n54,
  n22,
  n67,
  n21,
  n45,
  n87,
  n56,
  n52,
  n23,
  n29,
  n84,
  n92,
  n33,
  n487,
  n637,
  n635,
  n640,
  n634,
  n802,
  n799,
  n914,
  n940,
  n936,
  n939,
  n938,
  n942,
  n941,
  n937,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n75;output n35;output n54;output n22;output n67;output n21;output n45;output n87;output n56;output n52;output n23;output n29;output n84;output n92;output n33;output n487;output n637;output n635;output n640;output n634;output n802;output n799;output n914;output n940;output n936;output n939;output n938;output n942;output n941;output n937;
  wire n20;wire n24;wire n25;wire n26;wire n27;wire n28;wire n30;wire n31;wire n32;wire n34;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n53;wire n55;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n85;wire n86;wire n88;wire n89;wire n90;wire n91;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n636;wire n638;wire n639;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n800;wire n801;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyNOTWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyNOTWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n37,
    n6
  );


  not
  g1
  (
    n57,
    n2
  );


  not
  g2
  (
    n79,
    n18
  );


  not
  g3
  (
    n26,
    n15
  );


  not
  g4
  (
    n88,
    n16
  );


  not
  g5
  (
    n49,
    n12
  );


  buf
  g6
  (
    n74,
    n13
  );


  not
  g7
  (
    n80,
    n6
  );


  buf
  g8
  (
    n82,
    n10
  );


  not
  g9
  (
    n70,
    n7
  );


  not
  g10
  (
    n63,
    n1
  );


  not
  g11
  (
    n62,
    n11
  );


  not
  g12
  (
    n39,
    n19
  );


  not
  g13
  (
    n87,
    n7
  );


  buf
  g14
  (
    n34,
    n3
  );


  not
  g15
  (
    n89,
    n19
  );


  buf
  g16
  (
    n25,
    n14
  );


  not
  g17
  (
    KeyWire_0_10,
    n4
  );


  buf
  g18
  (
    n29,
    n8
  );


  buf
  g19
  (
    n85,
    n10
  );


  not
  g20
  (
    n51,
    n15
  );


  buf
  g21
  (
    n61,
    n13
  );


  not
  g22
  (
    n94,
    n9
  );


  not
  g23
  (
    n44,
    n19
  );


  buf
  g24
  (
    n90,
    n10
  );


  buf
  g25
  (
    n67,
    n15
  );


  buf
  g26
  (
    n35,
    n13
  );


  buf
  g27
  (
    n28,
    n17
  );


  not
  g28
  (
    n45,
    n5
  );


  not
  g29
  (
    n38,
    n9
  );


  not
  g30
  (
    n43,
    n16
  );


  not
  g31
  (
    n33,
    n7
  );


  buf
  g32
  (
    n55,
    n4
  );


  buf
  g33
  (
    n47,
    n18
  );


  buf
  g34
  (
    n32,
    n4
  );


  not
  g35
  (
    n66,
    n17
  );


  buf
  g36
  (
    n22,
    n11
  );


  buf
  g37
  (
    n54,
    n18
  );


  not
  g38
  (
    n72,
    n17
  );


  not
  g39
  (
    n50,
    n7
  );


  buf
  g40
  (
    n59,
    n1
  );


  buf
  g41
  (
    n24,
    n3
  );


  not
  g42
  (
    n42,
    n1
  );


  not
  g43
  (
    n91,
    n6
  );


  not
  g44
  (
    n36,
    n3
  );


  buf
  g45
  (
    n69,
    n12
  );


  not
  g46
  (
    n68,
    n14
  );


  not
  g47
  (
    n20,
    n10
  );


  not
  g48
  (
    n71,
    n14
  );


  not
  g49
  (
    n40,
    n8
  );


  not
  g50
  (
    n46,
    n3
  );


  not
  g51
  (
    n77,
    n16
  );


  buf
  g52
  (
    n75,
    n14
  );


  not
  g53
  (
    n53,
    n13
  );


  not
  g54
  (
    n81,
    n9
  );


  buf
  g55
  (
    n58,
    n16
  );


  not
  g56
  (
    n30,
    n18
  );


  not
  g57
  (
    n78,
    n1
  );


  not
  g58
  (
    n27,
    n11
  );


  buf
  g59
  (
    n56,
    n9
  );


  buf
  g60
  (
    n48,
    n17
  );


  buf
  g61
  (
    n60,
    n8
  );


  not
  g62
  (
    n76,
    n6
  );


  buf
  g63
  (
    n41,
    n12
  );


  not
  g64
  (
    KeyWire_0_26,
    n5
  );


  not
  g65
  (
    n65,
    n2
  );


  buf
  g66
  (
    n84,
    n2
  );


  buf
  g67
  (
    n52,
    n11
  );


  not
  g68
  (
    n86,
    n5
  );


  buf
  g69
  (
    n92,
    n8
  );


  not
  g70
  (
    n31,
    n2
  );


  buf
  g71
  (
    n83,
    n4
  );


  not
  g72
  (
    n64,
    n12
  );


  buf
  g73
  (
    n21,
    n5
  );


  not
  g74
  (
    n93,
    n15
  );


  not
  g75
  (
    n73,
    n19
  );


  buf
  g76
  (
    n161,
    n39
  );


  buf
  g77
  (
    KeyWire_0_24,
    n65
  );


  not
  g78
  (
    n267,
    n36
  );


  buf
  g79
  (
    n151,
    n26
  );


  not
  g80
  (
    n154,
    n36
  );


  buf
  g81
  (
    n218,
    n50
  );


  not
  g82
  (
    n129,
    n69
  );


  buf
  g83
  (
    n201,
    n39
  );


  not
  g84
  (
    n254,
    n29
  );


  not
  g85
  (
    n176,
    n63
  );


  buf
  g86
  (
    n114,
    n35
  );


  not
  g87
  (
    n204,
    n73
  );


  not
  g88
  (
    n236,
    n27
  );


  buf
  g89
  (
    n233,
    n36
  );


  buf
  g90
  (
    n131,
    n43
  );


  buf
  g91
  (
    n99,
    n71
  );


  not
  g92
  (
    n196,
    n53
  );


  buf
  g93
  (
    n211,
    n43
  );


  not
  g94
  (
    n110,
    n71
  );


  not
  g95
  (
    n147,
    n49
  );


  not
  g96
  (
    n266,
    n53
  );


  buf
  g97
  (
    n251,
    n46
  );


  buf
  g98
  (
    n222,
    n57
  );


  buf
  g99
  (
    n288,
    n41
  );


  not
  g100
  (
    n127,
    n73
  );


  not
  g101
  (
    n173,
    n46
  );


  not
  g102
  (
    n213,
    n66
  );


  not
  g103
  (
    n136,
    n53
  );


  buf
  g104
  (
    n121,
    n42
  );


  buf
  g105
  (
    n191,
    n32
  );


  not
  g106
  (
    n225,
    n55
  );


  buf
  g107
  (
    n111,
    n38
  );


  not
  g108
  (
    n192,
    n29
  );


  not
  g109
  (
    n115,
    n67
  );


  not
  g110
  (
    n123,
    n44
  );


  buf
  g111
  (
    n199,
    n27
  );


  not
  g112
  (
    n168,
    n61
  );


  not
  g113
  (
    n250,
    n56
  );


  buf
  g114
  (
    n295,
    n39
  );


  buf
  g115
  (
    n263,
    n52
  );


  buf
  g116
  (
    n108,
    n49
  );


  buf
  g117
  (
    n120,
    n30
  );


  buf
  g118
  (
    n239,
    n56
  );


  buf
  g119
  (
    n246,
    n52
  );


  buf
  g120
  (
    n112,
    n33
  );


  not
  g121
  (
    n142,
    n63
  );


  not
  g122
  (
    n242,
    n52
  );


  buf
  g123
  (
    n207,
    n31
  );


  not
  g124
  (
    n149,
    n71
  );


  not
  g125
  (
    n195,
    n23
  );


  buf
  g126
  (
    n96,
    n26
  );


  not
  g127
  (
    n128,
    n73
  );


  not
  g128
  (
    n103,
    n58
  );


  not
  g129
  (
    n274,
    n69
  );


  buf
  g130
  (
    n157,
    n65
  );


  not
  g131
  (
    n180,
    n30
  );


  not
  g132
  (
    n182,
    n27
  );


  not
  g133
  (
    n107,
    n35
  );


  not
  g134
  (
    n156,
    n67
  );


  buf
  g135
  (
    n163,
    n37
  );


  not
  g136
  (
    n208,
    n68
  );


  buf
  g137
  (
    n158,
    n29
  );


  buf
  g138
  (
    n134,
    n28
  );


  buf
  g139
  (
    n243,
    n41
  );


  not
  g140
  (
    n257,
    n48
  );


  not
  g141
  (
    n184,
    n23
  );


  not
  g142
  (
    n241,
    n33
  );


  buf
  g143
  (
    n290,
    n58
  );


  buf
  g144
  (
    n109,
    n54
  );


  buf
  g145
  (
    n200,
    n54
  );


  buf
  g146
  (
    n279,
    n51
  );


  buf
  g147
  (
    n193,
    n51
  );


  buf
  g148
  (
    n183,
    n69
  );


  buf
  g149
  (
    n268,
    n64
  );


  buf
  g150
  (
    KeyWire_0_4,
    n41
  );


  not
  g151
  (
    n140,
    n53
  );


  not
  g152
  (
    n169,
    n47
  );


  buf
  g153
  (
    n231,
    n37
  );


  buf
  g154
  (
    n247,
    n37
  );


  buf
  g155
  (
    n138,
    n46
  );


  buf
  g156
  (
    n178,
    n47
  );


  not
  g157
  (
    n287,
    n27
  );


  buf
  g158
  (
    n116,
    n50
  );


  not
  g159
  (
    n126,
    n60
  );


  buf
  g160
  (
    n118,
    n40
  );


  not
  g161
  (
    n276,
    n60
  );


  not
  g162
  (
    n152,
    n55
  );


  not
  g163
  (
    n113,
    n44
  );


  not
  g164
  (
    n235,
    n57
  );


  buf
  g165
  (
    n162,
    n33
  );


  not
  g166
  (
    n133,
    n48
  );


  not
  g167
  (
    n296,
    n67
  );


  buf
  g168
  (
    n175,
    n60
  );


  not
  g169
  (
    n124,
    n37
  );


  not
  g170
  (
    n212,
    n47
  );


  not
  g171
  (
    n214,
    n65
  );


  buf
  g172
  (
    n281,
    n66
  );


  buf
  g173
  (
    n260,
    n68
  );


  buf
  g174
  (
    n240,
    n72
  );


  not
  g175
  (
    n277,
    n30
  );


  buf
  g176
  (
    n269,
    n42
  );


  buf
  g177
  (
    n203,
    n41
  );


  buf
  g178
  (
    n285,
    n25
  );


  not
  g179
  (
    n186,
    n55
  );


  buf
  g180
  (
    n237,
    n48
  );


  not
  g181
  (
    n283,
    n73
  );


  buf
  g182
  (
    n153,
    n64
  );


  buf
  g183
  (
    n232,
    n67
  );


  not
  g184
  (
    n286,
    n46
  );


  buf
  g185
  (
    n137,
    n68
  );


  not
  g186
  (
    KeyWire_0_18,
    n45
  );


  buf
  g187
  (
    n171,
    n40
  );


  buf
  g188
  (
    n261,
    n62
  );


  buf
  g189
  (
    n229,
    n62
  );


  buf
  g190
  (
    n262,
    n59
  );


  buf
  g191
  (
    n284,
    n59
  );


  not
  g192
  (
    n282,
    n64
  );


  not
  g193
  (
    n275,
    n71
  );


  buf
  g194
  (
    n234,
    n32
  );


  not
  g195
  (
    n185,
    n44
  );


  buf
  g196
  (
    n172,
    n25
  );


  not
  g197
  (
    n294,
    n28
  );


  buf
  g198
  (
    n139,
    n52
  );


  buf
  g199
  (
    n228,
    n66
  );


  not
  g200
  (
    n141,
    n48
  );


  not
  g201
  (
    n219,
    n65
  );


  buf
  g202
  (
    n259,
    n45
  );


  buf
  g203
  (
    n217,
    n34
  );


  not
  g204
  (
    n272,
    n58
  );


  not
  g205
  (
    n170,
    n72
  );


  buf
  g206
  (
    n244,
    n63
  );


  not
  g207
  (
    n144,
    n20
  );


  buf
  g208
  (
    n252,
    n57
  );


  buf
  g209
  (
    n98,
    n69
  );


  buf
  g210
  (
    n164,
    n24
  );


  buf
  g211
  (
    n177,
    n51
  );


  buf
  g212
  (
    n206,
    n38
  );


  not
  g213
  (
    n155,
    n61
  );


  buf
  g214
  (
    n205,
    n68
  );


  not
  g215
  (
    n255,
    n47
  );


  not
  g216
  (
    n224,
    n50
  );


  buf
  g217
  (
    n181,
    n54
  );


  buf
  g218
  (
    n264,
    n44
  );


  buf
  g219
  (
    n245,
    n45
  );


  buf
  g220
  (
    n291,
    n31
  );


  not
  g221
  (
    n293,
    n72
  );


  not
  g222
  (
    n197,
    n58
  );


  not
  g223
  (
    n278,
    n32
  );


  not
  g224
  (
    n146,
    n43
  );


  buf
  g225
  (
    n117,
    n31
  );


  buf
  g226
  (
    n189,
    n49
  );


  buf
  g227
  (
    n179,
    n49
  );


  buf
  g228
  (
    n227,
    n21
  );


  buf
  g229
  (
    n194,
    n64
  );


  buf
  g230
  (
    n249,
    n40
  );


  buf
  g231
  (
    n150,
    n62
  );


  not
  g232
  (
    n166,
    n61
  );


  not
  g233
  (
    n265,
    n56
  );


  not
  g234
  (
    n148,
    n60
  );


  not
  g235
  (
    n105,
    n51
  );


  not
  g236
  (
    n216,
    n42
  );


  buf
  g237
  (
    n238,
    n24
  );


  not
  g238
  (
    n188,
    n34
  );


  buf
  g239
  (
    n165,
    n70
  );


  not
  g240
  (
    n273,
    n32
  );


  buf
  g241
  (
    n220,
    n70
  );


  buf
  g242
  (
    n190,
    n21
  );


  not
  g243
  (
    n292,
    n22
  );


  buf
  g244
  (
    n256,
    n22
  );


  buf
  g245
  (
    n270,
    n59
  );


  buf
  g246
  (
    n160,
    n34
  );


  buf
  g247
  (
    n106,
    n40
  );


  not
  g248
  (
    n122,
    n56
  );


  not
  g249
  (
    n215,
    n35
  );


  buf
  g250
  (
    n253,
    n62
  );


  not
  g251
  (
    n143,
    n31
  );


  buf
  g252
  (
    n125,
    n63
  );


  buf
  g253
  (
    n132,
    n38
  );


  buf
  g254
  (
    n101,
    n28
  );


  buf
  g255
  (
    n135,
    n29
  );


  not
  g256
  (
    n187,
    n61
  );


  not
  g257
  (
    n289,
    n66
  );


  buf
  g258
  (
    n159,
    n70
  );


  not
  g259
  (
    KeyWire_0_12,
    n59
  );


  not
  g260
  (
    n248,
    n43
  );


  buf
  g261
  (
    n258,
    n30
  );


  buf
  g262
  (
    n230,
    n34
  );


  not
  g263
  (
    n104,
    n35
  );


  not
  g264
  (
    n271,
    n28
  );


  not
  g265
  (
    n97,
    n39
  );


  not
  g266
  (
    n145,
    n36
  );


  not
  g267
  (
    n209,
    n57
  );


  not
  g268
  (
    n100,
    n50
  );


  not
  g269
  (
    n223,
    n54
  );


  not
  g270
  (
    n167,
    n42
  );


  buf
  g271
  (
    n210,
    n33
  );


  not
  g272
  (
    n202,
    n55
  );


  not
  g273
  (
    n198,
    n45
  );


  not
  g274
  (
    n226,
    n38
  );


  buf
  g275
  (
    n174,
    n72
  );


  not
  g276
  (
    n102,
    n70
  );


  not
  g277
  (
    n361,
    n231
  );


  buf
  g278
  (
    n511,
    n212
  );


  not
  g279
  (
    n478,
    n138
  );


  not
  g280
  (
    n335,
    n177
  );


  not
  g281
  (
    n494,
    n182
  );


  not
  g282
  (
    n540,
    n81
  );


  not
  g283
  (
    n325,
    n75
  );


  buf
  g284
  (
    n433,
    n83
  );


  not
  g285
  (
    n422,
    n260
  );


  buf
  g286
  (
    n405,
    n229
  );


  not
  g287
  (
    n340,
    n195
  );


  not
  g288
  (
    n376,
    n188
  );


  not
  g289
  (
    n455,
    n240
  );


  buf
  g290
  (
    n524,
    n263
  );


  not
  g291
  (
    n472,
    n262
  );


  buf
  g292
  (
    n582,
    n236
  );


  not
  g293
  (
    n305,
    n112
  );


  buf
  g294
  (
    n467,
    n223
  );


  buf
  g295
  (
    n375,
    n190
  );


  buf
  g296
  (
    n423,
    n187
  );


  buf
  g297
  (
    n513,
    n143
  );


  buf
  g298
  (
    n509,
    n88
  );


  buf
  g299
  (
    n410,
    n279
  );


  not
  g300
  (
    n548,
    n212
  );


  buf
  g301
  (
    n407,
    n91
  );


  not
  g302
  (
    n574,
    n224
  );


  not
  g303
  (
    n382,
    n75
  );


  buf
  g304
  (
    n420,
    n167
  );


  buf
  g305
  (
    n475,
    n170
  );


  buf
  g306
  (
    n299,
    n206
  );


  not
  g307
  (
    n387,
    n255
  );


  not
  g308
  (
    n326,
    n156
  );


  not
  g309
  (
    n590,
    n273
  );


  not
  g310
  (
    n490,
    n261
  );


  buf
  g311
  (
    n435,
    n104
  );


  not
  g312
  (
    n452,
    n152
  );


  not
  g313
  (
    n303,
    n127
  );


  buf
  g314
  (
    n512,
    n253
  );


  not
  g315
  (
    n364,
    n91
  );


  not
  g316
  (
    n487,
    n255
  );


  buf
  g317
  (
    n576,
    n101
  );


  buf
  g318
  (
    n496,
    n112
  );


  buf
  g319
  (
    n370,
    n165
  );


  not
  g320
  (
    n585,
    n141
  );


  buf
  g321
  (
    n533,
    n93
  );


  not
  g322
  (
    n308,
    n258
  );


  buf
  g323
  (
    n543,
    n265
  );


  buf
  g324
  (
    n411,
    n202
  );


  buf
  g325
  (
    n324,
    n263
  );


  not
  g326
  (
    n421,
    n85
  );


  not
  g327
  (
    n371,
    n79
  );


  buf
  g328
  (
    n347,
    n133
  );


  buf
  g329
  (
    n507,
    n184
  );


  not
  g330
  (
    n379,
    n203
  );


  not
  g331
  (
    n330,
    n276
  );


  not
  g332
  (
    n355,
    n254
  );


  not
  g333
  (
    n301,
    n246
  );


  buf
  g334
  (
    n541,
    n82
  );


  buf
  g335
  (
    n357,
    n243
  );


  buf
  g336
  (
    n395,
    n262
  );


  buf
  g337
  (
    n484,
    n148
  );


  not
  g338
  (
    n537,
    n80
  );


  not
  g339
  (
    n454,
    n200
  );


  buf
  g340
  (
    n529,
    n217
  );


  not
  g341
  (
    n327,
    n276
  );


  buf
  g342
  (
    n317,
    n187
  );


  not
  g343
  (
    n456,
    n266
  );


  buf
  g344
  (
    n432,
    n229
  );


  not
  g345
  (
    n604,
    n74
  );


  buf
  g346
  (
    n545,
    n140
  );


  not
  g347
  (
    n337,
    n151
  );


  not
  g348
  (
    n489,
    n117
  );


  not
  g349
  (
    n481,
    n77
  );


  not
  g350
  (
    n469,
    n124
  );


  buf
  g351
  (
    n413,
    n204
  );


  not
  g352
  (
    n431,
    n227
  );


  buf
  g353
  (
    n560,
    n205
  );


  buf
  g354
  (
    n448,
    n228
  );


  not
  g355
  (
    n390,
    n269
  );


  buf
  g356
  (
    n373,
    n253
  );


  buf
  g357
  (
    n600,
    n251
  );


  buf
  g358
  (
    n602,
    n114
  );


  buf
  g359
  (
    n446,
    n209
  );


  buf
  g360
  (
    n306,
    n160
  );


  buf
  g361
  (
    n599,
    n84
  );


  buf
  g362
  (
    n316,
    n193
  );


  buf
  g363
  (
    n417,
    n81
  );


  not
  g364
  (
    n346,
    n192
  );


  not
  g365
  (
    n447,
    n189
  );


  not
  g366
  (
    n596,
    n201
  );


  not
  g367
  (
    n384,
    n275
  );


  buf
  g368
  (
    KeyWire_0_13,
    n145
  );


  buf
  g369
  (
    KeyWire_0_9,
    n224
  );


  buf
  g370
  (
    n312,
    n267
  );


  buf
  g371
  (
    n441,
    n218
  );


  buf
  g372
  (
    n535,
    n204
  );


  buf
  g373
  (
    n424,
    n162
  );


  not
  g374
  (
    n597,
    n223
  );


  not
  g375
  (
    n608,
    n138
  );


  buf
  g376
  (
    n404,
    n266
  );


  buf
  g377
  (
    n366,
    n85
  );


  not
  g378
  (
    n434,
    n236
  );


  buf
  g379
  (
    n505,
    n216
  );


  not
  g380
  (
    n436,
    n213
  );


  not
  g381
  (
    n307,
    n221
  );


  buf
  g382
  (
    n315,
    n275
  );


  not
  g383
  (
    n297,
    n105
  );


  not
  g384
  (
    n348,
    n230
  );


  not
  g385
  (
    n464,
    n269
  );


  buf
  g386
  (
    n501,
    n226
  );


  buf
  g387
  (
    n443,
    n82
  );


  buf
  g388
  (
    n563,
    n240
  );


  not
  g389
  (
    n402,
    n227
  );


  not
  g390
  (
    n453,
    n189
  );


  not
  g391
  (
    n523,
    n242
  );


  not
  g392
  (
    KeyWire_0_7,
    n111
  );


  buf
  g393
  (
    n587,
    n221
  );


  not
  g394
  (
    n372,
    n258
  );


  buf
  g395
  (
    n525,
    n274
  );


  not
  g396
  (
    n569,
    n78
  );


  not
  g397
  (
    n396,
    n90
  );


  buf
  g398
  (
    n442,
    n273
  );


  buf
  g399
  (
    n439,
    n83
  );


  not
  g400
  (
    n437,
    n75
  );


  buf
  g401
  (
    n398,
    n204
  );


  not
  g402
  (
    n592,
    n212
  );


  not
  g403
  (
    n408,
    n252
  );


  buf
  g404
  (
    n532,
    n109
  );


  buf
  g405
  (
    n504,
    n131
  );


  buf
  g406
  (
    n440,
    n78
  );


  not
  g407
  (
    n580,
    n269
  );


  buf
  g408
  (
    n471,
    n260
  );


  buf
  g409
  (
    n333,
    n87
  );


  buf
  g410
  (
    n581,
    n245
  );


  not
  g411
  (
    n589,
    n209
  );


  not
  g412
  (
    n332,
    n117
  );


  buf
  g413
  (
    n329,
    n115
  );


  buf
  g414
  (
    n611,
    n105
  );


  buf
  g415
  (
    n538,
    n164
  );


  not
  g416
  (
    KeyWire_0_0,
    n231
  );


  buf
  g417
  (
    n528,
    n246
  );


  not
  g418
  (
    n601,
    n258
  );


  not
  g419
  (
    n531,
    n177
  );


  buf
  g420
  (
    n321,
    n172
  );


  buf
  g421
  (
    n350,
    n136
  );


  not
  g422
  (
    n362,
    n199
  );


  buf
  g423
  (
    n320,
    n132
  );


  not
  g424
  (
    n359,
    n153
  );


  not
  g425
  (
    n502,
    n140
  );


  buf
  g426
  (
    n377,
    n244
  );


  not
  g427
  (
    n520,
    n241
  );


  not
  g428
  (
    n342,
    n212
  );


  not
  g429
  (
    n383,
    n211
  );


  buf
  g430
  (
    n577,
    n268
  );


  buf
  g431
  (
    n415,
    n88
  );


  buf
  g432
  (
    n522,
    n205
  );


  buf
  g433
  (
    n555,
    n198
  );


  not
  g434
  (
    n483,
    n215
  );


  not
  g435
  (
    n336,
    n270
  );


  buf
  g436
  (
    n338,
    n86
  );


  not
  g437
  (
    n527,
    n116
  );


  not
  g438
  (
    KeyWire_0_19,
    n209
  );


  buf
  g439
  (
    n334,
    n77
  );


  buf
  g440
  (
    n603,
    n153
  );


  not
  g441
  (
    n341,
    n191
  );


  buf
  g442
  (
    n412,
    n215
  );


  buf
  g443
  (
    KeyWire_0_31,
    n235
  );


  buf
  g444
  (
    n488,
    n220
  );


  not
  g445
  (
    n530,
    n179
  );


  buf
  g446
  (
    n465,
    n123
  );


  not
  g447
  (
    n418,
    n206
  );


  buf
  g448
  (
    n473,
    n256
  );


  not
  g449
  (
    n610,
    n224
  );


  buf
  g450
  (
    n319,
    n147
  );


  not
  g451
  (
    KeyWire_0_23,
    n244
  );


  not
  g452
  (
    n500,
    n249
  );


  not
  g453
  (
    n598,
    n86
  );


  not
  g454
  (
    n539,
    n206
  );


  buf
  g455
  (
    n344,
    n195
  );


  buf
  g456
  (
    n356,
    n108
  );


  not
  g457
  (
    n367,
    n265
  );


  buf
  g458
  (
    n427,
    n237
  );


  not
  g459
  (
    n298,
    n166
  );


  not
  g460
  (
    n451,
    n256
  );


  not
  g461
  (
    n426,
    n275
  );


  buf
  g462
  (
    n514,
    n259
  );


  not
  g463
  (
    n479,
    n85
  );


  not
  g464
  (
    n595,
    n130
  );


  not
  g465
  (
    n491,
    n139
  );


  not
  g466
  (
    n572,
    n169
  );


  not
  g467
  (
    n605,
    n221
  );


  buf
  g468
  (
    n503,
    n163
  );


  buf
  g469
  (
    n445,
    n220
  );


  buf
  g470
  (
    n510,
    n93
  );


  not
  g471
  (
    n526,
    n133
  );


  not
  g472
  (
    n459,
    n149
  );


  buf
  g473
  (
    n518,
    n264
  );


  not
  g474
  (
    n463,
    n277
  );


  buf
  g475
  (
    KeyWire_0_20,
    n277
  );


  not
  g476
  (
    n461,
    n226
  );


  not
  g477
  (
    n575,
    n251
  );


  buf
  g478
  (
    n409,
    n136
  );


  buf
  g479
  (
    n568,
    n264
  );


  buf
  g480
  (
    n571,
    n239
  );


  not
  g481
  (
    n609,
    n231
  );


  buf
  g482
  (
    n552,
    n275
  );


  not
  g483
  (
    n358,
    n222
  );


  not
  g484
  (
    n517,
    n79
  );


  nor
  g485
  (
    n567,
    n84,
    n134,
    n250,
    n223
  );


  and
  g486
  (
    n542,
    n86,
    n164,
    n148,
    n183
  );


  and
  g487
  (
    n558,
    n247,
    n90,
    n232,
    n122
  );


  and
  g488
  (
    n345,
    n239,
    n80,
    n181,
    n193
  );


  and
  g489
  (
    n393,
    n128,
    n202,
    n248,
    n246
  );


  nor
  g490
  (
    n515,
    n255,
    n259,
    n192,
    n203
  );


  and
  g491
  (
    n388,
    n257,
    n107,
    n269,
    n173
  );


  nor
  g492
  (
    n492,
    n74,
    n197,
    n87,
    n178
  );


  nand
  g493
  (
    n425,
    n216,
    n194,
    n219,
    n218
  );


  nor
  g494
  (
    n544,
    n205,
    n232,
    n235,
    n265
  );


  xor
  g495
  (
    n462,
    n89,
    n274,
    n279,
    n187
  );


  and
  g496
  (
    n328,
    n185,
    n225,
    n219,
    n227
  );


  nand
  g497
  (
    n343,
    n276,
    n178,
    n271,
    n198
  );


  xnor
  g498
  (
    n360,
    n220,
    n214,
    n215,
    n155
  );


  xnor
  g499
  (
    n365,
    n200,
    n225,
    n75,
    n238
  );


  xor
  g500
  (
    n363,
    n268,
    n222,
    n99,
    n168
  );


  xor
  g501
  (
    KeyWire_0_22,
    n144,
    n217,
    n225,
    n243
  );


  nor
  g502
  (
    n476,
    n227,
    n247,
    n226,
    n81
  );


  xor
  g503
  (
    n564,
    n176,
    n274,
    n152,
    n100
  );


  and
  g504
  (
    n458,
    n214,
    n77,
    n271,
    n121
  );


  xor
  g505
  (
    n579,
    n278,
    n199,
    n229
  );


  and
  g506
  (
    n416,
    n256,
    n234,
    n161,
    n150
  );


  xor
  g507
  (
    KeyWire_0_28,
    n194,
    n141,
    n244,
    n193
  );


  nor
  g508
  (
    n583,
    n270,
    n266,
    n200,
    n163
  );


  xnor
  g509
  (
    n349,
    n254,
    n280,
    n113,
    n237
  );


  nand
  g510
  (
    n428,
    n250,
    n259,
    n268,
    n165
  );


  xnor
  g511
  (
    n309,
    n137,
    n93,
    n193,
    n249
  );


  xor
  g512
  (
    n606,
    n208,
    n232,
    n268,
    n180
  );


  and
  g513
  (
    n406,
    n252,
    n234,
    n98,
    n84
  );


  xor
  g514
  (
    n438,
    n191,
    n276,
    n187,
    n109
  );


  xnor
  g515
  (
    n485,
    n86,
    n88,
    n127,
    n211
  );


  nand
  g516
  (
    n313,
    n126,
    n248,
    n233,
    n207
  );


  nand
  g517
  (
    n553,
    n201,
    n78,
    n216,
    n245
  );


  nand
  g518
  (
    KeyWire_0_6,
    n201,
    n169,
    n188,
    n248
  );


  xnor
  g519
  (
    n497,
    n150,
    n90,
    n207,
    n215
  );


  nor
  g520
  (
    n351,
    n198,
    n256,
    n210
  );


  xor
  g521
  (
    n536,
    n239,
    n199,
    n196,
    n106
  );


  and
  g522
  (
    n323,
    n262,
    n245,
    n257,
    n144
  );


  or
  g523
  (
    n551,
    n97,
    n261,
    n175,
    n93
  );


  and
  g524
  (
    n399,
    n242,
    n214,
    n240,
    n196
  );


  nand
  g525
  (
    n310,
    n273,
    n211,
    n79,
    n198
  );


  xor
  g526
  (
    n403,
    n151,
    n263,
    n166,
    n106
  );


  nand
  g527
  (
    n554,
    n158,
    n242,
    n206,
    n222
  );


  and
  g528
  (
    n466,
    n274,
    n244,
    n161,
    n210
  );


  xor
  g529
  (
    n450,
    n88,
    n192,
    n80,
    n191
  );


  xnor
  g530
  (
    n419,
    n192,
    n254,
    n203,
    n189
  );


  nand
  g531
  (
    n392,
    n139,
    n252,
    n213,
    n271
  );


  xor
  g532
  (
    n397,
    n247,
    n76,
    n214,
    n101
  );


  xor
  g533
  (
    n588,
    n243,
    n156,
    n135,
    n186
  );


  xor
  g534
  (
    n322,
    n181,
    n87,
    n107,
    n154
  );


  xor
  g535
  (
    n547,
    n203,
    n119,
    n270,
    n84
  );


  xor
  g536
  (
    KeyWire_0_29,
    n226,
    n235,
    n257
  );


  and
  g537
  (
    n546,
    n185,
    n111,
    n80,
    n222
  );


  nand
  g538
  (
    n352,
    n110,
    n128,
    n265,
    n79
  );


  or
  g539
  (
    n369,
    n237,
    n242,
    n145,
    n238
  );


  xnor
  g540
  (
    n314,
    n182,
    n255,
    n186,
    n123
  );


  or
  g541
  (
    n486,
    n134,
    n132,
    n247,
    n92
  );


  nor
  g542
  (
    n444,
    n175,
    n102,
    n197,
    n146
  );


  and
  g543
  (
    n381,
    n82,
    n218,
    n76,
    n202
  );


  and
  g544
  (
    n353,
    n129,
    n125,
    n120,
    n238
  );


  xor
  g545
  (
    n430,
    n202,
    n216,
    n232,
    n149
  );


  or
  g546
  (
    n557,
    n208,
    n191,
    n159,
    n211
  );


  or
  g547
  (
    n562,
    n267,
    n267,
    n179,
    n218
  );


  xor
  g548
  (
    n449,
    n172,
    n262,
    n188,
    n104
  );


  xnor
  g549
  (
    n516,
    n121,
    n130,
    n190,
    n233
  );


  xor
  g550
  (
    n460,
    n273,
    n233,
    n230,
    n83
  );


  or
  g551
  (
    n561,
    n180,
    n157,
    n98,
    n260
  );


  or
  g552
  (
    n391,
    n260,
    n219,
    n110,
    n251
  );


  xnor
  g553
  (
    n591,
    n190,
    n170,
    n85,
    n272
  );


  xnor
  g554
  (
    n506,
    n108,
    n115,
    n280,
    n174
  );


  xor
  g555
  (
    n570,
    n238,
    n116,
    n125,
    n131
  );


  nor
  g556
  (
    n386,
    n261,
    n249,
    n272,
    n99
  );


  nand
  g557
  (
    n556,
    n82,
    n261,
    n246,
    n213
  );


  xnor
  g558
  (
    n474,
    n173,
    n230,
    n228,
    n97
  );


  xor
  g559
  (
    n401,
    n195,
    n168,
    n277,
    n91
  );


  or
  g560
  (
    n498,
    n230,
    n76,
    n279,
    n201
  );


  xor
  g561
  (
    n300,
    n167,
    n213,
    n81,
    n102
  );


  nor
  g562
  (
    n477,
    n92,
    n89,
    n229,
    n278
  );


  or
  g563
  (
    n468,
    n114,
    n135,
    n184,
    n272
  );


  nor
  g564
  (
    n549,
    n236,
    n188,
    n267,
    n77
  );


  and
  g565
  (
    n339,
    n118,
    n234,
    n159,
    n252
  );


  xor
  g566
  (
    n374,
    n245,
    n217,
    n209,
    n143
  );


  xor
  g567
  (
    KeyWire_0_30,
    n155,
    n189,
    n118,
    n237
  );


  nand
  g568
  (
    n578,
    n196,
    n147,
    n280,
    n266
  );


  xnor
  g569
  (
    n519,
    n194,
    n278,
    n91,
    n190
  );


  nor
  g570
  (
    n331,
    n90,
    n103,
    n83,
    n250
  );


  and
  g571
  (
    n573,
    n142,
    n142,
    n76,
    n250
  );


  xor
  g572
  (
    n304,
    n239,
    n241,
    n254,
    n89
  );


  or
  g573
  (
    n470,
    n176,
    n122,
    n87,
    n270
  );


  xnor
  g574
  (
    n368,
    n183,
    n234,
    n220,
    n92
  );


  nor
  g575
  (
    n400,
    n204,
    n74,
    n257,
    n263
  );


  xnor
  g576
  (
    n354,
    n233,
    n264,
    n208,
    n207
  );


  nor
  g577
  (
    n414,
    n74,
    n171,
    n224,
    n196
  );


  and
  g578
  (
    n593,
    n219,
    n113,
    n119,
    n280
  );


  or
  g579
  (
    n534,
    n207,
    n146,
    n228,
    n120
  );


  nor
  g580
  (
    n565,
    n137,
    n258,
    n249,
    n100
  );


  and
  g581
  (
    n495,
    n228,
    n200,
    n174,
    n154
  );


  or
  g582
  (
    n493,
    n194,
    n162,
    n89,
    n271
  );


  and
  g583
  (
    n378,
    n92,
    n129,
    n243,
    n205
  );


  nor
  g584
  (
    n302,
    n241,
    n231,
    n157,
    n197
  );


  xor
  g585
  (
    n311,
    n278,
    n171,
    n277,
    n253
  );


  xnor
  g586
  (
    KeyWire_0_17,
    n259,
    n210,
    n248,
    n225
  );


  and
  g587
  (
    n594,
    n236,
    n158,
    n124,
    n160
  );


  xor
  g588
  (
    n480,
    n217,
    n251,
    n195,
    n264
  );


  nand
  g589
  (
    n389,
    n253,
    n221,
    n223,
    n103
  );


  or
  g590
  (
    n521,
    n272,
    n78,
    n208,
    n240
  );


  nor
  g591
  (
    n586,
    n126,
    n279,
    n197,
    n241
  );


  not
  g592
  (
    n619,
    n309
  );


  not
  g593
  (
    n626,
    n301
  );


  buf
  g594
  (
    n623,
    n304
  );


  buf
  g595
  (
    n628,
    n323
  );


  buf
  g596
  (
    n621,
    n310
  );


  buf
  g597
  (
    n624,
    n319
  );


  buf
  g598
  (
    n616,
    n316
  );


  buf
  g599
  (
    n627,
    n298
  );


  buf
  g600
  (
    n614,
    n321
  );


  not
  g601
  (
    n625,
    n303
  );


  buf
  g602
  (
    KeyWire_0_2,
    n299
  );


  buf
  g603
  (
    n633,
    n313
  );


  not
  g604
  (
    n630,
    n314
  );


  buf
  g605
  (
    n632,
    n308
  );


  not
  g606
  (
    n618,
    n307
  );


  buf
  g607
  (
    n615,
    n312
  );


  buf
  g608
  (
    n617,
    n318
  );


  not
  g609
  (
    n620,
    n311
  );


  buf
  g610
  (
    n629,
    n300
  );


  not
  g611
  (
    n612,
    n315
  );


  nor
  g612
  (
    n631,
    n306,
    n325,
    n305,
    n324
  );


  nand
  g613
  (
    n622,
    n320,
    n317,
    n302,
    n322
  );


  xnor
  g614
  (
    n635,
    n625,
    n356,
    n331,
    n339
  );


  xor
  g615
  (
    n647,
    n335,
    n336,
    n355,
    n328
  );


  or
  g616
  (
    n636,
    n345,
    n326,
    n358,
    n334
  );


  nor
  g617
  (
    n643,
    n338,
    n350,
    n341,
    n621
  );


  nor
  g618
  (
    n641,
    n618,
    n615,
    n340,
    n333
  );


  and
  g619
  (
    n646,
    n361,
    n366,
    n351,
    n332
  );


  or
  g620
  (
    n638,
    n364,
    n349,
    n617,
    n363
  );


  or
  g621
  (
    n644,
    n616,
    n352,
    n614,
    n330
  );


  or
  g622
  (
    n642,
    n613,
    n622,
    n347,
    n362
  );


  nand
  g623
  (
    n637,
    n342,
    n348,
    n619,
    n343
  );


  or
  g624
  (
    n634,
    n329,
    n357,
    n354,
    n359
  );


  nand
  g625
  (
    n640,
    n367,
    n353,
    n337,
    n365
  );


  nand
  g626
  (
    n645,
    n612,
    n346,
    n620,
    n344
  );


  nor
  g627
  (
    n639,
    n624,
    n327,
    n360,
    n623
  );


  and
  g628
  (
    n654,
    n284,
    n283,
    n377,
    n642
  );


  nor
  g629
  (
    n651,
    n379,
    n370,
    n643,
    n281
  );


  nand
  g630
  (
    n657,
    n281,
    n641,
    n283,
    n376
  );


  or
  g631
  (
    n649,
    n371,
    n284,
    n283,
    n378
  );


  xnor
  g632
  (
    n653,
    n646,
    n647,
    n282,
    n283
  );


  xor
  g633
  (
    n656,
    n284,
    n281,
    n645,
    n373
  );


  xor
  g634
  (
    n655,
    n285,
    n369,
    n640,
    n282
  );


  and
  g635
  (
    n650,
    n282,
    n285,
    n281,
    n644
  );


  xnor
  g636
  (
    n648,
    n284,
    n638,
    n372,
    n282
  );


  xnor
  g637
  (
    KeyWire_0_11,
    n368,
    n639,
    n374,
    n375
  );


  not
  g638
  (
    n661,
    n388
  );


  buf
  g639
  (
    n658,
    n387
  );


  nand
  g640
  (
    n659,
    n649,
    n384
  );


  xnor
  g641
  (
    n662,
    n392,
    n386,
    n648,
    n383
  );


  nor
  g642
  (
    n664,
    n654,
    n385,
    n381,
    n653
  );


  nand
  g643
  (
    n660,
    n380,
    n391,
    n652,
    n651
  );


  or
  g644
  (
    n663,
    n389,
    n390,
    n650,
    n382
  );


  and
  g645
  (
    n665,
    n406,
    n660,
    n659,
    n428
  );


  or
  g646
  (
    n669,
    n417,
    n410,
    n403,
    n421
  );


  nand
  g647
  (
    n679,
    n661,
    n409,
    n402,
    n659
  );


  nor
  g648
  (
    KeyWire_0_8,
    n423,
    n405,
    n401,
    n659
  );


  or
  g649
  (
    n677,
    n437,
    n658,
    n418,
    n411
  );


  xor
  g650
  (
    n672,
    n661,
    n424,
    n658,
    n434
  );


  or
  g651
  (
    n671,
    n431,
    n432,
    n661,
    n659
  );


  nor
  g652
  (
    n678,
    n397,
    n414,
    n420,
    n660
  );


  or
  g653
  (
    n673,
    n419,
    n399,
    n661,
    n436
  );


  xor
  g654
  (
    n667,
    n662,
    n430,
    n407,
    n433
  );


  nor
  g655
  (
    n668,
    n413,
    n426,
    n394,
    n415
  );


  or
  g656
  (
    n670,
    n412,
    n396,
    n398,
    n422
  );


  xnor
  g657
  (
    n676,
    n395,
    n660,
    n425,
    n393
  );


  nand
  g658
  (
    n674,
    n400,
    n660,
    n427,
    n435
  );


  xor
  g659
  (
    n675,
    n404,
    n416,
    n429,
    n408
  );


  xor
  g660
  (
    n689,
    n285,
    n664,
    n667
  );


  nand
  g661
  (
    n693,
    n679,
    n628,
    n655,
    n666
  );


  and
  g662
  (
    n682,
    n678,
    n675,
    n676,
    n632
  );


  xnor
  g663
  (
    n681,
    n94,
    n288,
    n679,
    n626
  );


  xor
  g664
  (
    n686,
    n286,
    n440,
    n663,
    n629
  );


  nand
  g665
  (
    n695,
    n673,
    n630,
    n672,
    n288
  );


  nand
  g666
  (
    n683,
    n657,
    n663,
    n627,
    n662
  );


  or
  g667
  (
    n680,
    n289,
    n286,
    n438
  );


  or
  g668
  (
    n684,
    n671,
    n287,
    n285,
    n442
  );


  or
  g669
  (
    n694,
    n288,
    n289,
    n439
  );


  nand
  g670
  (
    n690,
    n286,
    n633,
    n631,
    n670
  );


  xor
  g671
  (
    n688,
    n287,
    n663,
    n664,
    n443
  );


  nand
  g672
  (
    n685,
    n665,
    n674,
    n287,
    n662
  );


  and
  g673
  (
    n691,
    n668,
    n287,
    n664,
    n669
  );


  nand
  g674
  (
    n687,
    n677,
    n656,
    n663,
    n94
  );


  nand
  g675
  (
    n692,
    n441,
    n289,
    n288,
    n662
  );


  not
  g676
  (
    n698,
    n680
  );


  buf
  g677
  (
    n718,
    n682
  );


  not
  g678
  (
    n707,
    n682
  );


  not
  g679
  (
    n699,
    n684
  );


  not
  g680
  (
    n710,
    n685
  );


  buf
  g681
  (
    n717,
    n685
  );


  not
  g682
  (
    n716,
    n684
  );


  not
  g683
  (
    n709,
    n684
  );


  buf
  g684
  (
    n702,
    n686
  );


  not
  g685
  (
    n711,
    n680
  );


  not
  g686
  (
    n703,
    n682
  );


  buf
  g687
  (
    n715,
    n686
  );


  not
  g688
  (
    n700,
    n683
  );


  buf
  g689
  (
    n704,
    n683
  );


  buf
  g690
  (
    n712,
    n683
  );


  not
  g691
  (
    n719,
    n684
  );


  not
  g692
  (
    n706,
    n681
  );


  buf
  g693
  (
    n701,
    n681
  );


  buf
  g694
  (
    n705,
    n685
  );


  buf
  g695
  (
    n708,
    n686
  );


  buf
  g696
  (
    n713,
    n683
  );


  not
  g697
  (
    n714,
    n682
  );


  not
  g698
  (
    n697,
    n685
  );


  buf
  g699
  (
    n696,
    n686
  );


  buf
  g700
  (
    n725,
    n697
  );


  buf
  g701
  (
    n727,
    n699
  );


  not
  g702
  (
    KeyWire_0_25,
    n698
  );


  buf
  g703
  (
    n726,
    n696
  );


  not
  g704
  (
    KeyWire_0_3,
    n687
  );


  not
  g705
  (
    n724,
    n700
  );


  xor
  g706
  (
    n720,
    n699,
    n687
  );


  nand
  g707
  (
    n729,
    n449,
    n697,
    n687,
    n698
  );


  nand
  g708
  (
    n723,
    n447,
    n448,
    n696,
    n445
  );


  xor
  g709
  (
    n722,
    n444,
    n446,
    n700,
    n687
  );


  not
  g710
  (
    n730,
    n720
  );


  xnor
  g711
  (
    n732,
    n701,
    n451,
    n454
  );


  and
  g712
  (
    n733,
    n721,
    n456,
    n450,
    n722
  );


  xnor
  g713
  (
    n731,
    n721,
    n453,
    n452,
    n455
  );


  buf
  g714
  (
    n740,
    n731
  );


  not
  g715
  (
    n736,
    n730
  );


  not
  g716
  (
    n738,
    n688
  );


  not
  g717
  (
    n735,
    n688
  );


  not
  g718
  (
    n737,
    n732
  );


  nand
  g719
  (
    n739,
    n689,
    n730,
    n731
  );


  and
  g720
  (
    n741,
    n732,
    n689,
    n731
  );


  xor
  g721
  (
    n734,
    n731,
    n688,
    n689
  );


  buf
  g722
  (
    n748,
    n741
  );


  buf
  g723
  (
    n745,
    n739
  );


  not
  g724
  (
    n743,
    n735
  );


  buf
  g725
  (
    n747,
    n741
  );


  buf
  g726
  (
    n750,
    n734
  );


  buf
  g727
  (
    n746,
    n737
  );


  buf
  g728
  (
    n749,
    n736
  );


  buf
  g729
  (
    n744,
    n738
  );


  nand
  g730
  (
    n742,
    n732,
    n740
  );


  nand
  g731
  (
    n777,
    n745,
    n712,
    n727,
    n716
  );


  or
  g732
  (
    n770,
    n742,
    n744,
    n458,
    n728
  );


  or
  g733
  (
    n758,
    n706,
    n746,
    n724
  );


  nand
  g734
  (
    n785,
    n722,
    n723,
    n705,
    n725
  );


  xor
  g735
  (
    n762,
    n729,
    n723,
    n702,
    n750
  );


  nor
  g736
  (
    n764,
    n722,
    n710,
    n723,
    n749
  );


  xnor
  g737
  (
    n759,
    n750,
    n750,
    n717,
    n713
  );


  xnor
  g738
  (
    n778,
    n728,
    n747,
    n290,
    n702
  );


  xnor
  g739
  (
    n771,
    n291,
    n709,
    n743,
    n742
  );


  or
  g740
  (
    KeyWire_0_14,
    n711,
    n711,
    n746,
    n712
  );


  xor
  g741
  (
    n765,
    n729,
    n716,
    n709,
    n727
  );


  or
  g742
  (
    n780,
    n457,
    n462,
    n722,
    n290
  );


  or
  g743
  (
    n784,
    n744,
    n715,
    n714,
    n725
  );


  xnor
  g744
  (
    n761,
    n742,
    n744,
    n711,
    n723
  );


  xnor
  g745
  (
    n753,
    n465,
    n466,
    n748,
    n706
  );


  xor
  g746
  (
    n782,
    n713,
    n708,
    n710,
    n742
  );


  or
  g747
  (
    n786,
    n709,
    n705,
    n715
  );


  and
  g748
  (
    n773,
    n726,
    n708,
    n707,
    n728
  );


  nand
  g749
  (
    n752,
    n710,
    n464,
    n714,
    n745
  );


  nor
  g750
  (
    n781,
    n704,
    n290,
    n712,
    n743
  );


  xnor
  g751
  (
    n760,
    n746,
    n749,
    n291,
    n463
  );


  xnor
  g752
  (
    n783,
    n726,
    n748,
    n706,
    n747
  );


  nand
  g753
  (
    KeyWire_0_5,
    n717,
    n744,
    n749,
    n707
  );


  xor
  g754
  (
    n755,
    n714,
    n710,
    n290,
    n717
  );


  and
  g755
  (
    n754,
    n291,
    n724,
    n715,
    n705
  );


  nand
  g756
  (
    n768,
    n727,
    n459,
    n743,
    n712
  );


  xor
  g757
  (
    n769,
    n749,
    n708,
    n745,
    n746
  );


  nand
  g758
  (
    n766,
    n715,
    n726,
    n748,
    n724
  );


  or
  g759
  (
    n763,
    n460,
    n725,
    n461,
    n709
  );


  xor
  g760
  (
    n775,
    n727,
    n703,
    n748,
    n729
  );


  xor
  g761
  (
    n757,
    n726,
    n716,
    n728,
    n713
  );


  nand
  g762
  (
    n774,
    n713,
    n706,
    n745,
    n708
  );


  xor
  g763
  (
    n779,
    n750,
    n704,
    n711,
    n729
  );


  xnor
  g764
  (
    n772,
    n716,
    n747,
    n714,
    n703
  );


  and
  g765
  (
    n751,
    n704,
    n743,
    n707,
    n701
  );


  and
  g766
  (
    n756,
    n747,
    n707,
    n704,
    n725
  );


  not
  g767
  (
    n789,
    n754
  );


  not
  g768
  (
    n793,
    n753
  );


  buf
  g769
  (
    n788,
    n754
  );


  buf
  g770
  (
    n792,
    n752
  );


  not
  g771
  (
    n795,
    n755
  );


  buf
  g772
  (
    n790,
    n751
  );


  buf
  g773
  (
    n791,
    n752
  );


  buf
  g774
  (
    n794,
    n755
  );


  not
  g775
  (
    n787,
    n753
  );


  not
  g776
  (
    n796,
    n751
  );


  xnor
  g777
  (
    n798,
    n474,
    n475,
    n477,
    n467
  );


  nand
  g778
  (
    n800,
    n468,
    n760,
    n476,
    n759
  );


  xnor
  g779
  (
    n799,
    n471,
    n760,
    n787,
    n473
  );


  nand
  g780
  (
    n801,
    n469,
    n472,
    n758,
    n757
  );


  nand
  g781
  (
    n802,
    n787,
    n787,
    n788,
    n756
  );


  and
  g782
  (
    n797,
    n756,
    n759,
    n758,
    n788
  );


  nand
  g783
  (
    n803,
    n757,
    n787,
    n470,
    n788
  );


  nor
  g784
  (
    n808,
    n690,
    n691,
    n692
  );


  xnor
  g785
  (
    n805,
    n802,
    n690,
    n692,
    n691
  );


  nor
  g786
  (
    n807,
    n788,
    n690,
    n799
  );


  xor
  g787
  (
    n804,
    n693,
    n691,
    n789,
    n803
  );


  xor
  g788
  (
    n806,
    n800,
    n801,
    n692
  );


  nor
  g789
  (
    n816,
    n762,
    n783,
    n775,
    n808
  );


  xnor
  g790
  (
    n822,
    n804,
    n782,
    n779,
    n766
  );


  xor
  g791
  (
    n812,
    n779,
    n806,
    n781,
    n763
  );


  xnor
  g792
  (
    n814,
    n783,
    n805,
    n807
  );


  xnor
  g793
  (
    n821,
    n806,
    n808,
    n769
  );


  nand
  g794
  (
    n826,
    n776,
    n774,
    n808,
    n806
  );


  or
  g795
  (
    n818,
    n808,
    n807,
    n766,
    n782
  );


  or
  g796
  (
    n823,
    n780,
    n765,
    n805,
    n778
  );


  nor
  g797
  (
    n810,
    n807,
    n768,
    n780,
    n763
  );


  nor
  g798
  (
    n811,
    n761,
    n768,
    n804,
    n771
  );


  nand
  g799
  (
    n824,
    n783,
    n770,
    n807,
    n775
  );


  xnor
  g800
  (
    n820,
    n764,
    n780,
    n762,
    n805
  );


  and
  g801
  (
    n815,
    n783,
    n776,
    n774,
    n771
  );


  or
  g802
  (
    n817,
    n806,
    n780,
    n772,
    n782
  );


  or
  g803
  (
    n819,
    n773,
    n777,
    n764,
    n767
  );


  xnor
  g804
  (
    n813,
    n765,
    n778,
    n773,
    n777
  );


  xnor
  g805
  (
    n825,
    n761,
    n772,
    n782,
    n767
  );


  xnor
  g806
  (
    n809,
    n770,
    n781
  );


  xor
  g807
  (
    n846,
    n816,
    n786,
    n823,
    n792
  );


  nand
  g808
  (
    n845,
    n789,
    n824,
    n794,
    n785
  );


  nor
  g809
  (
    n835,
    n789,
    n732,
    n785,
    n811
  );


  xnor
  g810
  (
    n828,
    n794,
    n791,
    n795
  );


  xor
  g811
  (
    n844,
    n790,
    n796,
    n821,
    n791
  );


  or
  g812
  (
    n827,
    n478,
    n95,
    n795,
    n792
  );


  nand
  g813
  (
    n847,
    n824,
    n820,
    n826,
    n789
  );


  and
  g814
  (
    n833,
    n796,
    n784,
    n794
  );


  xnor
  g815
  (
    n829,
    n718,
    n815,
    n793,
    n693
  );


  xnor
  g816
  (
    n841,
    n786,
    n793,
    n95,
    n826
  );


  nor
  g817
  (
    n830,
    n814,
    n785,
    n813,
    n733
  );


  nor
  g818
  (
    n838,
    n796,
    n479,
    n693,
    n784
  );


  nor
  g819
  (
    n849,
    n786,
    n94,
    n822
  );


  nor
  g820
  (
    n840,
    n733,
    n95,
    n693,
    n786
  );


  nor
  g821
  (
    n839,
    n809,
    n822,
    n718,
    n792
  );


  and
  g822
  (
    n850,
    n823,
    n821,
    n795,
    n733
  );


  nand
  g823
  (
    n832,
    n733,
    n718,
    n819,
    n694
  );


  xnor
  g824
  (
    n843,
    n717,
    n481,
    n718,
    n95
  );


  and
  g825
  (
    n831,
    n485,
    n791,
    n793,
    n790
  );


  or
  g826
  (
    n837,
    n794,
    n790,
    n817
  );


  and
  g827
  (
    n848,
    n484,
    n825,
    n818,
    n784
  );


  xor
  g828
  (
    n836,
    n812,
    n483,
    n810,
    n482
  );


  and
  g829
  (
    n842,
    n719,
    n480,
    n793,
    n791
  );


  nor
  g830
  (
    n834,
    n796,
    n792,
    n825,
    n785
  );


  or
  g831
  (
    n865,
    n845,
    n519,
    n573,
    n539
  );


  xor
  g832
  (
    n863,
    n526,
    n506,
    n491,
    n493
  );


  or
  g833
  (
    KeyWire_0_27,
    n546,
    n848,
    n495,
    n521
  );


  or
  g834
  (
    n881,
    n499,
    n515,
    n568,
    n848
  );


  and
  g835
  (
    n852,
    n842,
    n831,
    n516,
    n553
  );


  xor
  g836
  (
    n867,
    n517,
    n846,
    n534,
    n505
  );


  nor
  g837
  (
    n878,
    n508,
    n549,
    n528,
    n850
  );


  xnor
  g838
  (
    n851,
    n843,
    n532,
    n494,
    n844
  );


  and
  g839
  (
    n873,
    n522,
    n838,
    n525,
    n575
  );


  nor
  g840
  (
    n879,
    n832,
    n489,
    n510,
    n828
  );


  nand
  g841
  (
    n861,
    n847,
    n541,
    n574,
    n502
  );


  xor
  g842
  (
    n876,
    n488,
    n529,
    n840,
    n846
  );


  and
  g843
  (
    n869,
    n511,
    n538,
    n847,
    n556
  );


  xor
  g844
  (
    n857,
    n837,
    n567,
    n514,
    n554
  );


  xor
  g845
  (
    n859,
    n542,
    n512,
    n555,
    n503
  );


  nand
  g846
  (
    n854,
    n500,
    n490,
    n518,
    n536
  );


  and
  g847
  (
    n858,
    n835,
    n487,
    n513,
    n560
  );


  and
  g848
  (
    n868,
    n527,
    n545,
    n558,
    n486
  );


  nor
  g849
  (
    n880,
    n830,
    n829,
    n850,
    n572
  );


  nor
  g850
  (
    n855,
    n849,
    n523,
    n566,
    n497
  );


  or
  g851
  (
    n862,
    n827,
    n533,
    n509,
    n559
  );


  nor
  g852
  (
    n871,
    n548,
    n552,
    n520,
    n849
  );


  nand
  g853
  (
    n866,
    n577,
    n565,
    n547,
    n496
  );


  nor
  g854
  (
    n877,
    n564,
    n498,
    n845,
    n841
  );


  nand
  g855
  (
    KeyWire_0_15,
    n844,
    n543,
    n833,
    n569
  );


  xnor
  g856
  (
    n864,
    n836,
    n551,
    n507,
    n557
  );


  xor
  g857
  (
    KeyWire_0_16,
    n578,
    n540,
    n537,
    n501
  );


  or
  g858
  (
    n853,
    n530,
    n561,
    n504,
    n563
  );


  xor
  g859
  (
    n872,
    n492,
    n570,
    n535,
    n524
  );


  nor
  g860
  (
    n870,
    n562,
    n576,
    n531,
    n544
  );


  nor
  g861
  (
    n875,
    n839,
    n571,
    n834,
    n550
  );


  buf
  g862
  (
    n885,
    n857
  );


  not
  g863
  (
    n883,
    n856
  );


  buf
  g864
  (
    n882,
    n858
  );


  buf
  g865
  (
    n884,
    n855
  );


  not
  g866
  (
    n890,
    n866
  );


  not
  g867
  (
    n895,
    n883
  );


  buf
  g868
  (
    n888,
    n861
  );


  not
  g869
  (
    n886,
    n882
  );


  xor
  g870
  (
    n893,
    n864,
    n579,
    n585,
    n884
  );


  xor
  g871
  (
    n894,
    n883,
    n581,
    n862,
    n882
  );


  and
  g872
  (
    n887,
    n586,
    n884,
    n583,
    n582
  );


  xnor
  g873
  (
    n891,
    n867,
    n580,
    n882,
    n863
  );


  xnor
  g874
  (
    n889,
    n865,
    n860,
    n584,
    n882
  );


  and
  g875
  (
    n892,
    n859,
    n883,
    n587
  );


  xor
  g876
  (
    n908,
    n872,
    n888,
    n886,
    n876
  );


  or
  g877
  (
    n911,
    n886,
    n889
  );


  xor
  g878
  (
    n900,
    n890,
    n885,
    n879,
    n869
  );


  xnor
  g879
  (
    KeyWire_0_1,
    n889,
    n878,
    n887,
    n293
  );


  xor
  g880
  (
    n904,
    n295,
    n293,
    n888,
    n886
  );


  and
  g881
  (
    n896,
    n292,
    n873,
    n876,
    n293
  );


  nand
  g882
  (
    n902,
    n873,
    n872,
    n291,
    n887
  );


  xnor
  g883
  (
    n897,
    n294,
    n296,
    n867,
    n884
  );


  nor
  g884
  (
    n899,
    n889,
    n871,
    n294,
    n875
  );


  nand
  g885
  (
    n901,
    n294,
    n884,
    n878,
    n870
  );


  and
  g886
  (
    n910,
    n875,
    n888,
    n871,
    n885
  );


  nand
  g887
  (
    n907,
    n295,
    n890,
    n885,
    n292
  );


  or
  g888
  (
    n909,
    n885,
    n292,
    n296,
    n294
  );


  nor
  g889
  (
    n912,
    n888,
    n295,
    n874,
    n877
  );


  or
  g890
  (
    n905,
    n292,
    n887,
    n877
  );


  nand
  g891
  (
    n906,
    n293,
    n869,
    n296,
    n874
  );


  nand
  g892
  (
    n903,
    n868,
    n868,
    n870,
    n295
  );


  not
  g893
  (
    n913,
    n896
  );


  nor
  g894
  (
    n914,
    n880,
    n897,
    n879
  );


  or
  g895
  (
    n915,
    n914,
    n881,
    n880
  );


  nor
  g896
  (
    n917,
    n890,
    n915,
    n891
  );


  xor
  g897
  (
    n916,
    n892,
    n893,
    n915
  );


  or
  g898
  (
    n918,
    n892,
    n891
  );


  nor
  g899
  (
    n919,
    n915,
    n892,
    n893,
    n890
  );


  or
  g900
  (
    n925,
    n895,
    n903,
    n916,
    n917
  );


  xnor
  g901
  (
    n922,
    n591,
    n589,
    n919,
    n893
  );


  xor
  g902
  (
    n930,
    n609,
    n917,
    n608,
    n916
  );


  and
  g903
  (
    n928,
    n595,
    n895,
    n917,
    n893
  );


  or
  g904
  (
    n923,
    n603,
    n909,
    n592,
    n602
  );


  or
  g905
  (
    n927,
    n894,
    n901,
    n590,
    n604
  );


  nand
  g906
  (
    n934,
    n597,
    n904,
    n919,
    n900
  );


  xnor
  g907
  (
    n935,
    n912,
    n894,
    n593,
    n594
  );


  xnor
  g908
  (
    n924,
    n905,
    n898,
    n599,
    n600
  );


  nand
  g909
  (
    n932,
    n908,
    n899,
    n606,
    n919
  );


  xnor
  g910
  (
    n933,
    n918,
    n911,
    n588,
    n895
  );


  nor
  g911
  (
    n931,
    n916,
    n902,
    n601,
    n919
  );


  or
  g912
  (
    n929,
    n894,
    n907,
    n918,
    n906
  );


  nand
  g913
  (
    n920,
    n610,
    n598,
    n894,
    n916
  );


  and
  g914
  (
    n926,
    n596,
    n605,
    n918,
    n895
  );


  or
  g915
  (
    n921,
    n917,
    n910,
    n918,
    n607
  );


  or
  g916
  (
    n938,
    n695,
    n924,
    n935,
    n931
  );


  xnor
  g917
  (
    n939,
    n920,
    n694,
    n927
  );


  xor
  g918
  (
    n941,
    n611,
    n695,
    n921
  );


  and
  g919
  (
    n936,
    n719,
    n932,
    n933,
    n695
  );


  xor
  g920
  (
    n942,
    n928,
    n930,
    n926,
    n719
  );


  and
  g921
  (
    KeyWire_0_21,
    n925,
    n934,
    n923,
    n719
  );


  nor
  g922
  (
    n937,
    n694,
    n929,
    n296,
    n922
  );


  xor
  KeyGate_0_0
  (
    n457,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n898,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n613,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n728,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n130,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n776,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n429,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n566,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n666,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n385,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n23,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n652,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n221,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n499,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n767,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n856,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n860,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n550,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n119,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n318,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n380,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n940,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n394,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n508,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n280,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n721,
    keyIn_0_25,
    KeyWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n95,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n874,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n482,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n559,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n584,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n607,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule

