// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_322 written by SynthGen on 2021/04/05 11:24:15
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_3000_322 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n2756, n2798, n2787, n2805, n2775, n2799, n2802, n2788,
 n2807, n2808, n2796, n2801, n2777, n2783, n2779, n2791,
 n2789, n2792, n2784, n2782, n2786, n2804, n2778, n2800,
 n2785, n2809, n2780, n2793, n2790, n2803, n2906, n3032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n2756, n2798, n2787, n2805, n2775, n2799, n2802, n2788,
 n2807, n2808, n2796, n2801, n2777, n2783, n2779, n2791,
 n2789, n2792, n2784, n2782, n2786, n2804, n2778, n2800,
 n2785, n2809, n2780, n2793, n2790, n2803, n2906, n3032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n638, n639, n640,
 n641, n642, n643, n644, n645, n646, n647, n648,
 n649, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n668, n669, n670, n671, n672,
 n673, n674, n675, n676, n677, n678, n679, n680,
 n681, n682, n683, n684, n685, n686, n687, n688,
 n689, n690, n691, n692, n693, n694, n695, n696,
 n697, n698, n699, n700, n701, n702, n703, n704,
 n705, n706, n707, n708, n709, n710, n711, n712,
 n713, n714, n715, n716, n717, n718, n719, n720,
 n721, n722, n723, n724, n725, n726, n727, n728,
 n729, n730, n731, n732, n733, n734, n735, n736,
 n737, n738, n739, n740, n741, n742, n743, n744,
 n745, n746, n747, n748, n749, n750, n751, n752,
 n753, n754, n755, n756, n757, n758, n759, n760,
 n761, n762, n763, n764, n765, n766, n767, n768,
 n769, n770, n771, n772, n773, n774, n775, n776,
 n777, n778, n779, n780, n781, n782, n783, n784,
 n785, n786, n787, n788, n789, n790, n791, n792,
 n793, n794, n795, n796, n797, n798, n799, n800,
 n801, n802, n803, n804, n805, n806, n807, n808,
 n809, n810, n811, n812, n813, n814, n815, n816,
 n817, n818, n819, n820, n821, n822, n823, n824,
 n825, n826, n827, n828, n829, n830, n831, n832,
 n833, n834, n835, n836, n837, n838, n839, n840,
 n841, n842, n843, n844, n845, n846, n847, n848,
 n849, n850, n851, n852, n853, n854, n855, n856,
 n857, n858, n859, n860, n861, n862, n863, n864,
 n865, n866, n867, n868, n869, n870, n871, n872,
 n873, n874, n875, n876, n877, n878, n879, n880,
 n881, n882, n883, n884, n885, n886, n887, n888,
 n889, n890, n891, n892, n893, n894, n895, n896,
 n897, n898, n899, n900, n901, n902, n903, n904,
 n905, n906, n907, n908, n909, n910, n911, n912,
 n913, n914, n915, n916, n917, n918, n919, n920,
 n921, n922, n923, n924, n925, n926, n927, n928,
 n929, n930, n931, n932, n933, n934, n935, n936,
 n937, n938, n939, n940, n941, n942, n943, n944,
 n945, n946, n947, n948, n949, n950, n951, n952,
 n953, n954, n955, n956, n957, n958, n959, n960,
 n961, n962, n963, n964, n965, n966, n967, n968,
 n969, n970, n971, n972, n973, n974, n975, n976,
 n977, n978, n979, n980, n981, n982, n983, n984,
 n985, n986, n987, n988, n989, n990, n991, n992,
 n993, n994, n995, n996, n997, n998, n999, n1000,
 n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
 n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
 n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
 n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
 n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
 n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
 n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
 n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
 n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
 n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
 n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
 n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
 n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
 n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
 n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
 n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
 n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
 n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
 n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
 n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
 n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
 n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
 n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
 n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
 n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
 n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
 n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
 n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
 n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
 n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
 n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
 n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
 n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
 n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
 n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
 n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
 n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
 n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
 n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
 n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
 n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
 n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
 n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
 n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
 n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
 n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
 n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
 n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
 n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
 n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
 n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
 n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
 n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
 n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
 n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
 n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
 n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
 n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
 n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
 n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
 n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
 n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
 n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
 n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
 n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
 n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
 n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
 n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
 n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
 n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
 n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
 n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
 n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
 n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
 n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
 n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
 n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
 n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
 n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
 n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
 n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
 n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
 n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
 n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
 n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
 n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
 n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
 n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
 n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
 n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
 n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
 n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
 n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
 n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
 n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
 n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
 n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
 n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
 n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
 n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
 n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
 n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
 n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
 n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
 n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
 n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
 n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
 n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
 n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
 n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
 n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
 n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
 n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
 n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
 n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
 n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
 n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936,
 n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
 n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
 n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
 n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
 n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976,
 n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
 n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
 n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
 n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
 n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016,
 n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
 n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
 n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
 n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
 n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056,
 n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
 n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
 n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
 n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
 n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096,
 n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
 n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
 n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
 n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
 n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136,
 n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
 n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
 n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
 n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
 n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176,
 n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
 n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
 n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
 n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
 n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216,
 n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
 n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
 n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
 n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
 n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256,
 n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
 n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
 n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
 n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
 n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296,
 n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
 n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
 n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
 n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
 n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336,
 n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
 n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
 n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
 n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
 n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376,
 n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
 n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
 n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
 n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
 n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
 n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
 n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
 n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
 n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
 n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456,
 n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
 n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
 n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
 n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
 n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496,
 n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
 n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
 n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
 n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
 n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536,
 n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
 n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
 n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
 n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
 n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576,
 n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
 n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
 n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
 n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
 n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616,
 n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
 n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
 n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
 n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
 n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
 n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
 n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
 n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
 n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
 n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
 n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
 n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
 n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
 n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
 n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
 n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
 n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
 n2753, n2754, n2755, n2757, n2758, n2759, n2760, n2761,
 n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
 n2770, n2771, n2772, n2773, n2774, n2776, n2781, n2794,
 n2795, n2797, n2806, n2810, n2811, n2812, n2813, n2814,
 n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
 n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
 n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
 n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
 n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
 n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
 n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
 n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
 n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
 n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
 n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
 n2903, n2904, n2905, n2907, n2908, n2909, n2910, n2911,
 n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
 n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
 n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
 n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
 n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
 n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
 n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
 n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
 n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
 n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
 n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
 n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
 n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
 n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
 n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031;

not  g0 (n56, n22);
buf  g1 (n59, n11);
not  g2 (n125, n11);
not  g3 (n101, n18);
not  g4 (n81, n12);
buf  g5 (n94, n3);
buf  g6 (n39, n23);
buf  g7 (n96, n28);
buf  g8 (n70, n27);
buf  g9 (n83, n13);
buf  g10 (n119, n23);
buf  g11 (n54, n3);
not  g12 (n95, n21);
not  g13 (n82, n12);
not  g14 (n75, n13);
not  g15 (n86, n12);
buf  g16 (n131, n5);
buf  g17 (n51, n25);
buf  g18 (n110, n6);
buf  g19 (n53, n17);
buf  g20 (n106, n10);
not  g21 (n58, n4);
not  g22 (n60, n14);
buf  g23 (n73, n2);
not  g24 (n62, n25);
not  g25 (n111, n19);
buf  g26 (n118, n18);
not  g27 (n33, n3);
buf  g28 (n116, n27);
not  g29 (n115, n10);
buf  g30 (n55, n16);
not  g31 (n84, n14);
buf  g32 (n122, n11);
buf  g33 (n142, n21);
not  g34 (n132, n20);
buf  g35 (n77, n26);
buf  g36 (n105, n23);
not  g37 (n61, n5);
not  g38 (n103, n20);
not  g39 (n93, n23);
not  g40 (n92, n14);
buf  g41 (n44, n8);
not  g42 (n35, n8);
not  g43 (n138, n21);
not  g44 (n74, n27);
buf  g45 (n109, n28);
not  g46 (n48, n2);
buf  g47 (n99, n2);
not  g48 (n41, n24);
buf  g49 (n113, n7);
buf  g50 (n43, n25);
not  g51 (n45, n16);
buf  g52 (n78, n24);
not  g53 (n49, n15);
not  g54 (n69, n4);
buf  g55 (n141, n3);
not  g56 (n133, n15);
not  g57 (n80, n9);
not  g58 (n134, n28);
buf  g59 (n137, n1);
buf  g60 (n143, n5);
not  g61 (n104, n16);
buf  g62 (n34, n7);
not  g63 (n117, n27);
buf  g64 (n135, n12);
not  g65 (n64, n24);
buf  g66 (n140, n1);
buf  g67 (n102, n9);
buf  g68 (n114, n22);
buf  g69 (n139, n19);
not  g70 (n87, n13);
buf  g71 (n76, n11);
not  g72 (n36, n14);
buf  g73 (n124, n28);
not  g74 (n88, n22);
not  g75 (n50, n1);
buf  g76 (n68, n2);
not  g77 (n136, n7);
not  g78 (n40, n6);
buf  g79 (n90, n10);
buf  g80 (n127, n17);
buf  g81 (n121, n17);
buf  g82 (n52, n8);
buf  g83 (n72, n9);
buf  g84 (n91, n26);
not  g85 (n89, n20);
not  g86 (n144, n19);
buf  g87 (n65, n26);
buf  g88 (n98, n13);
not  g89 (n100, n15);
not  g90 (n120, n24);
buf  g91 (n123, n8);
not  g92 (n67, n6);
buf  g93 (n130, n25);
not  g94 (n71, n18);
buf  g95 (n128, n18);
not  g96 (n112, n10);
buf  g97 (n46, n1);
buf  g98 (n42, n4);
buf  g99 (n66, n4);
buf  g100 (n57, n17);
buf  g101 (n85, n6);
not  g102 (n79, n26);
not  g103 (n126, n22);
not  g104 (n63, n5);
buf  g105 (n97, n15);
not  g106 (n47, n9);
not  g107 (n37, n20);
buf  g108 (n107, n21);
buf  g109 (n38, n7);
buf  g110 (n129, n19);
buf  g111 (n108, n16);
not  g112 (n378, n124);
not  g113 (n261, n59);
buf  g114 (n552, n129);
buf  g115 (n197, n87);
not  g116 (n525, n45);
not  g117 (n463, n127);
buf  g118 (n510, n118);
buf  g119 (n461, n122);
not  g120 (n312, n85);
not  g121 (n392, n104);
buf  g122 (n405, n76);
buf  g123 (n207, n104);
buf  g124 (n333, n91);
not  g125 (n145, n132);
buf  g126 (n361, n142);
not  g127 (n176, n137);
not  g128 (n247, n41);
not  g129 (n239, n57);
buf  g130 (n534, n37);
buf  g131 (n386, n107);
buf  g132 (n523, n94);
not  g133 (n188, n119);
buf  g134 (n340, n63);
not  g135 (n388, n39);
not  g136 (n337, n142);
not  g137 (n230, n38);
not  g138 (n157, n57);
buf  g139 (n291, n123);
not  g140 (n183, n135);
not  g141 (n250, n75);
not  g142 (n406, n111);
buf  g143 (n258, n112);
buf  g144 (n536, n142);
not  g145 (n179, n83);
buf  g146 (n416, n93);
buf  g147 (n278, n40);
not  g148 (n351, n67);
buf  g149 (n509, n45);
not  g150 (n529, n123);
buf  g151 (n483, n55);
buf  g152 (n496, n120);
not  g153 (n297, n46);
not  g154 (n276, n116);
not  g155 (n399, n88);
not  g156 (n381, n36);
buf  g157 (n332, n43);
not  g158 (n253, n143);
buf  g159 (n477, n81);
not  g160 (n444, n139);
not  g161 (n453, n112);
not  g162 (n501, n91);
buf  g163 (n445, n85);
buf  g164 (n224, n67);
buf  g165 (n580, n125);
not  g166 (n262, n138);
not  g167 (n191, n105);
not  g168 (n284, n34);
not  g169 (n274, n41);
not  g170 (n317, n130);
buf  g171 (n216, n54);
not  g172 (n175, n135);
not  g173 (n422, n109);
not  g174 (n160, n70);
buf  g175 (n209, n141);
buf  g176 (n321, n61);
buf  g177 (n158, n51);
not  g178 (n283, n52);
buf  g179 (n478, n73);
buf  g180 (n513, n107);
not  g181 (n347, n51);
buf  g182 (n379, n101);
not  g183 (n555, n86);
not  g184 (n231, n53);
not  g185 (n561, n128);
not  g186 (n458, n48);
buf  g187 (n225, n129);
buf  g188 (n572, n89);
not  g189 (n193, n130);
buf  g190 (n409, n89);
not  g191 (n498, n47);
buf  g192 (n148, n93);
not  g193 (n526, n69);
not  g194 (n557, n74);
not  g195 (n192, n139);
not  g196 (n280, n112);
not  g197 (n485, n42);
not  g198 (n369, n110);
not  g199 (n189, n99);
buf  g200 (n232, n86);
buf  g201 (n475, n84);
buf  g202 (n168, n122);
not  g203 (n571, n79);
not  g204 (n431, n100);
not  g205 (n266, n47);
not  g206 (n420, n73);
buf  g207 (n376, n78);
buf  g208 (n447, n94);
not  g209 (n565, n35);
not  g210 (n546, n97);
buf  g211 (n588, n76);
not  g212 (n181, n90);
buf  g213 (n511, n109);
not  g214 (n198, n128);
buf  g215 (n357, n98);
not  g216 (n413, n127);
not  g217 (n150, n99);
not  g218 (n470, n143);
buf  g219 (n293, n69);
buf  g220 (n411, n106);
buf  g221 (n307, n40);
buf  g222 (n156, n81);
buf  g223 (n202, n91);
buf  g224 (n504, n37);
not  g225 (n305, n117);
buf  g226 (n272, n96);
buf  g227 (n449, n140);
not  g228 (n566, n94);
buf  g229 (n177, n94);
buf  g230 (n304, n34);
not  g231 (n573, n72);
buf  g232 (n185, n138);
not  g233 (n541, n128);
buf  g234 (n334, n87);
buf  g235 (n540, n102);
buf  g236 (n296, n63);
buf  g237 (n516, n67);
not  g238 (n348, n121);
buf  g239 (n371, n79);
not  g240 (n235, n103);
not  g241 (n178, n79);
buf  g242 (n290, n100);
buf  g243 (n465, n118);
not  g244 (n396, n60);
not  g245 (n473, n48);
buf  g246 (n295, n88);
buf  g247 (n173, n46);
not  g248 (n382, n35);
not  g249 (n389, n80);
buf  g250 (n315, n54);
buf  g251 (n339, n65);
buf  g252 (n490, n139);
buf  g253 (n301, n71);
not  g254 (n535, n88);
buf  g255 (n264, n123);
not  g256 (n578, n101);
buf  g257 (n481, n126);
not  g258 (n257, n143);
buf  g259 (n518, n48);
not  g260 (n414, n129);
not  g261 (n374, n41);
buf  g262 (n208, n104);
not  g263 (n433, n136);
not  g264 (n331, n140);
buf  g265 (n375, n44);
not  g266 (n244, n52);
buf  g267 (n352, n111);
buf  g268 (n459, n144);
not  g269 (n577, n84);
not  g270 (n243, n77);
buf  g271 (n538, n40);
buf  g272 (n583, n114);
not  g273 (n441, n126);
not  g274 (n214, n47);
not  g275 (n204, n103);
buf  g276 (n466, n70);
buf  g277 (n533, n116);
not  g278 (n424, n82);
buf  g279 (n165, n86);
buf  g280 (n575, n133);
buf  g281 (n520, n56);
not  g282 (n316, n60);
buf  g283 (n373, n134);
buf  g284 (n170, n85);
not  g285 (n328, n69);
buf  g286 (n454, n97);
buf  g287 (n482, n85);
buf  g288 (n237, n132);
not  g289 (n556, n139);
buf  g290 (n314, n83);
not  g291 (n545, n121);
not  g292 (n436, n119);
not  g293 (n497, n101);
buf  g294 (n443, n95);
not  g295 (n155, n38);
buf  g296 (n455, n55);
not  g297 (n159, n72);
not  g298 (n537, n86);
buf  g299 (n362, n39);
buf  g300 (n383, n110);
buf  g301 (n363, n98);
buf  g302 (n318, n119);
not  g303 (n323, n99);
buf  g304 (n452, n134);
not  g305 (n292, n90);
buf  g306 (n456, n124);
buf  g307 (n506, n112);
buf  g308 (n200, n87);
not  g309 (n223, n44);
not  g310 (n147, n113);
not  g311 (n408, n142);
not  g312 (n234, n124);
not  g313 (n169, n130);
not  g314 (n403, n58);
not  g315 (n367, n44);
buf  g316 (n270, n49);
not  g317 (n528, n111);
not  g318 (n310, n69);
buf  g319 (n275, n114);
not  g320 (n249, n84);
buf  g321 (n584, n56);
not  g322 (n587, n113);
buf  g323 (n218, n87);
not  g324 (n576, n143);
not  g325 (n279, n88);
buf  g326 (n567, n45);
not  g327 (n486, n46);
not  g328 (n222, n106);
not  g329 (n282, n37);
not  g330 (n564, n57);
not  g331 (n417, n40);
buf  g332 (n384, n60);
buf  g333 (n320, n140);
buf  g334 (n236, n108);
not  g335 (n400, n122);
buf  g336 (n263, n134);
not  g337 (n429, n120);
buf  g338 (n350, n61);
not  g339 (n586, n102);
not  g340 (n162, n50);
buf  g341 (n172, n33);
not  g342 (n194, n35);
buf  g343 (n560, n68);
buf  g344 (n402, n74);
buf  g345 (n472, n118);
not  g346 (n343, n47);
not  g347 (n495, n56);
buf  g348 (n558, n120);
buf  g349 (n353, n53);
not  g350 (n161, n98);
buf  g351 (n423, n58);
buf  g352 (n206, n107);
buf  g353 (n440, n42);
buf  g354 (n151, n33);
buf  g355 (n366, n80);
not  g356 (n233, n115);
buf  g357 (n269, n71);
buf  g358 (n248, n43);
buf  g359 (n539, n115);
buf  g360 (n471, n122);
buf  g361 (n356, n92);
not  g362 (n507, n131);
not  g363 (n568, n89);
buf  g364 (n460, n117);
buf  g365 (n585, n53);
not  g366 (n527, n127);
not  g367 (n322, n75);
not  g368 (n241, n109);
not  g369 (n186, n92);
buf  g370 (n574, n103);
buf  g371 (n238, n73);
not  g372 (n346, n141);
buf  g373 (n467, n73);
buf  g374 (n256, n42);
buf  g375 (n438, n74);
not  g376 (n450, n50);
not  g377 (n260, n80);
buf  g378 (n265, n115);
buf  g379 (n338, n81);
buf  g380 (n308, n108);
not  g381 (n427, n107);
buf  g382 (n474, n66);
buf  g383 (n149, n104);
not  g384 (n562, n95);
buf  g385 (n401, n34);
not  g386 (n294, n90);
buf  g387 (n268, n77);
buf  g388 (n152, n91);
not  g389 (n298, n72);
not  g390 (n434, n138);
not  g391 (n415, n113);
buf  g392 (n252, n34);
not  g393 (n324, n133);
not  g394 (n220, n39);
buf  g395 (n255, n134);
buf  g396 (n164, n55);
buf  g397 (n306, n68);
not  g398 (n184, n38);
not  g399 (n468, n39);
buf  g400 (n319, n78);
not  g401 (n563, n33);
buf  g402 (n211, n114);
buf  g403 (n311, n52);
not  g404 (n153, n41);
buf  g405 (n419, n111);
not  g406 (n227, n109);
not  g407 (n502, n137);
buf  g408 (n451, n138);
not  g409 (n421, n132);
buf  g410 (n457, n133);
buf  g411 (n508, n131);
not  g412 (n286, n93);
buf  g413 (n488, n65);
not  g414 (n245, n116);
buf  g415 (n554, n54);
buf  g416 (n167, n89);
buf  g417 (n480, n100);
buf  g418 (n242, n60);
not  g419 (n313, n129);
not  g420 (n418, n121);
buf  g421 (n462, n115);
buf  g422 (n358, n59);
not  g423 (n146, n92);
not  g424 (n364, n125);
buf  g425 (n385, n76);
not  g426 (n412, n43);
buf  g427 (n288, n106);
not  g428 (n330, n95);
buf  g429 (n309, n95);
buf  g430 (n469, n120);
buf  g431 (n489, n58);
not  g432 (n548, n49);
not  g433 (n300, n45);
buf  g434 (n163, n110);
not  g435 (n395, n132);
buf  g436 (n464, n52);
not  g437 (n182, n126);
not  g438 (n551, n59);
buf  g439 (n448, n61);
buf  g440 (n210, n108);
buf  g441 (n267, n75);
buf  g442 (n299, n62);
buf  g443 (n530, n99);
buf  g444 (n240, n108);
buf  g445 (n393, n72);
not  g446 (n212, n62);
buf  g447 (n277, n33);
not  g448 (n581, n137);
buf  g449 (n505, n67);
not  g450 (n215, n127);
buf  g451 (n582, n124);
not  g452 (n368, n97);
buf  g453 (n285, n105);
buf  g454 (n425, n121);
buf  g455 (n273, n102);
not  g456 (n171, n75);
not  g457 (n543, n106);
not  g458 (n589, n80);
not  g459 (n391, n114);
not  g460 (n326, n43);
buf  g461 (n404, n125);
buf  g462 (n335, n113);
not  g463 (n226, n131);
not  g464 (n387, n82);
not  g465 (n246, n130);
buf  g466 (n199, n50);
buf  g467 (n579, n68);
buf  g468 (n187, n49);
buf  g469 (n341, n116);
not  g470 (n345, n54);
buf  g471 (n336, n82);
buf  g472 (n360, n123);
not  g473 (n166, n71);
buf  g474 (n428, n62);
buf  g475 (n355, n70);
not  g476 (n550, n78);
buf  g477 (n514, n76);
buf  g478 (n435, n133);
buf  g479 (n519, n103);
not  g480 (n410, n97);
not  g481 (n476, n64);
buf  g482 (n377, n140);
buf  g483 (n397, n141);
not  g484 (n532, n141);
buf  g485 (n372, n42);
buf  g486 (n201, n110);
not  g487 (n570, n90);
buf  g488 (n205, n96);
not  g489 (n196, n58);
buf  g490 (n370, n65);
not  g491 (n432, n64);
not  g492 (n430, n63);
not  g493 (n544, n35);
buf  g494 (n491, n56);
not  g495 (n515, n53);
not  g496 (n380, n135);
buf  g497 (n549, n36);
buf  g498 (n344, n66);
not  g499 (n494, n66);
buf  g500 (n359, n135);
not  g501 (n190, n64);
not  g502 (n439, n68);
not  g503 (n327, n66);
not  g504 (n442, n102);
buf  g505 (n517, n36);
buf  g506 (n559, n100);
buf  g507 (n398, n51);
buf  g508 (n487, n136);
not  g509 (n289, n92);
buf  g510 (n569, n64);
not  g511 (n154, n119);
buf  g512 (n271, n50);
not  g513 (n394, n57);
buf  g514 (n521, n136);
not  g515 (n342, n131);
not  g516 (n228, n37);
not  g517 (n221, n105);
not  g518 (n547, n117);
buf  g519 (n390, n63);
not  g520 (n180, n101);
not  g521 (n281, n59);
buf  g522 (n354, n83);
not  g523 (n522, n105);
not  g524 (n365, n126);
not  g525 (n174, n125);
buf  g526 (n492, n93);
buf  g527 (n524, n77);
buf  g528 (n349, n36);
not  g529 (n303, n44);
not  g530 (n437, n78);
buf  g531 (n503, n137);
not  g532 (n499, n83);
buf  g533 (n251, n38);
buf  g534 (n302, n48);
buf  g535 (n446, n96);
not  g536 (n553, n61);
buf  g537 (n531, n79);
not  g538 (n213, n62);
not  g539 (n254, n98);
buf  g540 (n259, n118);
buf  g541 (n407, n136);
not  g542 (n195, n128);
not  g543 (n479, n65);
not  g544 (n542, n96);
buf  g545 (n325, n74);
not  g546 (n229, n46);
not  g547 (n329, n55);
not  g548 (n219, n117);
not  g549 (n493, n84);
buf  g550 (n426, n70);
buf  g551 (n512, n71);
buf  g552 (n500, n49);
buf  g553 (n203, n51);
buf  g554 (n217, n77);
buf  g555 (n484, n82);
buf  g556 (n287, n81);
buf  g557 (n1481, n470);
not  g558 (n1418, n239);
not  g559 (n1312, n516);
not  g560 (n1809, n538);
buf  g561 (n634, n332);
not  g562 (n1083, n514);
not  g563 (n866, n217);
buf  g564 (n659, n307);
not  g565 (n864, n334);
buf  g566 (n1104, n456);
buf  g567 (n1766, n229);
buf  g568 (n1718, n464);
buf  g569 (n1146, n510);
not  g570 (n654, n179);
buf  g571 (n1703, n262);
buf  g572 (n1195, n225);
buf  g573 (n712, n216);
not  g574 (n1080, n506);
not  g575 (n1183, n203);
not  g576 (n1212, n172);
buf  g577 (n1497, n313);
buf  g578 (n1675, n261);
buf  g579 (n1690, n450);
not  g580 (n1031, n453);
not  g581 (n1236, n406);
not  g582 (n964, n291);
buf  g583 (n1658, n214);
buf  g584 (n1492, n240);
buf  g585 (n1231, n176);
buf  g586 (n749, n451);
not  g587 (n899, n191);
buf  g588 (n1157, n321);
buf  g589 (n1523, n469);
buf  g590 (n775, n309);
buf  g591 (n1754, n306);
buf  g592 (n966, n509);
buf  g593 (n853, n443);
buf  g594 (n818, n448);
not  g595 (n1833, n469);
buf  g596 (n714, n531);
buf  g597 (n822, n301);
buf  g598 (n1151, n396);
buf  g599 (n1503, n354);
not  g600 (n1291, n417);
not  g601 (n1267, n365);
buf  g602 (n956, n425);
not  g603 (n1328, n214);
not  g604 (n989, n537);
not  g605 (n1731, n255);
buf  g606 (n1502, n472);
not  g607 (n1232, n184);
buf  g608 (n1223, n397);
not  g609 (n1780, n292);
not  g610 (n833, n431);
buf  g611 (n1471, n295);
buf  g612 (n856, n173);
not  g613 (n801, n440);
buf  g614 (n1821, n246);
buf  g615 (n1729, n222);
buf  g616 (n1327, n355);
not  g617 (n1406, n285);
not  g618 (n803, n420);
not  g619 (n1803, n278);
not  g620 (n1182, n367);
buf  g621 (n1525, n248);
not  g622 (n1558, n375);
not  g623 (n927, n426);
buf  g624 (n1679, n363);
not  g625 (n1217, n497);
not  g626 (n1113, n240);
not  g627 (n787, n170);
not  g628 (n1629, n434);
buf  g629 (n1022, n343);
buf  g630 (n1672, n515);
buf  g631 (n1135, n532);
not  g632 (n1596, n269);
buf  g633 (n1184, n319);
buf  g634 (n1448, n231);
not  g635 (n697, n415);
buf  g636 (n898, n382);
buf  g637 (n759, n510);
buf  g638 (n962, n405);
buf  g639 (n1190, n342);
not  g640 (n736, n175);
not  g641 (n1401, n396);
buf  g642 (n725, n283);
not  g643 (n1056, n289);
buf  g644 (n790, n359);
not  g645 (n1518, n406);
not  g646 (n1079, n335);
buf  g647 (n1815, n498);
not  g648 (n1255, n418);
not  g649 (n1608, n510);
not  g650 (n1588, n353);
not  g651 (n1090, n167);
buf  g652 (n999, n441);
buf  g653 (n1786, n453);
buf  g654 (n1379, n440);
not  g655 (n987, n448);
buf  g656 (n1823, n457);
buf  g657 (n1218, n430);
not  g658 (n1078, n220);
buf  g659 (n1553, n490);
not  g660 (n619, n258);
buf  g661 (n988, n426);
buf  g662 (n640, n264);
buf  g663 (n1562, n453);
not  g664 (n1038, n354);
not  g665 (n679, n303);
buf  g666 (n741, n410);
buf  g667 (n1094, n232);
not  g668 (n1433, n349);
not  g669 (n1572, n449);
not  g670 (n1004, n202);
buf  g671 (n1704, n265);
not  g672 (n1605, n440);
buf  g673 (n812, n388);
not  g674 (n844, n316);
not  g675 (n1213, n146);
not  g676 (n1555, n198);
not  g677 (n1033, n459);
buf  g678 (n636, n467);
not  g679 (n976, n363);
not  g680 (n1021, n329);
not  g681 (n707, n358);
not  g682 (n1480, n231);
not  g683 (n792, n151);
buf  g684 (n1771, n302);
not  g685 (n1606, n506);
not  g686 (n1086, n474);
not  g687 (n1561, n220);
buf  g688 (n832, n431);
buf  g689 (n1381, n266);
not  g690 (n1646, n381);
not  g691 (n1458, n325);
not  g692 (n1805, n314);
not  g693 (n1837, n424);
buf  g694 (n1622, n503);
buf  g695 (n1340, n495);
buf  g696 (n873, n224);
not  g697 (n931, n163);
not  g698 (n1246, n252);
not  g699 (n1466, n383);
not  g700 (n1493, n363);
buf  g701 (n862, n393);
buf  g702 (n648, n485);
buf  g703 (n1791, n410);
not  g704 (n609, n473);
not  g705 (n973, n213);
not  g706 (n1706, n239);
buf  g707 (n1166, n538);
buf  g708 (n1306, n337);
not  g709 (n1550, n211);
buf  g710 (n768, n263);
not  g711 (n1781, n535);
buf  g712 (n940, n379);
not  g713 (n932, n398);
not  g714 (n1334, n333);
not  g715 (n1478, n337);
not  g716 (n1724, n177);
buf  g717 (n1778, n159);
not  g718 (n1632, n294);
not  g719 (n1160, n372);
not  g720 (n1348, n436);
not  g721 (n1649, n362);
buf  g722 (n1573, n181);
buf  g723 (n817, n402);
buf  g724 (n903, n463);
not  g725 (n1095, n316);
not  g726 (n657, n434);
buf  g727 (n1473, n479);
buf  g728 (n891, n198);
buf  g729 (n724, n309);
not  g730 (n1536, n264);
not  g731 (n752, n289);
buf  g732 (n1100, n333);
not  g733 (n1696, n357);
buf  g734 (n1792, n323);
not  g735 (n1353, n463);
not  g736 (n594, n511);
buf  g737 (n793, n394);
not  g738 (n992, n504);
buf  g739 (n1013, n371);
not  g740 (n1584, n405);
not  g741 (n1419, n474);
not  g742 (n1272, n361);
not  g743 (n878, n183);
buf  g744 (n945, n494);
not  g745 (n690, n465);
buf  g746 (n951, n178);
not  g747 (n1585, n233);
not  g748 (n1730, n538);
not  g749 (n1609, n496);
not  g750 (n1633, n394);
not  g751 (n1621, n251);
not  g752 (n849, n255);
buf  g753 (n1126, n310);
not  g754 (n1544, n413);
not  g755 (n1738, n180);
buf  g756 (n1137, n153);
buf  g757 (n1671, n258);
not  g758 (n875, n328);
not  g759 (n1637, n249);
not  g760 (n1423, n299);
not  g761 (n614, n260);
buf  g762 (n895, n422);
not  g763 (n1265, n257);
buf  g764 (n1338, n220);
not  g765 (n715, n381);
buf  g766 (n1114, n193);
not  g767 (n1412, n194);
buf  g768 (n1198, n303);
buf  g769 (n1784, n441);
buf  g770 (n905, n402);
not  g771 (n1601, n214);
not  g772 (n857, n232);
not  g773 (n1131, n401);
not  g774 (n884, n294);
buf  g775 (n1054, n365);
buf  g776 (n1636, n287);
buf  g777 (n1717, n328);
buf  g778 (n991, n449);
not  g779 (n920, n498);
buf  g780 (n1832, n302);
not  g781 (n680, n469);
buf  g782 (n1297, n435);
not  g783 (n1436, n198);
not  g784 (n901, n452);
buf  g785 (n1688, n267);
not  g786 (n795, n337);
buf  g787 (n703, n304);
buf  g788 (n1354, n323);
not  g789 (n1304, n261);
not  g790 (n1856, n442);
not  g791 (n825, n497);
buf  g792 (n1529, n204);
not  g793 (n773, n332);
not  g794 (n1271, n218);
buf  g795 (n1479, n408);
not  g796 (n1089, n297);
buf  g797 (n985, n458);
buf  g798 (n1727, n185);
not  g799 (n671, n380);
not  g800 (n1101, n355);
not  g801 (n688, n284);
buf  g802 (n1644, n237);
buf  g803 (n1728, n348);
not  g804 (n603, n513);
buf  g805 (n1049, n266);
buf  g806 (n841, n451);
buf  g807 (n1852, n210);
not  g808 (n820, n487);
buf  g809 (n1611, n187);
buf  g810 (n1108, n215);
not  g811 (n859, n523);
buf  g812 (n1812, n523);
buf  g813 (n700, n341);
not  g814 (n1640, n454);
buf  g815 (n1323, n438);
not  g816 (n1247, n213);
not  g817 (n624, n482);
not  g818 (n942, n483);
buf  g819 (n1238, n291);
not  g820 (n1385, n219);
buf  g821 (n1000, n537);
buf  g822 (n1842, n533);
buf  g823 (n1783, n266);
not  g824 (n1158, n438);
buf  g825 (n963, n273);
not  g826 (n1491, n389);
not  g827 (n1026, n400);
buf  g828 (n1159, n357);
buf  g829 (n734, n156);
buf  g830 (n1439, n234);
buf  g831 (n1360, n229);
not  g832 (n1434, n455);
not  g833 (n1293, n378);
buf  g834 (n1219, n409);
not  g835 (n681, n201);
not  g836 (n1053, n499);
not  g837 (n746, n248);
not  g838 (n1251, n528);
buf  g839 (n1689, n270);
buf  g840 (n1590, n457);
not  g841 (n1639, n413);
not  g842 (n698, n464);
buf  g843 (n839, n272);
not  g844 (n914, n415);
not  g845 (n978, n452);
buf  g846 (n1041, n207);
buf  g847 (n1440, n247);
not  g848 (n1117, n433);
buf  g849 (n1035, n357);
not  g850 (n993, n245);
not  g851 (n865, n447);
buf  g852 (n913, n227);
buf  g853 (n1425, n358);
buf  g854 (n1206, n272);
buf  g855 (n1057, n364);
not  g856 (n1196, n155);
not  g857 (n1044, n500);
buf  g858 (n1377, n242);
not  g859 (n1844, n335);
not  g860 (n1741, n471);
not  g861 (n1779, n338);
buf  g862 (n1240, n409);
buf  g863 (n1282, n336);
buf  g864 (n627, n369);
not  g865 (n1472, n396);
not  g866 (n1432, n166);
buf  g867 (n767, n325);
not  g868 (n972, n306);
buf  g869 (n1563, n275);
buf  g870 (n1064, n261);
not  g871 (n1399, n163);
buf  g872 (n1192, n522);
buf  g873 (n804, n223);
buf  g874 (n1580, n498);
not  g875 (n1315, n291);
buf  g876 (n709, n473);
not  g877 (n1659, n319);
not  g878 (n1276, n417);
buf  g879 (n1853, n388);
not  g880 (n958, n349);
buf  g881 (n1726, n452);
not  g882 (n1515, n487);
not  g883 (n705, n312);
buf  g884 (n852, n289);
buf  g885 (n1662, n271);
buf  g886 (n821, n185);
buf  g887 (n830, n491);
buf  g888 (n1317, n466);
not  g889 (n1346, n206);
not  g890 (n1216, n292);
not  g891 (n1643, n344);
not  g892 (n1753, n160);
buf  g893 (n1801, n323);
not  g894 (n1344, n513);
buf  g895 (n1167, n316);
not  g896 (n883, n200);
buf  g897 (n843, n227);
buf  g898 (n922, n492);
buf  g899 (n1456, n215);
not  g900 (n1227, n238);
not  g901 (n1045, n351);
buf  g902 (n960, n165);
not  g903 (n1826, n480);
buf  g904 (n1693, n387);
not  g905 (n1337, n524);
not  g906 (n1663, n493);
buf  g907 (n969, n467);
buf  g908 (n994, n237);
not  g909 (n1405, n236);
not  g910 (n1604, n326);
not  g911 (n1150, n298);
buf  g912 (n1373, n273);
buf  g913 (n889, n459);
buf  g914 (n929, n210);
not  g915 (n1358, n503);
buf  g916 (n1397, n202);
buf  g917 (n1577, n514);
not  g918 (n1522, n254);
buf  g919 (n1178, n214);
not  g920 (n1626, n318);
not  g921 (n1464, n173);
buf  g922 (n601, n217);
not  g923 (n1645, n245);
buf  g924 (n1651, n419);
not  g925 (n984, n423);
buf  g926 (n1761, n456);
buf  g927 (n1093, n154);
not  g928 (n1156, n379);
not  g929 (n1191, n227);
not  g930 (n782, n397);
not  g931 (n1665, n250);
buf  g932 (n1488, n310);
not  g933 (n1283, n486);
not  g934 (n1711, n427);
not  g935 (n1618, n493);
buf  g936 (n1142, n360);
buf  g937 (n1591, n528);
not  g938 (n675, n358);
not  g939 (n823, n431);
buf  g940 (n1134, n505);
not  g941 (n761, n448);
not  g942 (n1285, n454);
buf  g943 (n590, n271);
buf  g944 (n1016, n298);
not  g945 (n1498, n325);
buf  g946 (n1593, n262);
not  g947 (n1084, n462);
not  g948 (n1258, n283);
not  g949 (n824, n522);
not  g950 (n1220, n264);
not  g951 (n1460, n437);
not  g952 (n1834, n370);
buf  g953 (n933, n494);
buf  g954 (n1313, n451);
buf  g955 (n1476, n280);
not  g956 (n1575, n242);
buf  g957 (n799, n311);
buf  g958 (n1003, n529);
not  g959 (n1830, n343);
not  g960 (n1598, n205);
not  g961 (n1389, n525);
buf  g962 (n798, n456);
buf  g963 (n1235, n276);
buf  g964 (n1303, n202);
buf  g965 (n780, n430);
buf  g966 (n1175, n207);
buf  g967 (n1650, n391);
not  g968 (n1787, n172);
not  g969 (n788, n500);
buf  g970 (n1597, n231);
not  g971 (n1748, n252);
not  g972 (n1806, n478);
not  g973 (n1200, n400);
not  g974 (n1164, n364);
buf  g975 (n1120, n427);
buf  g976 (n735, n300);
buf  g977 (n1708, n346);
buf  g978 (n794, n473);
buf  g979 (n1015, n505);
not  g980 (n626, n416);
not  g981 (n689, n518);
buf  g982 (n1660, n434);
buf  g983 (n1839, n347);
not  g984 (n1127, n238);
not  g985 (n1512, n290);
not  g986 (n1411, n209);
not  g987 (n663, n475);
buf  g988 (n776, n154);
buf  g989 (n1396, n485);
not  g990 (n954, n475);
not  g991 (n1775, n404);
buf  g992 (n1735, n538);
buf  g993 (n1287, n340);
buf  g994 (n778, n507);
buf  g995 (n732, n307);
buf  g996 (n1506, n283);
buf  g997 (n974, n419);
not  g998 (n1123, n256);
not  g999 (n1149, n445);
buf  g1000 (n702, n450);
not  g1001 (n1039, n205);
buf  g1002 (n1678, n239);
not  g1003 (n1071, n371);
not  g1004 (n622, n355);
not  g1005 (n796, n341);
buf  g1006 (n1023, n506);
not  g1007 (n944, n311);
buf  g1008 (n1530, n498);
buf  g1009 (n1500, n259);
not  g1010 (n1106, n293);
not  g1011 (n1122, n274);
buf  g1012 (n1484, n488);
not  g1013 (n965, n439);
buf  g1014 (n1228, n228);
buf  g1015 (n1459, n342);
not  g1016 (n1009, n378);
not  g1017 (n649, n241);
buf  g1018 (n1400, n295);
buf  g1019 (n658, n246);
buf  g1020 (n1091, n421);
not  g1021 (n831, n203);
buf  g1022 (n1239, n335);
not  g1023 (n757, n219);
buf  g1024 (n1420, n148);
buf  g1025 (n1413, n188);
not  g1026 (n1118, n514);
not  g1027 (n910, n487);
not  g1028 (n1571, n468);
not  g1029 (n1414, n189);
buf  g1030 (n630, n345);
buf  g1031 (n1513, n333);
buf  g1032 (n1132, n354);
buf  g1033 (n911, n356);
not  g1034 (n739, n332);
buf  g1035 (n633, n477);
buf  g1036 (n672, n373);
buf  g1037 (n1612, n418);
not  g1038 (n1615, n524);
buf  g1039 (n1817, n473);
buf  g1040 (n916, n300);
not  g1041 (n1368, n258);
not  g1042 (n1422, n521);
buf  g1043 (n1855, n267);
buf  g1044 (n1316, n509);
buf  g1045 (n1096, n258);
buf  g1046 (n1098, n324);
not  g1047 (n1332, n477);
buf  g1048 (n1286, n351);
buf  g1049 (n1557, n257);
buf  g1050 (n1827, n455);
buf  g1051 (n1301, n375);
not  g1052 (n1715, n206);
buf  g1053 (n1394, n376);
not  g1054 (n1005, n537);
buf  g1055 (n935, n247);
not  g1056 (n1578, n411);
not  g1057 (n677, n148);
buf  g1058 (n706, n508);
buf  g1059 (n1311, n182);
buf  g1060 (n1752, n464);
not  g1061 (n816, n197);
buf  g1062 (n897, n408);
buf  g1063 (n1595, n356);
not  g1064 (n892, n314);
buf  g1065 (n1350, n288);
buf  g1066 (n880, n383);
not  g1067 (n1048, n346);
buf  g1068 (n923, n304);
buf  g1069 (n961, n262);
buf  g1070 (n604, n436);
buf  g1071 (n1329, n529);
not  g1072 (n1508, n520);
not  g1073 (n691, n527);
buf  g1074 (n1374, n179);
buf  g1075 (n1416, n399);
buf  g1076 (n1161, n186);
buf  g1077 (n650, n407);
buf  g1078 (n731, n441);
not  g1079 (n879, n313);
buf  g1080 (n1443, n423);
not  g1081 (n926, n247);
buf  g1082 (n1770, n483);
not  g1083 (n1006, n221);
buf  g1084 (n1625, n275);
buf  g1085 (n1076, n512);
buf  g1086 (n1788, n310);
buf  g1087 (n1686, n540);
buf  g1088 (n1318, n365);
buf  g1089 (n1314, n488);
not  g1090 (n1296, n270);
buf  g1091 (n1514, n490);
buf  g1092 (n1468, n382);
buf  g1093 (n850, n535);
buf  g1094 (n1813, n208);
not  g1095 (n1321, n377);
not  g1096 (n1607, n311);
not  g1097 (n1260, n425);
buf  g1098 (n1060, n471);
not  g1099 (n1620, n526);
not  g1100 (n1720, n489);
not  g1101 (n1807, n253);
not  g1102 (n1362, n317);
not  g1103 (n1275, n502);
not  g1104 (n1461, n255);
not  g1105 (n1261, n307);
not  g1106 (n1387, n217);
not  g1107 (n753, n192);
not  g1108 (n1673, n523);
buf  g1109 (n1732, n235);
buf  g1110 (n1840, n422);
buf  g1111 (n611, n180);
not  g1112 (n1485, n398);
buf  g1113 (n1838, n187);
not  g1114 (n815, n276);
buf  g1115 (n1559, n320);
buf  g1116 (n1243, n504);
buf  g1117 (n1822, n183);
buf  g1118 (n1322, n380);
not  g1119 (n1777, n150);
buf  g1120 (n1366, n334);
not  g1121 (n1831, n243);
not  g1122 (n834, n280);
buf  g1123 (n743, n530);
buf  g1124 (n1204, n422);
not  g1125 (n858, n485);
buf  g1126 (n1066, n298);
not  g1127 (n623, n369);
not  g1128 (n1768, n332);
not  g1129 (n1451, n500);
not  g1130 (n1482, n429);
buf  g1131 (n1769, n327);
not  g1132 (n1630, n288);
buf  g1133 (n669, n324);
buf  g1134 (n1335, n472);
not  g1135 (n937, n478);
not  g1136 (n721, n528);
buf  g1137 (n1567, n292);
not  g1138 (n1483, n346);
buf  g1139 (n1359, n388);
buf  g1140 (n615, n484);
buf  g1141 (n1683, n207);
not  g1142 (n716, n257);
not  g1143 (n1361, n534);
buf  g1144 (n1203, n297);
buf  g1145 (n738, n375);
not  g1146 (n921, n532);
not  g1147 (n1654, n189);
not  g1148 (n1499, n401);
not  g1149 (n848, n186);
not  g1150 (n1429, n308);
not  g1151 (n592, n390);
not  g1152 (n1714, n223);
not  g1153 (n786, n393);
not  g1154 (n1767, n201);
buf  g1155 (n1020, n384);
buf  g1156 (n1656, n363);
buf  g1157 (n781, n322);
not  g1158 (n1288, n447);
buf  g1159 (n1325, n330);
not  g1160 (n837, n234);
not  g1161 (n1210, n311);
not  g1162 (n1165, n366);
buf  g1163 (n1037, n430);
buf  g1164 (n656, n159);
buf  g1165 (n1566, n151);
not  g1166 (n890, n347);
not  g1167 (n1018, n531);
buf  g1168 (n1189, n348);
not  g1169 (n1733, n457);
not  g1170 (n607, n251);
not  g1171 (n1666, n250);
buf  g1172 (n1507, n541);
buf  g1173 (n1776, n517);
not  g1174 (n1357, n190);
not  g1175 (n673, n187);
buf  g1176 (n1012, n396);
not  g1177 (n602, n384);
not  g1178 (n1351, n403);
not  g1179 (n1068, n338);
buf  g1180 (n1241, n244);
not  g1181 (n1713, n395);
buf  g1182 (n1040, n378);
not  g1183 (n1445, n467);
not  g1184 (n1772, n284);
buf  g1185 (n1176, n472);
not  g1186 (n1736, n489);
not  g1187 (n1829, n370);
buf  g1188 (n805, n344);
not  g1189 (n1367, n339);
buf  g1190 (n1782, n360);
buf  g1191 (n777, n324);
buf  g1192 (n997, n177);
buf  g1193 (n842, n432);
buf  g1194 (n1710, n319);
not  g1195 (n1462, n164);
not  g1196 (n750, n296);
not  g1197 (n810, n483);
not  g1198 (n1697, n497);
not  g1199 (n1211, n285);
not  g1200 (n1380, n187);
buf  g1201 (n696, n534);
buf  g1202 (n1143, n300);
buf  g1203 (n1737, n216);
not  g1204 (n807, n461);
buf  g1205 (n637, n285);
not  g1206 (n1130, n397);
buf  g1207 (n1430, n389);
buf  g1208 (n1799, n392);
buf  g1209 (n1551, n463);
buf  g1210 (n600, n439);
not  g1211 (n1734, n348);
not  g1212 (n967, n434);
not  g1213 (n789, n442);
buf  g1214 (n1001, n232);
not  g1215 (n1292, n249);
buf  g1216 (n1133, n215);
not  g1217 (n1616, n352);
buf  g1218 (n1682, n206);
buf  g1219 (n995, n524);
not  g1220 (n981, n277);
buf  g1221 (n1254, n448);
buf  g1222 (n1051, n303);
buf  g1223 (n670, n340);
buf  g1224 (n747, n313);
buf  g1225 (n1446, n409);
not  g1226 (n666, n433);
not  g1227 (n1568, n343);
not  g1228 (n1214, n443);
not  g1229 (n1309, n197);
not  g1230 (n1442, n478);
buf  g1231 (n941, n229);
buf  g1232 (n979, n183);
not  g1233 (n632, n226);
not  g1234 (n1407, n174);
buf  g1235 (n1221, n188);
not  g1236 (n693, n519);
not  g1237 (n1036, n530);
buf  g1238 (n1388, n331);
not  g1239 (n863, n230);
not  g1240 (n860, n440);
not  g1241 (n719, n374);
buf  g1242 (n1059, n485);
buf  g1243 (n730, n486);
buf  g1244 (n1319, n482);
not  g1245 (n774, n190);
not  g1246 (n1701, n443);
buf  g1247 (n1540, n499);
not  g1248 (n1810, n256);
buf  g1249 (n613, n181);
buf  g1250 (n1441, n321);
buf  g1251 (n740, n429);
buf  g1252 (n930, n345);
not  g1253 (n876, n344);
not  g1254 (n779, n167);
not  g1255 (n1215, n421);
not  g1256 (n996, n235);
buf  g1257 (n608, n186);
not  g1258 (n1740, n304);
buf  g1259 (n1670, n496);
not  g1260 (n1103, n386);
buf  g1261 (n1119, n246);
not  g1262 (n605, n415);
buf  g1263 (n1415, n284);
not  g1264 (n665, n392);
not  g1265 (n713, n280);
buf  g1266 (n1208, n350);
buf  g1267 (n797, n352);
buf  g1268 (n980, n224);
buf  g1269 (n887, n349);
buf  g1270 (n1789, n416);
buf  g1271 (n886, n526);
not  g1272 (n1613, n283);
not  g1273 (n711, n322);
not  g1274 (n1347, n490);
buf  g1275 (n1538, n381);
buf  g1276 (n1547, n437);
not  g1277 (n872, n458);
buf  g1278 (n1237, n484);
not  g1279 (n1569, n302);
not  g1280 (n695, n385);
buf  g1281 (n1531, n180);
buf  g1282 (n1721, n153);
not  g1283 (n1356, n386);
not  g1284 (n1138, n275);
not  g1285 (n1641, n306);
buf  g1286 (n639, n515);
not  g1287 (n646, n199);
not  g1288 (n1774, n350);
not  g1289 (n1274, n479);
buf  g1290 (n1075, n196);
buf  g1291 (n1707, n476);
buf  g1292 (n1341, n164);
buf  g1293 (n1505, n359);
not  g1294 (n1109, n245);
not  g1295 (n1188, n260);
buf  g1296 (n1764, n221);
buf  g1297 (n1841, n388);
not  g1298 (n950, n242);
not  g1299 (n1421, n157);
buf  g1300 (n1600, n454);
not  g1301 (n1438, n223);
buf  g1302 (n1193, n313);
not  g1303 (n1008, n468);
buf  g1304 (n1747, n369);
not  g1305 (n1082, n336);
not  g1306 (n1253, n344);
buf  g1307 (n1145, n408);
buf  g1308 (n1352, n250);
not  g1309 (n948, n499);
buf  g1310 (n1259, n287);
not  g1311 (n1264, n387);
not  g1312 (n1589, n254);
not  g1313 (n599, n401);
buf  g1314 (n1063, n433);
not  g1315 (n631, n329);
not  g1316 (n1128, n481);
buf  g1317 (n1371, n423);
not  g1318 (n1846, n424);
not  g1319 (n727, n465);
not  g1320 (n1092, n285);
buf  g1321 (n1107, n428);
not  g1322 (n1751, n405);
not  g1323 (n1564, n509);
not  g1324 (n662, n193);
buf  g1325 (n655, n314);
buf  g1326 (n867, n438);
not  g1327 (n827, n234);
not  g1328 (n610, n277);
not  g1329 (n1073, n271);
not  g1330 (n1676, n424);
not  g1331 (n813, n435);
buf  g1332 (n1234, n345);
not  g1333 (n667, n247);
not  g1334 (n1617, n291);
buf  g1335 (n1700, n495);
not  g1336 (n1386, n420);
buf  g1337 (n661, n181);
not  g1338 (n894, n233);
not  g1339 (n1331, n204);
buf  g1340 (n616, n493);
not  g1341 (n1757, n225);
not  g1342 (n1624, n432);
buf  g1343 (n1148, n395);
not  g1344 (n925, n391);
buf  g1345 (n882, n505);
buf  g1346 (n1121, n176);
buf  g1347 (n687, n482);
buf  g1348 (n1263, n507);
buf  g1349 (n1684, n210);
not  g1350 (n1171, n261);
not  g1351 (n1129, n350);
not  g1352 (n1105, n279);
not  g1353 (n1187, n466);
not  g1354 (n934, n171);
buf  g1355 (n1526, n275);
buf  g1356 (n718, n497);
not  g1357 (n1299, n474);
not  g1358 (n1278, n281);
buf  g1359 (n1739, n517);
not  g1360 (n1450, n282);
buf  g1361 (n1849, n253);
buf  g1362 (n811, n305);
not  g1363 (n1652, n189);
not  g1364 (n1543, n200);
not  g1365 (n829, n297);
buf  g1366 (n635, n156);
not  g1367 (n1687, n426);
buf  g1368 (n1449, n149);
not  g1369 (n1542, n371);
not  g1370 (n676, n385);
not  g1371 (n1742, n188);
buf  g1372 (n1570, n240);
not  g1373 (n733, n277);
buf  g1374 (n1242, n526);
buf  g1375 (n1648, n529);
buf  g1376 (n1029, n206);
buf  g1377 (n1019, n386);
buf  g1378 (n802, n165);
not  g1379 (n1222, n437);
not  g1380 (n1349, n481);
buf  g1381 (n1289, n338);
buf  g1382 (n1664, n536);
not  g1383 (n645, n169);
buf  g1384 (n1345, n437);
not  g1385 (n1410, n228);
not  g1386 (n1370, n458);
buf  g1387 (n1065, n449);
buf  g1388 (n908, n321);
not  g1389 (n800, n419);
buf  g1390 (n652, n219);
buf  g1391 (n1270, n530);
not  g1392 (n1115, n412);
buf  g1393 (n756, n384);
not  g1394 (n1229, n243);
not  g1395 (n729, n273);
buf  g1396 (n1268, n276);
not  g1397 (n717, n181);
not  g1398 (n1110, n400);
not  g1399 (n917, n178);
not  g1400 (n1520, n459);
not  g1401 (n755, n223);
not  g1402 (n1062, n424);
buf  g1403 (n1290, n278);
not  g1404 (n1205, n511);
buf  g1405 (n1355, n176);
buf  g1406 (n1716, n399);
not  g1407 (n1759, n414);
not  g1408 (n1404, n310);
not  g1409 (n1490, n483);
not  g1410 (n1011, n230);
not  g1411 (n1250, n460);
not  g1412 (n686, n520);
buf  g1413 (n1294, n490);
not  g1414 (n642, n231);
not  g1415 (n1081, n537);
buf  g1416 (n1230, n286);
buf  g1417 (n947, n540);
buf  g1418 (n606, n282);
buf  g1419 (n1527, n433);
not  g1420 (n1454, n296);
not  g1421 (n1489, n347);
buf  g1422 (n982, n506);
buf  g1423 (n1030, n446);
not  g1424 (n1136, n410);
buf  g1425 (n1760, n286);
not  g1426 (n1843, n241);
not  g1427 (n1378, n336);
not  g1428 (n1457, n215);
not  g1429 (n861, n242);
buf  g1430 (n1545, n465);
not  g1431 (n1592, n420);
not  g1432 (n1437, n320);
not  g1433 (n1552, n468);
buf  g1434 (n1463, n521);
not  g1435 (n597, n228);
buf  g1436 (n1685, n425);
buf  g1437 (n1816, n518);
not  g1438 (n1854, n300);
buf  g1439 (n828, n270);
buf  g1440 (n968, n212);
buf  g1441 (n1339, n539);
buf  g1442 (n1155, n208);
not  g1443 (n1072, n212);
buf  g1444 (n682, n436);
not  g1445 (n957, n204);
not  g1446 (n1383, n277);
buf  g1447 (n758, n178);
buf  g1448 (n742, n521);
not  g1449 (n1375, n504);
buf  g1450 (n836, n184);
not  g1451 (n769, n284);
buf  g1452 (n1042, n257);
buf  g1453 (n1116, n182);
not  g1454 (n668, n278);
buf  g1455 (n1070, n367);
not  g1456 (n1032, n254);
not  g1457 (n1695, n251);
not  g1458 (n1680, n308);
not  g1459 (n1047, n330);
buf  g1460 (n874, n444);
buf  g1461 (n1343, n269);
not  g1462 (n1517, n444);
buf  g1463 (n1447, n519);
buf  g1464 (n1280, n322);
buf  g1465 (n1384, n146);
not  g1466 (n1574, n190);
buf  g1467 (n1424, n404);
not  g1468 (n1539, n358);
buf  g1469 (n1034, n408);
not  g1470 (n1602, n281);
not  g1471 (n1667, n222);
not  g1472 (n970, n365);
not  g1473 (n1310, n307);
buf  g1474 (n1305, n337);
buf  g1475 (n1587, n268);
not  g1476 (n1342, n272);
buf  g1477 (n1623, n394);
not  g1478 (n1756, n326);
not  g1479 (n748, n535);
buf  g1480 (n909, n212);
buf  g1481 (n1835, n315);
buf  g1482 (n1668, n395);
buf  g1483 (n1702, n320);
not  g1484 (n1745, n464);
buf  g1485 (n1474, n270);
not  g1486 (n1112, n373);
not  g1487 (n1174, n372);
not  g1488 (n851, n248);
not  g1489 (n1694, n508);
not  g1490 (n1273, n462);
not  g1491 (n1581, n315);
not  g1492 (n737, n374);
buf  g1493 (n1444, n425);
not  g1494 (n664, n501);
not  g1495 (n1002, n299);
not  g1496 (n710, n472);
buf  g1497 (n1521, n466);
not  g1498 (n1548, n296);
not  g1499 (n1691, n340);
not  g1500 (n868, n210);
not  g1501 (n1692, n366);
buf  g1502 (n683, n457);
not  g1503 (n924, n501);
buf  g1504 (n1074, n356);
buf  g1505 (n1681, n286);
buf  g1506 (n1477, n375);
buf  g1507 (n1642, n501);
not  g1508 (n1487, n455);
not  g1509 (n846, n383);
buf  g1510 (n1376, n280);
not  g1511 (n1819, n426);
not  g1512 (n1435, n534);
not  g1513 (n1811, n252);
not  g1514 (n593, n292);
not  g1515 (n1565, n265);
buf  g1516 (n1043, n290);
not  g1517 (n625, n480);
not  g1518 (n1773, n303);
not  g1519 (n1194, n150);
not  g1520 (n1847, n225);
not  g1521 (n618, n305);
not  g1522 (n1392, n235);
not  g1523 (n1537, n539);
not  g1524 (n612, n475);
not  g1525 (n766, n219);
buf  g1526 (n1528, n370);
not  g1527 (n1124, n492);
not  g1528 (n1139, n355);
not  g1529 (n904, n523);
not  g1530 (n1808, n414);
buf  g1531 (n1028, n539);
not  g1532 (n1185, n245);
not  g1533 (n1698, n354);
not  g1534 (n1069, n166);
not  g1535 (n1393, n263);
not  g1536 (n1199, n512);
not  g1537 (n728, n184);
buf  g1538 (n617, n192);
buf  g1539 (n699, n158);
buf  g1540 (n1610, n486);
buf  g1541 (n1469, n417);
not  g1542 (n854, n236);
buf  g1543 (n784, n260);
buf  g1544 (n1509, n533);
not  g1545 (n763, n518);
not  g1546 (n1330, n360);
buf  g1547 (n1390, n339);
not  g1548 (n653, n373);
not  g1549 (n1586, n309);
buf  g1550 (n881, n228);
buf  g1551 (n1061, n318);
buf  g1552 (n651, n507);
buf  g1553 (n1402, n367);
buf  g1554 (n1147, n287);
not  g1555 (n1125, n168);
buf  g1556 (n1797, n382);
buf  g1557 (n1699, n463);
not  g1558 (n1284, n389);
not  g1559 (n893, n195);
buf  g1560 (n1556, n468);
buf  g1561 (n629, n194);
buf  g1562 (n855, n295);
not  g1563 (n1372, n269);
buf  g1564 (n1307, n315);
not  g1565 (n1281, n527);
not  g1566 (n1269, n204);
buf  g1567 (n1814, n478);
not  g1568 (n1825, n532);
buf  g1569 (n1850, n145);
buf  g1570 (n1661, n218);
not  g1571 (n1417, n477);
not  g1572 (n1455, n211);
not  g1573 (n870, n299);
buf  g1574 (n1226, n479);
not  g1575 (n1674, n525);
buf  g1576 (n692, n526);
buf  g1577 (n644, n194);
buf  g1578 (n1027, n353);
buf  g1579 (n1510, n174);
buf  g1580 (n1262, n400);
not  g1581 (n1511, n392);
not  g1582 (n906, n265);
not  g1583 (n1743, n306);
not  g1584 (n598, n340);
buf  g1585 (n1763, n446);
buf  g1586 (n1141, n227);
not  g1587 (n840, n282);
not  g1588 (n1179, n381);
not  g1589 (n647, n404);
not  g1590 (n1426, n175);
buf  g1591 (n1677, n385);
buf  g1592 (n1709, n494);
not  g1593 (n814, n447);
not  g1594 (n1828, n205);
buf  g1595 (n1762, n524);
not  g1596 (n1152, n203);
not  g1597 (n998, n492);
not  g1598 (n946, n268);
not  g1599 (n835, n402);
buf  g1600 (n1749, n361);
buf  g1601 (n1793, n244);
not  g1602 (n685, n168);
buf  g1603 (n1647, n200);
not  g1604 (n764, n250);
buf  g1605 (n1153, n312);
buf  g1606 (n1504, n385);
not  g1607 (n1007, n324);
buf  g1608 (n1170, n391);
not  g1609 (n918, n211);
not  g1610 (n1750, n465);
buf  g1611 (n1723, n193);
buf  g1612 (n704, n372);
buf  g1613 (n1207, n401);
not  g1614 (n959, n252);
buf  g1615 (n1249, n312);
not  g1616 (n949, n376);
buf  g1617 (n1785, n488);
not  g1618 (n1614, n266);
not  g1619 (n1765, n253);
not  g1620 (n1427, n221);
buf  g1621 (n1582, n342);
not  g1622 (n1818, n484);
not  g1623 (n1794, n395);
buf  g1624 (n1298, n380);
not  g1625 (n1758, n268);
buf  g1626 (n1795, n379);
not  g1627 (n1824, n314);
buf  g1628 (n943, n393);
not  g1629 (n595, n319);
buf  g1630 (n1144, n410);
buf  g1631 (n1501, n256);
not  g1632 (n1087, n321);
not  g1633 (n1295, n183);
not  g1634 (n990, n263);
buf  g1635 (n643, n335);
not  g1636 (n977, n439);
not  g1637 (n641, n249);
not  g1638 (n1050, n518);
not  g1639 (n744, n429);
buf  g1640 (n1746, n316);
buf  g1641 (n1798, n244);
not  g1642 (n1820, n378);
not  g1643 (n1364, n369);
not  g1644 (n845, n399);
buf  g1645 (n1836, n502);
buf  g1646 (n1619, n162);
not  g1647 (n1014, n500);
buf  g1648 (n1363, n508);
not  g1649 (n1010, n230);
buf  g1650 (n1225, n182);
not  g1651 (n1398, n233);
buf  g1652 (n1628, n387);
buf  g1653 (n1755, n197);
not  g1654 (n871, n444);
buf  g1655 (n896, n226);
not  g1656 (n726, n496);
not  g1657 (n638, n248);
buf  g1658 (n1494, n515);
buf  g1659 (n1172, n256);
buf  g1660 (n1277, n451);
buf  g1661 (n1365, n225);
not  g1662 (n1097, n470);
buf  g1663 (n701, n439);
not  g1664 (n1162, n213);
buf  g1665 (n1111, n173);
buf  g1666 (n1408, n197);
buf  g1667 (n1140, n447);
not  g1668 (n939, n470);
buf  g1669 (n986, n342);
not  g1670 (n1470, n360);
buf  g1671 (n1804, n471);
not  g1672 (n1168, n179);
not  g1673 (n1535, n536);
buf  g1674 (n722, n272);
not  g1675 (n1245, n217);
not  g1676 (n1266, n229);
not  g1677 (n1802, n377);
not  g1678 (n1324, n176);
buf  g1679 (n953, n274);
buf  g1680 (n1233, n331);
not  g1681 (n936, n460);
buf  g1682 (n907, n475);
buf  g1683 (n1516, n390);
not  g1684 (n1583, n510);
buf  g1685 (n1465, n413);
not  g1686 (n1052, n445);
buf  g1687 (n919, n515);
not  g1688 (n1725, n301);
buf  g1689 (n1163, n220);
buf  g1690 (n952, n368);
not  g1691 (n1257, n507);
buf  g1692 (n1627, n230);
not  g1693 (n1800, n348);
buf  g1694 (n877, n188);
buf  g1695 (n1669, n254);
not  g1696 (n1486, n308);
buf  g1697 (n1594, n322);
buf  g1698 (n975, n185);
not  g1699 (n1173, n237);
buf  g1700 (n1533, n407);
buf  g1701 (n628, n499);
not  g1702 (n1495, n222);
buf  g1703 (n915, n209);
buf  g1704 (n1154, n462);
not  g1705 (n1845, n199);
not  g1706 (n1197, n491);
buf  g1707 (n1403, n289);
buf  g1708 (n1244, n185);
not  g1709 (n1326, n182);
buf  g1710 (n751, n318);
buf  g1711 (n1579, n357);
not  g1712 (n888, n191);
buf  g1713 (n1655, n268);
not  g1714 (n1712, n325);
not  g1715 (n1705, n251);
buf  g1716 (n1085, n404);
not  g1717 (n1722, n531);
buf  g1718 (n1428, n177);
buf  g1719 (n1635, n328);
buf  g1720 (n1201, n450);
not  g1721 (n1099, n470);
not  g1722 (n1302, n519);
buf  g1723 (n955, n481);
not  g1724 (n1790, n305);
not  g1725 (n1209, n162);
not  g1726 (n1453, n487);
not  g1727 (n765, n403);
buf  g1728 (n900, n327);
buf  g1729 (n1467, n407);
not  g1730 (n708, n208);
buf  g1731 (n791, n202);
buf  g1732 (n1744, n412);
not  g1733 (n1719, n203);
buf  g1734 (n938, n147);
buf  g1735 (n1202, n328);
buf  g1736 (n928, n287);
and  g1737 (n1017, n241, n442, n149, n402);
xnor g1738 (n1524, n361, n480, n374, n190);
or   g1739 (n770, n411, n527, n406, n353);
nand g1740 (n1409, n394, n179, n418, n409);
or   g1741 (n1256, n391, n317, n195, n175);
and  g1742 (n808, n386, n198, n420, n170);
xnor g1743 (n1431, n246, n359, n366, n481);
nand g1744 (n745, n414, n372, n201, n233);
nor  g1745 (n720, n482, n349, n491, n323);
nor  g1746 (n596, n364, n290, n417, n456);
nand g1747 (n1077, n177, n298, n201, n488);
xor  g1748 (n1055, n157, n531, n509, n249);
or   g1749 (n1180, n450, n504, n514, n445);
xnor g1750 (n684, n459, n356, n260, n382);
xor  g1751 (n1382, n259, n236, n186, n371);
nand g1752 (n838, n454, n160, n453, n525);
xnor g1753 (n772, n334, n511, n452, n530);
xnor g1754 (n660, n302, n502, n377, n494);
nand g1755 (n1169, n423, n216, n516, n535);
nand g1756 (n1279, n155, n218, n341, n312);
and  g1757 (n1452, n320, n161, n432, n419);
xor  g1758 (n760, n436, n241, n399, n191);
nor  g1759 (n1336, n240, n267, n326);
and  g1760 (n819, n195, n393, n519, n259);
xor  g1761 (n1177, n353, n491, n195, n161);
nor  g1762 (n754, n235, n226, n327, n158);
xor  g1763 (n1851, n253, n218, n370, n207);
and  g1764 (n1067, n327, n501, n376, n520);
and  g1765 (n1546, n259, n492, n352, n496);
xor  g1766 (n1631, n411, n238, n397, n265);
xor  g1767 (n1519, n368, n421, n442, n281);
xor  g1768 (n771, n476, n359, n516, n221);
nor  g1769 (n826, n317, n389, n522, n290);
xnor g1770 (n1848, n517, n413, n539, n390);
or   g1771 (n885, n412, n152, n373, n278);
nand g1772 (n674, n416, n279, n293, n330);
and  g1773 (n902, n178, n305, n461, n403);
or   g1774 (n1576, n540, n361, n520, n403);
nor  g1775 (n847, n205, n301, n200, n368);
xor  g1776 (n1653, n438, n301, n238, n412);
xor  g1777 (n1300, n274, n414, n339, n479);
xnor g1778 (n1391, n199, n294, n226, n209);
nand g1779 (n620, n521, n428, n489, n345);
xnor g1780 (n1475, n374, n533, n503, n330);
xnor g1781 (n1046, n446, n294, n362, n304);
nor  g1782 (n762, n467, n513, n333, n366);
nand g1783 (n1088, n351, n152, n281, n466);
nor  g1784 (n723, n527, n237, n262, n528);
xor  g1785 (n678, n175, n318, n352, n383);
nand g1786 (n785, n263, n489, n279, n503);
nand g1787 (n1181, n474, n462, n392, n476);
xnor g1788 (n1308, n199, n338, n418, n297);
xor  g1789 (n591, n213, n367, n517, n435);
and  g1790 (n1224, n380, n196, n460, n276);
and  g1791 (n983, n476, n428, n477, n293);
nor  g1792 (n869, n331, n208, n172, n288);
nor  g1793 (n1638, n427, n529, n390, n189);
nor  g1794 (n1634, n484, n398, n296, n293);
nand g1795 (n1395, n444, n243, n379, n431);
nor  g1796 (n1186, n282, n376, n502, n295);
nor  g1797 (n1796, n274, n516, n368, n239);
xor  g1798 (n1554, n216, n512, n336, n346);
and  g1799 (n1549, n343, n232, n534, n243);
nor  g1800 (n1532, n415, n244, n405, n441);
xor  g1801 (n1496, n191, n432, n407, n192);
or   g1802 (n1333, n171, n194, n421, n536);
xnor g1803 (n694, n174, n222, n427, n331);
nor  g1804 (n1541, n279, n536, n493, n411);
nand g1805 (n1024, n234, n513, n326, n334);
nand g1806 (n621, n317, n212, n315, n308);
nor  g1807 (n1599, n511, n351, n384, n264);
xnor g1808 (n1102, n460, n458, n461, n416);
xor  g1809 (n1560, n455, n273, n288, n271);
or   g1810 (n971, n486, n445, n180, n147);
xnor g1811 (n1603, n362, n196, n540);
nor  g1812 (n1534, n522, n193, n443, n236);
xnor g1813 (n1248, n471, n329, n350, n430);
xnor g1814 (n783, n435, n184, n495, n145);
nand g1815 (n912, n299, n224, n209, n329);
or   g1816 (n1025, n364, n532, n446, n429);
xor  g1817 (n806, n398, n428, n377, n505);
xor  g1818 (n1058, n269, n286, n347, n533);
and  g1819 (n809, n469, n211, n362, n449);
nand g1820 (n1369, n169, n341, n224, n309);
nand g1821 (n1320, n495, n461, n480, n422);
nor  g1822 (n1657, n508, n255, n192, n512);
xor  g1823 (n1252, n339, n525, n387, n406);
not  g1824 (n2453, n912);
buf  g1825 (n1971, n1018);
buf  g1826 (n1915, n1626);
not  g1827 (n2307, n1164);
not  g1828 (n2115, n830);
buf  g1829 (n1967, n1075);
buf  g1830 (n2528, n1099);
not  g1831 (n1953, n1325);
not  g1832 (n2147, n792);
buf  g1833 (n1885, n1137);
buf  g1834 (n2174, n1551);
buf  g1835 (n2372, n743);
not  g1836 (n2095, n707);
buf  g1837 (n2218, n1565);
buf  g1838 (n2075, n1040);
not  g1839 (n2488, n1783);
not  g1840 (n2362, n1433);
buf  g1841 (n2469, n1665);
buf  g1842 (n1931, n941);
not  g1843 (n2149, n1733);
buf  g1844 (n2378, n756);
buf  g1845 (n2398, n1166);
not  g1846 (n2525, n1658);
not  g1847 (n2256, n883);
not  g1848 (n2046, n1214);
buf  g1849 (n2102, n1742);
buf  g1850 (n2294, n1158);
not  g1851 (n2053, n1464);
not  g1852 (n1927, n703);
buf  g1853 (n2047, n949);
buf  g1854 (n1928, n1380);
buf  g1855 (n2289, n1208);
not  g1856 (n2042, n921);
buf  g1857 (n1921, n881);
not  g1858 (n2076, n1429);
not  g1859 (n2198, n1476);
buf  g1860 (n2080, n1055);
not  g1861 (n2264, n812);
buf  g1862 (n2157, n801);
not  g1863 (n2441, n602);
buf  g1864 (n2404, n1178);
buf  g1865 (n2356, n1535);
not  g1866 (n2322, n1458);
buf  g1867 (n1952, n1531);
not  g1868 (n2317, n1226);
buf  g1869 (n2261, n718);
not  g1870 (n2146, n992);
buf  g1871 (n2339, n934);
not  g1872 (n2189, n1510);
not  g1873 (n2195, n956);
buf  g1874 (n2048, n1124);
buf  g1875 (n1973, n802);
buf  g1876 (n2170, n837);
buf  g1877 (n2492, n1582);
buf  g1878 (n1887, n1334);
buf  g1879 (n1898, n943);
buf  g1880 (n1934, n784);
buf  g1881 (n2277, n1797);
buf  g1882 (n2260, n1109);
buf  g1883 (n2502, n1631);
not  g1884 (n2238, n742);
buf  g1885 (n2055, n1475);
buf  g1886 (n1864, n1067);
buf  g1887 (n1869, n1484);
buf  g1888 (n2460, n854);
not  g1889 (n2024, n1022);
not  g1890 (n2282, n1690);
not  g1891 (n2463, n1161);
not  g1892 (n2414, n1561);
buf  g1893 (n2323, n1576);
buf  g1894 (n2171, n1533);
not  g1895 (n1970, n1388);
buf  g1896 (n2517, n1281);
buf  g1897 (n1888, n1257);
not  g1898 (n2311, n968);
buf  g1899 (n2522, n840);
not  g1900 (n1951, n1255);
not  g1901 (n2365, n1515);
not  g1902 (n2501, n1599);
buf  g1903 (n2001, n637);
buf  g1904 (n2196, n1605);
not  g1905 (n2192, n1627);
buf  g1906 (n2337, n795);
not  g1907 (n2380, n890);
not  g1908 (n1922, n1229);
not  g1909 (n1935, n872);
buf  g1910 (n2293, n1785);
buf  g1911 (n1948, n710);
not  g1912 (n2375, n1236);
buf  g1913 (n2406, n829);
buf  g1914 (n2142, n1344);
buf  g1915 (n2445, n744);
buf  g1916 (n2202, n1298);
not  g1917 (n2319, n925);
not  g1918 (n2205, n1125);
buf  g1919 (n2034, n1491);
buf  g1920 (n2318, n1691);
not  g1921 (n2310, n665);
buf  g1922 (n2231, n1374);
not  g1923 (n2420, n1736);
buf  g1924 (n2344, n951);
not  g1925 (n2506, n1655);
not  g1926 (n2464, n804);
not  g1927 (n2246, n1332);
buf  g1928 (n2043, n1778);
not  g1929 (n1914, n601);
not  g1930 (n2083, n936);
buf  g1931 (n2411, n1328);
buf  g1932 (n1996, n1267);
buf  g1933 (n1978, n1288);
buf  g1934 (n2104, n633);
buf  g1935 (n2345, n781);
buf  g1936 (n2148, n1552);
buf  g1937 (n2430, n1646);
buf  g1938 (n1926, n1722);
not  g1939 (n2392, n1301);
not  g1940 (n1897, n1580);
not  g1941 (n2094, n1549);
buf  g1942 (n2278, n858);
not  g1943 (n2128, n1472);
not  g1944 (n2340, n984);
not  g1945 (n2477, n961);
not  g1946 (n1865, n617);
buf  g1947 (n2520, n1442);
not  g1948 (n1959, n1280);
not  g1949 (n2435, n1718);
buf  g1950 (n2402, n1148);
not  g1951 (n2233, n708);
buf  g1952 (n1943, n1441);
buf  g1953 (n2090, n1139);
buf  g1954 (n2049, n928);
not  g1955 (n1920, n1727);
buf  g1956 (n2050, n679);
buf  g1957 (n2390, n977);
not  g1958 (n1916, n1575);
not  g1959 (n2212, n1322);
not  g1960 (n2440, n698);
not  g1961 (n2352, n1773);
buf  g1962 (n2133, n958);
not  g1963 (n2291, n1260);
not  g1964 (n2255, n1685);
buf  g1965 (n2244, n1493);
buf  g1966 (n1939, n1412);
buf  g1967 (n2391, n1543);
not  g1968 (n1861, n999);
not  g1969 (n2388, n729);
not  g1970 (n2286, n869);
not  g1971 (n2129, n1292);
buf  g1972 (n2208, n726);
not  g1973 (n2423, n1031);
not  g1974 (n2326, n1225);
buf  g1975 (n2251, n1324);
not  g1976 (n2155, n1248);
not  g1977 (n2029, n1023);
not  g1978 (n2138, n1370);
not  g1979 (n2107, n1251);
not  g1980 (n2037, n974);
buf  g1981 (n2065, n1024);
not  g1982 (n2331, n663);
not  g1983 (n2348, n931);
not  g1984 (n2439, n1348);
not  g1985 (n2203, n1762);
buf  g1986 (n2434, n1613);
not  g1987 (n2280, n1788);
buf  g1988 (n2006, n1306);
not  g1989 (n2227, n730);
not  g1990 (n2499, n774);
buf  g1991 (n1902, n866);
buf  g1992 (n2503, n782);
buf  g1993 (n1969, n1056);
not  g1994 (n2101, n1559);
buf  g1995 (n1965, n1309);
buf  g1996 (n2395, n1047);
not  g1997 (n2067, n1469);
buf  g1998 (n2369, n1446);
buf  g1999 (n2041, n1769);
not  g2000 (n1945, n1058);
buf  g2001 (n2105, n1327);
buf  g2002 (n1983, n1110);
not  g2003 (n2284, n759);
not  g2004 (n2346, n805);
buf  g2005 (n2073, n1457);
not  g2006 (n2304, n1030);
not  g2007 (n2514, n695);
not  g2008 (n2334, n1035);
not  g2009 (n2033, n1323);
buf  g2010 (n1932, n1761);
buf  g2011 (n2064, n1385);
buf  g2012 (n2308, n880);
not  g2013 (n2184, n794);
buf  g2014 (n2481, n1584);
buf  g2015 (n2089, n1610);
buf  g2016 (n1966, n739);
buf  g2017 (n2495, n1331);
not  g2018 (n1880, n966);
not  g2019 (n2511, n666);
not  g2020 (n2461, n1459);
not  g2021 (n2475, n902);
not  g2022 (n2131, n979);
buf  g2023 (n1947, n1617);
not  g2024 (n2152, n1714);
buf  g2025 (n2275, n1772);
buf  g2026 (n1918, n1573);
buf  g2027 (n2266, n1692);
buf  g2028 (n2421, n1059);
buf  g2029 (n2119, n1359);
buf  g2030 (n2169, n639);
buf  g2031 (n1950, n1500);
not  g2032 (n2446, n1244);
not  g2033 (n1879, n844);
not  g2034 (n2122, n990);
not  g2035 (n2281, n1767);
not  g2036 (n2168, n857);
buf  g2037 (n1929, n1707);
buf  g2038 (n2215, n1622);
buf  g2039 (n2058, n1735);
not  g2040 (n2342, n646);
not  g2041 (n2164, n605);
buf  g2042 (n2178, n1141);
not  g2043 (n1982, n910);
not  g2044 (n2267, n1273);
not  g2045 (n2336, n945);
not  g2046 (n2213, n1065);
not  g2047 (n2110, n1593);
buf  g2048 (n2400, n1641);
buf  g2049 (n2527, n1709);
buf  g2050 (n2015, n752);
buf  g2051 (n2002, n1317);
not  g2052 (n2222, n1302);
not  g2053 (n1911, n1032);
buf  g2054 (n1899, n1140);
not  g2055 (n2248, n1524);
buf  g2056 (n2470, n714);
buf  g2057 (n2262, n1223);
not  g2058 (n2523, n662);
buf  g2059 (n2223, n1405);
buf  g2060 (n2444, n915);
buf  g2061 (n2276, n621);
buf  g2062 (n2497, n705);
not  g2063 (n2139, n1016);
not  g2064 (n1938, n1759);
buf  g2065 (n2194, n1453);
buf  g2066 (n2399, n1277);
not  g2067 (n2478, n1061);
buf  g2068 (n1933, n1624);
not  g2069 (n2004, n1176);
buf  g2070 (n2023, n1497);
buf  g2071 (n1913, n1540);
not  g2072 (n2210, n959);
not  g2073 (n2166, n1054);
not  g2074 (n2158, n1670);
buf  g2075 (n1886, n1303);
not  g2076 (n2145, n1136);
buf  g2077 (n1930, n1057);
not  g2078 (n2224, n1452);
not  g2079 (n2088, n957);
not  g2080 (n2360, n594);
buf  g2081 (n2379, n1195);
buf  g2082 (n2341, n1642);
buf  g2083 (n2332, n1572);
not  g2084 (n2020, n1528);
not  g2085 (n2124, n723);
not  g2086 (n1906, n1525);
buf  g2087 (n2078, n1111);
buf  g2088 (n2269, n1606);
buf  g2089 (n2407, n1700);
not  g2090 (n2134, n894);
not  g2091 (n2112, n725);
buf  g2092 (n2381, n997);
buf  g2093 (n2253, n1723);
not  g2094 (n2199, n1364);
not  g2095 (n1997, n1038);
buf  g2096 (n2374, n711);
buf  g2097 (n2237, n942);
not  g2098 (n2144, n1211);
not  g2099 (n2358, n1747);
buf  g2100 (n2393, n1498);
buf  g2101 (n1995, n773);
buf  g2102 (n2303, n879);
buf  g2103 (n1993, n614);
buf  g2104 (n2486, n640);
buf  g2105 (n2016, n971);
buf  g2106 (n2132, n914);
not  g2107 (n2413, n724);
not  g2108 (n2193, n1034);
not  g2109 (n2455, n692);
not  g2110 (n2117, n1413);
not  g2111 (n2361, n810);
buf  g2112 (n1988, n803);
not  g2113 (n2257, n1679);
buf  g2114 (n2250, n1548);
buf  g2115 (n2239, n1463);
buf  g2116 (n2000, n1553);
buf  g2117 (n2180, n680);
buf  g2118 (n1984, n1122);
not  g2119 (n2396, n1644);
not  g2120 (n2507, n751);
buf  g2121 (n2359, n1435);
buf  g2122 (n2485, n1731);
not  g2123 (n1859, n793);
buf  g2124 (n2505, n1329);
not  g2125 (n2035, n1686);
not  g2126 (n2526, n906);
buf  g2127 (n2200, n1417);
buf  g2128 (n2209, n1340);
not  g2129 (n2312, n1155);
buf  g2130 (n1877, n1170);
not  g2131 (n2496, n838);
buf  g2132 (n1912, n1297);
not  g2133 (n2135, n1518);
not  g2134 (n1923, n1777);
buf  g2135 (n2099, n1085);
not  g2136 (n2241, n649);
not  g2137 (n2301, n1635);
not  g2138 (n2187, n892);
buf  g2139 (n2121, n888);
buf  g2140 (n1944, n1650);
buf  g2141 (n2462, n1365);
not  g2142 (n2274, n1204);
not  g2143 (n2040, n1760);
buf  g2144 (n2295, n1455);
buf  g2145 (n2007, n1082);
buf  g2146 (n2141, n1748);
not  g2147 (n1874, n1104);
buf  g2148 (n2039, n1647);
not  g2149 (n1925, n1490);
buf  g2150 (n2298, n1768);
not  g2151 (n2217, n1290);
not  g2152 (n2125, n1048);
buf  g2153 (n2529, n1120);
buf  g2154 (n1889, n1051);
not  g2155 (n1960, n1020);
buf  g2156 (n2242, n988);
not  g2157 (n2057, n1437);
buf  g2158 (n2324, n1710);
not  g2159 (n1868, n1357);
not  g2160 (n2181, n1604);
not  g2161 (n1871, n1237);
buf  g2162 (n1873, n731);
buf  g2163 (n2425, n1049);
not  g2164 (n2354, n1544);
not  g2165 (n2185, n1265);
not  g2166 (n1999, n918);
not  g2167 (n2188, n1132);
not  g2168 (n2401, n1218);
buf  g2169 (n2493, n1378);
not  g2170 (n2343, n632);
buf  g2171 (n2422, n1716);
buf  g2172 (n2367, n1473);
buf  g2173 (n2302, n1434);
not  g2174 (n2162, n1494);
buf  g2175 (n2447, n1060);
buf  g2176 (n2510, n1074);
buf  g2177 (n2027, n758);
buf  g2178 (n2418, n1330);
buf  g2179 (n2220, n1555);
buf  g2180 (n2032, n1001);
buf  g2181 (n2172, n1293);
not  g2182 (n1909, n1400);
not  g2183 (n2191, n1520);
not  g2184 (n2518, n1315);
buf  g2185 (n2426, n1172);
buf  g2186 (n2509, n653);
not  g2187 (n2448, n1162);
buf  g2188 (n1882, n1191);
buf  g2189 (n1892, n1144);
buf  g2190 (n2069, n764);
buf  g2191 (n2387, n1426);
not  g2192 (n2490, n1103);
buf  g2193 (n1900, n980);
not  g2194 (n2442, n789);
buf  g2195 (n2056, n668);
buf  g2196 (n1901, n1115);
not  g2197 (n2397, n950);
buf  g2198 (n2335, n1787);
buf  g2199 (n2459, n1007);
buf  g2200 (n2394, n852);
buf  g2201 (n1987, n1632);
buf  g2202 (n2279, n1749);
not  g2203 (n1980, n1246);
not  g2204 (n2092, n1420);
buf  g2205 (n2022, n1550);
not  g2206 (n2190, n832);
buf  g2207 (n2521, n1222);
buf  g2208 (n2176, n1129);
not  g2209 (n2074, n1356);
buf  g2210 (n2084, n613);
not  g2211 (n1858, n1369);
not  g2212 (n2216, n882);
buf  g2213 (n1875, n671);
buf  g2214 (n2285, n786);
not  g2215 (n2008, n1063);
not  g2216 (n2320, n940);
buf  g2217 (n2389, n704);
not  g2218 (n2467, n939);
buf  g2219 (n1919, n1095);
not  g2220 (n2366, n1093);
buf  g2221 (n2245, n1765);
buf  g2222 (n2091, n1382);
not  g2223 (n2179, n1758);
not  g2224 (n2156, n1377);
not  g2225 (n2066, n963);
buf  g2226 (n2230, n1003);
buf  g2227 (n2347, n741);
not  g2228 (n1895, n1102);
not  g2229 (n1942, n1568);
not  g2230 (n1955, n1687);
not  g2231 (n2159, n896);
buf  g2232 (n2173, n1431);
not  g2233 (n2283, n923);
not  g2234 (n1972, n1699);
buf  g2235 (n2026, n982);
buf  g2236 (n2265, n1416);
buf  g2237 (n2259, n1259);
not  g2238 (n2432, n828);
not  g2239 (n2480, n1563);
not  g2240 (n2063, n1702);
buf  g2241 (n1917, n985);
not  g2242 (n2045, n721);
buf  g2243 (n2315, n1542);
buf  g2244 (n2030, n1119);
not  g2245 (n1974, n1791);
buf  g2246 (n2059, n987);
buf  g2247 (n1964, n1284);
buf  g2248 (n2403, n1299);
not  g2249 (n2309, n702);
buf  g2250 (n2371, n611);
buf  g2251 (n2268, n1156);
buf  g2252 (n2232, n1167);
buf  g2253 (n2111, n1232);
buf  g2254 (n1860, n1680);
not  g2255 (n2012, n930);
buf  g2256 (n2410, n1419);
buf  g2257 (n2316, n661);
not  g2258 (n2126, n658);
buf  g2259 (n2087, n1675);
buf  g2260 (n2472, n604);
buf  g2261 (n1976, n1756);
not  g2262 (n1878, n1745);
not  g2263 (n2081, n1415);
buf  g2264 (n2140, n1053);
not  g2265 (n2482, n1445);
buf  g2266 (n2314, n1594);
not  g2267 (n2247, n1482);
not  g2268 (n2468, n927);
not  g2269 (n2270, n1252);
not  g2270 (n2513, n1752);
not  g2271 (n2385, n634);
not  g2272 (n2013, n1096);
buf  g2273 (n2098, n862);
buf  g2274 (n2384, n1728);
buf  g2275 (n2473, n924);
buf  g2276 (n2458, n1037);
not  g2277 (n2077, n899);
buf  g2278 (n1881, n1174);
not  g2279 (n1986, n656);
not  g2280 (n2226, n1402);
buf  g2281 (n2427, n1776);
not  g2282 (n1872, n1339);
buf  g2283 (n2221, n738);
buf  g2284 (n2054, n813);
buf  g2285 (n2086, n1502);
not  g2286 (n2009, n1373);
buf  g2287 (n2165, n1730);
buf  g2288 (n2382, n1487);
not  g2289 (n2498, n1375);
not  g2290 (n1890, n965);
buf  g2291 (n2504, n701);
not  g2292 (n2355, n1249);
buf  g2293 (n2219, n1354);
not  g2294 (n2431, n975);
buf  g2295 (n2031, n1283);
not  g2296 (n2429, n1509);
buf  g2297 (n2183, n1360);
buf  g2298 (n2457, n737);
not  g2299 (n1867, n1574);
not  g2300 (n2487, n1666);
not  g2301 (n1866, n1009);
buf  g2302 (n2153, n1304);
buf  g2303 (n1991, n1033);
buf  g2304 (n2363, n1189);
buf  g2305 (n2109, n850);
buf  g2306 (n1907, n1489);
buf  g2307 (n2258, n1697);
buf  g2308 (n2197, n1590);
buf  g2309 (n2186, n1614);
not  g2310 (n2018, n1300);
buf  g2311 (n2150, n1205);
not  g2312 (n2175, n1621);
buf  g2313 (n2305, n1786);
buf  g2314 (n2452, n1577);
buf  g2315 (n1979, n1186);
buf  g2316 (n2225, n967);
buf  g2317 (n2254, n1774);
not  g2318 (n2120, n1010);
nor  g2319 (n1876, n1462, n1083);
xnor g2320 (n2524, n1789, n1086, n685, n753);
xor  g2321 (n2214, n1750, n1106, n1268, n1333);
nor  g2322 (n2161, n856, n1097, n755, n827);
xnor g2323 (n2405, n1185, n1015, n1460, n1467);
nand g2324 (n2163, n1674, n1532, n1025, n1602);
xnor g2325 (n1896, n1401, n1628, n898, n678);
nor  g2326 (n2019, n1153, n627, n1101, n769);
xnor g2327 (n2516, n920, n749, n1438, n1570);
or   g2328 (n2349, n969, n1408, n1080, n809);
xnor g2329 (n2328, n740, n808, n807, n1775);
nand g2330 (n2451, n994, n1131, n1270, n1751);
or   g2331 (n1961, n922, n1571, n1234, n1276);
or   g2332 (n2234, n916, n1008, n820, n1689);
xnor g2333 (n2333, n1667, n745, n1505, n1150);
or   g2334 (n2137, n978, n1587, n822, n1200);
or   g2335 (n2300, n901, n1795, n1127, n635);
and  g2336 (n2325, n1084, n1243, n893, n989);
nor  g2337 (n2436, n1456, n1227, n1794, n1592);
xnor g2338 (n1941, n675, n1087, n1242, n1660);
and  g2339 (n2474, n775, n670, n624, n1712);
nor  g2340 (n1940, n1427, n843, n1607, n1028);
xnor g2341 (n1863, n732, n1603, n1050, n699);
xnor g2342 (n2005, n1654, n684, n700, n1444);
xnor g2343 (n1862, n791, n1046, n1261, n1608);
or   g2344 (n2479, n1175, n875, n1077, n762);
or   g2345 (n2484, n815, n1545, n638, n1230);
xnor g2346 (n2068, n1629, n1068, n895, n1041);
nor  g2347 (n1908, n1094, n1387, n1159, n1371);
xor  g2348 (n1957, n953, n696, n771, n831);
and  g2349 (n2377, n650, n1199, n1611, n1734);
xor  g2350 (n1963, n1744, n1741, n1305, n1521);
and  g2351 (n1962, n664, n1468, n907, n1719);
or   g2352 (n1958, n1423, n615, n1190, n1410);
xor  g2353 (n1883, n1729, n770, n715, n644);
and  g2354 (n1905, n1481, n612, n1285, n1683);
or   g2355 (n2465, n1743, n597, n1764, n851);
nand g2356 (n2428, n1508, n868, n636, n1656);
or   g2357 (n2449, n1335, n1790, n1254, n1755);
xnor g2358 (n2313, n811, n593, n1202, n874);
nor  g2359 (n2021, n1526, n1516, n1350, n1177);
and  g2360 (n2160, n608, n909, n859, n592);
or   g2361 (n2297, n1519, n860, n1351, n913);
nand g2362 (n2079, n1090, n1517, n677, n1383);
nor  g2363 (n2296, n1113, n1715, n1677, n1395);
nor  g2364 (n2287, n1554, n1321, n1362, n778);
nor  g2365 (n2272, n1036, n1355, n1341, n1358);
nand g2366 (n2412, n1536, n1366, n1005, n1514);
nand g2367 (n2386, n599, n1017, n1146, n669);
nand g2368 (n2093, n799, n1623, n1091, n1149);
nor  g2369 (n2415, n1636, n667, n1770, n1079);
xor  g2370 (n2271, n1678, n1062, n970, n1633);
xor  g2371 (n2290, n1217, n1396, n1296, n1737);
nand g2372 (n2103, n1027, n1583, n839, n1534);
xor  g2373 (n2025, n1154, n1002, n846, n1781);
or   g2374 (n2143, n1556, n780, n938, n825);
or   g2375 (n2417, n1615, n878, n929, n1701);
and  g2376 (n1884, n1338, n674, n1287, n849);
nor  g2377 (n1936, n1512, n1657, n1157, n1649);
or   g2378 (n2500, n1171, n1798, n797, n1363);
or   g2379 (n2450, n1698, n1000, n1663, n1209);
nor  g2380 (n2424, n1215, n1672, n1547, n1486);
nor  g2381 (n2249, n1275, n1316, n619, n676);
or   g2382 (n2443, n960, n1183, n955, n1703);
or   g2383 (n1954, n687, n911, n686, n1295);
xnor g2384 (n2338, n900, n1471, n1784, n1342);
or   g2385 (n2437, n986, n790, n1397, n1253);
xor  g2386 (n2206, n1754, n1695, n706, n1271);
nor  g2387 (n2376, n607, n1648, n722, n1188);
or   g2388 (n1975, n1392, n1376, n1589, n1081);
nand g2389 (n2014, n876, n1541, n870, n1414);
nor  g2390 (n2207, n693, n796, n954, n1326);
nand g2391 (n2028, n1337, n727, n1004, n1216);
xnor g2392 (n2329, n1238, n1522, n867, n1349);
and  g2393 (n2116, n1440, n1398, n772, n1108);
xnor g2394 (n2003, n886, n1428, n1078, n798);
nor  g2395 (n1870, n1245, n1272, n1352, n887);
nor  g2396 (n2273, n1274, n1588, n1506, n1021);
nand g2397 (n2357, n1262, n1618, n1105, n1263);
xor  g2398 (n2491, n660, n1432, n1310, n1461);
and  g2399 (n2085, n1477, n1114, n905, n853);
nand g2400 (n2235, n861, n1579, n1069, n761);
nand g2401 (n2100, n972, n596, n834, n1411);
nor  g2402 (n2011, n652, n1282, n1569, n1451);
or   g2403 (n1893, n683, n697, n1389, n1221);
or   g2404 (n2370, n1345, n1100, n1346, n1673);
or   g2405 (n2228, n1581, n1595, n1513, n735);
nor  g2406 (n2409, n835, n836, n1152, n800);
xor  g2407 (n2408, n651, n806, n1560, n908);
xnor g2408 (n2353, n1286, n1088, n788, n1527);
xnor g2409 (n2060, n919, n865, n628, n1121);
nand g2410 (n2070, n1126, n935, n1314, n952);
xor  g2411 (n2118, n1289, n1619, n1147, n877);
xor  g2412 (n2494, n1447, n1014, n1616, n983);
or   g2413 (n2530, n1198, n765, n1448, n1766);
xnor g2414 (n1904, n1092, n712, n1320, n1372);
xnor g2415 (n2010, n1567, n618, n736, n1220);
nand g2416 (n2419, n1347, n1682, n1193, n841);
and  g2417 (n1985, n1732, n1182, n643, n823);
or   g2418 (n2466, n897, n606, n1450, n1379);
nand g2419 (n2211, n728, n1160, n717, n1163);
xor  g2420 (n2052, n1598, n998, n819, n1187);
and  g2421 (n2483, n1566, n716, n1586, n595);
or   g2422 (n2113, n1757, n720, n747, n842);
xnor g2423 (n1977, n1384, n944, n1706, n1696);
xor  g2424 (n1903, n873, n1039, n1422, n1196);
and  g2425 (n1981, n1409, n690, n1089, n655);
and  g2426 (n2044, n1179, n1386, n1421, n1045);
xor  g2427 (n1857, n885, n1609, n814, n1042);
xnor g2428 (n2114, n672, n1138, n1436, n598);
xnor g2429 (n2201, n1044, n833, n630, n1117);
xor  g2430 (n2151, n1133, n817, n1643, n1499);
nor  g2431 (n1937, n1430, n1011, n620, n1381);
nor  g2432 (n2177, n1591, n891, n1652, n1792);
nor  g2433 (n2182, n1503, n1640, n1639, n625);
nand g2434 (n2240, n1278, n1194, n626, n1012);
nand g2435 (n2512, n1771, n648, n590, n694);
and  g2436 (n2123, n821, n713, n1597, n1501);
and  g2437 (n2051, n1312, n1072, n763, n1676);
nand g2438 (n2017, n1612, n1247, n1557, n1693);
xor  g2439 (n1891, n816, n1066, n1391, n622);
xnor g2440 (n2368, n1480, n1071, n937, n1367);
xor  g2441 (n1910, n1006, n623, n766, n926);
xor  g2442 (n2364, n682, n787, n1073, n1294);
nor  g2443 (n2167, n1307, n1763, n1135, n1130);
and  g2444 (n2416, n1393, n1479, n748, n1558);
nand g2445 (n1989, n1098, n600, n1235, n948);
or   g2446 (n2204, n750, n689, n1504, n932);
xor  g2447 (n2072, n933, n1782, n1669, n1168);
xor  g2448 (n2373, n1739, n1780, n1145, n1169);
xnor g2449 (n2454, n871, n681, n1076, n973);
xnor g2450 (n2321, n631, n962, n1256, n1488);
xnor g2451 (n2062, n1353, n1721, n1142, n757);
nand g2452 (n2136, n864, n1740, n824, n1779);
xor  g2453 (n2288, n946, n884, n688, n659);
xor  g2454 (n2351, n1684, n1052, n1705, n1578);
nor  g2455 (n2108, n1601, n1470, n1424, n616);
nand g2456 (n1968, n783, n1713, n1443, n1212);
xor  g2457 (n2292, n691, n1231, n1539, n1197);
nor  g2458 (n1894, n1793, n1449, n1224, n1026);
and  g2459 (n2096, n719, n964, n1478, n1291);
xor  g2460 (n2061, n1406, n1013, n1711, n591);
xnor g2461 (n2082, n1399, n1107, n1116, n1796);
and  g2462 (n2106, n848, n991, n847, n1368);
xor  g2463 (n2508, n1180, n785, n1266, n1753);
or   g2464 (n2476, n1717, n1390, n1634, n904);
xor  g2465 (n2097, n746, n1537, n1664, n1308);
nand g2466 (n2236, n976, n1313, n1070, n1661);
xor  g2467 (n1924, n654, n1343, n1662, n609);
and  g2468 (n2243, n1645, n1495, n1250, n1228);
nor  g2469 (n2383, n647, n610, n826, n1483);
and  g2470 (n2071, n1407, n995, n993, n1203);
nand g2471 (n2471, n768, n863, n1029, n1219);
xnor g2472 (n1946, n1184, n1492, n1264, n1319);
nand g2473 (n1998, n760, n1112, n1546, n1201);
xnor g2474 (n2350, n1403, n1233, n996, n1336);
or   g2475 (n2127, n603, n1439, n1620, n1585);
nor  g2476 (n2330, n1496, n673, n1724, n629);
or   g2477 (n1956, n1688, n1653, n889, n981);
nand g2478 (n2036, n642, n1523, n776, n1165);
nor  g2479 (n2154, n754, n1625, n1600, n845);
nand g2480 (n2515, n855, n1564, n1318, n779);
xor  g2481 (n2456, n1269, n733, n1418, n1681);
and  g2482 (n1992, n1361, n1466, n1143, n645);
nand g2483 (n2327, n709, n1694, n1507, n641);
and  g2484 (n2130, n1637, n1279, n1746, n1529);
or   g2485 (n1994, n1725, n1404, n1708, n1596);
or   g2486 (n2438, n1485, n767, n1241, n1538);
xnor g2487 (n2038, n1726, n818, n1530, n1192);
or   g2488 (n2519, n734, n1206, n903, n1638);
or   g2489 (n2433, n1454, n1630, n1213, n1651);
or   g2490 (n2489, n1134, n1659, n1181, n1425);
and  g2491 (n2252, n1668, n1311, n1394, n1151);
xnor g2492 (n2299, n1173, n1064, n1258, n1210);
xnor g2493 (n2229, n1511, n1704, n1043, n1562);
xnor g2494 (n2306, n917, n1128, n1240, n1465);
or   g2495 (n1990, n947, n657, n1738, n1474);
and  g2496 (n2263, n1720, n777, n1019, n1207);
nor  g2497 (n1949, n1239, n1118, n1123, n1671);
nand g2498 (n2629, n563, n565, n2174, n2358);
nand g2499 (n2633, n2142, n559, n1977, n575);
nand g2500 (n2665, n1996, n2357, n559, n2165);
or   g2501 (n2562, n2311, n2275, n562, n2396);
xor  g2502 (n2556, n2072, n559, n2324, n564);
xnor g2503 (n2674, n1920, n2267, n1929, n2272);
xnor g2504 (n2617, n2067, n2231, n2034, n567);
xor  g2505 (n2580, n2073, n2191, n1911, n2141);
xor  g2506 (n2635, n546, n2225, n571, n561);
nand g2507 (n2564, n2250, n1944, n2203, n2273);
and  g2508 (n2645, n2147, n1943, n2149, n2040);
or   g2509 (n2569, n553, n547, n2125, n2354);
and  g2510 (n2576, n2045, n550, n1912, n545);
nor  g2511 (n2626, n2253, n2195, n578, n557);
xnor g2512 (n2654, n570, n2279, n2115, n2332);
nand g2513 (n2701, n2265, n2200, n2021, n2098);
and  g2514 (n2608, n2158, n1997, n2005, n2113);
xor  g2515 (n2679, n2126, n1914, n2095, n2385);
and  g2516 (n2684, n2127, n2247, n2353, n2041);
xor  g2517 (n2656, n2164, n579, n2359, n1923);
xor  g2518 (n2581, n2026, n2116, n1922, n1936);
and  g2519 (n2660, n2001, n2157, n2341, n553);
or   g2520 (n2579, n2283, n577, n1859, n1862);
nor  g2521 (n2575, n552, n2317, n2376, n568);
or   g2522 (n2669, n2387, n576, n1891, n1909);
xnor g2523 (n2640, n1975, n1954, n1983, n2234);
xor  g2524 (n2676, n2068, n2096, n1988, n2289);
and  g2525 (n2698, n2349, n2137, n2258, n2352);
nand g2526 (n2616, n2333, n2082, n1999, n2107);
nor  g2527 (n2601, n546, n2084, n562, n542);
and  g2528 (n2583, n2066, n551, n2018, n2097);
xnor g2529 (n2655, n555, n2269, n547, n2009);
xnor g2530 (n2551, n1987, n2048, n2148, n2060);
or   g2531 (n2699, n2344, n1979, n1915, n2057);
xor  g2532 (n2696, n2185, n551, n2061, n560);
nand g2533 (n2653, n2364, n2198, n2199, n2375);
xnor g2534 (n2686, n541, n2189, n543, n2336);
xor  g2535 (n2599, n2188, n2103, n2215, n556);
and  g2536 (n2534, n2031, n547, n1888, n548);
or   g2537 (n2559, n2287, n554, n560, n1892);
xnor g2538 (n2615, n2080, n567, n579, n2160);
nor  g2539 (n2682, n2260, n2383, n1945, n2393);
and  g2540 (n2637, n1872, n2136, n1867, n576);
nor  g2541 (n2590, n561, n2134, n2105, n1857);
xor  g2542 (n2570, n558, n2327, n580, n564);
xor  g2543 (n2638, n2312, n2280, n2259, n555);
xnor g2544 (n2543, n2088, n567, n2322, n1890);
and  g2545 (n2602, n2184, n1952, n2384, n2294);
nor  g2546 (n2667, n2178, n2338, n1895, n2173);
xor  g2547 (n2649, n562, n1864, n2047, n2254);
nor  g2548 (n2659, n1972, n541, n1935, n1933);
or   g2549 (n2687, n2074, n2335, n2159, n2085);
nand g2550 (n2677, n2342, n2235, n1925, n1882);
and  g2551 (n2584, n2218, n2271, n2121, n1957);
and  g2552 (n2606, n1982, n1994, n2372, n2297);
xnor g2553 (n2619, n2326, n2181, n576, n2301);
nor  g2554 (n2612, n2270, n1889, n2024, n2256);
or   g2555 (n2571, n547, n2204, n2029, n2167);
xor  g2556 (n2572, n2140, n2340, n2062, n2243);
and  g2557 (n2681, n578, n2156, n2330, n552);
or   g2558 (n2651, n2089, n2076, n2263, n1955);
nand g2559 (n2690, n2039, n2374, n2362, n573);
nand g2560 (n2607, n1898, n2237, n2211, n2087);
nand g2561 (n2692, n2094, n1953, n2346, n2122);
nand g2562 (n2678, n1973, n566, n2251, n2356);
xnor g2563 (n2593, n2171, n2153, n2206, n2321);
xnor g2564 (n2549, n546, n1962, n2379, n572);
xor  g2565 (n2565, n2227, n1949, n2300, n2299);
xor  g2566 (n2548, n2197, n1976, n2224, n2007);
xor  g2567 (n2693, n2038, n2131, n1965, n549);
and  g2568 (n2623, n2023, n1913, n1861, n2310);
or   g2569 (n2618, n1879, n2304, n1971, n2130);
xor  g2570 (n2683, n2193, n2207, n1876, n559);
nor  g2571 (n2563, n2331, n2071, n574, n1897);
nand g2572 (n2634, n545, n549, n1937, n2285);
nand g2573 (n2545, n574, n1921, n2064, n2223);
xnor g2574 (n2624, n546, n1904, n2276, n2129);
nor  g2575 (n2537, n1991, n2182, n2216, n2296);
xnor g2576 (n2550, n2090, n1924, n1893, n2391);
nand g2577 (n2557, n572, n574, n1871);
xor  g2578 (n2688, n2004, n2124, n2264, n2170);
and  g2579 (n2621, n2081, n2006, n572, n2008);
nand g2580 (n2625, n1958, n2108, n2011, n1960);
nor  g2581 (n2695, n2120, n2106, n2086, n2220);
nand g2582 (n2700, n557, n1870, n561, n1927);
xor  g2583 (n2631, n571, n2161, n2282, n2014);
xor  g2584 (n2546, n1932, n2239, n564, n2030);
xor  g2585 (n2657, n2102, n1877, n1868, n551);
and  g2586 (n2611, n2051, n553, n1894, n550);
xnor g2587 (n2573, n2050, n1951, n2168, n2292);
xor  g2588 (n2630, n575, n1940, n571, n2183);
nor  g2589 (n2532, n2278, n1930, n2348, n565);
nor  g2590 (n2536, n1961, n2196, n2144, n1998);
and  g2591 (n2666, n2214, n2205, n568);
nor  g2592 (n2650, n2010, n2055, n2065, n2118);
and  g2593 (n2595, n1908, n2128, n560, n569);
xnor g2594 (n2597, n1978, n2132, n2143, n566);
or   g2595 (n2672, n2369, n2054, n2226, n1874);
or   g2596 (n2610, n2314, n2295, n1916, n1992);
xor  g2597 (n2636, n2133, n2303, n2163, n2036);
nor  g2598 (n2603, n1869, n2380, n2389, n1866);
or   g2599 (n2533, n567, n2366, n2392, n1950);
nor  g2600 (n2582, n2000, n2056, n573, n2192);
nor  g2601 (n2585, n569, n573, n2078, n1907);
xor  g2602 (n2591, n2365, n555, n1946, n2293);
xnor g2603 (n2689, n551, n2049, n2092, n2176);
and  g2604 (n2663, n568, n2252, n543, n1974);
nand g2605 (n2567, n563, n2210, n569, n549);
nand g2606 (n2558, n2249, n2079, n2248, n2025);
nor  g2607 (n2553, n563, n561, n2244, n2347);
and  g2608 (n2703, n2135, n2395, n2329, n570);
nor  g2609 (n2628, n1881, n2394, n1956, n2228);
xor  g2610 (n2578, n580, n2212, n2268, n2177);
xor  g2611 (n2671, n1995, n579, n549, n1964);
xnor g2612 (n2588, n2172, n2016, n1928, n577);
xnor g2613 (n2541, n577, n2242, n1918, n2052);
xnor g2614 (n2566, n556, n556, n2077, n2233);
nor  g2615 (n2648, n2377, n1875, n2033, n2281);
and  g2616 (n2586, n2319, n2044, n2138, n2187);
nor  g2617 (n2577, n2230, n1858, n1917, n2217);
xnor g2618 (n2641, n2219, n2111, n2179, n2307);
or   g2619 (n2531, n558, n2070, n1880, n548);
nor  g2620 (n2555, n557, n1990, n2020, n1887);
and  g2621 (n2661, n1860, n575, n2334, n552);
xnor g2622 (n2627, n576, n2104, n2325, n1910);
xor  g2623 (n2604, n2069, n2154, n580, n2110);
nor  g2624 (n2668, n554, n2345, n2240, n2305);
and  g2625 (n2544, n2190, n2246, n2241, n2180);
nor  g2626 (n2574, n578, n1903, n2063, n2355);
nand g2627 (n2552, n2361, n2284, n2277, n2290);
and  g2628 (n2594, n2155, n1984, n2043, n2302);
nand g2629 (n2673, n2012, n1947, n575, n2288);
or   g2630 (n2664, n572, n2274, n542, n2022);
xor  g2631 (n2694, n2222, n2313, n550, n1963);
nor  g2632 (n2704, n2245, n566, n2397, n2286);
and  g2633 (n2568, n2208, n2037, n571, n2058);
or   g2634 (n2658, n2053, n558, n2367, n1948);
nor  g2635 (n2596, n2019, n2145, n2386, n1865);
or   g2636 (n2600, n2101, n2027, n1980, n2059);
xor  g2637 (n2620, n2209, n2151, n2360, n2042);
or   g2638 (n2685, n1985, n2368, n1934, n565);
nor  g2639 (n2675, n2236, n2337, n2261, n1959);
and  g2640 (n2560, n1886, n2162, n2150, n1986);
xor  g2641 (n2632, n558, n2112, n2083, n2238);
or   g2642 (n2642, n2099, n560, n1938, n2175);
nand g2643 (n2539, n2306, n2093, n2032, n2318);
nor  g2644 (n2547, n542, n2035, n1970, n1941);
nor  g2645 (n2691, n1969, n2309, n544, n2186);
and  g2646 (n2589, n2262, n2255, n1926, n2351);
xnor g2647 (n2647, n1905, n542, n564, n2291);
xor  g2648 (n2670, n2013, n2152, n2339, n1989);
nand g2649 (n2644, n579, n545, n1878, n543);
nand g2650 (n2652, n2316, n570, n2381, n1968);
or   g2651 (n2561, n2370, n1942, n545, n2169);
xor  g2652 (n2613, n569, n2194, n566, n2109);
or   g2653 (n2587, n2100, n2117, n552, n1939);
xor  g2654 (n2680, n2323, n562, n2046, n2075);
nor  g2655 (n2605, n2266, n570, n2015, n1902);
nor  g2656 (n2598, n1966, n2017, n548, n557);
nor  g2657 (n2540, n1873, n573, n2308, n2028);
or   g2658 (n2542, n1919, n1981, n2373, n543);
and  g2659 (n2697, n2315, n1900, n554, n2213);
xor  g2660 (n2554, n1899, n1896, n556, n2146);
nand g2661 (n2614, n544, n2166, n2139, n1901);
nor  g2662 (n2646, n2257, n1906, n1885, n1931);
and  g2663 (n2639, n580, n548, n2221, n2003);
nor  g2664 (n2592, n2229, n2201, n1863, n2343);
xnor g2665 (n2622, n565, n578, n554, n2320);
or   g2666 (n2643, n555, n1883, n2232, n2298);
and  g2667 (n2702, n2002, n2388, n2119, n2091);
xor  g2668 (n2535, n2378, n563, n2371, n544);
or   g2669 (n2705, n550, n577, n2123, n2114);
nor  g2670 (n2662, n544, n2390, n2202, n1884);
xor  g2671 (n2609, n2350, n1967, n541, n553);
nor  g2672 (n2538, n2328, n1993, n2382, n2363);
buf  g2673 (n2710, n2559);
buf  g2674 (n2722, n2534);
buf  g2675 (n2712, n2542);
buf  g2676 (n2727, n2537);
not  g2677 (n2719, n2547);
not  g2678 (n2732, n2548);
buf  g2679 (n2717, n2533);
not  g2680 (n2726, n2554);
buf  g2681 (n2714, n2532);
not  g2682 (n2725, n2541);
not  g2683 (n2734, n2550);
buf  g2684 (n2721, n2561);
not  g2685 (n2730, n2535);
not  g2686 (n2731, n2558);
buf  g2687 (n2728, n2540);
buf  g2688 (n2706, n2545);
buf  g2689 (n2713, n2539);
not  g2690 (n2708, n2557);
buf  g2691 (n2716, n2556);
buf  g2692 (n2736, n2549);
not  g2693 (n2715, n2536);
not  g2694 (n2707, n2555);
not  g2695 (n2709, n2553);
buf  g2696 (n2718, n2560);
not  g2697 (n2737, n2551);
buf  g2698 (n2733, n2552);
not  g2699 (n2711, n2544);
buf  g2700 (n2724, n2546);
not  g2701 (n2723, n2538);
buf  g2702 (n2735, n2562);
not  g2703 (n2720, n2543);
not  g2704 (n2729, n2531);
nand g2705 (n2745, n2709, n2429, n581, n2403);
xnor g2706 (n2752, n2439, n2416, n2706, n2402);
xor  g2707 (n2747, n2709, n2418, n2400, n2398);
nor  g2708 (n2750, n2708, n2708, n2427, n2399);
xor  g2709 (n2740, n2407, n2423, n2443, n2708);
xor  g2710 (n2748, n2417, n2709, n2708, n2401);
xnor g2711 (n2739, n2436, n2415, n2442, n2437);
xor  g2712 (n2743, n2426, n2706, n2434, n2707);
nor  g2713 (n2742, n2420, n2409, n2440, n2435);
xor  g2714 (n2744, n2411, n2706, n2441, n2438);
xnor g2715 (n2746, n2410, n2413, n2707, n2424);
and  g2716 (n2741, n2706, n2414, n2404, n2422);
nor  g2717 (n2749, n2412, n2408, n2405, n581);
or   g2718 (n2753, n2707, n2430, n2433, n2431);
and  g2719 (n2738, n2709, n2419, n2421, n2428);
xor  g2720 (n2751, n2425, n2707, n2406, n2432);
xnor g2721 (n2755, n1806, n1801, n1803, n1810);
nand g2722 (n2757, n2739, n2740, n2738, n1807);
and  g2723 (n2756, n1805, n1804, n1808, n2741);
xor  g2724 (n2754, n1802, n1799, n1800, n1809);
or   g2725 (n2760, n2757, n2450, n2755, n2448);
or   g2726 (n2759, n2449, n2452, n2444, n2445);
and  g2727 (n2758, n2756, n2447, n2446, n2451);
not  g2728 (n2768, n2760);
not  g2729 (n2765, n2565);
buf  g2730 (n2771, n2581);
buf  g2731 (n2772, n2566);
and  g2732 (n2767, n2567, n2760, n2577, n2586);
and  g2733 (n2769, n2563, n2759, n2583);
nor  g2734 (n2766, n2570, n2760, n2758, n2572);
nor  g2735 (n2762, n2582, n2758, n2584);
nand g2736 (n2770, n2574, n2564, n2580, n2573);
nand g2737 (n2761, n2758, n2569, n2571, n2760);
xnor g2738 (n2764, n2576, n2585, n2575, n2759);
nand g2739 (n2763, n2579, n2568, n2759, n2578);
and  g2740 (n2775, n581, n2728, n2725, n2712);
nor  g2741 (n2808, n2719, n2768, n583);
and  g2742 (n2796, n2761, n584, n2456, n2718);
xor  g2743 (n2777, n2761, n2724, n2770, n2716);
and  g2744 (n2809, n2717, n30, n2725, n2721);
xor  g2745 (n2802, n32, n581, n583, n2727);
nor  g2746 (n2793, n2767, n2766, n584, n30);
nand g2747 (n2784, n2724, n2721, n2765, n584);
xor  g2748 (n2801, n2722, n2722, n2764, n2767);
and  g2749 (n2776, n2765, n2721, n2766, n2723);
xor  g2750 (n2794, n2454, n2769, n2726, n2717);
or   g2751 (n2806, n2764, n2720, n2713, n2725);
xnor g2752 (n2778, n31, n2453, n2761, n2718);
xor  g2753 (n2779, n2711, n2716, n2722, n2720);
or   g2754 (n2788, n2711, n29, n2713, n32);
and  g2755 (n2789, n2762, n2762, n583, n2769);
xor  g2756 (n2780, n2726, n582, n2763, n585);
xnor g2757 (n2797, n2767, n2726, n2710, n2727);
nor  g2758 (n2790, n2721, n2714, n2715, n2710);
nand g2759 (n2799, n2716, n2724, n30, n2719);
or   g2760 (n2805, n2720, n582, n2717, n2712);
and  g2761 (n2774, n32, n2714, n2711, n29);
and  g2762 (n2798, n2713, n2455, n2712, n32);
xnor g2763 (n2773, n2723, n2764, n2768, n2724);
or   g2764 (n2787, n2727, n2720, n31, n2726);
xnor g2765 (n2804, n2723, n2763, n2718, n2728);
nor  g2766 (n2800, n2716, n2710, n29, n2763);
nand g2767 (n2807, n2761, n2766, n2713, n30);
xnor g2768 (n2782, n2766, n2711, n2719, n2765);
xnor g2769 (n2803, n2763, n2764, n2717, n2767);
and  g2770 (n2792, n2710, n2728, n2762, n582);
xnor g2771 (n2795, n584, n2769, n585, n29);
or   g2772 (n2781, n2768, n2762, n31, n2725);
and  g2773 (n2783, n2715, n2718, n2719, n2727);
nor  g2774 (n2791, n2715, n2723, n2722, n583);
xnor g2775 (n2786, n2712, n2715, n2714);
and  g2776 (n2785, n31, n582, n2769, n2765);
not  g2777 (n2811, n2802);
not  g2778 (n2810, n2803);
xnor g2779 (n2815, n588, n587, n586);
nor  g2780 (n2812, n586, n2810, n587, n585);
and  g2781 (n2814, n2810, n2810, n586, n587);
nor  g2782 (n2813, n588, n585, n586, n2810);
nand g2783 (n2821, n1825, n1815, n1827, n1833);
and  g2784 (n2818, n2815, n1823, n1834, n1819);
and  g2785 (n2822, n2812, n1822, n1829, n1831);
nor  g2786 (n2817, n2813, n1811, n1824, n1830);
nand g2787 (n2816, n1820, n1832, n2814, n1813);
and  g2788 (n2819, n1816, n1814, n1812, n2814);
xor  g2789 (n2823, n1828, n1818, n1817, n2813);
or   g2790 (n2820, n1821, n1826, n2815, n2812);
not  g2791 (n2824, n2822);
buf  g2792 (n2825, n2462);
buf  g2793 (n2826, n2820);
buf  g2794 (n2832, n2821);
not  g2795 (n2831, n2816);
not  g2796 (n2833, n2822);
buf  g2797 (n2830, n2457);
buf  g2798 (n2827, n2459);
xor  g2799 (n2829, n2461, n2820, n2821, n2817);
xor  g2800 (n2828, n2460, n2818, n2458, n2819);
and  g2801 (n2834, n2589, n2592, n2824, n2591);
xnor g2802 (n2835, n2590, n2824, n2587, n2588);
nor  g2803 (n2840, n2734, n2835, n2730, n2729);
and  g2804 (n2843, n2731, n2835, n2733, n2730);
nor  g2805 (n2838, n2834, n2730, n2734);
nand g2806 (n2842, n2834, n2732);
and  g2807 (n2837, n2732, n2834, n2729, n2733);
and  g2808 (n2841, n2733, n2732, n2730, n2835);
or   g2809 (n2839, n2729, n2835, n2731, n2733);
nor  g2810 (n2836, n2731, n2731, n2728, n2729);
buf  g2811 (n2873, n2828);
not  g2812 (n2848, n2474);
not  g2813 (n2871, n2843);
xor  g2814 (n2854, n2735, n2829, n2836, n2831);
nor  g2815 (n2847, n2829, n2838, n1842, n2826);
xor  g2816 (n2844, n2468, n2748, n2839, n2832);
xnor g2817 (n2865, n2842, n2827, n1837, n2832);
nand g2818 (n2858, n2752, n1849, n2838, n2833);
nand g2819 (n2870, n1844, n2842, n2464, n2476);
nor  g2820 (n2849, n2735, n2843, n2841, n2833);
nor  g2821 (n2856, n2840, n2839, n2826);
nand g2822 (n2866, n2745, n2828, n2469, n1839);
xnor g2823 (n2874, n1846, n2827, n2825, n2475);
and  g2824 (n2864, n2753, n1841, n2841, n2840);
nor  g2825 (n2850, n2463, n2751, n2843, n2735);
nand g2826 (n2857, n2842, n2824, n1847, n1836);
nand g2827 (n2859, n2746, n2472, n2838, n1848);
or   g2828 (n2852, n2840, n1845, n2837);
nor  g2829 (n2853, n2832, n2465, n1838, n2828);
or   g2830 (n2868, n2842, n2825, n2829, n2827);
xnor g2831 (n2867, n2743, n2827, n2830, n2747);
nor  g2832 (n2846, n2836, n2471, n2466, n1840);
or   g2833 (n2851, n2744, n2839, n2829, n2828);
nand g2834 (n2862, n2830, n2839, n2831, n2841);
nand g2835 (n2860, n1843, n2734, n2838, n2831);
or   g2836 (n2869, n2841, n2832, n2837, n2843);
nand g2837 (n2863, n2826, n144, n1835);
nor  g2838 (n2875, n2837, n2473, n2830, n2467);
or   g2839 (n2845, n2831, n2824, n2836);
and  g2840 (n2861, n2825, n144, n2833, n2830);
nand g2841 (n2855, n2825, n2750, n2749, n2742);
xnor g2842 (n2872, n2735, n2840, n2833, n2470);
not  g2843 (n2879, n2844);
not  g2844 (n2877, n2844);
not  g2845 (n2878, n2844);
buf  g2846 (n2876, n2844);
buf  g2847 (n2881, n2876);
not  g2848 (n2880, n2876);
xor  g2849 (n2882, n2771, n2479, n2482, n2772);
nand g2850 (n2888, n2481, n2771, n2483, n2770);
and  g2851 (n2883, n2770, n2772, n2881);
nand g2852 (n2886, n2484, n2485, n2880, n2772);
xnor g2853 (n2884, n2478, n2771, n2772, n2880);
nand g2854 (n2885, n2480, n2477, n2880);
nand g2855 (n2887, n2770, n2486, n2881, n2771);
or   g2856 (n2890, n2600, n2882, n2888, n2596);
or   g2857 (n2892, n2604, n2888, n2605, n2808);
xnor g2858 (n2896, n2609, n2599, n2884, n2593);
or   g2859 (n2895, n2607, n2610, n2608, n2809);
xnor g2860 (n2894, n2805, n2806, n2606, n2594);
xnor g2861 (n2893, n2597, n2886, n2595, n2807);
and  g2862 (n2889, n2883, n2804, n2598, n2887);
and  g2863 (n2891, n2602, n2603, n2601, n2885);
not  g2864 (n2900, n2811);
buf  g2865 (n2898, n2811);
buf  g2866 (n2897, n2890);
nor  g2867 (n2899, n2891, n2889);
nor  g2868 (n2901, n2889, n2811, n2890);
and  g2869 (n2905, n2489, n589, n588, n1850);
nor  g2870 (n2904, n2488, n2493, n2494, n588);
nor  g2871 (n2902, n2487, n2897, n2492);
or   g2872 (n2903, n2490, n2491, n2897);
xnor g2873 (n2906, n2902, n2881, n1854, n2905);
xnor g2874 (n2908, n2495, n1855, n2823, n2496);
or   g2875 (n2907, n2903, n1856, n1852, n2497);
xnor g2876 (n2909, n1853, n2904, n1851, n2823);
not  g2877 (n2911, n2909);
buf  g2878 (n2910, n2907);
buf  g2879 (n2912, n2908);
nand g2880 (n2923, n2510, n2894, n2503, n2896);
or   g2881 (n2916, n2611, n2893, n2910, n2896);
nor  g2882 (n2914, n2912, n2910, n2896);
nor  g2883 (n2921, n2499, n2912, n2612, n2891);
nor  g2884 (n2920, n2511, n2895, n2892, n2500);
nand g2885 (n2915, n2894, n2504, n2895, n2498);
nor  g2886 (n2917, n2505, n2911, n2512, n2912);
nor  g2887 (n2922, n2893, n2911, n2506);
and  g2888 (n2918, n2911, n2613, n2892, n2508);
nor  g2889 (n2913, n2894, n2509, n2895, n2501);
nand g2890 (n2919, n2502, n2893, n2912, n2507);
or   g2891 (n2935, n2692, n2621, n2679, n2899);
xor  g2892 (n2961, n2918, n2899, n2901, n2634);
or   g2893 (n2926, n2668, n2922, n2920, n2648);
and  g2894 (n2960, n2650, n2671, n2667, n2919);
nor  g2895 (n2951, n2654, n2915, n2917, n2900);
xor  g2896 (n2945, n2694, n2651, n2690, n2693);
and  g2897 (n2942, n2919, n2915, n2736, n2917);
and  g2898 (n2936, n2663, n2918, n2687, n2914);
nor  g2899 (n2948, n2921, n2657, n2697, n2631);
nand g2900 (n2941, n589, n2659, n2636, n2653);
or   g2901 (n2959, n2900, n2630, n2704, n2678);
nand g2902 (n2949, n2736, n2618, n2898, n2617);
xnor g2903 (n2962, n2699, n2691, n2898, n2649);
nand g2904 (n2939, n2705, n2637, n2661, n2642);
nor  g2905 (n2943, n2700, n2899, n2921, n2914);
and  g2906 (n2950, n2920, n2645, n2673, n2923);
nor  g2907 (n2940, n2914, n2695, n2913, n2646);
and  g2908 (n2947, n2628, n2647, n2737, n2660);
xor  g2909 (n2955, n2641, n2917, n2698, n2737);
or   g2910 (n2933, n2916, n2624, n2702, n2899);
xnor g2911 (n2927, n2898, n2696, n2652, n2629);
or   g2912 (n2954, n2701, n2901, n2680, n2913);
nand g2913 (n2932, n2913, n2620, n2915, n2632);
xnor g2914 (n2953, n2922, n2640, n2643, n2616);
or   g2915 (n2925, n2916, n2619, n2914, n2918);
xor  g2916 (n2930, n2669, n2677, n2676, n2625);
nand g2917 (n2944, n2919, n2684, n2623, n2670);
or   g2918 (n2956, n2922, n2675, n2900, n2664);
xor  g2919 (n2937, n2672, n2686, n2674, n589);
nand g2920 (n2958, n2918, n2615, n2627, n2682);
nor  g2921 (n2929, n2683, n2658, n2614, n2703);
xor  g2922 (n2957, n2622, n2921, n2737);
nor  g2923 (n2946, n2635, n2633, n2662, n2901);
xnor g2924 (n2928, n2639, n2688, n2920, n2736);
or   g2925 (n2938, n2666, n2638, n2685, n2655);
or   g2926 (n2931, n2898, n2736, n2916, n2665);
xor  g2927 (n2963, n2681, n2922, n2689, n2916);
nand g2928 (n2924, n2656, n2901, n2920, n2915);
xor  g2929 (n2934, n2644, n2737, n2900, n2626);
nand g2930 (n2952, n2919, n2513, n2917, n589);
nand g2931 (n2984, n2863, n2952, n2848, n2959);
xnor g2932 (n2976, n2847, n2852, n2864, n2858);
or   g2933 (n2989, n2948, n2963, n2850, n2855);
and  g2934 (n2994, n2857, n2866, n2862);
and  g2935 (n2991, n2872, n2864, n2855, n2865);
or   g2936 (n2999, n2931, n2962, n2864, n2851);
xor  g2937 (n2980, n2872, n2848, n2947, n2949);
nor  g2938 (n2996, n2846, n2521, n2861, n2522);
or   g2939 (n2971, n2871, n2853, n2924, n2941);
xnor g2940 (n2977, n2811, n2853, n2845);
xnor g2941 (n3004, n2870, n2854, n2945, n2861);
or   g2942 (n2992, n2862, n2868, n2961, n2525);
or   g2943 (n2998, n2860, n2865, n2847, n2871);
nor  g2944 (n2967, n2851, n2872, n2849, n2867);
xnor g2945 (n2974, n2862, n2515, n2854, n2939);
xnor g2946 (n2970, n2852, n2960, n2858, n2868);
nand g2947 (n3003, n2875, n2858, n2955, n2860);
nor  g2948 (n2972, n2850, n2850, n2518, n2528);
nand g2949 (n3002, n2940, n2869, n2953, n2849);
nand g2950 (n2985, n2936, n2861, n2865, n2526);
nand g2951 (n2981, n2960, n2519, n2856, n2848);
or   g2952 (n2995, n2856, n2926, n2857, n2871);
xor  g2953 (n3009, n2871, n2845, n2872, n2867);
nor  g2954 (n3000, n2946, n2864, n2846);
xnor g2955 (n2965, n2856, n2962, n2859);
xnor g2956 (n3006, n2851, n2875, n2870, n2849);
nand g2957 (n2986, n2853, n2957, n2874, n2867);
xnor g2958 (n2978, n2958, n2870, n2516, n2851);
xor  g2959 (n2966, n2846, n2933, n2959, n2847);
xnor g2960 (n2973, n2866, n2958, n2858, n2930);
xor  g2961 (n2982, n2857, n2855, n2874, n2873);
xnor g2962 (n2969, n2956, n2868, n2944);
or   g2963 (n2964, n2523, n2855, n2954, n2928);
or   g2964 (n2997, n2860, n2524, n2932, n2861);
xnor g2965 (n2987, n2852, n2963, n2867, n2961);
xnor g2966 (n2968, n2934, n2869, n2854, n2957);
xor  g2967 (n2983, n2873, n2935, n2527, n2929);
and  g2968 (n3005, n2950, n2845, n2874, n2859);
nand g2969 (n3011, n2865, n2937, n2875, n2955);
xor  g2970 (n2990, n2860, n2954, n2873, n2856);
or   g2971 (n3007, n2956, n2870, n2927, n2869);
and  g2972 (n2979, n2854, n2863, n2514, n2849);
or   g2973 (n2988, n2866, n2853, n2859, n2520);
and  g2974 (n2975, n2857, n2873, n2847, n2925);
and  g2975 (n3008, n2850, n2530, n2863, n2938);
xnor g2976 (n2993, n2852, n2848, n2942, n2529);
and  g2977 (n3010, n2869, n2951, n2517, n2874);
and  g2978 (n3001, n2875, n2943, n2863, n2866);
and  g2979 (n3012, n2982, n2977, n3006, n2970);
xor  g2980 (n3022, n2978, n2997, n2995, n2985);
xnor g2981 (n3024, n2969, n2989, n2879, n2877);
xnor g2982 (n3020, n2967, n3007, n3000, n2876);
xnor g2983 (n3014, n2879, n2879, n2976, n2972);
xor  g2984 (n3021, n2878, n2878, n2971, n2994);
xor  g2985 (n3013, n2878, n2964, n3010, n2993);
xor  g2986 (n3017, n2980, n2973, n2877, n2966);
or   g2987 (n3023, n2879, n2986, n2923);
and  g2988 (n3026, n2923, n3002, n2878, n3001);
or   g2989 (n3016, n2987, n2996, n2991, n3003);
and  g2990 (n3015, n3009, n2965, n3004, n2999);
and  g2991 (n3025, n3008, n2990, n2968, n2992);
nor  g2992 (n3027, n2984, n2988, n2983, n2998);
xnor g2993 (n3019, n2981, n2877, n3011, n2974);
or   g2994 (n3018, n2979, n2975, n3005, n2877);
xnor g2995 (n3030, n3023, n3020, n3017, n3016);
xnor g2996 (n3028, n3025, n3019, n3013, n3015);
nand g2997 (n3031, n3014, n3027, n3012, n3024);
or   g2998 (n3029, n3018, n3021, n3022, n3026);
nand g2999 (n3032, n3030, n3031, n3028, n3029);
endmodule
