// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_157 written by SynthGen on 2021/04/05 11:08:35
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_157 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n638, n733, n759, n753, n778, n775, n768, n748,
 n758, n779, n754, n750, n734, n751, n745, n762,
 n771, n767, n776, n747, n740, n756, n798, n1032,
 n1027, n1024, n1025, n1030, n1026, n1028, n1029, n1031);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n638, n733, n759, n753, n778, n775, n768, n748,
 n758, n779, n754, n750, n734, n751, n745, n762,
 n771, n767, n776, n747, n740, n756, n798, n1032,
 n1027, n1024, n1025, n1030, n1026, n1028, n1029, n1031;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n616,
 n617, n618, n619, n620, n621, n622, n623, n624,
 n625, n626, n627, n628, n629, n630, n631, n632,
 n633, n634, n635, n636, n637, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n735, n736, n737, n738, n739,
 n741, n742, n743, n744, n746, n749, n752, n755,
 n757, n760, n761, n763, n764, n765, n766, n769,
 n770, n772, n773, n774, n777, n780, n781, n782,
 n783, n784, n785, n786, n787, n788, n789, n790,
 n791, n792, n793, n794, n795, n796, n797, n799,
 n800, n801, n802, n803, n804, n805, n806, n807,
 n808, n809, n810, n811, n812, n813, n814, n815,
 n816, n817, n818, n819, n820, n821, n822, n823,
 n824, n825, n826, n827, n828, n829, n830, n831,
 n832, n833, n834, n835, n836, n837, n838, n839,
 n840, n841, n842, n843, n844, n845, n846, n847,
 n848, n849, n850, n851, n852, n853, n854, n855,
 n856, n857, n858, n859, n860, n861, n862, n863,
 n864, n865, n866, n867, n868, n869, n870, n871,
 n872, n873, n874, n875, n876, n877, n878, n879,
 n880, n881, n882, n883, n884, n885, n886, n887,
 n888, n889, n890, n891, n892, n893, n894, n895,
 n896, n897, n898, n899, n900, n901, n902, n903,
 n904, n905, n906, n907, n908, n909, n910, n911,
 n912, n913, n914, n915, n916, n917, n918, n919,
 n920, n921, n922, n923, n924, n925, n926, n927,
 n928, n929, n930, n931, n932, n933, n934, n935,
 n936, n937, n938, n939, n940, n941, n942, n943,
 n944, n945, n946, n947, n948, n949, n950, n951,
 n952, n953, n954, n955, n956, n957, n958, n959,
 n960, n961, n962, n963, n964, n965, n966, n967,
 n968, n969, n970, n971, n972, n973, n974, n975,
 n976, n977, n978, n979, n980, n981, n982, n983,
 n984, n985, n986, n987, n988, n989, n990, n991,
 n992, n993, n994, n995, n996, n997, n998, n999,
 n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
 n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
 n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;

not  g0 (n50, n13);
buf  g1 (n69, n11);
not  g2 (n86, n20);
buf  g3 (n84, n17);
not  g4 (n37, n21);
buf  g5 (n43, n4);
not  g6 (n115, n7);
not  g7 (n49, n14);
not  g8 (n88, n17);
buf  g9 (n100, n16);
buf  g10 (n98, n19);
buf  g11 (n44, n10);
buf  g12 (n63, n4);
buf  g13 (n87, n16);
buf  g14 (n108, n7);
buf  g15 (n111, n7);
not  g16 (n104, n16);
not  g17 (n67, n13);
buf  g18 (n113, n22);
not  g19 (n70, n2);
buf  g20 (n106, n3);
not  g21 (n81, n12);
not  g22 (n38, n9);
buf  g23 (n91, n6);
buf  g24 (n55, n18);
not  g25 (n33, n8);
buf  g26 (n90, n5);
not  g27 (n85, n9);
not  g28 (n116, n20);
buf  g29 (n41, n21);
buf  g30 (n114, n3);
buf  g31 (n34, n12);
buf  g32 (n53, n2);
buf  g33 (n93, n10);
not  g34 (n71, n6);
buf  g35 (n51, n10);
buf  g36 (n79, n14);
buf  g37 (n110, n7);
not  g38 (n74, n1);
buf  g39 (n54, n21);
not  g40 (n95, n14);
buf  g41 (n82, n18);
buf  g42 (n105, n3);
not  g43 (n39, n13);
not  g44 (n59, n1);
buf  g45 (n47, n15);
buf  g46 (n76, n1);
buf  g47 (n60, n19);
buf  g48 (n75, n20);
buf  g49 (n64, n18);
not  g50 (n102, n17);
not  g51 (n89, n12);
buf  g52 (n118, n19);
buf  g53 (n48, n11);
buf  g54 (n40, n8);
buf  g55 (n107, n22);
buf  g56 (n112, n6);
buf  g57 (n78, n9);
not  g58 (n72, n11);
not  g59 (n36, n12);
not  g60 (n97, n5);
not  g61 (n80, n8);
not  g62 (n109, n1);
not  g63 (n57, n2);
buf  g64 (n52, n3);
buf  g65 (n73, n18);
buf  g66 (n68, n14);
not  g67 (n42, n5);
buf  g68 (n46, n20);
not  g69 (n83, n8);
buf  g70 (n56, n2);
not  g71 (n94, n6);
not  g72 (n45, n4);
buf  g73 (n66, n16);
buf  g74 (n101, n15);
not  g75 (n58, n15);
buf  g76 (n35, n5);
not  g77 (n62, n9);
buf  g78 (n61, n19);
buf  g79 (n77, n15);
buf  g80 (n99, n21);
not  g81 (n65, n4);
buf  g82 (n92, n11);
buf  g83 (n96, n13);
not  g84 (n117, n17);
not  g85 (n103, n10);
not  g86 (n163, n72);
not  g87 (n172, n49);
buf  g88 (n150, n70);
not  g89 (n209, n39);
not  g90 (n169, n46);
buf  g91 (n242, n48);
not  g92 (n282, n46);
not  g93 (n141, n34);
not  g94 (n243, n62);
not  g95 (n137, n68);
not  g96 (n232, n35);
not  g97 (n143, n63);
buf  g98 (n193, n57);
not  g99 (n170, n62);
not  g100 (n192, n55);
buf  g101 (n124, n55);
not  g102 (n203, n43);
buf  g103 (n182, n36);
not  g104 (n119, n47);
buf  g105 (n228, n40);
not  g106 (n259, n73);
buf  g107 (n175, n63);
buf  g108 (n186, n53);
buf  g109 (n146, n50);
buf  g110 (n256, n74);
not  g111 (n204, n41);
buf  g112 (n248, n48);
buf  g113 (n247, n64);
not  g114 (n158, n69);
buf  g115 (n178, n74);
not  g116 (n221, n71);
buf  g117 (n196, n74);
buf  g118 (n128, n57);
buf  g119 (n260, n59);
not  g120 (n273, n66);
buf  g121 (n162, n45);
not  g122 (n250, n43);
buf  g123 (n263, n75);
not  g124 (n153, n67);
not  g125 (n202, n75);
buf  g126 (n223, n35);
not  g127 (n244, n38);
not  g128 (n293, n42);
buf  g129 (n218, n56);
not  g130 (n165, n37);
not  g131 (n206, n34);
not  g132 (n281, n40);
buf  g133 (n227, n44);
not  g134 (n230, n36);
buf  g135 (n171, n53);
buf  g136 (n144, n77);
not  g137 (n274, n42);
not  g138 (n145, n71);
not  g139 (n164, n63);
not  g140 (n131, n39);
not  g141 (n139, n72);
not  g142 (n138, n65);
buf  g143 (n199, n72);
not  g144 (n268, n45);
not  g145 (n147, n48);
not  g146 (n253, n46);
buf  g147 (n200, n47);
not  g148 (n127, n36);
buf  g149 (n246, n49);
buf  g150 (n217, n69);
buf  g151 (n135, n69);
not  g152 (n180, n38);
buf  g153 (n160, n52);
buf  g154 (n213, n47);
buf  g155 (n215, n54);
buf  g156 (n264, n65);
not  g157 (n185, n53);
buf  g158 (n262, n33);
not  g159 (n129, n68);
buf  g160 (n208, n61);
not  g161 (n212, n58);
buf  g162 (n149, n38);
not  g163 (n234, n45);
buf  g164 (n177, n50);
not  g165 (n214, n57);
not  g166 (n152, n46);
not  g167 (n132, n73);
buf  g168 (n181, n34);
not  g169 (n183, n74);
buf  g170 (n220, n34);
buf  g171 (n276, n40);
buf  g172 (n292, n63);
buf  g173 (n222, n49);
buf  g174 (n151, n33);
buf  g175 (n252, n56);
not  g176 (n195, n70);
not  g177 (n184, n76);
buf  g178 (n142, n60);
buf  g179 (n155, n61);
not  g180 (n122, n54);
buf  g181 (n271, n41);
not  g182 (n156, n65);
buf  g183 (n189, n39);
buf  g184 (n159, n72);
not  g185 (n279, n53);
not  g186 (n236, n44);
buf  g187 (n261, n51);
buf  g188 (n266, n44);
not  g189 (n201, n52);
buf  g190 (n205, n76);
not  g191 (n283, n66);
buf  g192 (n255, n37);
buf  g193 (n297, n50);
not  g194 (n290, n62);
not  g195 (n207, n71);
buf  g196 (n120, n35);
not  g197 (n284, n70);
buf  g198 (n148, n42);
buf  g199 (n157, n70);
not  g200 (n133, n51);
not  g201 (n278, n65);
not  g202 (n167, n60);
not  g203 (n211, n61);
not  g204 (n254, n66);
not  g205 (n225, n71);
buf  g206 (n123, n59);
buf  g207 (n229, n58);
buf  g208 (n237, n76);
not  g209 (n191, n66);
not  g210 (n251, n56);
buf  g211 (n277, n52);
not  g212 (n289, n77);
not  g213 (n187, n33);
not  g214 (n291, n55);
buf  g215 (n296, n36);
not  g216 (n197, n37);
not  g217 (n176, n51);
not  g218 (n241, n76);
buf  g219 (n219, n45);
not  g220 (n154, n57);
buf  g221 (n245, n50);
buf  g222 (n125, n59);
buf  g223 (n216, n60);
not  g224 (n161, n48);
not  g225 (n286, n75);
not  g226 (n280, n35);
buf  g227 (n269, n69);
buf  g228 (n121, n64);
not  g229 (n168, n42);
not  g230 (n249, n60);
buf  g231 (n258, n62);
buf  g232 (n194, n52);
buf  g233 (n265, n73);
buf  g234 (n130, n47);
buf  g235 (n136, n67);
buf  g236 (n173, n77);
buf  g237 (n275, n68);
not  g238 (n285, n55);
not  g239 (n235, n33);
not  g240 (n174, n58);
not  g241 (n287, n58);
not  g242 (n179, n56);
not  g243 (n190, n39);
buf  g244 (n233, n54);
not  g245 (n231, n64);
not  g246 (n267, n43);
not  g247 (n240, n61);
buf  g248 (n126, n73);
buf  g249 (n210, n41);
not  g250 (n295, n59);
not  g251 (n188, n37);
not  g252 (n272, n49);
not  g253 (n226, n40);
buf  g254 (n288, n43);
buf  g255 (n239, n41);
not  g256 (n294, n64);
not  g257 (n257, n75);
not  g258 (n270, n67);
buf  g259 (n166, n38);
buf  g260 (n140, n51);
buf  g261 (n224, n44);
buf  g262 (n134, n67);
not  g263 (n198, n54);
buf  g264 (n238, n68);
not  g265 (n302, n259);
not  g266 (n555, n160);
not  g267 (n316, n274);
not  g268 (n315, n166);
not  g269 (n359, n264);
not  g270 (n496, n194);
buf  g271 (n367, n261);
not  g272 (n509, n266);
buf  g273 (n401, n267);
buf  g274 (n567, n193);
not  g275 (n545, n174);
not  g276 (n331, n199);
not  g277 (n422, n213);
buf  g278 (n395, n263);
not  g279 (n369, n204);
not  g280 (n341, n276);
buf  g281 (n488, n264);
buf  g282 (n404, n219);
not  g283 (n571, n291);
buf  g284 (n343, n274);
buf  g285 (n423, n158);
buf  g286 (n410, n272);
buf  g287 (n531, n287);
not  g288 (n564, n292);
not  g289 (n500, n257);
not  g290 (n476, n273);
not  g291 (n510, n275);
buf  g292 (n480, n136);
not  g293 (n419, n138);
not  g294 (n346, n133);
not  g295 (n335, n269);
buf  g296 (n308, n134);
not  g297 (n319, n152);
buf  g298 (n578, n225);
not  g299 (n378, n263);
not  g300 (n455, n151);
not  g301 (n396, n256);
buf  g302 (n458, n271);
not  g303 (n533, n241);
buf  g304 (n324, n272);
buf  g305 (n390, n279);
buf  g306 (n358, n275);
not  g307 (n537, n263);
not  g308 (n575, n146);
not  g309 (n362, n248);
not  g310 (n321, n282);
buf  g311 (n393, n282);
buf  g312 (n377, n234);
not  g313 (n303, n252);
buf  g314 (n546, n232);
not  g315 (n351, n226);
not  g316 (n439, n171);
buf  g317 (n498, n282);
not  g318 (n322, n266);
buf  g319 (n492, n127);
buf  g320 (n364, n290);
not  g321 (n443, n242);
not  g322 (n317, n292);
buf  g323 (n483, n277);
buf  g324 (n549, n126);
not  g325 (n415, n235);
buf  g326 (n334, n164);
not  g327 (n327, n256);
not  g328 (n421, n265);
buf  g329 (n428, n150);
not  g330 (n583, n208);
not  g331 (n576, n195);
not  g332 (n445, n184);
not  g333 (n389, n285);
not  g334 (n543, n182);
not  g335 (n298, n200);
not  g336 (n536, n254);
buf  g337 (n357, n132);
not  g338 (n526, n217);
not  g339 (n552, n255);
not  g340 (n484, n287);
not  g341 (n352, n272);
buf  g342 (n407, n270);
buf  g343 (n425, n190);
not  g344 (n568, n220);
not  g345 (n508, n269);
not  g346 (n414, n264);
not  g347 (n538, n212);
buf  g348 (n311, n288);
buf  g349 (n363, n180);
not  g350 (n465, n163);
not  g351 (n519, n144);
not  g352 (n332, n291);
buf  g353 (n547, n266);
not  g354 (n548, n250);
not  g355 (n350, n161);
buf  g356 (n456, n211);
not  g357 (n444, n222);
not  g358 (n386, n279);
not  g359 (n562, n268);
not  g360 (n521, n280);
buf  g361 (n482, n267);
buf  g362 (n345, n215);
not  g363 (n307, n276);
buf  g364 (n540, n196);
buf  g365 (n323, n145);
buf  g366 (n494, n187);
buf  g367 (n318, n256);
not  g368 (n513, n272);
not  g369 (n541, n261);
buf  g370 (n398, n262);
not  g371 (n330, n246);
buf  g372 (n372, n262);
not  g373 (n581, n261);
buf  g374 (n418, n277);
buf  g375 (n512, n287);
buf  g376 (n473, n269);
buf  g377 (n557, n273);
buf  g378 (n577, n256);
not  g379 (n544, n153);
not  g380 (n355, n178);
not  g381 (n515, n276);
buf  g382 (n388, n189);
not  g383 (n551, n277);
buf  g384 (n329, n121);
buf  g385 (n374, n125);
not  g386 (n481, n279);
not  g387 (n313, n289);
buf  g388 (n520, n282);
not  g389 (n559, n259);
buf  g390 (n470, n284);
not  g391 (n522, n147);
not  g392 (n493, n257);
buf  g393 (n347, n175);
not  g394 (n572, n283);
not  g395 (n495, n201);
buf  g396 (n530, n293);
buf  g397 (n447, n188);
not  g398 (n527, n286);
buf  g399 (n382, n271);
buf  g400 (n349, n244);
not  g401 (n460, n284);
buf  g402 (n457, n142);
not  g403 (n504, n274);
not  g404 (n475, n286);
not  g405 (n365, n270);
buf  g406 (n429, n139);
buf  g407 (n535, n224);
not  g408 (n394, n245);
not  g409 (n333, n261);
not  g410 (n477, n249);
buf  g411 (n400, n230);
buf  g412 (n406, n185);
buf  g413 (n381, n172);
not  g414 (n342, n258);
not  g415 (n437, n262);
buf  g416 (n325, n165);
not  g417 (n405, n198);
not  g418 (n353, n280);
buf  g419 (n474, n216);
buf  g420 (n497, n238);
buf  g421 (n573, n169);
not  g422 (n397, n237);
not  g423 (n556, n258);
not  g424 (n517, n260);
not  g425 (n542, n271);
not  g426 (n469, n168);
buf  g427 (n301, n278);
not  g428 (n448, n281);
buf  g429 (n574, n275);
not  g430 (n501, n271);
not  g431 (n487, n285);
not  g432 (n340, n289);
not  g433 (n507, n130);
buf  g434 (n503, n197);
buf  g435 (n464, n231);
not  g436 (n408, n119);
buf  g437 (n385, n257);
not  g438 (n499, n131);
buf  g439 (n360, n278);
buf  g440 (n413, n183);
not  g441 (n454, n154);
not  g442 (n471, n203);
buf  g443 (n561, n283);
buf  g444 (n361, n287);
not  g445 (n433, n290);
not  g446 (n304, n291);
buf  g447 (n514, n124);
buf  g448 (n370, n273);
buf  g449 (n441, n157);
buf  g450 (n305, n240);
not  g451 (n534, n191);
not  g452 (n384, n265);
not  g453 (n339, n275);
buf  g454 (n468, n283);
not  g455 (n579, n202);
buf  g456 (n452, n258);
buf  g457 (n326, n260);
buf  g458 (n449, n159);
buf  g459 (n336, n292);
buf  g460 (n434, n262);
not  g461 (n344, n143);
buf  g462 (n430, n268);
not  g463 (n461, n278);
not  g464 (n417, n288);
buf  g465 (n320, n284);
not  g466 (n442, n274);
buf  g467 (n523, n167);
not  g468 (n467, n277);
buf  g469 (n354, n290);
buf  g470 (n424, n279);
not  g471 (n565, n264);
buf  g472 (n314, n156);
not  g473 (n373, n267);
buf  g474 (n511, n290);
not  g475 (n462, n206);
not  g476 (n582, n192);
buf  g477 (n516, n283);
buf  g478 (n402, n268);
not  g479 (n554, n135);
not  g480 (n356, n181);
buf  g481 (n309, n276);
not  g482 (n485, n247);
not  g483 (n478, n236);
buf  g484 (n506, n269);
not  g485 (n420, n259);
buf  g486 (n306, n148);
buf  g487 (n524, n260);
buf  g488 (n532, n289);
not  g489 (n489, n278);
buf  g490 (n399, n288);
buf  g491 (n529, n284);
not  g492 (n463, n141);
buf  g493 (n392, n286);
not  g494 (n375, n285);
buf  g495 (n348, n162);
not  g496 (n432, n122);
buf  g497 (n438, n265);
buf  g498 (n376, n267);
buf  g499 (n558, n209);
not  g500 (n436, n258);
not  g501 (n440, n280);
not  g502 (n391, n289);
not  g503 (n379, n292);
not  g504 (n337, n229);
not  g505 (n409, n155);
buf  g506 (n371, n228);
not  g507 (n310, n129);
not  g508 (n490, n281);
buf  g509 (n380, n173);
buf  g510 (n412, n281);
buf  g511 (n569, n207);
not  g512 (n387, n280);
not  g513 (n560, n281);
buf  g514 (n426, n218);
buf  g515 (n472, n286);
not  g516 (n505, n273);
buf  g517 (n580, n239);
buf  g518 (n416, n214);
not  g519 (n466, n243);
buf  g520 (n525, n137);
not  g521 (n563, n170);
not  g522 (n450, n266);
buf  g523 (n431, n186);
buf  g524 (n312, n140);
buf  g525 (n479, n223);
buf  g526 (n553, n288);
not  g527 (n486, n179);
not  g528 (n491, n128);
buf  g529 (n459, n265);
buf  g530 (n453, n268);
not  g531 (n566, n285);
not  g532 (n338, n221);
buf  g533 (n299, n176);
buf  g534 (n427, n233);
not  g535 (n502, n270);
not  g536 (n328, n263);
not  g537 (n518, n251);
not  g538 (n383, n177);
buf  g539 (n528, n253);
not  g540 (n368, n259);
buf  g541 (n435, n227);
buf  g542 (n451, n120);
buf  g543 (n403, n270);
buf  g544 (n570, n205);
not  g545 (n300, n149);
buf  g546 (n550, n260);
buf  g547 (n366, n210);
not  g548 (n539, n291);
buf  g549 (n411, n123);
buf  g550 (n446, n257);
buf  g551 (n616, n333);
buf  g552 (n609, n308);
buf  g553 (n624, n327);
not  g554 (n618, n348);
buf  g555 (n645, n359);
not  g556 (n593, n331);
buf  g557 (n622, n324);
buf  g558 (n617, n311);
not  g559 (n628, n319);
not  g560 (n646, n316);
not  g561 (n637, n332);
buf  g562 (n640, n361);
buf  g563 (n607, n306);
not  g564 (n601, n350);
buf  g565 (n627, n337);
buf  g566 (n610, n339);
not  g567 (n633, n307);
buf  g568 (n625, n347);
not  g569 (n634, n355);
buf  g570 (n591, n360);
buf  g571 (n600, n330);
buf  g572 (n619, n349);
not  g573 (n636, n321);
buf  g574 (n613, n336);
buf  g575 (n629, n303);
not  g576 (n635, n342);
buf  g577 (n588, n343);
not  g578 (n596, n313);
buf  g579 (n595, n358);
not  g580 (n602, n299);
not  g581 (n639, n312);
buf  g582 (n586, n325);
buf  g583 (n604, n329);
not  g584 (n620, n300);
not  g585 (n585, n326);
buf  g586 (n611, n310);
not  g587 (n608, n314);
not  g588 (n597, n335);
buf  g589 (n647, n315);
not  g590 (n642, n340);
buf  g591 (n598, n352);
buf  g592 (n615, n346);
buf  g593 (n641, n338);
buf  g594 (n612, n357);
not  g595 (n631, n341);
not  g596 (n594, n328);
buf  g597 (n643, n317);
buf  g598 (n606, n334);
buf  g599 (n605, n304);
buf  g600 (n590, n351);
buf  g601 (n587, n322);
buf  g602 (n603, n305);
not  g603 (n638, n318);
not  g604 (n584, n301);
buf  g605 (n626, n354);
buf  g606 (n592, n345);
not  g607 (n599, n356);
buf  g608 (n621, n298);
buf  g609 (n614, n320);
buf  g610 (n630, n323);
buf  g611 (n623, n344);
not  g612 (n644, n353);
buf  g613 (n589, n309);
buf  g614 (n632, n302);
buf  g615 (n658, n587);
not  g616 (n659, n599);
not  g617 (n650, n597);
not  g618 (n674, n599);
not  g619 (n649, n591);
buf  g620 (n666, n597);
not  g621 (n667, n592);
buf  g622 (n648, n593);
buf  g623 (n668, n584);
not  g624 (n677, n596);
not  g625 (n665, n585);
buf  g626 (n669, n598);
not  g627 (n673, n595);
buf  g628 (n661, n596);
buf  g629 (n652, n597);
buf  g630 (n664, n597);
not  g631 (n670, n589);
not  g632 (n662, n586);
buf  g633 (n653, n599);
buf  g634 (n654, n600);
not  g635 (n671, n595);
not  g636 (n663, n588);
not  g637 (n675, n599);
not  g638 (n655, n598);
buf  g639 (n676, n598);
not  g640 (n651, n596);
not  g641 (n656, n590);
not  g642 (n672, n598);
buf  g643 (n657, n594);
buf  g644 (n660, n596);
nor  g645 (n729, n26, n398, n458, n441);
and  g646 (n683, n365, n380, n651, n409);
nor  g647 (n687, n482, n454, n384, n455);
and  g648 (n726, n30, n665, n25, n666);
or   g649 (n696, n435, n28, n29, n432);
nor  g650 (n711, n464, n427, n470, n367);
and  g651 (n698, n658, n481, n668, n394);
nor  g652 (n715, n667, n376, n418, n26);
xor  g653 (n704, n32, n450, n392, n404);
or   g654 (n721, n661, n662, n421, n461);
or   g655 (n731, n28, n370, n456, n663);
or   g656 (n682, n467, n665, n438, n22);
or   g657 (n680, n476, n660, n24, n433);
and  g658 (n679, n420, n668, n452, n661);
xnor g659 (n690, n480, n664, n24, n31);
and  g660 (n697, n652, n32, n414, n25);
nor  g661 (n691, n664, n663, n406, n373);
or   g662 (n727, n666, n419, n29, n483);
nor  g663 (n725, n366, n449, n402, n408);
or   g664 (n681, n473, n29, n665, n417);
xor  g665 (n706, n428, n23, n386, n375);
nor  g666 (n700, n654, n478, n383, n405);
or   g667 (n699, n388, n451, n660, n391);
xor  g668 (n730, n400, n393, n649, n474);
xnor g669 (n689, n442, n443, n410, n378);
nor  g670 (n684, n379, n371, n377, n466);
nand g671 (n707, n436, n31, n656, n445);
and  g672 (n716, n662, n413, n660, n430);
and  g673 (n724, n30, n477, n440, n23);
nand g674 (n723, n659, n664, n25, n471);
xnor g675 (n694, n653, n395, n23, n368);
nand g676 (n710, n479, n668, n27, n667);
and  g677 (n693, n661, n28, n659, n24);
nor  g678 (n718, n658, n22, n27, n659);
xor  g679 (n695, n389, n364, n472, n484);
xnor g680 (n678, n469, n666, n667, n363);
nor  g681 (n701, n403, n439, n385, n663);
nand g682 (n708, n669, n666, n659, n457);
and  g683 (n709, n663, n369, n426, n30);
or   g684 (n686, n423, n669, n650, n381);
xor  g685 (n728, n668, n416, n429, n434);
nand g686 (n720, n27, n655, n397, n453);
or   g687 (n703, n372, n660, n648, n448);
xor  g688 (n722, n28, n669, n657, n437);
and  g689 (n688, n665, n412, n465, n459);
xor  g690 (n713, n444, n390, n431, n382);
nand g691 (n732, n387, n475, n26, n463);
xnor g692 (n705, n23, n32, n30);
nor  g693 (n719, n462, n399, n31, n446);
xor  g694 (n717, n407, n29, n422, n662);
and  g695 (n714, n26, n25, n460, n425);
xnor g696 (n702, n415, n661, n447, n662);
nand g697 (n712, n664, n27, n411, n401);
nor  g698 (n685, n424, n24, n396, n362);
or   g699 (n692, n468, n31, n667, n374);
nand g700 (n775, n97, n95, n81, n688);
nand g701 (n748, n702, n86, n687, n689);
xor  g702 (n759, n697, n90, n95, n91);
and  g703 (n747, n708, n707, n98, n700);
xor  g704 (n740, n85, n90, n698, n94);
or   g705 (n767, n678, n698, n79, n687);
nand g706 (n769, n699, n96, n98, n707);
or   g707 (n754, n78, n694, n686, n89);
xnor g708 (n749, n92, n81, n701, n686);
xnor g709 (n772, n697, n692, n79, n91);
nor  g710 (n771, n693, n696, n79, n94);
nor  g711 (n745, n693, n92, n94, n690);
or   g712 (n739, n97, n695, n91, n77);
xor  g713 (n742, n82, n691, n80, n81);
and  g714 (n757, n699, n84, n86, n691);
xor  g715 (n744, n687, n82, n696, n87);
or   g716 (n773, n81, n704, n705, n91);
or   g717 (n750, n97, n689, n86, n679);
or   g718 (n763, n700, n87, n685, n705);
nand g719 (n761, n705, n80, n89);
and  g720 (n743, n92, n97, n98, n84);
xnor g721 (n736, n85, n706, n80, n695);
or   g722 (n776, n701, n90, n96, n694);
xor  g723 (n779, n86, n88, n691, n702);
xnor g724 (n778, n696, n78, n84, n682);
or   g725 (n735, n90, n83, n708, n87);
nand g726 (n738, n88, n702, n706, n701);
xor  g727 (n777, n95, n95, n87, n93);
xnor g728 (n770, n697, n78, n703, n93);
nand g729 (n768, n685, n693, n692, n707);
or   g730 (n766, n690, n79, n93, n695);
nand g731 (n774, n690, n89, n684, n85);
xnor g732 (n746, n88, n680, n699, n85);
xor  g733 (n737, n704, n88, n688, n701);
or   g734 (n758, n707, n94, n697, n693);
or   g735 (n752, n99, n686, n690, n96);
nand g736 (n762, n600, n696, n703, n93);
xor  g737 (n760, n83, n84, n82, n78);
xor  g738 (n741, n83, n699, n689, n698);
and  g739 (n755, n687, n691, n703, n688);
or   g740 (n753, n99, n689, n694, n82);
xor  g741 (n734, n692, n700, n704, n703);
nor  g742 (n756, n694, n681, n695, n692);
nor  g743 (n765, n83, n92, n706, n96);
or   g744 (n733, n702, n686, n698, n704);
and  g745 (n751, n705, n688, n89, n706);
xnor g746 (n764, n683, n700, n98, n600);
xor  g747 (n787, n605, n607, n604, n601);
nand g748 (n783, n763, n293, n760);
xor  g749 (n790, n297, n607, n709, n766);
xnor g750 (n797, n770, n602, n710, n295);
xnor g751 (n794, n601, n709, n710, n711);
nand g752 (n789, n755, n294, n606, n602);
xor  g753 (n798, n294, n709, n711, n603);
xor  g754 (n799, n757, n294, n710);
xor  g755 (n781, n762, n295, n603, n605);
or   g756 (n786, n297, n296, n604, n772);
and  g757 (n785, n605, n708, n754, n709);
and  g758 (n793, n603, n293, n296, n602);
or   g759 (n780, n765, n761, n297, n759);
nor  g760 (n791, n602, n601, n603, n771);
or   g761 (n792, n296, n604, n756, n295);
and  g762 (n788, n606, n604, n601, n758);
nor  g763 (n796, n296, n768, n764, n773);
nand g764 (n795, n769, n605, n295, n607);
and  g765 (n784, n600, n294, n607, n708);
xnor g766 (n782, n606, n606, n297, n767);
xnor g767 (n802, n549, n555, n792, n783);
and  g768 (n807, n560, n541, n556, n531);
nor  g769 (n801, n559, n505, n519, n523);
and  g770 (n819, n506, n542, n500, n522);
or   g771 (n820, n503, n543, n711, n547);
or   g772 (n806, n791, n540, n784, n495);
nand g773 (n817, n497, n535, n537, n780);
nor  g774 (n800, n538, n533, n510, n790);
xor  g775 (n815, n791, n554, n485, n496);
nand g776 (n824, n498, n787, n504, n552);
xor  g777 (n803, n544, n507, n527, n550);
nor  g778 (n805, n539, n509, n789, n516);
and  g779 (n812, n524, n532, n515, n790);
xor  g780 (n825, n488, n712, n781, n526);
xor  g781 (n810, n513, n521, n551, n512);
or   g782 (n811, n490, n782, n712, n557);
or   g783 (n809, n502, n530, n786, n514);
nor  g784 (n826, n791, n499, n493, n789);
nand g785 (n823, n791, n790, n789, n494);
xnor g786 (n822, n788, n487, n711, n534);
xnor g787 (n813, n545, n520, n792, n536);
xnor g788 (n816, n712, n787, n528, n788);
nor  g789 (n821, n789, n501, n517, n529);
xnor g790 (n804, n792, n548, n492, n558);
and  g791 (n814, n491, n790, n792, n525);
and  g792 (n818, n553, n486, n511, n785);
or   g793 (n808, n546, n508, n489, n518);
not  g794 (n830, n818);
buf  g795 (n836, n608);
not  g796 (n840, n609);
buf  g797 (n847, n812);
not  g798 (n835, n806);
buf  g799 (n833, n805);
not  g800 (n828, n807);
not  g801 (n832, n813);
buf  g802 (n827, n610);
buf  g803 (n846, n815);
not  g804 (n850, n822);
buf  g805 (n838, n816);
buf  g806 (n843, n811);
buf  g807 (n837, n810);
buf  g808 (n829, n801);
buf  g809 (n848, n610);
not  g810 (n842, n809);
buf  g811 (n839, n608);
buf  g812 (n845, n808);
buf  g813 (n841, n814);
and  g814 (n834, n610, n802, n817, n803);
or   g815 (n844, n610, n823, n804, n820);
and  g816 (n849, n819, n821, n608, n609);
nand g817 (n831, n800, n608, n609);
xor  g818 (n858, n566, n721);
and  g819 (n852, n612, n564);
nor  g820 (n936, n612, n836, n832, n619);
or   g821 (n902, n639, n848, n614, n846);
xnor g822 (n938, n840, n634, n847, n844);
or   g823 (n914, n794, n632, n672, n842);
xor  g824 (n860, n568, n799, n716, n640);
xnor g825 (n886, n799, n616, n674, n719);
xor  g826 (n923, n831, n828, n625, n633);
and  g827 (n911, n622, n716, n844, n717);
xnor g828 (n888, n614, n673, n675, n616);
xor  g829 (n865, n798, n574, n577, n718);
nand g830 (n929, n623, n619, n632, n725);
nand g831 (n855, n629, n715, n621, n620);
or   g832 (n916, n837, n635, n638, n726);
and  g833 (n900, n615, n846, n628, n834);
xnor g834 (n935, n831, n674, n620, n617);
and  g835 (n862, n845, n836, n674, n614);
nor  g836 (n878, n724, n570, n841, n670);
xor  g837 (n875, n846, n794, n676, n848);
xor  g838 (n895, n843, n840, n617, n572);
xor  g839 (n925, n828, n845, n576, n847);
nor  g840 (n941, n578, n672, n842, n675);
xnor g841 (n937, n641, n631, n848, n629);
xor  g842 (n861, n631, n830, n718, n617);
or   g843 (n920, n842, n611, n672, n563);
xnor g844 (n879, n630, n720, n799, n562);
xnor g845 (n898, n627, n835, n722, n828);
xnor g846 (n868, n712, n793, n637, n721);
xnor g847 (n896, n674, n832, n833, n713);
or   g848 (n870, n101, n671, n835);
xor  g849 (n921, n677, n621, n633, n640);
and  g850 (n857, n841, n841, n613, n845);
nor  g851 (n871, n722, n627, n673, n677);
nand g852 (n910, n834, n642, n717, n845);
or   g853 (n851, n638, n796, n636, n613);
nand g854 (n881, n617, n793, n641, n796);
or   g855 (n872, n624, n638, n726, n794);
and  g856 (n905, n628, n838, n626, n621);
nor  g857 (n913, n673, n846, n832, n100);
and  g858 (n931, n632, n633, n628, n840);
xnor g859 (n928, n839, n641, n636, n642);
or   g860 (n891, n616, n848, n724, n676);
nor  g861 (n934, n834, n722, n843, n828);
nand g862 (n932, n839, n714, n670, n720);
nor  g863 (n899, n844, n626, n723, n575);
xnor g864 (n924, n849, n795, n671, n639);
or   g865 (n893, n623, n796, n850, n673);
nand g866 (n880, n718, n615, n849, n619);
xor  g867 (n892, n637, n795, n831, n99);
and  g868 (n942, n677, n850, n720, n582);
nor  g869 (n853, n672, n621, n849, n797);
xnor g870 (n890, n629, n640, n571, n624);
and  g871 (n906, n622, n631, n794, n625);
nor  g872 (n856, n716, n723, n626, n847);
and  g873 (n922, n837, n618, n713, n714);
xor  g874 (n926, n727, n642, n849, n829);
nor  g875 (n907, n716, n629, n721, n623);
nor  g876 (n854, n714, n634, n630, n622);
xor  g877 (n915, n625, n635, n638, n723);
nor  g878 (n864, n715, n834, n827, n632);
xor  g879 (n877, n833, n639, n724, n827);
and  g880 (n882, n830, n613, n796, n618);
xor  g881 (n889, n713, n99, n850, n630);
and  g882 (n919, n798, n832, n623, n634);
nor  g883 (n887, n627, n569, n714, n612);
or   g884 (n912, n831, n611, n615, n850);
and  g885 (n930, n625, n612, n100, n627);
xor  g886 (n908, n836, n719, n830, n725);
nor  g887 (n944, n833, n622, n829, n100);
nor  g888 (n918, n641, n726, n626, n573);
and  g889 (n939, n636, n567, n799, n797);
nor  g890 (n897, n620, n624, n671, n615);
or   g891 (n884, n634, n793, n677, n636);
xnor g892 (n866, n725, n620, n727, n675);
or   g893 (n909, n829, n842, n843, n635);
and  g894 (n885, n639, n613, n713, n725);
xor  g895 (n943, n637, n841, n721, n840);
or   g896 (n883, n793, n628, n611, n614);
nand g897 (n933, n797, n795, n836, n838);
and  g898 (n901, n724, n676, n795, n835);
and  g899 (n940, n839, n833, n581, n637);
and  g900 (n863, n838, n669, n797, n642);
nor  g901 (n917, n726, n670, n830, n619);
or   g902 (n859, n565, n618, n640, n722);
and  g903 (n873, n670, n847, n839, n837);
or   g904 (n903, n838, n843, n844, n580);
xor  g905 (n869, n100, n676, n719, n723);
and  g906 (n927, n616, n618, n837, n579);
or   g907 (n876, n718, n631, n715, n624);
xnor g908 (n904, n798, n630, n675, n829);
or   g909 (n874, n720, n717, n633, n719);
nor  g910 (n867, n611, n635, n717, n101);
and  g911 (n894, n798, n715, n561, n835);
not  g912 (n945, n858);
buf  g913 (n946, n854);
not  g914 (n954, n727);
buf  g915 (n947, n855);
buf  g916 (n950, n859);
buf  g917 (n948, n852);
buf  g918 (n953, n857);
not  g919 (n951, n727);
not  g920 (n952, n856);
xnor g921 (n949, n860, n851, n853);
nor  g922 (n966, n645, n947, n730, n946);
xnor g923 (n974, n644, n110, n105, n108);
xnor g924 (n973, n729, n117, n105, n948);
xor  g925 (n981, n730, n103, n107, n104);
nor  g926 (n979, n950, n107, n949, n948);
or   g927 (n989, n115, n111, n950, n103);
nand g928 (n983, n728, n646, n949, n643);
nor  g929 (n955, n102, n104, n113);
nor  g930 (n991, n108, n106, n643, n647);
or   g931 (n980, n118, n112, n111, n946);
xor  g932 (n984, n948, n117, n107, n728);
nor  g933 (n960, n953, n102, n644);
xnor g934 (n978, n646, n949, n116);
nor  g935 (n965, n646, n947, n729, n775);
nand g936 (n971, n105, n107, n948, n952);
or   g937 (n987, n777, n950, n114, n104);
or   g938 (n957, n954, n109, n108, n952);
xor  g939 (n962, n645, n111, n114, n947);
nand g940 (n990, n106, n951, n731);
nand g941 (n982, n731, n113, n103, n952);
nand g942 (n967, n774, n954, n946, n729);
nand g943 (n970, n945, n111, n731, n112);
xor  g944 (n988, n647, n118, n779, n953);
or   g945 (n969, n116, n108, n106, n101);
xor  g946 (n976, n110, n728, n117, n954);
or   g947 (n985, n115, n110, n101, n949);
xnor g948 (n968, n954, n730, n109, n118);
nand g949 (n986, n113, n730, n112, n109);
or   g950 (n959, n953, n114, n946, n646);
xor  g951 (n964, n114, n109, n729, n644);
and  g952 (n977, n110, n643, n951, n947);
nand g953 (n956, n102, n103, n644, n113);
xor  g954 (n961, n950, n952, n117, n778);
or   g955 (n972, n105, n106, n115);
xnor g956 (n963, n116, n112, n953, n643);
xor  g957 (n958, n645, n951, n776, n731);
nor  g958 (n975, n645, n647, n728);
xor  g959 (n996, n732, n975, n960, n963);
xor  g960 (n992, n912, n900, n932, n918);
or   g961 (n1013, n902, n940, n890, n982);
xor  g962 (n1006, n898, n882, n583, n961);
or   g963 (n1017, n732, n910, n985, n892);
xnor g964 (n1011, n916, n894, n964, n974);
xnor g965 (n1018, n965, n938, n939, n906);
nand g966 (n1010, n970, n862, n891, n986);
nand g967 (n1009, n929, n958, n887, n903);
and  g968 (n1005, n899, n914, n959, n927);
nor  g969 (n999, n880, n989, n864, n981);
nor  g970 (n1020, n878, n926, n913, n941);
or   g971 (n1012, n978, n872, n943, n922);
nor  g972 (n1004, n583, n920, n930, n935);
xnor g973 (n1021, n869, n988, n921, n861);
xor  g974 (n998, n908, n917, n972, n934);
and  g975 (n1016, n968, n889, n937, n990);
xnor g976 (n993, n911, n886, n871, n944);
nand g977 (n1002, n969, n732, n919, n987);
nor  g978 (n1003, n883, n955, n866, n976);
nor  g979 (n994, n973, n896, n925, n881);
nor  g980 (n1007, n909, n924, n991, n867);
xnor g981 (n1015, n983, n868, n984, n876);
nor  g982 (n1001, n732, n865, n888, n933);
nor  g983 (n997, n863, n956, n877, n875);
or   g984 (n1000, n879, n923, n897, n971);
or   g985 (n1014, n870, n967, n901, n966);
and  g986 (n1008, n942, n907, n931, n118);
or   g987 (n1022, n928, n905, n979, n873);
xnor g988 (n1023, n915, n895, n962, n893);
nor  g989 (n995, n874, n980, n904, n936);
nand g990 (n1019, n884, n885, n957, n977);
xor  g991 (n1027, n1012, n995, n826, n1020);
xnor g992 (n1032, n1008, n1010, n997, n1004);
nor  g993 (n1024, n1009, n1015, n1000, n1023);
nor  g994 (n1030, n1016, n993, n1007, n1021);
xor  g995 (n1029, n1014, n998, n1017, n1006);
and  g996 (n1028, n1001, n1018, n1002, n1005);
or   g997 (n1026, n1003, n826, n1011, n994);
nand g998 (n1031, n996, n992, n1019, n1013);
xnor g999 (n1025, n825, n999, n1022, n824);
endmodule
