// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_102 written by SynthGen on 2021/04/05 11:08:33
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_102 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n497, n1009, n1032, n1007, n1003, n1010, n1013, n1011,
 n1028, n1025, n1005, n1016, n1031, n1012, n1015, n1027,
 n1019, n1014, n1023, n1020, n1002, n1008, n1024, n1029,
 n1021, n1004, n1022, n1017, n1006, n1026, n1018, n1030);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n497, n1009, n1032, n1007, n1003, n1010, n1013, n1011,
 n1028, n1025, n1005, n1016, n1031, n1012, n1015, n1027,
 n1019, n1014, n1023, n1020, n1002, n1008, n1024, n1029,
 n1021, n1004, n1022, n1017, n1006, n1026, n1018, n1030;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001;

buf  g0 (n69, n12);
not  g1 (n49, n16);
buf  g2 (n39, n14);
buf  g3 (n33, n22);
not  g4 (n59, n12);
buf  g5 (n53, n17);
not  g6 (n48, n20);
not  g7 (n63, n25);
not  g8 (n74, n8);
buf  g9 (n52, n7);
not  g10 (n76, n28);
buf  g11 (n41, n25);
buf  g12 (n62, n11);
buf  g13 (n46, n6);
not  g14 (n60, n30);
buf  g15 (n64, n24);
buf  g16 (n58, n7);
not  g17 (n75, n18);
not  g18 (n40, n23);
not  g19 (n35, n26);
not  g20 (n54, n27);
not  g21 (n34, n23);
buf  g22 (n37, n19);
buf  g23 (n51, n25);
not  g24 (n86, n28);
buf  g25 (n47, n30);
buf  g26 (n77, n3);
not  g27 (n85, n9);
not  g28 (n50, n19);
buf  g29 (n42, n10);
buf  g30 (n72, n14);
and  g31 (n71, n21, n24);
or   g32 (n65, n1, n26, n13);
nor  g33 (n83, n3, n20, n16, n18);
xor  g34 (n68, n6, n14, n21, n17);
and  g35 (n43, n27, n20, n13);
or   g36 (n56, n29, n7);
xor  g37 (n78, n26, n15, n18);
xor  g38 (n55, n17, n20, n26, n10);
xor  g39 (n38, n16, n22, n14, n12);
xor  g40 (n61, n8, n1, n30, n16);
xor  g41 (n36, n8, n4, n5);
xnor g42 (n67, n2, n3, n29, n4);
xor  g43 (n84, n1, n23, n29, n5);
nand g44 (n66, n12, n24, n18, n15);
or   g45 (n44, n4, n10, n19, n2);
and  g46 (n70, n11, n22, n8, n28);
xor  g47 (n82, n22, n15, n23, n28);
nand g48 (n81, n6, n6, n9, n1);
nor  g49 (n80, n5, n31, n11, n21);
xnor g50 (n73, n10, n27, n19, n9);
xnor g51 (n45, n11, n27, n17, n21);
nor  g52 (n79, n25, n24, n2, n9);
xnor g53 (n57, n3, n2, n4, n30);
buf  g54 (n92, n70);
buf  g55 (n136, n61);
buf  g56 (n222, n81);
buf  g57 (n232, n59);
not  g58 (n87, n66);
not  g59 (n124, n62);
buf  g60 (n211, n39);
buf  g61 (n158, n63);
buf  g62 (n190, n65);
buf  g63 (n157, n50);
buf  g64 (n116, n43);
not  g65 (n128, n68);
buf  g66 (n105, n69);
not  g67 (n97, n64);
not  g68 (n206, n77);
not  g69 (n208, n64);
not  g70 (n242, n63);
buf  g71 (n171, n74);
not  g72 (n160, n80);
buf  g73 (n189, n86);
not  g74 (n145, n82);
not  g75 (n112, n62);
buf  g76 (n235, n39);
buf  g77 (n108, n75);
not  g78 (n229, n74);
not  g79 (n178, n41);
buf  g80 (n238, n41);
buf  g81 (n88, n36);
buf  g82 (n103, n65);
buf  g83 (n164, n76);
not  g84 (n91, n35);
buf  g85 (n197, n44);
buf  g86 (n114, n59);
not  g87 (n90, n53);
not  g88 (n224, n80);
buf  g89 (n153, n57);
buf  g90 (n241, n44);
not  g91 (n95, n83);
not  g92 (n161, n62);
buf  g93 (n111, n44);
not  g94 (n94, n73);
buf  g95 (n188, n49);
buf  g96 (n155, n56);
not  g97 (n173, n52);
not  g98 (n228, n84);
buf  g99 (n148, n31);
buf  g100 (n202, n60);
buf  g101 (n130, n60);
buf  g102 (n89, n85);
not  g103 (n193, n55);
not  g104 (n126, n45);
buf  g105 (n101, n53);
not  g106 (n156, n55);
not  g107 (n205, n84);
not  g108 (n107, n80);
buf  g109 (n175, n71);
buf  g110 (n100, n78);
not  g111 (n187, n50);
buf  g112 (n249, n69);
buf  g113 (n123, n37);
not  g114 (n110, n56);
buf  g115 (n137, n48);
not  g116 (n220, n33);
not  g117 (n98, n31);
not  g118 (n198, n72);
not  g119 (n201, n46);
buf  g120 (n106, n33);
buf  g121 (n217, n85);
buf  g122 (n183, n59);
not  g123 (n179, n83);
not  g124 (n247, n37);
buf  g125 (n199, n35);
buf  g126 (n237, n55);
not  g127 (n104, n67);
not  g128 (n162, n67);
not  g129 (n109, n54);
buf  g130 (n163, n54);
buf  g131 (n218, n38);
buf  g132 (n236, n41);
buf  g133 (n144, n86);
not  g134 (n172, n84);
not  g135 (n125, n82);
not  g136 (n233, n61);
buf  g137 (n182, n67);
buf  g138 (n200, n51);
buf  g139 (n150, n47);
buf  g140 (n196, n79);
buf  g141 (n239, n68);
buf  g142 (n133, n65);
not  g143 (n119, n42);
not  g144 (n118, n34);
buf  g145 (n165, n53);
buf  g146 (n231, n56);
not  g147 (n115, n70);
buf  g148 (n230, n71);
buf  g149 (n140, n57);
buf  g150 (n176, n79);
buf  g151 (n210, n71);
buf  g152 (n243, n76);
not  g153 (n121, n48);
not  g154 (n99, n69);
not  g155 (n143, n77);
buf  g156 (n141, n69);
not  g157 (n147, n82);
not  g158 (n240, n38);
not  g159 (n191, n54);
buf  g160 (n209, n37);
buf  g161 (n168, n79);
not  g162 (n127, n66);
buf  g163 (n154, n83);
buf  g164 (n120, n61);
buf  g165 (n135, n81);
buf  g166 (n223, n49);
buf  g167 (n166, n71);
buf  g168 (n177, n48);
not  g169 (n93, n38);
buf  g170 (n227, n81);
not  g171 (n169, n60);
buf  g172 (n134, n62);
not  g173 (n234, n51);
buf  g174 (n113, n55);
not  g175 (n167, n47);
not  g176 (n213, n52);
buf  g177 (n244, n48);
not  g178 (n152, n32);
buf  g179 (n203, n57);
buf  g180 (n159, n35);
buf  g181 (n151, n60);
not  g182 (n207, n34);
not  g183 (n214, n36);
not  g184 (n181, n72);
buf  g185 (n146, n38);
buf  g186 (n184, n64);
buf  g187 (n138, n42);
not  g188 (n132, n85);
buf  g189 (n250, n51);
buf  g190 (n245, n67);
buf  g191 (n225, n39);
buf  g192 (n221, n73);
buf  g193 (n129, n47);
buf  g194 (n212, n58);
not  g195 (n117, n58);
buf  g196 (n219, n75);
not  g197 (n246, n73);
not  g198 (n186, n31);
xnor g199 (n174, n82, n34);
and  g200 (n122, n61, n33, n74, n41);
xor  g201 (n192, n50, n75, n81, n46);
or   g202 (n194, n77, n43, n64, n54);
or   g203 (n149, n45, n70, n50, n85);
or   g204 (n226, n63, n35, n72, n68);
and  g205 (n180, n77, n57, n65, n74);
xnor g206 (n216, n43, n36, n66, n40);
and  g207 (n96, n52, n46, n49, n42);
nor  g208 (n248, n44, n40, n53, n80);
or   g209 (n195, n59, n49, n75, n39);
xnor g210 (n131, n52, n40, n66);
or   g211 (n215, n78, n37, n70, n51);
nor  g212 (n139, n72, n83, n36, n43);
and  g213 (n142, n76, n42, n56, n73);
xor  g214 (n102, n76, n46, n68, n34);
nor  g215 (n170, n84, n78, n47);
xor  g216 (n204, n33, n58, n45);
or   g217 (n185, n79, n32, n63, n58);
nor  g218 (n399, n193, n161, n247, n195);
or   g219 (n298, n232, n198, n87, n228);
xor  g220 (n326, n88, n239, n173, n102);
nor  g221 (n392, n206, n180, n170, n150);
nor  g222 (n322, n101, n91, n104, n135);
or   g223 (n373, n93, n198, n138, n112);
xnor g224 (n334, n182, n227, n194, n196);
xnor g225 (n343, n140, n109, n169, n166);
nand g226 (n308, n144, n243, n129, n200);
nand g227 (n385, n169, n153, n109, n171);
and  g228 (n380, n240, n222, n172, n221);
nand g229 (n402, n178, n143, n134, n162);
or   g230 (n258, n131, n247, n229, n250);
and  g231 (n286, n140, n116, n94, n168);
xor  g232 (n302, n200, n239, n181, n110);
xnor g233 (n328, n103, n97, n161, n186);
nand g234 (n362, n87, n229, n194, n242);
nand g235 (n271, n117, n184, n123, n165);
and  g236 (n301, n152, n116, n210, n158);
xnor g237 (n382, n125, n223, n233, n93);
xor  g238 (n337, n148, n214, n221, n175);
and  g239 (n253, n168, n107, n106, n144);
xor  g240 (n381, n246, n228, n143, n107);
xnor g241 (n356, n220, n90, n186, n207);
xnor g242 (n281, n167, n193, n95, n222);
nor  g243 (n318, n230, n239, n96, n100);
and  g244 (n325, n243, n231, n146, n242);
nor  g245 (n376, n146, n122, n242, n185);
xor  g246 (n379, n169, n139, n244, n245);
xor  g247 (n341, n137, n108, n102, n148);
and  g248 (n393, n163, n209, n245, n89);
xor  g249 (n375, n196, n196, n226, n106);
nor  g250 (n378, n118, n185, n190, n184);
nor  g251 (n377, n111, n249, n116, n105);
xnor g252 (n278, n153, n202, n147, n241);
and  g253 (n383, n211, n222, n158, n164);
or   g254 (n303, n157, n125, n122, n206);
xnor g255 (n305, n98, n207, n117, n120);
and  g256 (n400, n218, n86, n141, n110);
and  g257 (n285, n225, n88, n206, n97);
xnor g258 (n269, n160, n95, n93, n205);
or   g259 (n273, n147, n236, n249, n179);
xnor g260 (n256, n101, n114, n167, n171);
nand g261 (n394, n133, n134, n201, n154);
or   g262 (n335, n238, n118, n191, n129);
or   g263 (n361, n115, n137, n197, n180);
nand g264 (n374, n126, n124, n232, n230);
nor  g265 (n327, n217, n147, n118, n183);
nor  g266 (n370, n213, n136, n233, n113);
and  g267 (n268, n166, n109, n205, n176);
nor  g268 (n355, n150, n141, n223, n134);
and  g269 (n396, n142, n154, n210, n132);
nand g270 (n364, n178, n121, n250);
nand g271 (n288, n231, n193, n234, n215);
and  g272 (n330, n143, n149, n120, n240);
xnor g273 (n295, n134, n160, n120, n147);
nand g274 (n290, n194, n241, n247, n96);
xnor g275 (n255, n208, n104, n131, n212);
and  g276 (n357, n174, n170, n187, n103);
xnor g277 (n340, n110, n119, n145, n131);
nor  g278 (n321, n168, n204, n189, n224);
xnor g279 (n350, n212, n230, n135, n227);
or   g280 (n367, n195, n102, n215, n132);
nand g281 (n409, n240, n228, n123, n152);
nand g282 (n289, n201, n208, n164, n227);
or   g283 (n304, n241, n170, n231, n202);
or   g284 (n311, n145, n192, n172, n86);
xor  g285 (n401, n87, n181, n185, n209);
or   g286 (n263, n111, n211, n234, n202);
or   g287 (n358, n128, n190, n96, n127);
nand g288 (n389, n201, n235, n177, n221);
and  g289 (n299, n154, n125, n236, n191);
and  g290 (n296, n239, n90, n170, n151);
nor  g291 (n313, n138, n112, n250, n179);
nand g292 (n413, n87, n101, n114, n189);
xor  g293 (n336, n244, n166, n218, n95);
nor  g294 (n411, n167, n158, n217, n122);
nand g295 (n363, n144, n194, n130, n159);
nor  g296 (n410, n219, n199, n90, n152);
nor  g297 (n282, n246, n184, n238, n117);
or   g298 (n293, n199, n213, n165, n161);
xor  g299 (n387, n95, n132, n92, n219);
xor  g300 (n384, n91, n218, n225, n205);
xor  g301 (n338, n235, n176, n232, n200);
or   g302 (n372, n154, n238, n151, n123);
xor  g303 (n307, n113, n98, n32, n192);
nand g304 (n397, n119, n136, n203, n247);
xor  g305 (n407, n206, n126, n197, n90);
and  g306 (n300, n248, n188, n157, n217);
or   g307 (n398, n229, n145, n204, n135);
nor  g308 (n406, n171, n195, n105, n137);
and  g309 (n395, n233, n98, n207, n127);
and  g310 (n405, n164, n186, n169, n191);
or   g311 (n316, n188, n132, n180, n229);
and  g312 (n348, n234, n198, n181, n94);
nor  g313 (n324, n209, n248, n223, n240);
xnor g314 (n339, n232, n88, n102, n159);
or   g315 (n319, n135, n163, n127, n145);
xor  g316 (n264, n153, n220, n211, n197);
xor  g317 (n314, n183, n121, n107, n214);
or   g318 (n315, n179, n123, n221, n186);
or   g319 (n403, n245, n216, n115, n173);
xnor g320 (n279, n156, n159, n127, n100);
nor  g321 (n317, n183, n88, n155, n103);
or   g322 (n412, n173, n129, n160, n246);
or   g323 (n292, n104, n248, n141, n168);
or   g324 (n366, n215, n185, n99, n165);
nand g325 (n323, n209, n199, n228, n226);
nor  g326 (n257, n150, n100, n241, n161);
nor  g327 (n365, n105, n100, n178, n126);
nand g328 (n267, n207, n224, n243, n94);
or   g329 (n254, n237, n182, n106, n136);
nand g330 (n353, n112, n142, n97, n133);
and  g331 (n404, n128, n236, n113, n163);
xor  g332 (n354, n188, n139, n142, n203);
xnor g333 (n260, n148, n173, n174, n235);
or   g334 (n306, n136, n198, n151, n141);
and  g335 (n276, n126, n172, n219, n212);
and  g336 (n275, n158, n149, n156, n174);
xor  g337 (n344, n152, n217, n142, n146);
or   g338 (n369, n226, n156, n111, n248);
xnor g339 (n414, n138, n249, n130, n211);
xor  g340 (n320, n242, n213, n92, n93);
xnor g341 (n270, n110, n224, n202, n130);
xnor g342 (n272, n103, n91, n214, n223);
xor  g343 (n351, n188, n113, n164, n203);
nor  g344 (n408, n187, n216, n124, n99);
xor  g345 (n360, n96, n208, n143, n249);
nand g346 (n352, n153, n204, n192, n244);
or   g347 (n332, n212, n176, n97, n216);
nand g348 (n349, n162, n183, n233, n177);
xnor g349 (n342, n104, n167, n245, n191);
nand g350 (n262, n150, n105, n237);
nand g351 (n386, n114, n187, n157, n155);
or   g352 (n309, n231, n182, n177, n148);
nor  g353 (n283, n89, n244, n200, n179);
or   g354 (n294, n187, n108, n32, n131);
nor  g355 (n388, n189, n190, n106, n162);
or   g356 (n251, n122, n204, n130, n144);
xor  g357 (n310, n119, n128, n190, n138);
xnor g358 (n297, n177, n195, n220, n184);
xnor g359 (n390, n140, n92, n175, n91);
xnor g360 (n265, n189, n149, n176);
or   g361 (n331, n213, n171, n133, n99);
nand g362 (n368, n124, n181, n120, n230);
xor  g363 (n261, n218, n175, n140, n89);
and  g364 (n259, n159, n243, n208, n128);
nor  g365 (n333, n115, n155, n124, n116);
nor  g366 (n359, n197, n234, n193, n101);
xnor g367 (n252, n220, n199, n151, n178);
xor  g368 (n280, n205, n119, n219, n201);
nor  g369 (n329, n112, n114, n236, n115);
and  g370 (n346, n139, n108, n203, n107);
nor  g371 (n266, n210, n174, n108, n117);
or   g372 (n347, n214, n180, n192, n250);
or   g373 (n284, n163, n99, n121, n156);
nand g374 (n371, n139, n225, n210, n238);
xor  g375 (n277, n146, n225, n175, n196);
xor  g376 (n274, n216, n111, n227, n129);
xor  g377 (n312, n172, n246, n94, n155);
xnor g378 (n287, n235, n160, n89, n109);
or   g379 (n415, n118, n133, n166, n215);
xnor g380 (n391, n125, n224, n222, n226);
nand g381 (n291, n165, n92, n98, n162);
nand g382 (n345, n137, n237, n157, n182);
and  g383 (n485, n306, n265, n259, n296);
nor  g384 (n426, n323, n321, n268, n284);
or   g385 (n441, n253, n313, n300, n325);
and  g386 (n461, n272, n294, n304, n300);
and  g387 (n428, n272, n256, n308, n265);
and  g388 (n488, n258, n312, n301, n270);
and  g389 (n483, n315, n251, n311, n303);
and  g390 (n453, n308, n273, n326, n307);
xor  g391 (n477, n314, n272, n269, n327);
xnor g392 (n425, n306, n263, n320, n278);
xnor g393 (n474, n312, n321, n274);
or   g394 (n439, n315, n271, n301, n262);
or   g395 (n492, n310, n276, n291, n257);
nor  g396 (n478, n304, n304, n295, n310);
nor  g397 (n434, n263, n314, n277, n305);
and  g398 (n486, n284, n251, n275, n307);
xnor g399 (n448, n325, n267, n311, n299);
nor  g400 (n460, n296, n323, n310, n322);
nand g401 (n479, n293, n270, n318, n277);
or   g402 (n480, n253, n322, n270, n319);
or   g403 (n451, n282, n286, n252, n328);
and  g404 (n469, n260, n293, n263, n303);
xor  g405 (n455, n252, n293, n284, n256);
xor  g406 (n420, n267, n302, n283, n318);
xnor g407 (n417, n319, n283, n302, n309);
xnor g408 (n430, n296, n274, n266, n307);
nor  g409 (n429, n315, n272, n305, n280);
xnor g410 (n467, n275, n328, n309, n290);
nor  g411 (n491, n267, n319, n282, n279);
or   g412 (n435, n270, n327, n297, n281);
xor  g413 (n463, n305, n278, n324, n268);
or   g414 (n432, n323, n251, n310, n289);
or   g415 (n482, n271, n297, n255, n257);
xnor g416 (n431, n264, n260, n279, n262);
xor  g417 (n484, n287, n274, n279, n322);
xor  g418 (n447, n262, n292, n261, n256);
nand g419 (n468, n275, n291, n263, n285);
nand g420 (n481, n318, n320, n266, n328);
nand g421 (n424, n294, n267, n317, n262);
xnor g422 (n422, n277, n288, n278, n307);
nand g423 (n475, n326, n323, n327, n266);
or   g424 (n456, n290, n283, n287, n293);
nand g425 (n449, n261, n321, n324, n313);
and  g426 (n446, n257, n264, n320, n268);
xnor g427 (n457, n261, n286, n264, n285);
or   g428 (n436, n276, n300, n281, n254);
nor  g429 (n493, n289, n288, n253, n286);
xnor g430 (n466, n328, n302, n259, n278);
xor  g431 (n423, n260, n294, n287, n281);
nor  g432 (n489, n269, n324, n299, n317);
nor  g433 (n443, n301, n255, n287, n261);
nand g434 (n458, n259, n281, n292, n321);
nand g435 (n465, n273, n285, n282, n296);
or   g436 (n440, n298, n309, n302, n254);
or   g437 (n471, n269, n275, n292, n314);
or   g438 (n437, n291, n290, n301, n297);
nor  g439 (n419, n297, n316, n257, n326);
and  g440 (n473, n308, n271, n286, n280);
and  g441 (n438, n290, n292, n322, n311);
xor  g442 (n444, n258, n303, n300, n319);
xor  g443 (n418, n325, n316, n265, n289);
xnor g444 (n450, n325, n266, n265, n298);
or   g445 (n421, n252, n308, n317, n311);
and  g446 (n464, n285, n315, n289, n255);
xor  g447 (n490, n299, n318, n312, n280);
nor  g448 (n459, n298, n273, n280, n312);
xor  g449 (n462, n258, n320, n288, n295);
or   g450 (n472, n306, n251, n295, n324);
xnor g451 (n445, n284, n277, n295, n253);
or   g452 (n476, n291, n314, n255, n252);
or   g453 (n433, n313, n316, n269, n304);
and  g454 (n442, n283, n299, n313, n264);
nand g455 (n487, n271, n288, n276, n256);
nor  g456 (n470, n276, n298, n327, n305);
and  g457 (n452, n303, n260, n254, n268);
nor  g458 (n416, n306, n294, n279, n316);
and  g459 (n454, n326, n282, n259, n273);
nand g460 (n427, n309, n254, n258, n317);
not  g461 (n499, n424);
not  g462 (n509, n420);
not  g463 (n505, n421);
buf  g464 (n504, n416);
buf  g465 (n522, n428);
not  g466 (n513, n419);
not  g467 (n520, n417);
buf  g468 (n501, n418);
not  g469 (n496, n417);
not  g470 (n497, n419);
buf  g471 (n515, n424);
not  g472 (n507, n428);
buf  g473 (n506, n420);
buf  g474 (n503, n427);
not  g475 (n514, n416);
not  g476 (n510, n426);
buf  g477 (n500, n423);
not  g478 (n512, n429);
nor  g479 (n519, n426, n421);
xnor g480 (n502, n420, n416);
and  g481 (n494, n428, n420, n421, n418);
xnor g482 (n508, n429, n425, n427, n418);
or   g483 (n516, n426, n422, n418, n417);
and  g484 (n517, n423, n429, n422);
nor  g485 (n498, n430, n423, n419, n422);
nor  g486 (n511, n428, n421, n423, n425);
xnor g487 (n495, n422, n426, n427, n425);
or   g488 (n521, n425, n424, n417, n427);
nor  g489 (n518, n419, n430, n416, n424);
xor  g490 (n615, n432, n357, n334, n502);
xnor g491 (n556, n351, n504, n349, n519);
xor  g492 (n596, n507, n434, n501, n503);
nor  g493 (n551, n516, n348, n453, n467);
nor  g494 (n563, n332, n335, n513, n454);
and  g495 (n555, n512, n329, n440, n507);
and  g496 (n540, n357, n342, n368, n364);
xnor g497 (n548, n341, n440, n463, n466);
nand g498 (n625, n329, n445, n351, n364);
xor  g499 (n568, n435, n335, n436, n466);
or   g500 (n547, n456, n462, n435, n496);
or   g501 (n589, n442, n439, n367, n346);
nor  g502 (n583, n520, n462, n365, n500);
nor  g503 (n605, n520, n363, n508, n515);
nand g504 (n533, n459, n340, n331);
nand g505 (n591, n444, n440, n336, n455);
xnor g506 (n576, n447, n465, n452, n436);
or   g507 (n586, n504, n446, n441, n442);
xnor g508 (n617, n348, n457, n347, n361);
xnor g509 (n580, n459, n442, n454, n503);
xnor g510 (n590, n501, n504, n453, n337);
nor  g511 (n543, n508, n443, n504, n439);
xor  g512 (n539, n518, n342, n451, n336);
nand g513 (n569, n360, n437, n337, n451);
nand g514 (n624, n438, n338, n362, n357);
xor  g515 (n595, n335, n469, n467, n347);
nor  g516 (n558, n461, n467, n468, n343);
xnor g517 (n573, n500, n498, n463, n457);
nor  g518 (n571, n517, n502, n447, n366);
and  g519 (n544, n464, n445, n439, n330);
and  g520 (n623, n351, n444, n449, n505);
and  g521 (n626, n510, n347, n453, n340);
xor  g522 (n554, n468, n369, n511, n350);
xor  g523 (n582, n364, n367, n458, n443);
xnor g524 (n535, n444, n512, n431, n338);
and  g525 (n600, n446, n365, n517, n514);
nand g526 (n621, n498, n499, n348, n452);
nor  g527 (n545, n451, n450, n515, n341);
xor  g528 (n541, n342, n447, n430, n515);
nor  g529 (n561, n508, n498, n462, n331);
or   g530 (n592, n521, n441, n455, n506);
xnor g531 (n581, n332, n511, n502, n460);
and  g532 (n538, n517, n512, n457, n514);
xnor g533 (n526, n362, n441, n333, n451);
and  g534 (n577, n456, n511, n501, n333);
xor  g535 (n601, n438, n360, n363, n522);
and  g536 (n528, n518, n505, n438, n503);
xor  g537 (n542, n509, n436, n461, n363);
and  g538 (n552, n349, n349, n445, n334);
nor  g539 (n565, n467, n495, n443, n338);
xnor g540 (n629, n341, n352, n496, n516);
and  g541 (n611, n464, n515, n499, n367);
xnor g542 (n578, n433, n438, n458, n343);
and  g543 (n598, n461, n510, n450, n351);
nor  g544 (n608, n452, n506, n344, n512);
and  g545 (n531, n329, n366, n353, n434);
xor  g546 (n614, n360, n500, n457, n448);
nor  g547 (n562, n340, n510, n436, n333);
or   g548 (n525, n352, n366, n465, n461);
nor  g549 (n534, n454, n516, n502);
xor  g550 (n619, n339, n346, n435, n433);
or   g551 (n570, n503, n433, n353, n464);
nand g552 (n628, n443, n431, n333, n495);
nor  g553 (n567, n446, n334, n513, n355);
or   g554 (n584, n444, n434, n353, n361);
xor  g555 (n527, n509, n356, n332, n460);
xor  g556 (n557, n346, n511, n356, n330);
nand g557 (n618, n522, n498, n494, n345);
xor  g558 (n575, n508, n363, n466, n495);
or   g559 (n607, n350, n339, n495, n365);
xor  g560 (n579, n466, n507, n344, n343);
nand g561 (n546, n433, n340, n344, n501);
nor  g562 (n550, n361, n354, n519, n449);
nor  g563 (n532, n432, n339, n519, n500);
nand g564 (n574, n362, n458, n355, n369);
xor  g565 (n620, n437, n368, n445, n447);
or   g566 (n599, n346, n345, n455, n449);
xnor g567 (n609, n359, n448, n356, n468);
or   g568 (n549, n519, n434, n330, n442);
xnor g569 (n560, n456, n455, n331, n462);
xor  g570 (n594, n448, n337, n496, n509);
or   g571 (n616, n345, n464, n497, n446);
xnor g572 (n530, n496, n448, n463, n518);
nand g573 (n564, n522, n522, n468, n334);
nor  g574 (n536, n338, n432, n359, n350);
and  g575 (n603, n453, n359, n505, n459);
nand g576 (n610, n341, n456, n499, n345);
or   g577 (n627, n521, n460, n431, n358);
or   g578 (n630, n332, n518, n367, n459);
nand g579 (n606, n352, n497, n521, n342);
xor  g580 (n593, n353, n336, n449, n362);
or   g581 (n587, n369, n450, n514, n505);
or   g582 (n622, n344, n513, n359, n360);
or   g583 (n529, n347, n354, n465, n509);
or   g584 (n524, n465, n458, n435, n450);
nand g585 (n572, n507, n339, n349, n432);
nor  g586 (n585, n354, n520, n329, n356);
or   g587 (n612, n521, n364, n439, n369);
xnor g588 (n553, n514, n454, n348, n352);
or   g589 (n602, n330, n355, n460);
nand g590 (n566, n497, n506, n431, n358);
nand g591 (n597, n452, n365, n337, n361);
xor  g592 (n588, n350, n335, n368, n440);
and  g593 (n604, n358, n368, n354, n441);
or   g594 (n559, n358, n343, n463, n366);
nand g595 (n613, n336, n437, n497);
xnor g596 (n537, n517, n506, n510, n520);
xor  g597 (n523, n499, n357, n513, n430);
xor  g598 (n658, n617, n409, n479, n606);
nor  g599 (n678, n619, n604, n484, n605);
nand g600 (n742, n586, n535, n393, n475);
xnor g601 (n646, n477, n626, n376, n615);
nor  g602 (n642, n599, n386, n380, n485);
xor  g603 (n656, n611, n600, n627, n618);
or   g604 (n677, n552, n492, n372, n493);
xor  g605 (n744, n613, n381, n626, n409);
nor  g606 (n699, n476, n623, n384, n403);
and  g607 (n633, n392, n555, n379, n370);
nor  g608 (n640, n598, n479, n411, n388);
and  g609 (n696, n594, n624, n400, n380);
or   g610 (n670, n539, n382, n625, n581);
and  g611 (n664, n620, n472, n408, n414);
and  g612 (n737, n576, n381, n615, n600);
and  g613 (n695, n536, n411, n571, n378);
nand g614 (n648, n575, n408, n578, n613);
xnor g615 (n724, n616, n596, n597, n614);
xnor g616 (n647, n394, n630, n403, n550);
nor  g617 (n644, n628, n607, n485, n483);
or   g618 (n703, n390, n613, n406, n381);
xnor g619 (n727, n492, n399, n480, n379);
and  g620 (n746, n478, n610, n412, n386);
or   g621 (n717, n477, n413, n470, n606);
nand g622 (n721, n569, n629, n618, n378);
xor  g623 (n665, n398, n469, n406, n568);
and  g624 (n728, n389, n380, n600, n624);
nor  g625 (n729, n612, n626, n401, n481);
or   g626 (n751, n485, n414, n376, n484);
and  g627 (n711, n629, n387, n388, n384);
nand g628 (n649, n606, n615, n413, n381);
nand g629 (n693, n566, n617, n478, n533);
xnor g630 (n679, n493, n474, n623, n407);
xor  g631 (n716, n372, n402, n593, n391);
xor  g632 (n705, n492, n388, n384, n375);
and  g633 (n682, n415, n481, n405, n630);
or   g634 (n689, n574, n616, n470, n397);
xor  g635 (n754, n493, n394, n610, n573);
nor  g636 (n710, n486, n376, n371, n563);
nor  g637 (n674, n547, n627, n617, n628);
or   g638 (n708, n542, n482, n372, n612);
and  g639 (n735, n409, n469, n391, n615);
nor  g640 (n733, n614, n480, n383, n396);
nor  g641 (n666, n376, n476, n485, n382);
or   g642 (n720, n486, n604, n411, n389);
nand g643 (n655, n608, n628, n597, n605);
xor  g644 (n707, n582, n469, n371, n471);
nand g645 (n697, n391, n415, n407, n383);
or   g646 (n688, n609, n408, n401, n375);
nand g647 (n676, n385, n373, n405, n413);
nor  g648 (n726, n621, n487, n393, n560);
nor  g649 (n706, n597, n395, n540, n532);
xnor g650 (n718, n612, n375, n413, n588);
or   g651 (n631, n478, n407, n487, n383);
nor  g652 (n651, n412, n412, n478, n579);
xor  g653 (n650, n396, n608, n598, n541);
nand g654 (n681, n479, n558, n553, n623);
xor  g655 (n654, n409, n587, n549, n392);
xnor g656 (n741, n380, n527, n481, n604);
or   g657 (n734, n622, n475, n483, n406);
nand g658 (n672, n378, n472, n548, n374);
xnor g659 (n709, n404, n392, n414, n477);
nor  g660 (n645, n484, n609, n590, n410);
xor  g661 (n698, n402, n405, n412, n370);
and  g662 (n700, n608, n408, n414, n609);
or   g663 (n669, n620, n611, n395, n604);
xnor g664 (n714, n370, n371, n559, n477);
nor  g665 (n661, n601, n393, n405, n398);
xnor g666 (n752, n383, n395, n482, n398);
and  g667 (n635, n609, n374, n493, n373);
nand g668 (n634, n584, n603, n472, n602);
nor  g669 (n738, n474, n373, n398, n607);
xor  g670 (n639, n538, n470, n489, n622);
or   g671 (n750, n396, n402, n530, n523);
nand g672 (n660, n601, n531, n545, n386);
nand g673 (n691, n602, n618, n625);
xnor g674 (n659, n394, n387, n489, n490);
xnor g675 (n662, n621, n374, n399, n480);
nand g676 (n657, n606, n537, n596, n619);
xnor g677 (n704, n583, n620, n387, n404);
or   g678 (n638, n628, n410, n475, n476);
and  g679 (n736, n611, n618, n492, n473);
xnor g680 (n686, n395, n612, n377, n630);
xor  g681 (n653, n602, n603, n599, n565);
nor  g682 (n692, n610, n474, n484, n377);
or   g683 (n731, n473, n389, n399, n402);
xnor g684 (n701, n483, n482, n597, n544);
nor  g685 (n685, n629, n397, n624, n603);
or   g686 (n632, n475, n567, n614, n561);
or   g687 (n643, n490, n490, n410, n385);
or   g688 (n636, n603, n572, n371, n525);
and  g689 (n694, n379, n589, n621, n382);
xnor g690 (n723, n400, n403, n471, n619);
or   g691 (n732, n392, n616, n486, n526);
and  g692 (n667, n591, n375, n543, n622);
nand g693 (n719, n599, n610, n470, n614);
or   g694 (n702, n483, n389, n487, n397);
xor  g695 (n753, n488, n387, n607, n474);
xor  g696 (n673, n601, n393, n399, n415);
nand g697 (n713, n601, n528, n407, n390);
xor  g698 (n739, n476, n620, n556, n564);
nor  g699 (n740, n491, n627, n570, n384);
and  g700 (n652, n473, n599, n374, n390);
xnor g701 (n687, n619, n400, n415, n382);
nand g702 (n749, n406, n397, n373, n372);
and  g703 (n745, n488, n396, n401, n491);
nand g704 (n722, n481, n629, n400, n630);
xor  g705 (n683, n489, n613, n404, n473);
xnor g706 (n748, n472, n627, n595, n471);
or   g707 (n747, n546, n377, n580);
and  g708 (n725, n482, n602, n534, n611);
xnor g709 (n637, n385, n608, n625, n605);
xor  g710 (n671, n596, n404, n621, n551);
xnor g711 (n663, n598, n471, n491, n401);
nor  g712 (n641, n390, n486, n598, n626);
xor  g713 (n675, n386, n487, n623, n562);
nor  g714 (n680, n607, n596, n617, n624);
xnor g715 (n743, n616, n394, n577, n600);
nor  g716 (n668, n391, n378, n489, n410);
nand g717 (n715, n491, n622, n370, n385);
xnor g718 (n712, n557, n592, n490, n488);
xor  g719 (n684, n480, n479, n411, n605);
nand g720 (n730, n488, n379, n585, n388);
xnor g721 (n690, n524, n554, n529, n403);
or   g722 (n779, n638, n738, n742, n721);
nor  g723 (n855, n751, n642, n670, n716);
or   g724 (n762, n738, n636, n637, n694);
xnor g725 (n764, n724, n745, n741, n715);
nor  g726 (n827, n732, n694, n704, n664);
xnor g727 (n765, n712, n739, n699, n696);
xor  g728 (n858, n687, n675, n719, n720);
or   g729 (n826, n636, n692, n632, n701);
xor  g730 (n776, n702, n703, n676, n697);
xor  g731 (n841, n672, n733, n681, n674);
nor  g732 (n781, n748, n691, n650, n692);
nand g733 (n824, n722, n659, n665, n634);
and  g734 (n840, n741, n713, n660, n661);
or   g735 (n773, n668, n706, n725, n710);
xor  g736 (n852, n736, n646, n683, n636);
nor  g737 (n847, n660, n723, n662, n717);
or   g738 (n843, n737, n635, n637, n711);
and  g739 (n784, n664, n649, n731, n729);
xor  g740 (n875, n732, n699, n750, n647);
and  g741 (n821, n641, n730, n675, n705);
xor  g742 (n857, n652, n732, n681, n673);
xnor g743 (n872, n747, n737, n724, n712);
or   g744 (n778, n741, n727, n702, n664);
or   g745 (n863, n711, n681, n721, n753);
nor  g746 (n864, n727, n689, n717, n680);
nor  g747 (n805, n669, n719, n650, n656);
nand g748 (n814, n701, n745, n668, n656);
nor  g749 (n804, n703, n753, n659, n700);
and  g750 (n758, n730, n682, n674, n658);
nor  g751 (n761, n634, n751, n647, n633);
xnor g752 (n763, n725, n673, n644, n651);
xor  g753 (n819, n710, n749, n745, n666);
or   g754 (n759, n649, n736, n715, n717);
nor  g755 (n799, n738, n739, n727, n719);
nand g756 (n795, n689, n748, n688, n746);
xnor g757 (n823, n733, n646, n720, n647);
nand g758 (n856, n748, n703, n683, n678);
nand g759 (n772, n666, n709, n713, n705);
nor  g760 (n791, n655, n735, n646, n719);
xnor g761 (n801, n752, n631, n721, n706);
and  g762 (n831, n667, n644, n632, n671);
and  g763 (n783, n656, n641, n708, n734);
and  g764 (n782, n722, n694, n687, n643);
nor  g765 (n822, n645, n749, n708, n686);
or   g766 (n755, n707, n653, n654, n677);
nor  g767 (n833, n684, n700, n641, n656);
or   g768 (n839, n711, n668, n669, n718);
or   g769 (n853, n648, n659, n733, n676);
and  g770 (n849, n697, n700, n735, n657);
and  g771 (n792, n704, n734, n710, n644);
nor  g772 (n766, n722, n651, n720, n730);
or   g773 (n850, n746, n740, n708, n679);
nor  g774 (n777, n676, n726, n741, n728);
nand g775 (n867, n638, n673, n702, n700);
xor  g776 (n793, n711, n736, n639, n672);
and  g777 (n859, n652, n640, n750, n679);
xor  g778 (n780, n720, n747, n652, n636);
nor  g779 (n870, n632, n663, n697, n729);
nand g780 (n806, n717, n690, n683, n731);
or   g781 (n790, n747, n645, n678, n665);
and  g782 (n811, n696, n635, n731, n680);
xnor g783 (n861, n736, n635, n726, n685);
and  g784 (n774, n665, n680, n690, n637);
or   g785 (n800, n726, n721, n715, n647);
xor  g786 (n771, n658, n723, n638, n714);
xnor g787 (n810, n686, n702, n657, n716);
nand g788 (n812, n678, n715, n701, n728);
and  g789 (n865, n642, n648, n633, n706);
and  g790 (n816, n648, n751, n642, n696);
nor  g791 (n842, n654, n685, n695, n634);
nand g792 (n851, n692, n701, n714, n725);
nand g793 (n770, n641, n743, n655, n643);
or   g794 (n846, n674, n735, n749, n710);
or   g795 (n798, n646, n675, n740, n684);
nor  g796 (n788, n743, n671, n752, n753);
xnor g797 (n796, n648, n696, n709, n698);
nand g798 (n768, n687, n677, n733, n639);
nor  g799 (n808, n635, n740, n653, n668);
or   g800 (n874, n737, n691, n750, n669);
xor  g801 (n838, n731, n750, n709, n714);
xor  g802 (n835, n737, n723, n697, n661);
or   g803 (n802, n640, n734, n639, n671);
nor  g804 (n862, n732, n742, n643, n674);
or   g805 (n866, n752, n640, n662, n713);
xnor g806 (n803, n693, n665, n673, n688);
xor  g807 (n871, n693, n724, n638, n723);
and  g808 (n868, n667, n657, n653, n705);
or   g809 (n775, n713, n689, n640, n631);
xor  g810 (n767, n726, n667, n722, n712);
and  g811 (n820, n658, n727, n676, n663);
xor  g812 (n813, n655, n684, n670, n650);
nand g813 (n844, n728, n747, n671, n695);
xnor g814 (n830, n718, n746, n735, n692);
nand g815 (n785, n730, n681, n661, n645);
or   g816 (n769, n724, n657, n675, n651);
and  g817 (n877, n695, n698, n688, n691);
xor  g818 (n845, n643, n740, n716, n695);
nand g819 (n807, n684, n743, n633, n661);
xnor g820 (n834, n744, n631, n679, n654);
and  g821 (n873, n752, n679, n729, n682);
and  g822 (n828, n670, n699, n734, n739);
or   g823 (n836, n685, n660, n729);
xor  g824 (n815, n693, n716, n698, n653);
xor  g825 (n876, n748, n677, n633, n662);
nor  g826 (n869, n709, n642, n686, n663);
xor  g827 (n760, n662, n705, n718, n706);
nand g828 (n818, n637, n683, n707, n686);
nand g829 (n848, n689, n714, n670, n744);
nor  g830 (n854, n651, n738, n703, n739);
xor  g831 (n832, n685, n687, n688, n744);
xnor g832 (n794, n655, n677, n753, n669);
xor  g833 (n829, n672, n649, n742);
nor  g834 (n825, n704, n690, n751, n694);
or   g835 (n817, n728, n743, n712, n708);
xor  g836 (n860, n663, n749, n659, n645);
xnor g837 (n786, n745, n639, n654, n644);
or   g838 (n797, n682, n744, n693, n707);
xor  g839 (n789, n682, n650, n698, n718);
xnor g840 (n756, n725, n632, n680, n707);
xor  g841 (n809, n667, n699, n666);
or   g842 (n787, n631, n691, n672, n664);
and  g843 (n837, n742, n678, n690, n704);
nand g844 (n757, n652, n634, n746, n658);
nand g845 (n896, n790, n761, n868, n763);
xor  g846 (n911, n832, n835, n767, n756);
xnor g847 (n930, n809, n756, n754, n797);
nand g848 (n880, n839, n768, n872, n821);
or   g849 (n981, n803, n797, n790);
nor  g850 (n914, n825, n817, n863, n764);
and  g851 (n993, n875, n843, n814, n798);
nor  g852 (n907, n873, n846, n762, n776);
nor  g853 (n982, n828, n847, n839, n773);
nand g854 (n1000, n817, n841, n779, n850);
nand g855 (n970, n765, n858, n802, n792);
and  g856 (n901, n852, n810, n862, n782);
or   g857 (n919, n764, n834, n794, n835);
nand g858 (n902, n820, n768, n803, n845);
and  g859 (n897, n875, n861, n827, n772);
xnor g860 (n947, n817, n869, n786, n840);
nor  g861 (n965, n786, n795, n761, n876);
and  g862 (n985, n770, n807, n857, n837);
xnor g863 (n898, n812, n870, n864, n869);
and  g864 (n974, n874, n794, n848, n787);
xor  g865 (n953, n777, n844, n823, n780);
xor  g866 (n950, n869, n835, n823, n848);
xnor g867 (n881, n800, n772, n846, n872);
nor  g868 (n926, n834, n854, n877, n814);
or   g869 (n928, n809, n840, n855, n839);
xnor g870 (n975, n764, n791, n789, n841);
and  g871 (n987, n779, n811, n849, n760);
xor  g872 (n972, n862, n818, n809, n829);
nor  g873 (n929, n831, n780, n863, n769);
nand g874 (n989, n774, n819, n876, n824);
xor  g875 (n969, n860, n840, n825, n784);
or   g876 (n962, n767, n792, n868, n811);
or   g877 (n984, n851, n851, n858, n795);
or   g878 (n948, n875, n865, n774, n848);
xor  g879 (n899, n844, n820, n850, n792);
nor  g880 (n994, n873, n826, n860, n857);
or   g881 (n976, n761, n769, n804, n863);
xor  g882 (n908, n868, n837, n826, n852);
or   g883 (n913, n769, n757, n760, n755);
or   g884 (n954, n808, n822, n866, n832);
xnor g885 (n966, n806, n761, n781, n785);
and  g886 (n963, n770, n778, n805, n768);
xor  g887 (n1001, n762, n774, n862, n872);
xnor g888 (n891, n856, n868, n760, n855);
xnor g889 (n951, n822, n866, n816, n796);
nor  g890 (n910, n788, n812, n838, n772);
nor  g891 (n973, n859, n764, n857, n876);
xnor g892 (n932, n831, n812, n815, n872);
nor  g893 (n923, n793, n849, n844, n836);
or   g894 (n939, n755, n874, n833, n864);
nand g895 (n904, n813, n818, n804, n877);
xor  g896 (n958, n841, n869, n788, n854);
xor  g897 (n905, n830, n852, n805, n871);
xnor g898 (n884, n758, n824, n784, n794);
nor  g899 (n921, n775, n847, n856, n854);
or   g900 (n931, n846, n860, n780);
xor  g901 (n894, n792, n790, n773, n800);
or   g902 (n955, n801, n757, n805, n802);
xor  g903 (n906, n824, n831, n837, n804);
or   g904 (n886, n785, n819, n833, n807);
nand g905 (n887, n820, n773, n776, n799);
or   g906 (n878, n842, n754, n785, n841);
xor  g907 (n980, n844, n859, n786, n832);
xnor g908 (n917, n877, n871, n796, n822);
or   g909 (n888, n865, n791, n776, n830);
xnor g910 (n938, n789, n827, n774, n788);
nor  g911 (n885, n781, n832, n830, n823);
nand g912 (n960, n772, n793, n815, n758);
xnor g913 (n988, n810, n762, n797, n801);
xnor g914 (n952, n858, n777, n829, n873);
nor  g915 (n942, n766, n855, n842, n798);
xnor g916 (n998, n775, n817, n785, n776);
nor  g917 (n990, n819, n847, n859, n813);
xor  g918 (n892, n862, n851, n799, n867);
and  g919 (n895, n847, n777, n806, n796);
xnor g920 (n915, n791, n851, n797, n861);
nor  g921 (n959, n765, n770, n784, n826);
and  g922 (n900, n864, n867, n782, n857);
xor  g923 (n890, n827, n754, n777, n765);
xor  g924 (n968, n809, n763, n759, n873);
nand g925 (n943, n811, n757, n838, n849);
xor  g926 (n893, n798, n766, n839, n775);
nor  g927 (n912, n816, n866, n778, n853);
and  g928 (n967, n843, n846, n860, n816);
and  g929 (n934, n803, n871, n816, n789);
nand g930 (n978, n814, n822, n799, n831);
nor  g931 (n922, n829, n782, n783, n815);
and  g932 (n889, n850, n850, n854, n863);
xor  g933 (n937, n836, n824, n825, n758);
nand g934 (n949, n826, n783, n788);
xnor g935 (n916, n833, n802, n756, n877);
and  g936 (n925, n767, n843, n821, n836);
xor  g937 (n991, n755, n875, n775, n815);
and  g938 (n996, n829, n864, n767, n805);
nand g939 (n924, n845, n766, n853, n778);
xor  g940 (n961, n810, n823, n827, n861);
and  g941 (n979, n795, n843, n811, n821);
xor  g942 (n956, n791, n825, n866, n849);
and  g943 (n882, n798, n758, n837, n801);
nand g944 (n940, n842, n830, n803, n779);
nor  g945 (n941, n793, n865, n794, n795);
nand g946 (n997, n768, n865, n876, n870);
nand g947 (n927, n778, n757, n871, n804);
nor  g948 (n920, n861, n820, n874, n853);
xor  g949 (n936, n760, n799, n771, n858);
or   g950 (n964, n765, n852, n870, n818);
xor  g951 (n903, n759, n771, n808, n786);
or   g952 (n971, n796, n819, n754, n834);
or   g953 (n918, n802, n800, n807, n845);
xnor g954 (n935, n756, n814, n833, n867);
and  g955 (n946, n828, n755, n834, n840);
and  g956 (n999, n771, n766, n808, n787);
nand g957 (n909, n779, n763, n874, n838);
nand g958 (n933, n793, n838, n770, n789);
and  g959 (n945, n781, n769, n859, n787);
or   g960 (n883, n842, n781, n821, n806);
nor  g961 (n992, n759, n759, n813, n856);
xnor g962 (n977, n807, n806, n813, n828);
nand g963 (n995, n773, n818, n762, n835);
nand g964 (n957, n800, n812, n836, n808);
xnor g965 (n879, n801, n828, n783, n853);
nand g966 (n983, n855, n784, n771, n856);
xnor g967 (n986, n787, n845, n848, n867);
or   g968 (n944, n763, n782, n870, n810);
xnor g969 (n1019, n897, n985, n953, n921);
nor  g970 (n1011, n976, n916, n883, n955);
xor  g971 (n1024, n885, n931, n881, n882);
xor  g972 (n1004, n986, n908, n989, n929);
or   g973 (n1007, n951, n879, n926, n966);
nor  g974 (n1027, n889, n997, n992, n972);
or   g975 (n1028, n937, n924, n944, n995);
nand g976 (n1016, n984, n918, n957, n896);
xor  g977 (n1005, n941, n880, n969, n909);
nor  g978 (n1030, n893, n978, n934, n884);
nand g979 (n1015, n900, n952, n903, n938);
xnor g980 (n1020, n901, n996, n940, n967);
xnor g981 (n1002, n922, n878, n974, n962);
xnor g982 (n1032, n894, n988, n927, n963);
nand g983 (n1025, n888, n971, n948, n975);
xor  g984 (n1014, n935, n961, n959, n915);
xnor g985 (n1031, n942, n950, n980, n917);
nand g986 (n1010, n973, n936, n949, n920);
and  g987 (n1023, n965, n905, n891, n930);
xnor g988 (n1018, n943, n1000, n914, n958);
xnor g989 (n1003, n983, n939, n933, n902);
nor  g990 (n1022, n970, n911, n904, n993);
nand g991 (n1008, n923, n925, n910, n977);
and  g992 (n1009, n932, n928, n991, n898);
or   g993 (n1006, n890, n999, n912, n907);
nand g994 (n1017, n892, n987, n982, n906);
xor  g995 (n1026, n887, n979, n960, n998);
nor  g996 (n1029, n945, n981, n964, n954);
nand g997 (n1012, n1001, n886, n968, n994);
nor  g998 (n1013, n956, n919, n946, n913);
xor  g999 (n1021, n899, n990, n895, n947);
endmodule
