

module Stat_2000_311
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n892,
  n886,
  n877,
  n890,
  n870,
  n880,
  n872,
  n884,
  n871,
  n883,
  n881,
  n869,
  n891,
  n873,
  n887,
  n882,
  n866,
  n1953,
  n2028,
  n2023,
  n2022,
  n2020,
  n2027,
  n2031,
  n2029,
  n2025,
  n2030,
  n2021,
  n2019,
  n2026,
  n2032,
  n2024,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n892;output n886;output n877;output n890;output n870;output n880;output n872;output n884;output n871;output n883;output n881;output n869;output n891;output n873;output n887;output n882;output n866;output n1953;output n2028;output n2023;output n2022;output n2020;output n2027;output n2031;output n2029;output n2025;output n2030;output n2021;output n2019;output n2026;output n2032;output n2024;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n867;wire n868;wire n874;wire n875;wire n876;wire n878;wire n879;wire n885;wire n888;wire n889;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n61,
    n24
  );


  buf
  g1
  (
    n52,
    n20
  );


  buf
  g2
  (
    n143,
    n29
  );


  not
  g3
  (
    n50,
    n18
  );


  not
  g4
  (
    n56,
    n9
  );


  buf
  g5
  (
    n126,
    n19
  );


  not
  g6
  (
    n131,
    n29
  );


  not
  g7
  (
    n39,
    n13
  );


  buf
  g8
  (
    n93,
    n11
  );


  buf
  g9
  (
    n70,
    n25
  );


  not
  g10
  (
    n103,
    n31
  );


  buf
  g11
  (
    n65,
    n12
  );


  not
  g12
  (
    n62,
    n7
  );


  not
  g13
  (
    n134,
    n27
  );


  not
  g14
  (
    n66,
    n23
  );


  buf
  g15
  (
    n35,
    n27
  );


  not
  g16
  (
    n105,
    n7
  );


  buf
  g17
  (
    n40,
    n18
  );


  not
  g18
  (
    n112,
    n7
  );


  buf
  g19
  (
    n140,
    n30
  );


  buf
  g20
  (
    n33,
    n3
  );


  not
  g21
  (
    n94,
    n1
  );


  buf
  g22
  (
    n67,
    n22
  );


  not
  g23
  (
    n37,
    n19
  );


  buf
  g24
  (
    n92,
    n20
  );


  not
  g25
  (
    n108,
    n30
  );


  not
  g26
  (
    n144,
    n13
  );


  not
  g27
  (
    n88,
    n16
  );


  not
  g28
  (
    n129,
    n3
  );


  not
  g29
  (
    n46,
    n15
  );


  buf
  g30
  (
    n136,
    n25
  );


  buf
  g31
  (
    n47,
    n6
  );


  buf
  g32
  (
    n45,
    n12
  );


  not
  g33
  (
    n49,
    n7
  );


  buf
  g34
  (
    n118,
    n9
  );


  buf
  g35
  (
    n121,
    n29
  );


  not
  g36
  (
    n34,
    n28
  );


  not
  g37
  (
    n78,
    n13
  );


  not
  g38
  (
    n132,
    n13
  );


  buf
  g39
  (
    n122,
    n28
  );


  not
  g40
  (
    n135,
    n26
  );


  buf
  g41
  (
    n97,
    n23
  );


  buf
  g42
  (
    n74,
    n8
  );


  buf
  g43
  (
    n128,
    n26
  );


  not
  g44
  (
    n130,
    n4
  );


  buf
  g45
  (
    n58,
    n1
  );


  buf
  g46
  (
    n107,
    n17
  );


  buf
  g47
  (
    n53,
    n14
  );


  buf
  g48
  (
    n63,
    n17
  );


  buf
  g49
  (
    n96,
    n6
  );


  buf
  g50
  (
    n42,
    n21
  );


  not
  g51
  (
    n113,
    n8
  );


  buf
  g52
  (
    n119,
    n15
  );


  not
  g53
  (
    n44,
    n29
  );


  not
  g54
  (
    n87,
    n11
  );


  buf
  g55
  (
    n84,
    n5
  );


  not
  g56
  (
    n55,
    n3
  );


  not
  g57
  (
    n137,
    n5
  );


  not
  g58
  (
    n139,
    n9
  );


  buf
  g59
  (
    n141,
    n27
  );


  not
  g60
  (
    n138,
    n23
  );


  buf
  g61
  (
    n100,
    n8
  );


  buf
  g62
  (
    n101,
    n14
  );


  not
  g63
  (
    n69,
    n2
  );


  not
  g64
  (
    n77,
    n26
  );


  not
  g65
  (
    n115,
    n24
  );


  not
  g66
  (
    n83,
    n20
  );


  not
  g67
  (
    n89,
    n18
  );


  buf
  g68
  (
    n81,
    n1
  );


  buf
  g69
  (
    n124,
    n16
  );


  buf
  g70
  (
    n57,
    n24
  );


  not
  g71
  (
    n82,
    n22
  );


  not
  g72
  (
    n111,
    n26
  );


  not
  g73
  (
    n99,
    n2
  );


  not
  g74
  (
    n106,
    n12
  );


  buf
  g75
  (
    n114,
    n4
  );


  not
  g76
  (
    n117,
    n9
  );


  buf
  g77
  (
    n68,
    n23
  );


  buf
  g78
  (
    n120,
    n10
  );


  not
  g79
  (
    n38,
    n14
  );


  not
  g80
  (
    n133,
    n16
  );


  not
  g81
  (
    n95,
    n19
  );


  buf
  g82
  (
    n125,
    n18
  );


  not
  g83
  (
    n147,
    n25
  );


  not
  g84
  (
    n64,
    n10
  );


  buf
  g85
  (
    n109,
    n28
  );


  not
  g86
  (
    n54,
    n10
  );


  buf
  g87
  (
    n60,
    n17
  );


  buf
  g88
  (
    n91,
    n22
  );


  buf
  g89
  (
    n80,
    n8
  );


  buf
  g90
  (
    n59,
    n21
  );


  not
  g91
  (
    n98,
    n4
  );


  buf
  g92
  (
    n127,
    n5
  );


  not
  g93
  (
    n110,
    n21
  );


  buf
  g94
  (
    n48,
    n11
  );


  not
  g95
  (
    n43,
    n21
  );


  not
  g96
  (
    n145,
    n30
  );


  buf
  g97
  (
    n142,
    n6
  );


  not
  g98
  (
    n51,
    n22
  );


  not
  g99
  (
    n72,
    n14
  );


  not
  g100
  (
    n148,
    n30
  );


  not
  g101
  (
    n79,
    n16
  );


  not
  g102
  (
    n90,
    n6
  );


  not
  g103
  (
    n123,
    n24
  );


  buf
  g104
  (
    n86,
    n2
  );


  not
  g105
  (
    n75,
    n28
  );


  buf
  g106
  (
    n102,
    n17
  );


  not
  g107
  (
    n73,
    n27
  );


  not
  g108
  (
    n85,
    n12
  );


  buf
  g109
  (
    n41,
    n15
  );


  buf
  g110
  (
    n116,
    n11
  );


  not
  g111
  (
    n76,
    n25
  );


  buf
  g112
  (
    n104,
    n15
  );


  not
  g113
  (
    n71,
    n19
  );


  not
  g114
  (
    n146,
    n20
  );


  buf
  g115
  (
    n36,
    n10
  );


  not
  g116
  (
    n446,
    n98
  );


  buf
  g117
  (
    n292,
    n48
  );


  not
  g118
  (
    n387,
    n85
  );


  not
  g119
  (
    n463,
    n35
  );


  not
  g120
  (
    n383,
    n66
  );


  buf
  g121
  (
    n343,
    n111
  );


  not
  g122
  (
    n376,
    n48
  );


  not
  g123
  (
    n169,
    n97
  );


  buf
  g124
  (
    n166,
    n72
  );


  not
  g125
  (
    n335,
    n88
  );


  not
  g126
  (
    n431,
    n49
  );


  buf
  g127
  (
    n175,
    n36
  );


  not
  g128
  (
    n185,
    n44
  );


  not
  g129
  (
    n274,
    n49
  );


  not
  g130
  (
    n237,
    n91
  );


  buf
  g131
  (
    n219,
    n113
  );


  buf
  g132
  (
    n440,
    n42
  );


  not
  g133
  (
    n295,
    n68
  );


  not
  g134
  (
    n331,
    n92
  );


  buf
  g135
  (
    n277,
    n54
  );


  not
  g136
  (
    n281,
    n87
  );


  not
  g137
  (
    n485,
    n114
  );


  buf
  g138
  (
    n260,
    n94
  );


  not
  g139
  (
    n241,
    n73
  );


  buf
  g140
  (
    n452,
    n37
  );


  not
  g141
  (
    n242,
    n79
  );


  not
  g142
  (
    n300,
    n92
  );


  buf
  g143
  (
    n430,
    n52
  );


  buf
  g144
  (
    n276,
    n87
  );


  buf
  g145
  (
    n438,
    n89
  );


  buf
  g146
  (
    n416,
    n101
  );


  not
  g147
  (
    n244,
    n45
  );


  not
  g148
  (
    n384,
    n101
  );


  buf
  g149
  (
    n428,
    n104
  );


  not
  g150
  (
    n195,
    n69
  );


  buf
  g151
  (
    n330,
    n82
  );


  buf
  g152
  (
    n378,
    n86
  );


  not
  g153
  (
    n153,
    n68
  );


  buf
  g154
  (
    n163,
    n58
  );


  buf
  g155
  (
    n196,
    n65
  );


  not
  g156
  (
    n471,
    n112
  );


  not
  g157
  (
    n298,
    n60
  );


  buf
  g158
  (
    n389,
    n74
  );


  not
  g159
  (
    n417,
    n112
  );


  not
  g160
  (
    n272,
    n41
  );


  not
  g161
  (
    n412,
    n68
  );


  buf
  g162
  (
    n315,
    n104
  );


  not
  g163
  (
    n204,
    n50
  );


  buf
  g164
  (
    n225,
    n116
  );


  buf
  g165
  (
    n290,
    n117
  );


  buf
  g166
  (
    n210,
    n84
  );


  buf
  g167
  (
    n309,
    n100
  );


  not
  g168
  (
    n443,
    n90
  );


  not
  g169
  (
    n406,
    n63
  );


  not
  g170
  (
    n371,
    n72
  );


  not
  g171
  (
    n402,
    n77
  );


  buf
  g172
  (
    n350,
    n114
  );


  buf
  g173
  (
    n296,
    n77
  );


  buf
  g174
  (
    n477,
    n44
  );


  buf
  g175
  (
    n271,
    n85
  );


  buf
  g176
  (
    n338,
    n108
  );


  buf
  g177
  (
    n181,
    n65
  );


  buf
  g178
  (
    n340,
    n89
  );


  buf
  g179
  (
    n474,
    n115
  );


  buf
  g180
  (
    n313,
    n71
  );


  not
  g181
  (
    n191,
    n37
  );


  buf
  g182
  (
    n388,
    n50
  );


  buf
  g183
  (
    n461,
    n68
  );


  buf
  g184
  (
    n421,
    n93
  );


  not
  g185
  (
    n304,
    n38
  );


  not
  g186
  (
    n324,
    n106
  );


  buf
  g187
  (
    n186,
    n70
  );


  buf
  g188
  (
    n256,
    n73
  );


  not
  g189
  (
    n162,
    n66
  );


  buf
  g190
  (
    n483,
    n106
  );


  not
  g191
  (
    n265,
    n88
  );


  buf
  g192
  (
    n280,
    n89
  );


  not
  g193
  (
    n258,
    n33
  );


  not
  g194
  (
    n359,
    n70
  );


  not
  g195
  (
    n426,
    n115
  );


  buf
  g196
  (
    n355,
    n110
  );


  buf
  g197
  (
    n167,
    n52
  );


  buf
  g198
  (
    n165,
    n39
  );


  buf
  g199
  (
    n467,
    n64
  );


  buf
  g200
  (
    n328,
    n83
  );


  not
  g201
  (
    n423,
    n56
  );


  not
  g202
  (
    n158,
    n77
  );


  not
  g203
  (
    n351,
    n71
  );


  not
  g204
  (
    n202,
    n56
  );


  buf
  g205
  (
    n332,
    n51
  );


  buf
  g206
  (
    n220,
    n74
  );


  not
  g207
  (
    n170,
    n66
  );


  not
  g208
  (
    n369,
    n95
  );


  not
  g209
  (
    n187,
    n111
  );


  not
  g210
  (
    n222,
    n85
  );


  buf
  g211
  (
    n236,
    n38
  );


  not
  g212
  (
    n311,
    n35
  );


  not
  g213
  (
    n490,
    n98
  );


  not
  g214
  (
    n229,
    n57
  );


  not
  g215
  (
    n278,
    n102
  );


  not
  g216
  (
    n156,
    n104
  );


  buf
  g217
  (
    n245,
    n81
  );


  buf
  g218
  (
    n396,
    n49
  );


  not
  g219
  (
    n329,
    n62
  );


  not
  g220
  (
    n414,
    n97
  );


  not
  g221
  (
    n447,
    n95
  );


  buf
  g222
  (
    n385,
    n106
  );


  buf
  g223
  (
    n390,
    n90
  );


  not
  g224
  (
    n294,
    n54
  );


  not
  g225
  (
    n234,
    n62
  );


  buf
  g226
  (
    n442,
    n96
  );


  not
  g227
  (
    n363,
    n34
  );


  not
  g228
  (
    n424,
    n67
  );


  not
  g229
  (
    n221,
    n33
  );


  not
  g230
  (
    n445,
    n39
  );


  buf
  g231
  (
    n218,
    n61
  );


  not
  g232
  (
    n200,
    n62
  );


  not
  g233
  (
    n183,
    n72
  );


  not
  g234
  (
    n392,
    n69
  );


  not
  g235
  (
    n365,
    n80
  );


  not
  g236
  (
    n456,
    n100
  );


  buf
  g237
  (
    n382,
    n105
  );


  buf
  g238
  (
    n320,
    n39
  );


  not
  g239
  (
    n429,
    n38
  );


  buf
  g240
  (
    n246,
    n64
  );


  not
  g241
  (
    n238,
    n115
  );


  not
  g242
  (
    n268,
    n60
  );


  not
  g243
  (
    n286,
    n54
  );


  not
  g244
  (
    n302,
    n113
  );


  not
  g245
  (
    n386,
    n34
  );


  buf
  g246
  (
    n336,
    n116
  );


  not
  g247
  (
    n345,
    n112
  );


  not
  g248
  (
    n160,
    n47
  );


  not
  g249
  (
    n251,
    n63
  );


  not
  g250
  (
    n151,
    n41
  );


  buf
  g251
  (
    n189,
    n53
  );


  buf
  g252
  (
    n168,
    n55
  );


  not
  g253
  (
    n287,
    n61
  );


  not
  g254
  (
    n283,
    n61
  );


  not
  g255
  (
    n341,
    n73
  );


  buf
  g256
  (
    n269,
    n35
  );


  not
  g257
  (
    n481,
    n41
  );


  buf
  g258
  (
    n157,
    n72
  );


  buf
  g259
  (
    n472,
    n39
  );


  not
  g260
  (
    n205,
    n99
  );


  buf
  g261
  (
    n449,
    n116
  );


  buf
  g262
  (
    n319,
    n107
  );


  not
  g263
  (
    n325,
    n60
  );


  not
  g264
  (
    n337,
    n90
  );


  buf
  g265
  (
    n487,
    n61
  );


  not
  g266
  (
    n259,
    n69
  );


  not
  g267
  (
    n391,
    n75
  );


  not
  g268
  (
    n398,
    n55
  );


  not
  g269
  (
    n179,
    n103
  );


  not
  g270
  (
    n413,
    n76
  );


  buf
  g271
  (
    n275,
    n94
  );


  not
  g272
  (
    n357,
    n96
  );


  not
  g273
  (
    n354,
    n52
  );


  not
  g274
  (
    n239,
    n76
  );


  not
  g275
  (
    n451,
    n65
  );


  not
  g276
  (
    n240,
    n59
  );


  buf
  g277
  (
    n203,
    n44
  );


  buf
  g278
  (
    n489,
    n46
  );


  not
  g279
  (
    n444,
    n97
  );


  not
  g280
  (
    n448,
    n40
  );


  not
  g281
  (
    n310,
    n55
  );


  not
  g282
  (
    n347,
    n107
  );


  not
  g283
  (
    n194,
    n101
  );


  not
  g284
  (
    n235,
    n93
  );


  not
  g285
  (
    n326,
    n63
  );


  buf
  g286
  (
    n373,
    n94
  );


  buf
  g287
  (
    n411,
    n91
  );


  buf
  g288
  (
    n314,
    n73
  );


  not
  g289
  (
    n291,
    n64
  );


  not
  g290
  (
    n334,
    n104
  );


  buf
  g291
  (
    n395,
    n64
  );


  not
  g292
  (
    n257,
    n99
  );


  buf
  g293
  (
    n217,
    n46
  );


  buf
  g294
  (
    n261,
    n52
  );


  buf
  g295
  (
    n409,
    n118
  );


  not
  g296
  (
    n255,
    n98
  );


  buf
  g297
  (
    n422,
    n110
  );


  not
  g298
  (
    n484,
    n91
  );


  buf
  g299
  (
    n214,
    n37
  );


  not
  g300
  (
    n273,
    n92
  );


  not
  g301
  (
    n228,
    n83
  );


  not
  g302
  (
    n152,
    n109
  );


  buf
  g303
  (
    n394,
    n38
  );


  not
  g304
  (
    n420,
    n96
  );


  not
  g305
  (
    n410,
    n51
  );


  not
  g306
  (
    n178,
    n99
  );


  not
  g307
  (
    n397,
    n80
  );


  not
  g308
  (
    n342,
    n54
  );


  buf
  g309
  (
    n208,
    n53
  );


  not
  g310
  (
    n233,
    n117
  );


  buf
  g311
  (
    n486,
    n76
  );


  not
  g312
  (
    n379,
    n93
  );


  buf
  g313
  (
    n209,
    n114
  );


  buf
  g314
  (
    n358,
    n78
  );


  buf
  g315
  (
    n321,
    n111
  );


  buf
  g316
  (
    n375,
    n33
  );


  buf
  g317
  (
    n457,
    n50
  );


  not
  g318
  (
    n348,
    n71
  );


  buf
  g319
  (
    n279,
    n60
  );


  not
  g320
  (
    n333,
    n92
  );


  not
  g321
  (
    n466,
    n70
  );


  not
  g322
  (
    n403,
    n67
  );


  buf
  g323
  (
    n212,
    n108
  );


  buf
  g324
  (
    n380,
    n95
  );


  not
  g325
  (
    n254,
    n46
  );


  buf
  g326
  (
    n437,
    n43
  );


  buf
  g327
  (
    n289,
    n35
  );


  buf
  g328
  (
    n312,
    n70
  );


  buf
  g329
  (
    n188,
    n99
  );


  buf
  g330
  (
    n197,
    n115
  );


  buf
  g331
  (
    n364,
    n100
  );


  buf
  g332
  (
    n404,
    n67
  );


  buf
  g333
  (
    n308,
    n106
  );


  buf
  g334
  (
    n473,
    n59
  );


  not
  g335
  (
    n339,
    n102
  );


  buf
  g336
  (
    n370,
    n65
  );


  buf
  g337
  (
    n253,
    n78
  );


  buf
  g338
  (
    n267,
    n34
  );


  buf
  g339
  (
    n482,
    n109
  );


  buf
  g340
  (
    n478,
    n77
  );


  buf
  g341
  (
    n182,
    n48
  );


  buf
  g342
  (
    n177,
    n57
  );


  not
  g343
  (
    n206,
    n86
  );


  not
  g344
  (
    n207,
    n113
  );


  not
  g345
  (
    n401,
    n82
  );


  buf
  g346
  (
    n159,
    n84
  );


  buf
  g347
  (
    n353,
    n66
  );


  buf
  g348
  (
    n262,
    n43
  );


  buf
  g349
  (
    n465,
    n105
  );


  not
  g350
  (
    n322,
    n78
  );


  buf
  g351
  (
    n476,
    n59
  );


  buf
  g352
  (
    n367,
    n83
  );


  buf
  g353
  (
    n434,
    n85
  );


  buf
  g354
  (
    n211,
    n102
  );


  not
  g355
  (
    n480,
    n103
  );


  not
  g356
  (
    n264,
    n105
  );


  not
  g357
  (
    n180,
    n78
  );


  buf
  g358
  (
    n366,
    n58
  );


  not
  g359
  (
    n469,
    n80
  );


  not
  g360
  (
    n393,
    n40
  );


  buf
  g361
  (
    n432,
    n86
  );


  not
  g362
  (
    n154,
    n76
  );


  not
  g363
  (
    n293,
    n91
  );


  buf
  g364
  (
    n149,
    n107
  );


  not
  g365
  (
    n226,
    n113
  );


  not
  g366
  (
    n468,
    n88
  );


  not
  g367
  (
    n305,
    n87
  );


  buf
  g368
  (
    n352,
    n79
  );


  buf
  g369
  (
    n303,
    n58
  );


  not
  g370
  (
    n318,
    n59
  );


  not
  g371
  (
    n462,
    n40
  );


  not
  g372
  (
    n356,
    n43
  );


  buf
  g373
  (
    n323,
    n51
  );


  not
  g374
  (
    n361,
    n41
  );


  not
  g375
  (
    n231,
    n40
  );


  not
  g376
  (
    n427,
    n67
  );


  not
  g377
  (
    n285,
    n56
  );


  buf
  g378
  (
    n435,
    n44
  );


  not
  g379
  (
    n150,
    n58
  );


  buf
  g380
  (
    n266,
    n82
  );


  not
  g381
  (
    n458,
    n79
  );


  not
  g382
  (
    n450,
    n57
  );


  buf
  g383
  (
    n176,
    n80
  );


  not
  g384
  (
    n299,
    n101
  );


  buf
  g385
  (
    n232,
    n88
  );


  buf
  g386
  (
    n263,
    n87
  );


  buf
  g387
  (
    n199,
    n57
  );


  buf
  g388
  (
    n174,
    n75
  );


  buf
  g389
  (
    n190,
    n84
  );


  buf
  g390
  (
    n297,
    n74
  );


  buf
  g391
  (
    n164,
    n84
  );


  not
  g392
  (
    n243,
    n69
  );


  buf
  g393
  (
    n455,
    n42
  );


  buf
  g394
  (
    n368,
    n33
  );


  not
  g395
  (
    n247,
    n117
  );


  buf
  g396
  (
    n439,
    n111
  );


  buf
  g397
  (
    n216,
    n48
  );


  not
  g398
  (
    n327,
    n45
  );


  not
  g399
  (
    n193,
    n96
  );


  not
  g400
  (
    n400,
    n110
  );


  buf
  g401
  (
    n184,
    n36
  );


  buf
  g402
  (
    n415,
    n83
  );


  buf
  g403
  (
    n374,
    n117
  );


  not
  g404
  (
    n282,
    n36
  );


  buf
  g405
  (
    n192,
    n98
  );


  buf
  g406
  (
    n418,
    n79
  );


  not
  g407
  (
    n230,
    n51
  );


  buf
  g408
  (
    n201,
    n108
  );


  buf
  g409
  (
    n213,
    n36
  );


  buf
  g410
  (
    n307,
    n100
  );


  not
  g411
  (
    n464,
    n102
  );


  buf
  g412
  (
    n407,
    n103
  );


  buf
  g413
  (
    n284,
    n93
  );


  buf
  g414
  (
    n316,
    n97
  );


  buf
  g415
  (
    n408,
    n45
  );


  not
  g416
  (
    n173,
    n55
  );


  buf
  g417
  (
    n249,
    n81
  );


  not
  g418
  (
    n362,
    n47
  );


  not
  g419
  (
    n215,
    n43
  );


  buf
  g420
  (
    n224,
    n49
  );


  not
  g421
  (
    n317,
    n90
  );


  not
  g422
  (
    n453,
    n103
  );


  not
  g423
  (
    n475,
    n86
  );


  not
  g424
  (
    n288,
    n109
  );


  buf
  g425
  (
    n433,
    n89
  );


  not
  g426
  (
    n372,
    n114
  );


  not
  g427
  (
    n399,
    n105
  );


  buf
  g428
  (
    n155,
    n74
  );


  not
  g429
  (
    n425,
    n53
  );


  buf
  g430
  (
    n470,
    n116
  );


  buf
  g431
  (
    n248,
    n63
  );


  buf
  g432
  (
    n360,
    n81
  );


  buf
  g433
  (
    n301,
    n118
  );


  not
  g434
  (
    n223,
    n108
  );


  buf
  g435
  (
    n381,
    n62
  );


  not
  g436
  (
    n488,
    n95
  );


  not
  g437
  (
    n171,
    n109
  );


  not
  g438
  (
    n270,
    n45
  );


  not
  g439
  (
    n227,
    n46
  );


  not
  g440
  (
    n454,
    n110
  );


  buf
  g441
  (
    n349,
    n42
  );


  not
  g442
  (
    n436,
    n50
  );


  buf
  g443
  (
    n479,
    n81
  );


  not
  g444
  (
    n198,
    n42
  );


  buf
  g445
  (
    n344,
    n37
  );


  buf
  g446
  (
    n419,
    n71
  );


  not
  g447
  (
    n306,
    n75
  );


  not
  g448
  (
    n161,
    n47
  );


  buf
  g449
  (
    n252,
    n56
  );


  not
  g450
  (
    n346,
    n107
  );


  not
  g451
  (
    n441,
    n112
  );


  not
  g452
  (
    n405,
    n94
  );


  not
  g453
  (
    n172,
    n47
  );


  not
  g454
  (
    n460,
    n53
  );


  buf
  g455
  (
    n459,
    n34
  );


  not
  g456
  (
    n377,
    n82
  );


  not
  g457
  (
    n250,
    n75
  );


  buf
  g458
  (
    n733,
    n289
  );


  buf
  g459
  (
    n575,
    n410
  );


  not
  g460
  (
    n594,
    n402
  );


  not
  g461
  (
    n516,
    n463
  );


  not
  g462
  (
    n623,
    n207
  );


  buf
  g463
  (
    n504,
    n231
  );


  buf
  g464
  (
    n546,
    n279
  );


  not
  g465
  (
    n551,
    n309
  );


  not
  g466
  (
    n672,
    n130
  );


  buf
  g467
  (
    n579,
    n165
  );


  not
  g468
  (
    n835,
    n418
  );


  not
  g469
  (
    n804,
    n328
  );


  buf
  g470
  (
    n653,
    n194
  );


  not
  g471
  (
    n659,
    n402
  );


  nor
  g472
  (
    n669,
    n176,
    n126,
    n311
  );


  nand
  g473
  (
    n513,
    n128,
    n405,
    n457,
    n390
  );


  or
  g474
  (
    n693,
    n227,
    n296,
    n418,
    n123
  );


  xnor
  g475
  (
    n825,
    n392,
    n378,
    n454,
    n443
  );


  nand
  g476
  (
    n592,
    n365,
    n374,
    n123,
    n342
  );


  xnor
  g477
  (
    n599,
    n379,
    n347,
    n415,
    n307
  );


  nor
  g478
  (
    n701,
    n431,
    n399,
    n345,
    n448
  );


  and
  g479
  (
    n529,
    n364,
    n263,
    n273,
    n217
  );


  or
  g480
  (
    n823,
    n250,
    n423,
    n449,
    n317
  );


  xor
  g481
  (
    n614,
    n243,
    n185,
    n222
  );


  nand
  g482
  (
    n637,
    n354,
    n280,
    n306,
    n409
  );


  nand
  g483
  (
    n617,
    n191,
    n142,
    n366,
    n160
  );


  and
  g484
  (
    n729,
    n437,
    n351,
    n320,
    n173
  );


  nand
  g485
  (
    n814,
    n184,
    n292,
    n275,
    n437
  );


  and
  g486
  (
    n709,
    n319,
    n410,
    n364,
    n421
  );


  nor
  g487
  (
    n522,
    n295,
    n137,
    n315,
    n455
  );


  nand
  g488
  (
    n569,
    n250,
    n188,
    n285,
    n284
  );


  xnor
  g489
  (
    n827,
    n150,
    n243,
    n184,
    n219
  );


  xnor
  g490
  (
    n536,
    n357,
    n324,
    n318,
    n287
  );


  and
  g491
  (
    n773,
    n211,
    n189,
    n456,
    n438
  );


  and
  g492
  (
    n567,
    n333,
    n215,
    n442,
    n163
  );


  and
  g493
  (
    n717,
    n369,
    n178,
    n459,
    n157
  );


  or
  g494
  (
    n721,
    n162,
    n372,
    n390,
    n376
  );


  xor
  g495
  (
    n616,
    n240,
    n340,
    n439,
    n453
  );


  and
  g496
  (
    n683,
    n275,
    n191,
    n452,
    n264
  );


  nor
  g497
  (
    n707,
    n127,
    n328,
    n318,
    n383
  );


  xor
  g498
  (
    n784,
    n119,
    n337,
    n359,
    n238
  );


  and
  g499
  (
    n615,
    n135,
    n385,
    n198,
    n159
  );


  and
  g500
  (
    n754,
    n237,
    n237,
    n138,
    n290
  );


  nor
  g501
  (
    n788,
    n360,
    n128,
    n219,
    n427
  );


  nor
  g502
  (
    n743,
    n197,
    n327,
    n408,
    n236
  );


  and
  g503
  (
    n571,
    n284,
    n204,
    n308,
    n235
  );


  nor
  g504
  (
    n620,
    n258,
    n198,
    n323,
    n281
  );


  and
  g505
  (
    n787,
    n310,
    n371,
    n386,
    n425
  );


  nand
  g506
  (
    n570,
    n454,
    n318,
    n333,
    n194
  );


  nand
  g507
  (
    n770,
    n374,
    n195,
    n142,
    n332
  );


  xnor
  g508
  (
    n526,
    n264,
    n316,
    n393,
    n372
  );


  or
  g509
  (
    n532,
    n351,
    n141,
    n275,
    n211
  );


  nand
  g510
  (
    n728,
    n261,
    n225,
    n449,
    n424
  );


  nand
  g511
  (
    n818,
    n290,
    n234,
    n356,
    n179
  );


  nand
  g512
  (
    n587,
    n234,
    n282,
    n176
  );


  xor
  g513
  (
    n657,
    n157,
    n184,
    n457,
    n188
  );


  xor
  g514
  (
    n673,
    n170,
    n165,
    n127,
    n432
  );


  or
  g515
  (
    n793,
    n314,
    n181,
    n174,
    n198
  );


  nand
  g516
  (
    n760,
    n441,
    n328,
    n370,
    n353
  );


  and
  g517
  (
    n766,
    n229,
    n344,
    n345,
    n442
  );


  nand
  g518
  (
    n745,
    n216,
    n444,
    n355,
    n323
  );


  and
  g519
  (
    n639,
    n316,
    n143,
    n420,
    n336
  );


  nor
  g520
  (
    n635,
    n153,
    n119,
    n461,
    n267
  );


  nand
  g521
  (
    n552,
    n406,
    n457,
    n318,
    n411
  );


  or
  g522
  (
    n736,
    n245,
    n426,
    n371,
    n374
  );


  xnor
  g523
  (
    n803,
    n317,
    n261,
    n395,
    n170
  );


  nand
  g524
  (
    n660,
    n288,
    n224,
    n451,
    n363
  );


  xor
  g525
  (
    n514,
    n139,
    n397,
    n272,
    n136
  );


  xor
  g526
  (
    n842,
    n426,
    n256,
    n189,
    n201
  );


  and
  g527
  (
    n578,
    n460,
    n358,
    n298,
    n151
  );


  nand
  g528
  (
    n649,
    n302,
    n356,
    n369,
    n403
  );


  nand
  g529
  (
    n624,
    n422,
    n245,
    n300,
    n215
  );


  xor
  g530
  (
    n663,
    n451,
    n316,
    n245,
    n186
  );


  nor
  g531
  (
    n506,
    n408,
    n163,
    n140,
    n173
  );


  xnor
  g532
  (
    n491,
    n254,
    n269,
    n443,
    n382
  );


  xnor
  g533
  (
    n824,
    n214,
    n136,
    n352,
    n181
  );


  or
  g534
  (
    n661,
    n226,
    n226,
    n258,
    n425
  );


  and
  g535
  (
    n613,
    n298,
    n158,
    n341,
    n230
  );


  xor
  g536
  (
    n518,
    n217,
    n393,
    n435,
    n200
  );


  nor
  g537
  (
    n610,
    n387,
    n459,
    n211,
    n413
  );


  nand
  g538
  (
    n727,
    n240,
    n259,
    n249,
    n357
  );


  xor
  g539
  (
    n688,
    n385,
    n369,
    n163,
    n306
  );


  xor
  g540
  (
    n495,
    n187,
    n131,
    n448,
    n168
  );


  nand
  g541
  (
    n682,
    n444,
    n436,
    n311,
    n297
  );


  or
  g542
  (
    n550,
    n461,
    n181,
    n367,
    n334
  );


  nor
  g543
  (
    n791,
    n263,
    n128,
    n347,
    n305
  );


  xnor
  g544
  (
    n515,
    n429,
    n445,
    n122,
    n359
  );


  xnor
  g545
  (
    n609,
    n127,
    n283,
    n321,
    n217
  );


  and
  g546
  (
    n805,
    n439,
    n438,
    n128,
    n252
  );


  nor
  g547
  (
    n564,
    n186,
    n391,
    n201,
    n250
  );


  and
  g548
  (
    n723,
    n334,
    n294,
    n420,
    n207
  );


  nand
  g549
  (
    n598,
    n149,
    n371,
    n377,
    n429
  );


  and
  g550
  (
    n815,
    n382,
    n229,
    n396,
    n418
  );


  and
  g551
  (
    n519,
    n327,
    n120,
    n313,
    n345
  );


  and
  g552
  (
    n811,
    n400,
    n160,
    n152
  );


  xnor
  g553
  (
    n744,
    n405,
    n313,
    n400,
    n459
  );


  xnor
  g554
  (
    n801,
    n139,
    n459,
    n264,
    n460
  );


  nand
  g555
  (
    n679,
    n305,
    n338,
    n381,
    n375
  );


  and
  g556
  (
    n535,
    n450,
    n405,
    n169,
    n232
  );


  nand
  g557
  (
    n528,
    n252,
    n143,
    n140,
    n441
  );


  xnor
  g558
  (
    n580,
    n219,
    n223,
    n398,
    n379
  );


  and
  g559
  (
    n530,
    n417,
    n322,
    n131,
    n151
  );


  or
  g560
  (
    n658,
    n337,
    n430,
    n413,
    n278
  );


  and
  g561
  (
    n525,
    n319,
    n298,
    n237,
    n150
  );


  xor
  g562
  (
    n700,
    n194,
    n289,
    n173,
    n221
  );


  xor
  g563
  (
    n675,
    n291,
    n453,
    n266,
    n153
  );


  xor
  g564
  (
    n554,
    n372,
    n121,
    n203,
    n355
  );


  and
  g565
  (
    n618,
    n224,
    n260,
    n390,
    n174
  );


  nand
  g566
  (
    n666,
    n263,
    n363,
    n376,
    n321
  );


  nand
  g567
  (
    n588,
    n379,
    n156,
    n266,
    n376
  );


  and
  g568
  (
    n605,
    n270,
    n416,
    n401,
    n463
  );


  or
  g569
  (
    n668,
    n320,
    n299,
    n350,
    n272
  );


  and
  g570
  (
    n544,
    n319,
    n416,
    n387,
    n126
  );


  or
  g571
  (
    n769,
    n388,
    n346,
    n368,
    n389
  );


  xnor
  g572
  (
    n708,
    n248,
    n269,
    n320,
    n296
  );


  or
  g573
  (
    n547,
    n229,
    n368,
    n389,
    n167
  );


  xor
  g574
  (
    n549,
    n449,
    n347,
    n161,
    n215
  );


  and
  g575
  (
    n589,
    n202,
    n361,
    n253,
    n404
  );


  and
  g576
  (
    n566,
    n431,
    n291,
    n362,
    n283
  );


  and
  g577
  (
    n630,
    n182,
    n154,
    n407,
    n163
  );


  nand
  g578
  (
    n507,
    n243,
    n296,
    n378,
    n452
  );


  nand
  g579
  (
    n795,
    n174,
    n299,
    n213,
    n232
  );


  nor
  g580
  (
    n565,
    n196,
    n274,
    n187,
    n289
  );


  xor
  g581
  (
    n493,
    n461,
    n204,
    n230,
    n450
  );


  xnor
  g582
  (
    n828,
    n150,
    n434,
    n346,
    n212
  );


  nor
  g583
  (
    n636,
    n412,
    n134,
    n439,
    n301
  );


  and
  g584
  (
    n541,
    n152,
    n206,
    n351,
    n155
  );


  and
  g585
  (
    n762,
    n352,
    n120,
    n341,
    n382
  );


  xnor
  g586
  (
    n687,
    n303,
    n187,
    n140,
    n449
  );


  xnor
  g587
  (
    n799,
    n236,
    n388,
    n189,
    n363
  );


  xor
  g588
  (
    n591,
    n122,
    n404,
    n217,
    n222
  );


  or
  g589
  (
    n523,
    n252,
    n322,
    n422,
    n291
  );


  or
  g590
  (
    n832,
    n370,
    n360,
    n129,
    n440
  );


  nand
  g591
  (
    n511,
    n279,
    n339,
    n314,
    n286
  );


  nor
  g592
  (
    n557,
    n266,
    n435,
    n279,
    n228
  );


  xnor
  g593
  (
    n582,
    n402,
    n244,
    n255,
    n311
  );


  nand
  g594
  (
    n713,
    n280,
    n190,
    n357,
    n287
  );


  and
  g595
  (
    n667,
    n407,
    n218,
    n221,
    n377
  );


  and
  g596
  (
    n711,
    n268,
    n313,
    n336,
    n462
  );


  and
  g597
  (
    n619,
    n342,
    n303,
    n204,
    n247
  );


  nand
  g598
  (
    n771,
    n141,
    n285,
    n200,
    n359
  );


  xor
  g599
  (
    n735,
    n338,
    n192,
    n406,
    n314
  );


  or
  g600
  (
    n689,
    n118,
    n423,
    n246,
    n260
  );


  xor
  g601
  (
    n696,
    n229,
    n430,
    n325,
    n349
  );


  and
  g602
  (
    n739,
    n200,
    n271,
    n144,
    n391
  );


  xor
  g603
  (
    n524,
    n219,
    n171,
    n391,
    n142
  );


  xor
  g604
  (
    n782,
    n189,
    n282,
    n187,
    n417
  );


  xor
  g605
  (
    n819,
    n193,
    n237,
    n225,
    n197
  );


  xnor
  g606
  (
    n656,
    n133,
    n232,
    n284,
    n412
  );


  xnor
  g607
  (
    n662,
    n394,
    n253,
    n170,
    n368
  );


  xnor
  g608
  (
    n652,
    n243,
    n132,
    n302,
    n195
  );


  nor
  g609
  (
    n645,
    n268,
    n227,
    n425,
    n166
  );


  nand
  g610
  (
    n840,
    n144,
    n415,
    n262,
    n276
  );


  and
  g611
  (
    n545,
    n440,
    n438,
    n166,
    n124
  );


  xnor
  g612
  (
    n562,
    n337,
    n168,
    n336,
    n210
  );


  or
  g613
  (
    n703,
    n339,
    n373,
    n392,
    n435
  );


  nor
  g614
  (
    n521,
    n433,
    n335,
    n201,
    n209
  );


  or
  g615
  (
    n698,
    n216,
    n423,
    n279,
    n383
  );


  nor
  g616
  (
    n633,
    n350,
    n261,
    n445,
    n253
  );


  and
  g617
  (
    n642,
    n155,
    n238,
    n314,
    n276
  );


  nor
  g618
  (
    n671,
    n215,
    n218,
    n278,
    n349
  );


  or
  g619
  (
    n500,
    n142,
    n188,
    n307,
    n248
  );


  xor
  g620
  (
    n681,
    n131,
    n406,
    n185,
    n329
  );


  nand
  g621
  (
    n759,
    n292,
    n418,
    n207,
    n428
  );


  nand
  g622
  (
    n830,
    n285,
    n305,
    n458,
    n380
  );


  xnor
  g623
  (
    n699,
    n348,
    n190,
    n233,
    n331
  );


  and
  g624
  (
    n563,
    n366,
    n358,
    n143,
    n132
  );


  xnor
  g625
  (
    n680,
    n119,
    n233,
    n230,
    n201
  );


  xor
  g626
  (
    n691,
    n133,
    n289,
    n386,
    n188
  );


  and
  g627
  (
    n765,
    n427,
    n293,
    n316,
    n436
  );


  xnor
  g628
  (
    n593,
    n393,
    n387,
    n450,
    n180
  );


  and
  g629
  (
    n806,
    n137,
    n294,
    n267,
    n446
  );


  nand
  g630
  (
    n737,
    n307,
    n420,
    n228,
    n421
  );


  nand
  g631
  (
    n749,
    n424,
    n456,
    n249,
    n395
  );


  xnor
  g632
  (
    n585,
    n342,
    n238,
    n358,
    n183
  );


  nor
  g633
  (
    n790,
    n356,
    n406,
    n265,
    n330
  );


  xor
  g634
  (
    n738,
    n277,
    n247,
    n137,
    n203
  );


  nor
  g635
  (
    n752,
    n234,
    n305,
    n399,
    n304
  );


  or
  g636
  (
    n651,
    n259,
    n296,
    n138,
    n199
  );


  xnor
  g637
  (
    n779,
    n306,
    n145,
    n401,
    n235
  );


  xnor
  g638
  (
    n692,
    n422,
    n274,
    n239,
    n151
  );


  xnor
  g639
  (
    n503,
    n281,
    n361,
    n440,
    n400
  );


  nand
  g640
  (
    n785,
    n267,
    n455,
    n249,
    n248
  );


  nand
  g641
  (
    n542,
    n177,
    n274,
    n303,
    n162
  );


  and
  g642
  (
    n494,
    n401,
    n149,
    n389,
    n276
  );


  xnor
  g643
  (
    n750,
    n231,
    n213,
    n355,
    n170
  );


  and
  g644
  (
    n686,
    n343,
    n433,
    n425,
    n302
  );


  xnor
  g645
  (
    n628,
    n233,
    n417,
    n414,
    n180
  );


  xor
  g646
  (
    n600,
    n335,
    n412,
    n210,
    n132
  );


  or
  g647
  (
    n757,
    n384,
    n202,
    n339,
    n319
  );


  nor
  g648
  (
    n724,
    n443,
    n178,
    n144,
    n411
  );


  nor
  g649
  (
    n556,
    n227,
    n295,
    n446,
    n152
  );


  nor
  g650
  (
    n577,
    n438,
    n277,
    n445,
    n169
  );


  nand
  g651
  (
    n809,
    n285,
    n356,
    n302,
    n138
  );


  nand
  g652
  (
    n626,
    n192,
    n136,
    n159,
    n221
  );


  xnor
  g653
  (
    n670,
    n360,
    n327,
    n220,
    n136
  );


  xor
  g654
  (
    n751,
    n254,
    n365,
    n336,
    n157
  );


  nor
  g655
  (
    n621,
    n323,
    n268,
    n368,
    n446
  );


  and
  g656
  (
    n798,
    n190,
    n197,
    n378,
    n431
  );


  nand
  g657
  (
    n706,
    n282,
    n326,
    n392,
    n145
  );


  and
  g658
  (
    n810,
    n442,
    n258,
    n447,
    n451
  );


  nor
  g659
  (
    n820,
    n390,
    n123,
    n154,
    n360
  );


  nor
  g660
  (
    n634,
    n294,
    n396,
    n301,
    n175
  );


  nor
  g661
  (
    n789,
    n329,
    n309,
    n444,
    n455
  );


  or
  g662
  (
    n539,
    n304,
    n265,
    n164,
    n172
  );


  or
  g663
  (
    n627,
    n426,
    n135,
    n242,
    n140
  );


  and
  g664
  (
    n641,
    n199,
    n165,
    n378,
    n206
  );


  xor
  g665
  (
    n838,
    n286,
    n387,
    n416,
    n220
  );


  nor
  g666
  (
    n796,
    n269,
    n408,
    n162,
    n153
  );


  xnor
  g667
  (
    n677,
    n317,
    n295,
    n236,
    n332
  );


  and
  g668
  (
    n829,
    n263,
    n343,
    n240,
    n130
  );


  xnor
  g669
  (
    n761,
    n386,
    n315,
    n311,
    n177
  );


  xnor
  g670
  (
    n568,
    n164,
    n251,
    n185,
    n376
  );


  or
  g671
  (
    n697,
    n396,
    n177,
    n432,
    n191
  );


  nor
  g672
  (
    n548,
    n179,
    n431,
    n380,
    n423
  );


  nand
  g673
  (
    n501,
    n242,
    n195,
    n340,
    n450
  );


  nor
  g674
  (
    n678,
    n238,
    n380,
    n293,
    n176
  );


  nor
  g675
  (
    n802,
    n297,
    n435,
    n426,
    n456
  );


  or
  g676
  (
    n543,
    n324,
    n172,
    n458,
    n270
  );


  nand
  g677
  (
    n538,
    n228,
    n404,
    n299,
    n150
  );


  and
  g678
  (
    n684,
    n299,
    n278,
    n403,
    n375
  );


  nor
  g679
  (
    n622,
    n358,
    n329,
    n132,
    n137
  );


  nor
  g680
  (
    n775,
    n224,
    n326,
    n381,
    n421
  );


  xnor
  g681
  (
    n643,
    n239,
    n331,
    n246,
    n380
  );


  and
  g682
  (
    n772,
    n462,
    n312,
    n382,
    n164
  );


  and
  g683
  (
    n517,
    n166,
    n354,
    n208,
    n452
  );


  or
  g684
  (
    n734,
    n300,
    n199,
    n192,
    n256
  );


  xor
  g685
  (
    n647,
    n151,
    n121,
    n347,
    n286
  );


  nor
  g686
  (
    n822,
    n171,
    n153,
    n265,
    n428
  );


  nor
  g687
  (
    n755,
    n293,
    n182,
    n350,
    n255
  );


  and
  g688
  (
    n590,
    n275,
    n271,
    n283,
    n396
  );


  or
  g689
  (
    n774,
    n362,
    n144,
    n260,
    n127
  );


  or
  g690
  (
    n581,
    n287,
    n309,
    n308,
    n220
  );


  nor
  g691
  (
    n715,
    n301,
    n264,
    n257,
    n134
  );


  nor
  g692
  (
    n797,
    n191,
    n421,
    n135,
    n366
  );


  xor
  g693
  (
    n502,
    n444,
    n304,
    n303,
    n167
  );


  and
  g694
  (
    n595,
    n411,
    n443,
    n227,
    n448
  );


  nor
  g695
  (
    n586,
    n291,
    n436,
    n241,
    n442
  );


  xnor
  g696
  (
    n654,
    n205,
    n175,
    n255,
    n218
  );


  xnor
  g697
  (
    n740,
    n301,
    n209,
    n258,
    n414
  );


  nor
  g698
  (
    n821,
    n293,
    n331,
    n326,
    n129
  );


  xnor
  g699
  (
    n718,
    n274,
    n413,
    n174,
    n180
  );


  xor
  g700
  (
    n836,
    n175,
    n181,
    n462,
    n411
  );


  and
  g701
  (
    n533,
    n412,
    n131,
    n461,
    n306
  );


  nand
  g702
  (
    n510,
    n246,
    n397,
    n434,
    n367
  );


  and
  g703
  (
    n674,
    n122,
    n119,
    n143,
    n460
  );


  nor
  g704
  (
    n492,
    n394,
    n139,
    n255,
    n428
  );


  nor
  g705
  (
    n572,
    n185,
    n300,
    n216,
    n434
  );


  xnor
  g706
  (
    n531,
    n180,
    n308,
    n122,
    n254
  );


  nor
  g707
  (
    n534,
    n231,
    n224,
    n353,
    n197
  );


  xor
  g708
  (
    n690,
    n251,
    n310,
    n177,
    n343
  );


  nor
  g709
  (
    n527,
    n451,
    n196,
    n292,
    n322
  );


  nor
  g710
  (
    n640,
    n400,
    n226,
    n337,
    n329
  );


  nor
  g711
  (
    n625,
    n300,
    n212,
    n354,
    n343
  );


  xnor
  g712
  (
    n509,
    n242,
    n398,
    n183,
    n440
  );


  xor
  g713
  (
    n747,
    n424,
    n458,
    n355,
    n262
  );


  nand
  g714
  (
    n753,
    n365,
    n298,
    n159,
    n161
  );


  nor
  g715
  (
    n608,
    n167,
    n156,
    n335,
    n130
  );


  or
  g716
  (
    n748,
    n214,
    n330,
    n223,
    n362
  );


  nor
  g717
  (
    n646,
    n193,
    n322,
    n377
  );


  or
  g718
  (
    n732,
    n138,
    n182,
    n341,
    n348
  );


  nor
  g719
  (
    n596,
    n383,
    n272,
    n453,
    n164
  );


  nor
  g720
  (
    n722,
    n231,
    n371,
    n359,
    n269
  );


  nand
  g721
  (
    n758,
    n346,
    n447,
    n179,
    n169
  );


  or
  g722
  (
    n720,
    n251,
    n364,
    n385,
    n367
  );


  and
  g723
  (
    n574,
    n419,
    n309,
    n134,
    n233
  );


  xnor
  g724
  (
    n655,
    n208,
    n384,
    n325,
    n157
  );


  or
  g725
  (
    n555,
    n235,
    n453,
    n141,
    n308
  );


  nand
  g726
  (
    n781,
    n253,
    n324,
    n391,
    n272
  );


  xor
  g727
  (
    n611,
    n121,
    n340,
    n433,
    n152
  );


  and
  g728
  (
    n560,
    n344,
    n349,
    n433,
    n333
  );


  xnor
  g729
  (
    n764,
    n247,
    n288,
    n419
  );


  nand
  g730
  (
    n712,
    n161,
    n245,
    n198,
    n430
  );


  and
  g731
  (
    n583,
    n381,
    n210,
    n256,
    n211
  );


  xnor
  g732
  (
    n710,
    n458,
    n385,
    n464,
    n193
  );


  xor
  g733
  (
    n606,
    n402,
    n405,
    n196,
    n214
  );


  and
  g734
  (
    n794,
    n234,
    n203,
    n373,
    n429
  );


  xor
  g735
  (
    n508,
    n280,
    n206,
    n168,
    n395
  );


  nand
  g736
  (
    n792,
    n236,
    n447,
    n248,
    n249
  );


  or
  g737
  (
    n839,
    n434,
    n124,
    n246,
    n325
  );


  and
  g738
  (
    n786,
    n394,
    n221,
    n125,
    n213
  );


  xnor
  g739
  (
    n714,
    n223,
    n171,
    n257,
    n375
  );


  nor
  g740
  (
    n597,
    n353,
    n313,
    n158,
    n321
  );


  nand
  g741
  (
    n837,
    n126,
    n262,
    n348,
    n195
  );


  xor
  g742
  (
    n576,
    n184,
    n398,
    n222,
    n339
  );


  xnor
  g743
  (
    n780,
    n410,
    n183,
    n186,
    n407
  );


  nor
  g744
  (
    n665,
    n439,
    n284,
    n280,
    n134
  );


  xor
  g745
  (
    n612,
    n330,
    n327,
    n403,
    n125
  );


  nor
  g746
  (
    n632,
    n244,
    n352,
    n315,
    n172
  );


  xnor
  g747
  (
    n741,
    n341,
    n230,
    n190,
    n204
  );


  xor
  g748
  (
    n763,
    n383,
    n205,
    n266,
    n323
  );


  xor
  g749
  (
    n843,
    n178,
    n139,
    n363,
    n398
  );


  xnor
  g750
  (
    n498,
    n273,
    n209,
    n457,
    n365
  );


  nor
  g751
  (
    n584,
    n235,
    n123,
    n321,
    n373
  );


  xnor
  g752
  (
    n685,
    n239,
    n155,
    n388,
    n214
  );


  xnor
  g753
  (
    n631,
    n397,
    n463,
    n349,
    n270
  );


  nand
  g754
  (
    n812,
    n312,
    n294,
    n257,
    n125
  );


  and
  g755
  (
    n676,
    n283,
    n118,
    n361,
    n352
  );


  nor
  g756
  (
    n834,
    n166,
    n307,
    n448,
    n346
  );


  or
  g757
  (
    n813,
    n158,
    n437,
    n415,
    n121
  );


  nor
  g758
  (
    n704,
    n392,
    n129,
    n428
  );


  and
  g759
  (
    n520,
    n460,
    n193,
    n455,
    n281
  );


  xnor
  g760
  (
    n831,
    n397,
    n270,
    n427
  );


  xnor
  g761
  (
    n817,
    n202,
    n286,
    n271,
    n209
  );


  nor
  g762
  (
    n731,
    n162,
    n159,
    n141,
    n218
  );


  nand
  g763
  (
    n730,
    n432,
    n277,
    n344,
    n192
  );


  xnor
  g764
  (
    n756,
    n429,
    n273,
    n216,
    n342
  );


  nand
  g765
  (
    n768,
    n384,
    n331,
    n401,
    n315
  );


  nand
  g766
  (
    n783,
    n364,
    n271,
    n292,
    n223
  );


  nor
  g767
  (
    n650,
    n367,
    n208,
    n145,
    n415
  );


  xor
  g768
  (
    n629,
    n332,
    n156,
    n297,
    n247
  );


  nand
  g769
  (
    n702,
    n165,
    n374,
    n437,
    n179
  );


  nor
  g770
  (
    n499,
    n244,
    n409,
    n447,
    n175
  );


  or
  g771
  (
    n833,
    n194,
    n454,
    n261,
    n370
  );


  xor
  g772
  (
    n776,
    n333,
    n332,
    n133,
    n203
  );


  xnor
  g773
  (
    n694,
    n196,
    n155,
    n372,
    n254
  );


  or
  g774
  (
    n644,
    n259,
    n420,
    n220,
    n265
  );


  nor
  g775
  (
    n767,
    n357,
    n369,
    n171,
    n409
  );


  xnor
  g776
  (
    n559,
    n176,
    n242,
    n154,
    n133
  );


  and
  g777
  (
    n725,
    n256,
    n225,
    n407,
    n317
  );


  nand
  g778
  (
    n726,
    n335,
    n403,
    n430,
    n172
  );


  xnor
  g779
  (
    n777,
    n169,
    n257,
    n158,
    n324
  );


  nor
  g780
  (
    n778,
    n202,
    n240,
    n445,
    n409
  );


  xor
  g781
  (
    n601,
    n239,
    n441,
    n334,
    n379
  );


  xnor
  g782
  (
    n603,
    n416,
    n161,
    n232,
    n168
  );


  xnor
  g783
  (
    n496,
    n373,
    n205,
    n199,
    n226
  );


  xor
  g784
  (
    n540,
    n208,
    n393,
    n320,
    n399
  );


  nand
  g785
  (
    n695,
    n381,
    n395,
    n375,
    n135
  );


  nor
  g786
  (
    n742,
    n250,
    n419,
    n212,
    n326
  );


  or
  g787
  (
    n841,
    n340,
    n278,
    n334,
    n251
  );


  xor
  g788
  (
    n573,
    n344,
    n312,
    n244,
    n384
  );


  xor
  g789
  (
    n561,
    n210,
    n160,
    n124,
    n297
  );


  or
  g790
  (
    n719,
    n178,
    n173,
    n432,
    n441
  );


  xor
  g791
  (
    n602,
    n312,
    n125,
    n213,
    n281
  );


  nor
  g792
  (
    n553,
    n345,
    n295,
    n354,
    n462
  );


  or
  g793
  (
    n558,
    n205,
    n225,
    n328,
    n304
  );


  xor
  g794
  (
    n807,
    n290,
    n414,
    n241,
    n386
  );


  nor
  g795
  (
    n648,
    n463,
    n273,
    n353,
    n351
  );


  nor
  g796
  (
    n607,
    n424,
    n130,
    n241,
    n389
  );


  and
  g797
  (
    n826,
    n370,
    n446,
    n252,
    n408
  );


  xor
  g798
  (
    n800,
    n456,
    n212,
    n413,
    n330
  );


  nor
  g799
  (
    n664,
    n149,
    n350,
    n325,
    n419
  );


  nand
  g800
  (
    n705,
    n156,
    n200,
    n338,
    n120
  );


  and
  g801
  (
    n746,
    n366,
    n126,
    n267,
    n186
  );


  xor
  g802
  (
    n497,
    n404,
    n436,
    n277,
    n310
  );


  nand
  g803
  (
    n808,
    n290,
    n454,
    n259,
    n452
  );


  xnor
  g804
  (
    n816,
    n120,
    n417,
    n414,
    n348
  );


  nand
  g805
  (
    n604,
    n228,
    n310,
    n394,
    n422
  );


  and
  g806
  (
    n512,
    n207,
    n287,
    n268,
    n399
  );


  and
  g807
  (
    n537,
    n260,
    n167,
    n288,
    n241
  );


  or
  g808
  (
    n505,
    n182,
    n124,
    n338,
    n410
  );


  nand
  g809
  (
    n716,
    n262,
    n276,
    n183,
    n388
  );


  and
  g810
  (
    n638,
    n154,
    n362,
    n206,
    n361
  );


  not
  g811
  (
    n846,
    n495
  );


  not
  g812
  (
    n854,
    n493
  );


  not
  g813
  (
    n853,
    n492
  );


  not
  g814
  (
    n855,
    n147
  );


  not
  g815
  (
    n848,
    n496
  );


  buf
  g816
  (
    n852,
    n494
  );


  and
  g817
  (
    n850,
    n146,
    n145
  );


  xnor
  g818
  (
    n845,
    n146,
    n146,
    n492,
    n491
  );


  nand
  g819
  (
    n851,
    n494,
    n146,
    n491
  );


  or
  g820
  (
    n849,
    n494,
    n495,
    n491,
    n493
  );


  xnor
  g821
  (
    n847,
    n493,
    n495,
    n494,
    n147
  );


  nand
  g822
  (
    n844,
    n492,
    n492,
    n493,
    n495
  );


  buf
  g823
  (
    n857,
    n844
  );


  not
  g824
  (
    n856,
    n844
  );


  or
  g825
  (
    n865,
    n496,
    n501,
    n499,
    n857
  );


  xnor
  g826
  (
    n864,
    n857,
    n497,
    n500,
    n501
  );


  nor
  g827
  (
    n862,
    n856,
    n498,
    n499
  );


  xnor
  g828
  (
    n859,
    n502,
    n501,
    n857,
    n856
  );


  and
  g829
  (
    n863,
    n497,
    n499,
    n857,
    n500
  );


  nor
  g830
  (
    n860,
    n497,
    n499,
    n501,
    n496
  );


  or
  g831
  (
    n861,
    n500,
    n497,
    n498
  );


  nor
  g832
  (
    n858,
    n500,
    n856,
    n496
  );


  nand
  g833
  (
    n869,
    n863,
    n466,
    n862,
    n470
  );


  nor
  g834
  (
    n880,
    n477,
    n480,
    n861,
    n482
  );


  nor
  g835
  (
    n876,
    n465,
    n476,
    n472
  );


  xor
  g836
  (
    n885,
    n474,
    n479,
    n470,
    n859
  );


  xnor
  g837
  (
    n867,
    n860,
    n844,
    n476,
    n467
  );


  and
  g838
  (
    n878,
    n859,
    n477,
    n863,
    n464
  );


  xnor
  g839
  (
    n870,
    n466,
    n465,
    n481,
    n464
  );


  xnor
  g840
  (
    n872,
    n478,
    n473,
    n845,
    n468
  );


  and
  g841
  (
    n881,
    n469,
    n478,
    n473,
    n863
  );


  xnor
  g842
  (
    n891,
    n474,
    n860,
    n479,
    n862
  );


  and
  g843
  (
    n879,
    n471,
    n475,
    n858,
    n478
  );


  and
  g844
  (
    n887,
    n481,
    n468,
    n861,
    n471
  );


  xor
  g845
  (
    n888,
    n480,
    n858,
    n470,
    n859
  );


  and
  g846
  (
    n875,
    n863,
    n469,
    n478
  );


  or
  g847
  (
    n877,
    n467,
    n858,
    n862,
    n469
  );


  nand
  g848
  (
    n874,
    n481,
    n468,
    n472,
    n473
  );


  nor
  g849
  (
    AntiSAT_key_wire,
    n466,
    n480,
    n471,
    n864
  );


  xnor
  g850
  (
    n883,
    n846,
    n465,
    n482,
    n858
  );


  and
  g851
  (
    n889,
    n859,
    n477,
    n860,
    n861
  );


  or
  g852
  (
    n884,
    n845,
    n475,
    n481,
    n476
  );


  xnor
  g853
  (
    n868,
    n864,
    n482,
    n475,
    n474
  );


  nor
  g854
  (
    n890,
    n466,
    n482,
    n479,
    n477
  );


  xor
  g855
  (
    n886,
    n861,
    n471,
    n845,
    n480
  );


  xor
  g856
  (
    n871,
    n472,
    n475,
    n465,
    n470
  );


  nor
  g857
  (
    n866,
    n479,
    n472,
    n860,
    n464
  );


  nor
  g858
  (
    n892,
    n473,
    n474,
    n467
  );


  or
  g859
  (
    n873,
    n862,
    n468,
    n845,
    n864
  );


  xor
  g860
  (
    n893,
    n504,
    n502,
    n503
  );


  nand
  g861
  (
    n896,
    n886,
    n883,
    n503,
    n502
  );


  nand
  g862
  (
    n895,
    n505,
    n503,
    n884,
    n504
  );


  or
  g863
  (
    n894,
    n885,
    n504,
    n502
  );


  xor
  g864
  (
    n911,
    n507,
    n895,
    n511,
    n847
  );


  and
  g865
  (
    n898,
    n893,
    n509,
    n505,
    n510
  );


  xnor
  g866
  (
    n900,
    n508,
    n513,
    n864,
    n846
  );


  or
  g867
  (
    n906,
    n893,
    n512,
    n894
  );


  xor
  g868
  (
    n901,
    n509,
    n508,
    n506,
    n896
  );


  nand
  g869
  (
    n910,
    n511,
    n847,
    n512,
    n846
  );


  and
  g870
  (
    n899,
    n508,
    n507,
    n505,
    n895
  );


  and
  g871
  (
    n897,
    n894,
    n896,
    n847,
    n506
  );


  or
  g872
  (
    n907,
    n846,
    n894,
    n847
  );


  and
  g873
  (
    n905,
    n509,
    n506,
    n514,
    n513
  );


  or
  g874
  (
    n909,
    n510,
    n893,
    n512,
    n895
  );


  nor
  g875
  (
    n902,
    n513,
    n895,
    n509,
    n507
  );


  nor
  g876
  (
    n908,
    n893,
    n896,
    n505,
    n510
  );


  and
  g877
  (
    n903,
    n511,
    n510,
    n508,
    n507
  );


  xnor
  g878
  (
    n904,
    n514,
    n513,
    n511,
    n506
  );


  or
  g879
  (
    n916,
    n515,
    n517,
    n514
  );


  xnor
  g880
  (
    n917,
    n515,
    n518,
    n899
  );


  nand
  g881
  (
    n912,
    n901,
    n515,
    n516,
    n902
  );


  nand
  g882
  (
    n915,
    n515,
    n516,
    n900,
    n518
  );


  xnor
  g883
  (
    n914,
    n517,
    n516,
    n518,
    n898
  );


  nor
  g884
  (
    n913,
    n517,
    n897,
    n516,
    n514
  );


  not
  g885
  (
    n919,
    n915
  );


  not
  g886
  (
    n918,
    n913
  );


  buf
  g887
  (
    n920,
    n914
  );


  not
  g888
  (
    n921,
    n915
  );


  not
  g889
  (
    n922,
    n919
  );


  not
  g890
  (
    n932,
    n907
  );


  buf
  g891
  (
    n928,
    n921
  );


  not
  g892
  (
    n924,
    n918
  );


  buf
  g893
  (
    n923,
    n848
  );


  buf
  g894
  (
    n936,
    n920
  );


  or
  g895
  (
    n930,
    n904,
    n865
  );


  nor
  g896
  (
    n933,
    n908,
    n920
  );


  or
  g897
  (
    n935,
    n849,
    n918,
    n865,
    n919
  );


  nor
  g898
  (
    n934,
    n921,
    n919,
    n848,
    n905
  );


  xor
  g899
  (
    n931,
    n887,
    n889,
    n920,
    n921
  );


  nor
  g900
  (
    n925,
    n910,
    n888,
    n849,
    n918
  );


  xnor
  g901
  (
    n926,
    n919,
    n918,
    n850,
    n849
  );


  nor
  g902
  (
    n927,
    n890,
    n909,
    n891,
    n921
  );


  xor
  g903
  (
    n937,
    n920,
    n906,
    n865,
    n850
  );


  or
  g904
  (
    n929,
    n849,
    n903,
    n848
  );


  buf
  g905
  (
    n941,
    n923
  );


  not
  g906
  (
    n939,
    n922
  );


  not
  g907
  (
    n940,
    n922
  );


  buf
  g908
  (
    n942,
    n922
  );


  not
  g909
  (
    n938,
    n923
  );


  xnor
  g910
  (
    n943,
    n922,
    n519,
    n916
  );


  not
  g911
  (
    n946,
    n911
  );


  not
  g912
  (
    n958,
    n923
  );


  buf
  g913
  (
    n947,
    n943
  );


  buf
  g914
  (
    n957,
    n850
  );


  buf
  g915
  (
    n952,
    n939
  );


  buf
  g916
  (
    n955,
    n924
  );


  not
  g917
  (
    n950,
    n943
  );


  not
  g918
  (
    n949,
    n519
  );


  not
  g919
  (
    n954,
    n940
  );


  not
  g920
  (
    n948,
    n938
  );


  buf
  g921
  (
    n951,
    n940
  );


  nand
  g922
  (
    n944,
    n520,
    n942,
    n943
  );


  nand
  g923
  (
    n953,
    n911,
    n923,
    n942,
    n943
  );


  nand
  g924
  (
    n956,
    n939,
    n942,
    n941
  );


  nand
  g925
  (
    n945,
    n924,
    n519,
    n942
  );


  nor
  g926
  (
    n961,
    n927,
    n945,
    n924,
    n926
  );


  xor
  g927
  (
    n959,
    n928,
    n944,
    n926
  );


  nor
  g928
  (
    n963,
    n944,
    n925,
    n927
  );


  and
  g929
  (
    n960,
    n924,
    n925,
    n927
  );


  xnor
  g930
  (
    n962,
    n926,
    n944,
    n927
  );


  nor
  g931
  (
    n968,
    n961,
    n865,
    n948,
    n960
  );


  nand
  g932
  (
    n969,
    n962,
    n950,
    n951
  );


  and
  g933
  (
    n967,
    n947,
    n916,
    n946,
    n960
  );


  xor
  g934
  (
    n966,
    n950,
    n945,
    n949,
    n962
  );


  nor
  g935
  (
    n964,
    n950,
    n948,
    n961,
    n949
  );


  nand
  g936
  (
    n972,
    n945,
    n946,
    n948,
    n949
  );


  nand
  g937
  (
    n965,
    n951,
    n945,
    n946
  );


  xor
  g938
  (
    n970,
    n959,
    n947,
    n963
  );


  and
  g939
  (
    n971,
    n949,
    n947,
    n948
  );


  not
  g940
  (
    n981,
    n968
  );


  buf
  g941
  (
    n978,
    n967
  );


  not
  g942
  (
    n974,
    n970
  );


  not
  g943
  (
    n983,
    n929
  );


  not
  g944
  (
    n982,
    n969
  );


  not
  g945
  (
    n980,
    n970
  );


  not
  g946
  (
    n984,
    n928
  );


  buf
  g947
  (
    n979,
    n929
  );


  not
  g948
  (
    n976,
    n964
  );


  buf
  g949
  (
    n977,
    n971
  );


  or
  g950
  (
    n975,
    n968,
    n965,
    n969,
    n966
  );


  xnor
  g951
  (
    n973,
    n929,
    n967,
    n928
  );


  nor
  g952
  (
    n985,
    n929,
    n973
  );


  xnor
  g953
  (
    n986,
    n951,
    n985,
    n952
  );


  nand
  g954
  (
    n987,
    n985,
    n951,
    n520
  );


  nand
  g955
  (
    n988,
    n523,
    n973,
    n987,
    n520
  );


  xnor
  g956
  (
    n989,
    n987,
    n522,
    n523
  );


  nor
  g957
  (
    n990,
    n973,
    n522,
    n986,
    n521
  );


  or
  g958
  (
    n992,
    n986,
    n521,
    n987
  );


  xor
  g959
  (
    n991,
    n523,
    n521,
    n522
  );


  xnor
  g960
  (
    n993,
    n486,
    n988,
    n990,
    n485
  );


  nor
  g961
  (
    n1010,
    n990,
    n483,
    n992,
    n991
  );


  and
  g962
  (
    n1002,
    n486,
    n853,
    n483,
    n992
  );


  nand
  g963
  (
    n1006,
    n992,
    n524,
    n852,
    n952
  );


  xnor
  g964
  (
    n1007,
    n989,
    n954,
    n953,
    n486
  );


  and
  g965
  (
    n995,
    n988,
    n525,
    n524
  );


  or
  g966
  (
    n998,
    n991,
    n972,
    n483,
    n851
  );


  nand
  g967
  (
    n999,
    n991,
    n990,
    n852,
    n954
  );


  nor
  g968
  (
    n1004,
    n954,
    n991,
    n483,
    n525
  );


  nand
  g969
  (
    n996,
    n992,
    n972,
    n484,
    n853
  );


  nor
  g970
  (
    n1003,
    n851,
    n989,
    n853,
    n525
  );


  nor
  g971
  (
    n1008,
    n955,
    n955,
    n852,
    n953
  );


  xor
  g972
  (
    n1001,
    n989,
    n988,
    n485,
    n851
  );


  xnor
  g973
  (
    n1000,
    n990,
    n851,
    n486,
    n954
  );


  nor
  g974
  (
    n994,
    n484,
    n526,
    n485,
    n524
  );


  nor
  g975
  (
    n1005,
    n484,
    n526,
    n953,
    n853
  );


  nand
  g976
  (
    n1009,
    n953,
    n952,
    n971,
    n485
  );


  nor
  g977
  (
    n997,
    n852,
    n524,
    n850,
    n484
  );


  nand
  g978
  (
    n1014,
    n527,
    n529,
    n993
  );


  or
  g979
  (
    n1012,
    n529,
    n526,
    n993
  );


  nand
  g980
  (
    n1011,
    n994,
    n528,
    n526
  );


  and
  g981
  (
    n1013,
    n993,
    n528,
    n530,
    n527
  );


  xnor
  g982
  (
    n1015,
    n528,
    n527,
    n529
  );


  buf
  g983
  (
    n1019,
    n1012
  );


  buf
  g984
  (
    n1017,
    n1012
  );


  not
  g985
  (
    n1022,
    n1011
  );


  buf
  g986
  (
    n1020,
    n1011
  );


  buf
  g987
  (
    n1016,
    n1013
  );


  buf
  g988
  (
    n1024,
    n1011
  );


  buf
  g989
  (
    n1023,
    n1011
  );


  not
  g990
  (
    n1025,
    n1012
  );


  not
  g991
  (
    n1018,
    n1013
  );


  not
  g992
  (
    n1021,
    n1012
  );


  xor
  g993
  (
    n1060,
    n981,
    n1018,
    n973,
    n1023
  );


  xor
  g994
  (
    n1036,
    n981,
    n855,
    n930,
    n999
  );


  or
  g995
  (
    n1050,
    n530,
    n1024,
    n930,
    n892
  );


  or
  g996
  (
    n1044,
    n1022,
    n999,
    n933,
    n1019
  );


  nor
  g997
  (
    n1032,
    n996,
    n855,
    n931
  );


  xnor
  g998
  (
    n1042,
    n1022,
    n975,
    n1021,
    n1025
  );


  xnor
  g999
  (
    n1045,
    n1025,
    n1023,
    n958
  );


  xnor
  g1000
  (
    n1029,
    n1001,
    n1000,
    n977,
    n998
  );


  xor
  g1001
  (
    n1039,
    n1022,
    n979,
    n1002,
    n1020
  );


  xor
  g1002
  (
    n1049,
    n958,
    n531,
    n1018,
    n1021
  );


  or
  g1003
  (
    n1048,
    n930,
    n957,
    n1017,
    n532
  );


  nand
  g1004
  (
    n1038,
    n854,
    n995,
    n974,
    n1016
  );


  xnor
  g1005
  (
    n1056,
    n1023,
    n933,
    n995,
    n1024
  );


  nor
  g1006
  (
    n1055,
    n994,
    n981,
    n1021,
    n1016
  );


  nand
  g1007
  (
    n1062,
    n979,
    n976,
    n1021,
    n1000
  );


  nand
  g1008
  (
    n1059,
    n956,
    n854,
    n955,
    n979
  );


  or
  g1009
  (
    n1026,
    n974,
    n956,
    n996
  );


  xor
  g1010
  (
    n1065,
    n1024,
    n1025,
    n1018,
    n531
  );


  nand
  g1011
  (
    n1061,
    n1020,
    n1024,
    n854,
    n979
  );


  xnor
  g1012
  (
    n1052,
    n932,
    n1017,
    n976,
    n854
  );


  xor
  g1013
  (
    n1040,
    n982,
    n931,
    n932,
    n955
  );


  nand
  g1014
  (
    n1027,
    n933,
    n855,
    n996,
    n1000
  );


  and
  g1015
  (
    n1033,
    n1020,
    n995,
    n994,
    n1022
  );


  xor
  g1016
  (
    n1053,
    n999,
    n999,
    n930,
    n980
  );


  nor
  g1017
  (
    n1051,
    n996,
    n530,
    n974,
    n531
  );


  and
  g1018
  (
    n1030,
    n998,
    n978,
    n1016,
    n1019
  );


  nand
  g1019
  (
    n1046,
    n980,
    n975,
    n997,
    n994
  );


  xnor
  g1020
  (
    n1054,
    n1001,
    n956,
    n1017,
    n976
  );


  nor
  g1021
  (
    n1063,
    n958,
    n934,
    n998,
    n957
  );


  xnor
  g1022
  (
    n1047,
    n1018,
    n980,
    n977,
    n997
  );


  xnor
  g1023
  (
    n1058,
    n933,
    n1000,
    n980,
    n995
  );


  xnor
  g1024
  (
    n1043,
    n975,
    n997,
    n532,
    n982
  );


  nor
  g1025
  (
    n1064,
    n1001,
    n1017,
    n977,
    n533
  );


  nand
  g1026
  (
    n1037,
    n530,
    n531,
    n1020,
    n982
  );


  and
  g1027
  (
    n1041,
    n855,
    n977,
    n532,
    n978
  );


  or
  g1028
  (
    n1035,
    n1025,
    n932,
    n974
  );


  or
  g1029
  (
    n1028,
    n978,
    n1019,
    n998,
    n1001
  );


  or
  g1030
  (
    n1031,
    n997,
    n976,
    n978,
    n981
  );


  nand
  g1031
  (
    n1034,
    n1019,
    n957,
    n931,
    n975
  );


  xnor
  g1032
  (
    n1057,
    n957,
    n1016,
    n532,
    n958
  );


  xnor
  g1033
  (
    n1132,
    n626,
    n579,
    n561,
    n615
  );


  nor
  g1034
  (
    n1190,
    n594,
    n629,
    n628,
    n566
  );


  or
  g1035
  (
    n1177,
    n592,
    n1033,
    n553,
    n620
  );


  xnor
  g1036
  (
    n1102,
    n549,
    n567,
    n1064,
    n1036
  );


  nor
  g1037
  (
    n1166,
    n628,
    n1063,
    n590,
    n1014
  );


  xnor
  g1038
  (
    n1208,
    n650,
    n1026,
    n541,
    n619
  );


  xor
  g1039
  (
    n1113,
    n533,
    n646,
    n540,
    n1061
  );


  and
  g1040
  (
    n1117,
    n1034,
    n577,
    n580,
    n1055
  );


  and
  g1041
  (
    n1187,
    n643,
    n554,
    n577,
    n589
  );


  nor
  g1042
  (
    n1186,
    n1030,
    n624,
    n646,
    n1028
  );


  xor
  g1043
  (
    n1211,
    n620,
    n623,
    n595,
    n597
  );


  xor
  g1044
  (
    n1179,
    n1043,
    n1047,
    n600,
    n599
  );


  xor
  g1045
  (
    n1076,
    n1047,
    n543,
    n1043,
    n1044
  );


  and
  g1046
  (
    n1189,
    n1032,
    n583,
    n1061,
    n636
  );


  xor
  g1047
  (
    n1141,
    n626,
    n568,
    n566,
    n585
  );


  nor
  g1048
  (
    n1171,
    n617,
    n639,
    n583,
    n550
  );


  or
  g1049
  (
    n1140,
    n534,
    n589,
    n598,
    n1063
  );


  and
  g1050
  (
    n1180,
    n1041,
    n577,
    n636,
    n641
  );


  xor
  g1051
  (
    n1134,
    n643,
    n1059,
    n594,
    n631
  );


  nor
  g1052
  (
    n1108,
    n638,
    n622,
    n572,
    n551
  );


  and
  g1053
  (
    n1198,
    n536,
    n571,
    n1062,
    n1057
  );


  nor
  g1054
  (
    n1195,
    n627,
    n535,
    n583,
    n602
  );


  nand
  g1055
  (
    n1105,
    n621,
    n552,
    n605
  );


  xnor
  g1056
  (
    n1178,
    n633,
    n582,
    n646,
    n1042
  );


  and
  g1057
  (
    n1082,
    n586,
    n643,
    n648,
    n1028
  );


  nand
  g1058
  (
    n1212,
    n610,
    n564,
    n635,
    n585
  );


  xor
  g1059
  (
    n1191,
    n645,
    n534,
    n567,
    n1035
  );


  or
  g1060
  (
    n1217,
    n572,
    n1063,
    n555,
    n595
  );


  xnor
  g1061
  (
    n1072,
    n584,
    n535,
    n591,
    n574
  );


  nor
  g1062
  (
    n1090,
    n1030,
    n563,
    n1038,
    n568
  );


  nand
  g1063
  (
    n1078,
    n581,
    n649,
    n611,
    n637
  );


  xor
  g1064
  (
    n1183,
    n1059,
    n613,
    n1036,
    n600
  );


  nor
  g1065
  (
    n1074,
    n627,
    n543,
    n1053,
    n592
  );


  and
  g1066
  (
    n1207,
    n587,
    n1063,
    n584,
    n1052
  );


  and
  g1067
  (
    n1147,
    n574,
    n1052,
    n606,
    n578
  );


  nor
  g1068
  (
    n1167,
    n632,
    n1048,
    n600,
    n619
  );


  nor
  g1069
  (
    n1160,
    n563,
    n555,
    n595,
    n621
  );


  nand
  g1070
  (
    n1094,
    n630,
    n1057,
    n1031,
    n538
  );


  nor
  g1071
  (
    n1158,
    n1026,
    n590,
    n606,
    n638
  );


  nand
  g1072
  (
    n1081,
    n596,
    n983,
    n577,
    n555
  );


  nor
  g1073
  (
    n1069,
    n982,
    n544,
    n576,
    n627
  );


  or
  g1074
  (
    n1223,
    n614,
    n590,
    n1039,
    n559
  );


  xnor
  g1075
  (
    n1083,
    n648,
    n617,
    n1036,
    n643
  );


  xor
  g1076
  (
    n1116,
    n1013,
    n618,
    n1064,
    n1033
  );


  xnor
  g1077
  (
    n1123,
    n1058,
    n1064,
    n588,
    n642
  );


  xnor
  g1078
  (
    n1193,
    n1039,
    n556,
    n575,
    n1035
  );


  and
  g1079
  (
    n1219,
    n625,
    n568,
    n615,
    n1058
  );


  xnor
  g1080
  (
    n1203,
    n544,
    n603,
    n606,
    n632
  );


  nor
  g1081
  (
    n1168,
    n1048,
    n605,
    n580,
    n564
  );


  nand
  g1082
  (
    n1104,
    n605,
    n639,
    n1037,
    n549
  );


  xnor
  g1083
  (
    n1096,
    n1050,
    n565,
    n1028,
    n597
  );


  nand
  g1084
  (
    n1111,
    n1031,
    n1053,
    n1027,
    n576
  );


  or
  g1085
  (
    n1201,
    n600,
    n570,
    n611,
    n1041
  );


  nand
  g1086
  (
    n1097,
    n541,
    n557,
    n1059,
    n1046
  );


  or
  g1087
  (
    n1086,
    n571,
    n536,
    n1026,
    n579
  );


  nor
  g1088
  (
    n1109,
    n641,
    n558,
    n618,
    n648
  );


  nand
  g1089
  (
    n1070,
    n588,
    n597,
    n1051,
    n573
  );


  or
  g1090
  (
    n1080,
    n571,
    n591,
    n597,
    n544
  );


  nand
  g1091
  (
    n1133,
    n623,
    n585,
    n596,
    n603
  );


  and
  g1092
  (
    n1143,
    n1047,
    n612,
    n616,
    n618
  );


  nand
  g1093
  (
    n1126,
    n604,
    n645,
    n633,
    n649
  );


  or
  g1094
  (
    n1206,
    n539,
    n1034,
    n595,
    n583
  );


  xnor
  g1095
  (
    n1200,
    n1065,
    n602,
    n1064,
    n537
  );


  or
  g1096
  (
    n1192,
    n564,
    n543,
    n1037,
    n558
  );


  and
  g1097
  (
    n1176,
    n593,
    n533,
    n549,
    n608
  );


  or
  g1098
  (
    n1066,
    n609,
    n551,
    n1052,
    n1040
  );


  or
  g1099
  (
    n1152,
    n1046,
    n615,
    n562,
    n645
  );


  and
  g1100
  (
    n1071,
    n1034,
    n983,
    n601,
    n630
  );


  xor
  g1101
  (
    n1087,
    n579,
    n561,
    n637,
    n567
  );


  xor
  g1102
  (
    n1222,
    n560,
    n1054,
    n645,
    n650
  );


  or
  g1103
  (
    n1121,
    n574,
    n1044,
    n538,
    n613
  );


  xnor
  g1104
  (
    n1079,
    n602,
    n539,
    n584,
    n618
  );


  nor
  g1105
  (
    n1091,
    n544,
    n1027,
    n647,
    n598
  );


  and
  g1106
  (
    n1225,
    n555,
    n550,
    n537,
    n566
  );


  nor
  g1107
  (
    n1196,
    n1050,
    n1035,
    n548,
    n617
  );


  or
  g1108
  (
    n1088,
    n1055,
    n538,
    n599,
    n1035
  );


  nand
  g1109
  (
    n1202,
    n536,
    n622,
    n533,
    n1043
  );


  xor
  g1110
  (
    n1153,
    n1040,
    n559,
    n610,
    n1061
  );


  nor
  g1111
  (
    n1095,
    n1028,
    n1040,
    n1041,
    n1045
  );


  xor
  g1112
  (
    n1101,
    n545,
    n559,
    n1031,
    n622
  );


  and
  g1113
  (
    n1213,
    n539,
    n542,
    n1014
  );


  xor
  g1114
  (
    n1214,
    n1029,
    n564,
    n625,
    n575
  );


  or
  g1115
  (
    n1172,
    n983,
    n546,
    n1058,
    n642
  );


  or
  g1116
  (
    n1130,
    n568,
    n623,
    n647,
    n586
  );


  or
  g1117
  (
    n1098,
    n1037,
    n1014,
    n586,
    n546
  );


  and
  g1118
  (
    n1077,
    n641,
    n628,
    n581,
    n629
  );


  nand
  g1119
  (
    n1136,
    n553,
    n552,
    n649,
    n579
  );


  xor
  g1120
  (
    n1085,
    n570,
    n538,
    n569,
    n1039
  );


  and
  g1121
  (
    n1159,
    n562,
    n634,
    n609,
    n607
  );


  or
  g1122
  (
    n1120,
    n1049,
    n630,
    n1048,
    n626
  );


  nor
  g1123
  (
    n1182,
    n601,
    n614,
    n615,
    n619
  );


  xnor
  g1124
  (
    n1115,
    n984,
    n554,
    n644,
    n563
  );


  nand
  g1125
  (
    n1119,
    n553,
    n566,
    n638,
    n1049
  );


  nor
  g1126
  (
    n1110,
    n593,
    n598,
    n1044,
    n535
  );


  xnor
  g1127
  (
    n1092,
    n1034,
    n1065,
    n644,
    n587
  );


  xor
  g1128
  (
    n1164,
    n545,
    n541,
    n1049,
    n638
  );


  xnor
  g1129
  (
    n1199,
    n640,
    n1057,
    n548,
    n1038
  );


  nand
  g1130
  (
    n1138,
    n560,
    n644,
    n610,
    n604
  );


  nand
  g1131
  (
    n1156,
    n606,
    n570,
    n599,
    n1056
  );


  xor
  g1132
  (
    n1100,
    n649,
    n619,
    n610,
    n546
  );


  xnor
  g1133
  (
    n1181,
    n648,
    n547,
    n554,
    n562
  );


  or
  g1134
  (
    n1220,
    n537,
    n616,
    n621,
    n634
  );


  and
  g1135
  (
    n1129,
    n536,
    n1060,
    n1045,
    n594
  );


  nor
  g1136
  (
    n1224,
    n644,
    n631,
    n614,
    n635
  );


  and
  g1137
  (
    n1089,
    n558,
    n572,
    n1056,
    n588
  );


  nand
  g1138
  (
    n1154,
    n624,
    n636,
    n574,
    n569
  );


  xor
  g1139
  (
    n1197,
    n551,
    n1043,
    n603,
    n642
  );


  and
  g1140
  (
    n1099,
    n633,
    n573,
    n545,
    n604
  );


  nand
  g1141
  (
    n1209,
    n563,
    n983,
    n560,
    n559
  );


  xor
  g1142
  (
    n1163,
    n557,
    n635,
    n592,
    n625
  );


  nand
  g1143
  (
    n1075,
    n565,
    n628,
    n560,
    n1058
  );


  or
  g1144
  (
    n1205,
    n575,
    n588,
    n591,
    n1050
  );


  nor
  g1145
  (
    n1204,
    n534,
    n1039,
    n1054,
    n1046
  );


  and
  g1146
  (
    n1218,
    n541,
    n552,
    n1030,
    n569
  );


  or
  g1147
  (
    n1073,
    n556,
    n624,
    n547,
    n551
  );


  or
  g1148
  (
    n1107,
    n1062,
    n621,
    n585,
    n608
  );


  nor
  g1149
  (
    n1174,
    n591,
    n1030,
    n625,
    n1029
  );


  nor
  g1150
  (
    n1103,
    n1045,
    n612,
    n594,
    n578
  );


  xor
  g1151
  (
    n1106,
    n548,
    n608,
    n590,
    n547
  );


  nor
  g1152
  (
    n1165,
    n1033,
    n601,
    n1051,
    n1061
  );


  and
  g1153
  (
    n1145,
    n1053,
    n540,
    n1032,
    n640
  );


  xor
  g1154
  (
    n1142,
    n534,
    n1065,
    n1056,
    n582
  );


  nand
  g1155
  (
    n1149,
    n626,
    n586,
    n1050,
    n578
  );


  nor
  g1156
  (
    n1148,
    n604,
    n554,
    n647,
    n587
  );


  nand
  g1157
  (
    n1114,
    n1040,
    n1054,
    n1038,
    n631
  );


  xnor
  g1158
  (
    n1068,
    n570,
    n1013,
    n1047,
    n1060
  );


  xor
  g1159
  (
    n1215,
    n1051,
    n569,
    n624,
    n1045
  );


  nor
  g1160
  (
    n1124,
    n633,
    n1046,
    n640,
    n607
  );


  and
  g1161
  (
    n1210,
    n539,
    n632,
    n1029,
    n614
  );


  xor
  g1162
  (
    n1162,
    n616,
    n593,
    n634
  );


  xor
  g1163
  (
    n1150,
    n576,
    n608,
    n1036,
    n646
  );


  nor
  g1164
  (
    n1137,
    n580,
    n542,
    n1056,
    n556
  );


  nand
  g1165
  (
    n1146,
    n1060,
    n596,
    n553,
    n545
  );


  nor
  g1166
  (
    n1131,
    n1049,
    n601,
    n1053,
    n578
  );


  nand
  g1167
  (
    n1194,
    n612,
    n582,
    n1062,
    n639
  );


  nand
  g1168
  (
    n1184,
    n589,
    n1065,
    n609,
    n622
  );


  xor
  g1169
  (
    n1157,
    n581,
    n557,
    n641,
    n1060
  );


  xor
  g1170
  (
    n1175,
    n1052,
    n1062,
    n613,
    n598
  );


  xor
  g1171
  (
    n1155,
    n587,
    n548,
    n635,
    n1027
  );


  and
  g1172
  (
    n1161,
    n582,
    n1026,
    n639,
    n556
  );


  and
  g1173
  (
    n1170,
    n567,
    n617,
    n640,
    n565
  );


  nor
  g1174
  (
    n1173,
    n1037,
    n636,
    n596,
    n607
  );


  nand
  g1175
  (
    n1144,
    n573,
    n543,
    n642,
    n613
  );


  nand
  g1176
  (
    n1169,
    n557,
    n1054,
    n647,
    n542
  );


  xor
  g1177
  (
    n1216,
    n1042,
    n571,
    n581,
    n609
  );


  and
  g1178
  (
    n1188,
    n620,
    n630,
    n552,
    n623
  );


  nor
  g1179
  (
    n1093,
    n1032,
    n561,
    n1027,
    n607
  );


  nand
  g1180
  (
    n1122,
    n540,
    n562,
    n637,
    n1041
  );


  xnor
  g1181
  (
    n1067,
    n572,
    n629,
    n627,
    n573
  );


  and
  g1182
  (
    n1151,
    n592,
    n611,
    n1044,
    n1048
  );


  xnor
  g1183
  (
    n1118,
    n589,
    n580,
    n602,
    n561
  );


  nor
  g1184
  (
    n1139,
    n565,
    n550,
    n603,
    n549
  );


  and
  g1185
  (
    n1125,
    n1038,
    n599,
    n1031,
    n540
  );


  xnor
  g1186
  (
    n1128,
    n1029,
    n1032,
    n558,
    n1057
  );


  or
  g1187
  (
    n1135,
    n1055,
    n550,
    n584,
    n612
  );


  and
  g1188
  (
    n1084,
    n616,
    n547,
    n632,
    n1059
  );


  nand
  g1189
  (
    n1127,
    n593,
    n546,
    n537,
    n575
  );


  nor
  g1190
  (
    n1221,
    n576,
    n1051,
    n637,
    n1033
  );


  xor
  g1191
  (
    n1112,
    n620,
    n631,
    n1042,
    n535
  );


  nand
  g1192
  (
    n1185,
    n611,
    n1055,
    n629,
    n1042
  );


  buf
  g1193
  (
    n1316,
    n1090
  );


  nor
  g1194
  (
    n1273,
    n1125,
    n1004,
    n1148,
    n1167
  );


  xor
  g1195
  (
    n1305,
    n1145,
    n1163,
    n1157,
    n1138
  );


  nor
  g1196
  (
    n1302,
    n1107,
    n1141,
    n1156,
    n1115
  );


  xnor
  g1197
  (
    n1262,
    n1173,
    n1119,
    n1176,
    n1136
  );


  nand
  g1198
  (
    n1301,
    n1141,
    n1175,
    n1131,
    n1125
  );


  nand
  g1199
  (
    n1279,
    n1077,
    n1173,
    n1106,
    n1005
  );


  xnor
  g1200
  (
    n1339,
    n1098,
    n1002,
    n1140,
    n1183
  );


  and
  g1201
  (
    n1315,
    n937,
    n1180,
    n1096,
    n1112
  );


  and
  g1202
  (
    n1296,
    n1148,
    n1070,
    n1143,
    n1134
  );


  or
  g1203
  (
    n1360,
    n1086,
    n1153,
    n1143,
    n1145
  );


  and
  g1204
  (
    n1270,
    n1080,
    n1153,
    n1167,
    n1083
  );


  xnor
  g1205
  (
    n1240,
    n1068,
    n1098,
    n1114,
    n1095
  );


  nor
  g1206
  (
    n1234,
    n1126,
    n1072,
    n1087,
    n1170
  );


  xor
  g1207
  (
    n1300,
    n1184,
    n1141,
    n1079,
    n1144
  );


  nand
  g1208
  (
    n1338,
    n1111,
    n1149,
    n1123,
    n1182
  );


  xnor
  g1209
  (
    n1285,
    n1132,
    n1005,
    n1181,
    n1155
  );


  xor
  g1210
  (
    n1310,
    n1179,
    n1138,
    n651,
    n1078
  );


  nor
  g1211
  (
    n1352,
    n1106,
    n1148,
    n1083,
    n1072
  );


  xnor
  g1212
  (
    n1344,
    n1083,
    n1181,
    n1087,
    n1102
  );


  xnor
  g1213
  (
    n1243,
    n1099,
    n1124,
    n935,
    n1111
  );


  and
  g1214
  (
    n1246,
    n935,
    n1158,
    n1005,
    n1160
  );


  or
  g1215
  (
    n1331,
    n1172,
    n1089,
    n1140,
    n1125
  );


  nand
  g1216
  (
    n1256,
    n1113,
    n1073,
    n1142,
    n1162
  );


  xor
  g1217
  (
    n1321,
    n1166,
    n1185,
    n1089,
    n1076
  );


  or
  g1218
  (
    n1238,
    n1103,
    n1181,
    n1154,
    n1010
  );


  nand
  g1219
  (
    n1319,
    n1118,
    n1007,
    n1176,
    n1159
  );


  nor
  g1220
  (
    n1280,
    n1101,
    n1074,
    n1153,
    n1069
  );


  or
  g1221
  (
    n1332,
    n1118,
    n1093,
    n1128,
    n1117
  );


  xor
  g1222
  (
    n1269,
    n1086,
    n1104,
    n1068,
    n1174
  );


  xnor
  g1223
  (
    n1288,
    n1168,
    n1163,
    n1113,
    n1104
  );


  nor
  g1224
  (
    n1231,
    n1097,
    n1154,
    n1098,
    n1089
  );


  or
  g1225
  (
    n1320,
    n1073,
    n1099,
    n1002,
    n1104
  );


  xnor
  g1226
  (
    n1295,
    n1178,
    n1133,
    n1107,
    n934
  );


  nor
  g1227
  (
    n1325,
    n652,
    n1138,
    n1172,
    n1105
  );


  nand
  g1228
  (
    n1260,
    n1112,
    n1120,
    n1184,
    n1178
  );


  nand
  g1229
  (
    n1244,
    n1117,
    n1082,
    n1120,
    n1173
  );


  or
  g1230
  (
    n1329,
    n1159,
    n1183,
    n1116,
    n1142
  );


  nand
  g1231
  (
    n1347,
    n1082,
    n1143,
    n1066,
    n1115
  );


  or
  g1232
  (
    n1290,
    n1129,
    n1174,
    n1086,
    n1156
  );


  nand
  g1233
  (
    n1228,
    n1110,
    n1183,
    n1138,
    n1100
  );


  xnor
  g1234
  (
    n1335,
    n1140,
    n1080,
    n1114,
    n1177
  );


  and
  g1235
  (
    n1277,
    n1133,
    n1152,
    n1173,
    n1135
  );


  xor
  g1236
  (
    n1237,
    n1094,
    n1073,
    n1147,
    n1137
  );


  nand
  g1237
  (
    n1275,
    n1132,
    n1175,
    n1135,
    n1078
  );


  and
  g1238
  (
    n1272,
    n1125,
    n1171,
    n1110,
    n1127
  );


  xor
  g1239
  (
    n1333,
    n1109,
    n1110,
    n1162,
    n1123
  );


  or
  g1240
  (
    n1309,
    n1144,
    n1185,
    n1102,
    n937
  );


  nand
  g1241
  (
    n1343,
    n1097,
    n1003,
    n1160,
    n1112
  );


  or
  g1242
  (
    n1322,
    n1124,
    n1180,
    n1127,
    n1179
  );


  nand
  g1243
  (
    n1304,
    n1159,
    n1115,
    n1161,
    n1153
  );


  or
  g1244
  (
    n1266,
    n1091,
    n1164,
    n1069,
    n1093
  );


  or
  g1245
  (
    n1247,
    n1131,
    n1120,
    n1091,
    n1006
  );


  xnor
  g1246
  (
    n1251,
    n1166,
    n1136,
    n1112,
    n652
  );


  nand
  g1247
  (
    n1351,
    n1004,
    n1077,
    n1009,
    n1161
  );


  xnor
  g1248
  (
    n1263,
    n1146,
    n1128,
    n1168,
    n1157
  );


  xor
  g1249
  (
    n1233,
    n1009,
    n1121,
    n1094,
    n1171
  );


  or
  g1250
  (
    n1291,
    n1072,
    n1102,
    n1085
  );


  xnor
  g1251
  (
    n1307,
    n1096,
    n1150,
    n1007,
    n1161
  );


  and
  g1252
  (
    n1271,
    n1130,
    n1123,
    n1088,
    n1167
  );


  nor
  g1253
  (
    n1337,
    n1148,
    n1079,
    n935,
    n1074
  );


  and
  g1254
  (
    n1357,
    n1069,
    n1149,
    n1113,
    n1123
  );


  nor
  g1255
  (
    n1254,
    n1067,
    n1151,
    n1164,
    n1106
  );


  nand
  g1256
  (
    n1283,
    n1139,
    n1068,
    n1119,
    n1135
  );


  nor
  g1257
  (
    n1226,
    n1103,
    n1120,
    n1006,
    n1132
  );


  nand
  g1258
  (
    n1232,
    n1099,
    n1111,
    n1119,
    n1133
  );


  xor
  g1259
  (
    n1249,
    n1094,
    n1071,
    n1119,
    n1155
  );


  xor
  g1260
  (
    n1359,
    n1091,
    n1092,
    n1166,
    n1003
  );


  xor
  g1261
  (
    n1230,
    n1085,
    n1166,
    n1122,
    n1150
  );


  nor
  g1262
  (
    n1278,
    n1151,
    n1006,
    n1134,
    n1146
  );


  or
  g1263
  (
    n1354,
    n1115,
    n1156,
    n1005,
    n1144
  );


  and
  g1264
  (
    n1350,
    n937,
    n936,
    n1086,
    n1091
  );


  nor
  g1265
  (
    n1340,
    n1186,
    n1126,
    n1010,
    n1142
  );


  nand
  g1266
  (
    n1252,
    n1163,
    n1108,
    n1146,
    n1179
  );


  or
  g1267
  (
    n1314,
    n1117,
    n1164,
    n1137,
    n1067
  );


  xnor
  g1268
  (
    n1242,
    n1150,
    n1097,
    n1139,
    n1146
  );


  or
  g1269
  (
    n1348,
    n1070,
    n1010,
    n1143,
    n1109
  );


  nor
  g1270
  (
    n1346,
    n1176,
    n1067,
    n934,
    n1170
  );


  and
  g1271
  (
    n1324,
    n1003,
    n917,
    n1007,
    n1172
  );


  nand
  g1272
  (
    n1236,
    n1095,
    n1157,
    n1078,
    n1177
  );


  and
  g1273
  (
    n1265,
    n650,
    n1155,
    n1008,
    n1088
  );


  nand
  g1274
  (
    n1361,
    n1075,
    n650,
    n1182,
    n1087
  );


  and
  g1275
  (
    n1345,
    n1080,
    n1110,
    n1002,
    n1089
  );


  xnor
  g1276
  (
    n1358,
    n1082,
    n1073,
    n1128,
    n1066
  );


  nor
  g1277
  (
    n1289,
    n1163,
    n1136,
    n1066,
    n1124
  );


  nor
  g1278
  (
    n1286,
    n1066,
    n1128,
    n651,
    n1183
  );


  nor
  g1279
  (
    n1239,
    n1152,
    n1095,
    n1116,
    n1177
  );


  nor
  g1280
  (
    n1284,
    n1114,
    n1004,
    n1116,
    n1177
  );


  nand
  g1281
  (
    n1330,
    n1075,
    n1184,
    n1084,
    n1150
  );


  nor
  g1282
  (
    n1313,
    n1130,
    n1105,
    n1118,
    n1077
  );


  xnor
  g1283
  (
    n1274,
    n1084,
    n1116,
    n1076,
    n1137
  );


  nor
  g1284
  (
    n1312,
    n1127,
    n1081,
    n1090,
    n1170
  );


  nand
  g1285
  (
    n1258,
    n1152,
    n1165,
    n1092,
    n1080
  );


  nand
  g1286
  (
    n1299,
    n1109,
    n1147,
    n652,
    n1136
  );


  or
  g1287
  (
    n1298,
    n1105,
    n1126,
    n1129,
    n1006
  );


  nor
  g1288
  (
    n1327,
    n1165,
    n1100,
    n1180,
    n936
  );


  nand
  g1289
  (
    n1318,
    n1145,
    n1097,
    n935,
    n1176
  );


  nand
  g1290
  (
    n1227,
    n1092,
    n1100,
    n1185,
    n1008
  );


  nand
  g1291
  (
    n1276,
    n1149,
    n1101,
    n1157,
    n1121
  );


  nand
  g1292
  (
    n1326,
    n1104,
    n1167,
    n1132,
    n1168
  );


  xor
  g1293
  (
    n1336,
    n1094,
    n1181,
    n1141,
    n1071
  );


  nand
  g1294
  (
    n1323,
    n1103,
    n1084,
    n1008,
    n1168
  );


  or
  g1295
  (
    n1341,
    n1078,
    n1008,
    n651,
    n1079
  );


  and
  g1296
  (
    n1334,
    n1071,
    n1129,
    n1079,
    n1170
  );


  nand
  g1297
  (
    n1306,
    n1131,
    n1130,
    n1108,
    n1178
  );


  or
  g1298
  (
    n1297,
    n1135,
    n1144,
    n1122,
    n1121
  );


  xor
  g1299
  (
    n1287,
    n1169,
    n1075,
    n1149,
    n1070
  );


  and
  g1300
  (
    n1267,
    n1004,
    n1175,
    n1172,
    n1165
  );


  and
  g1301
  (
    n1248,
    n1105,
    n1070,
    n1162,
    n1185
  );


  nand
  g1302
  (
    n1342,
    n1130,
    n1169,
    n1122,
    n1108
  );


  and
  g1303
  (
    n1235,
    n1109,
    n1075,
    n1152,
    n1118
  );


  xor
  g1304
  (
    n1253,
    n1142,
    n1139,
    n1129,
    n1154
  );


  xor
  g1305
  (
    n1241,
    n1090,
    n1133,
    n1147,
    n936
  );


  xor
  g1306
  (
    n1250,
    n1074,
    n1147,
    n1140,
    n1082
  );


  xor
  g1307
  (
    n1311,
    n1111,
    n917,
    n1067,
    n936
  );


  and
  g1308
  (
    n1261,
    n1117,
    n1159,
    n1179,
    n1093
  );


  xor
  g1309
  (
    n1294,
    n1081,
    n1180,
    n1162,
    n1093
  );


  nand
  g1310
  (
    n1293,
    n1174,
    n1009,
    n1158,
    n1077
  );


  xnor
  g1311
  (
    n1259,
    n1154,
    n1076,
    n1161
  );


  xor
  g1312
  (
    n1281,
    n1092,
    n1099,
    n1100,
    n1158
  );


  xnor
  g1313
  (
    n1264,
    n1081,
    n1124,
    n1178,
    n1088
  );


  or
  g1314
  (
    n1356,
    n1101,
    n1083,
    n1113,
    n1102
  );


  xor
  g1315
  (
    n1257,
    n1098,
    n1160,
    n1169,
    n1175
  );


  nand
  g1316
  (
    n1255,
    n1139,
    n1010,
    n1085,
    n1088
  );


  xor
  g1317
  (
    n1292,
    n1107,
    n1156,
    n1072,
    n1122
  );


  nor
  g1318
  (
    n1268,
    n1007,
    n1069,
    n1127,
    n1169
  );


  and
  g1319
  (
    n1282,
    n934,
    n1174,
    n1103,
    n1160
  );


  or
  g1320
  (
    n1303,
    n1095,
    n1090,
    n1151,
    n651
  );


  xor
  g1321
  (
    n1328,
    n1151,
    n1074,
    n1096
  );


  and
  g1322
  (
    n1349,
    n1126,
    n1009,
    n1155,
    n1068
  );


  xnor
  g1323
  (
    n1353,
    n1114,
    n1171,
    n1134
  );


  nor
  g1324
  (
    n1245,
    n1158,
    n1101,
    n1107,
    n1165
  );


  or
  g1325
  (
    n1229,
    n1182,
    n1071,
    n1164,
    n1003
  );


  or
  g1326
  (
    n1317,
    n1145,
    n1087,
    n1108,
    n1106
  );


  xnor
  g1327
  (
    n1355,
    n1171,
    n1084,
    n1131,
    n1182
  );


  and
  g1328
  (
    n1308,
    n1184,
    n1137,
    n1121,
    n1081
  );


  and
  g1329
  (
    n1677,
    n1292,
    n717,
    n780,
    n1360
  );


  xnor
  g1330
  (
    n1493,
    n1223,
    n1259,
    n1245,
    n728
  );


  or
  g1331
  (
    n1590,
    n786,
    n695,
    n1293,
    n1283
  );


  and
  g1332
  (
    n1514,
    n1345,
    n1253,
    n753
  );


  and
  g1333
  (
    n1520,
    n682,
    n828,
    n1191,
    n1310
  );


  nand
  g1334
  (
    n1592,
    n837,
    n1253,
    n697,
    n1265
  );


  xor
  g1335
  (
    n1704,
    n1318,
    n739,
    n1252,
    n662
  );


  and
  g1336
  (
    n1474,
    n715,
    n1346,
    n1289,
    n1360
  );


  or
  g1337
  (
    n1699,
    n715,
    n1243,
    n1221,
    n812
  );


  xor
  g1338
  (
    n1568,
    n676,
    n832,
    n662,
    n1314
  );


  xnor
  g1339
  (
    n1503,
    n655,
    n1323,
    n839,
    n1297
  );


  nand
  g1340
  (
    n1484,
    n827,
    n1243,
    n1322,
    n1213
  );


  or
  g1341
  (
    n1475,
    n712,
    n782,
    n490,
    n1230
  );


  and
  g1342
  (
    n1695,
    n840,
    n749,
    n832,
    n1298
  );


  or
  g1343
  (
    n1429,
    n1226,
    n801,
    n1237,
    n1015
  );


  xor
  g1344
  (
    n1521,
    n774,
    n670,
    n747,
    n1342
  );


  xor
  g1345
  (
    n1727,
    n1276,
    n1347,
    n1241,
    n1295
  );


  nand
  g1346
  (
    n1606,
    n1285,
    n1277,
    n821,
    n1219
  );


  nor
  g1347
  (
    n1389,
    n790,
    n761,
    n742,
    n1236
  );


  xor
  g1348
  (
    n1731,
    n826,
    n1339,
    n1343,
    n1313
  );


  xor
  g1349
  (
    n1670,
    n792,
    n1236,
    n1298,
    n751
  );


  and
  g1350
  (
    n1630,
    n1314,
    n694,
    n1223,
    n771
  );


  xnor
  g1351
  (
    n1644,
    n1208,
    n729,
    n1237,
    n673
  );


  or
  g1352
  (
    n1496,
    n1214,
    n1192,
    n757,
    n843
  );


  xor
  g1353
  (
    n1689,
    n726,
    n1251,
    n736,
    n1352
  );


  nor
  g1354
  (
    n1382,
    n1187,
    n1361,
    n1291,
    n689
  );


  nor
  g1355
  (
    n1435,
    n719,
    n1329,
    n1296,
    n807
  );


  xor
  g1356
  (
    n1684,
    n1239,
    n1262,
    n705,
    n822
  );


  xnor
  g1357
  (
    n1585,
    n699,
    n746,
    n689,
    n1242
  );


  xnor
  g1358
  (
    n1694,
    n811,
    n836,
    n1199,
    n1222
  );


  nand
  g1359
  (
    n1528,
    n1198,
    n1209,
    n710,
    n1317
  );


  nand
  g1360
  (
    n1519,
    n811,
    n841,
    n1331,
    n742
  );


  nor
  g1361
  (
    n1634,
    n1305,
    n1335,
    n1256,
    n699
  );


  nor
  g1362
  (
    n1525,
    n1330,
    n838,
    n666,
    n671
  );


  and
  g1363
  (
    n1579,
    n811,
    n727,
    n825,
    n1294
  );


  and
  g1364
  (
    n1556,
    n767,
    n825,
    n812,
    n1194
  );


  nand
  g1365
  (
    n1529,
    n1250,
    n753,
    n1356,
    n729
  );


  xor
  g1366
  (
    n1413,
    n1223,
    n715,
    n769,
    n694
  );


  nand
  g1367
  (
    n1444,
    n1202,
    n795,
    n685,
    n1217
  );


  xor
  g1368
  (
    n1646,
    n1243,
    n817,
    n839,
    n1214
  );


  xor
  g1369
  (
    n1708,
    n681,
    n743,
    n1211,
    n816
  );


  xnor
  g1370
  (
    n1460,
    n808,
    n740,
    n1263,
    n697
  );


  xnor
  g1371
  (
    n1669,
    n1322,
    n658,
    n653,
    n762
  );


  xnor
  g1372
  (
    n1485,
    n1205,
    n771,
    n1194,
    n674
  );


  nand
  g1373
  (
    n1655,
    n1276,
    n707,
    n1271,
    n1351
  );


  or
  g1374
  (
    n1392,
    n734,
    n1300,
    n1257,
    n758
  );


  and
  g1375
  (
    n1407,
    n1267,
    n1270,
    n745,
    n1315
  );


  or
  g1376
  (
    n1645,
    n728,
    n770,
    n691,
    n725
  );


  and
  g1377
  (
    n1406,
    n685,
    n770,
    n714,
    n814
  );


  xor
  g1378
  (
    n1458,
    n837,
    n677,
    n1299,
    n1272
  );


  nor
  g1379
  (
    n1553,
    n758,
    n793,
    n832,
    n764
  );


  and
  g1380
  (
    n1540,
    n775,
    n1261,
    n782,
    n700
  );


  nand
  g1381
  (
    n1633,
    n1316,
    n822,
    n716,
    n756
  );


  xnor
  g1382
  (
    n1650,
    n819,
    n718,
    n1329,
    n1288
  );


  xor
  g1383
  (
    n1602,
    n788,
    n789,
    n719,
    n1204
  );


  xor
  g1384
  (
    n1608,
    n1312,
    n669,
    n1309,
    n819
  );


  nand
  g1385
  (
    n1533,
    n750,
    n1306,
    n653,
    n746
  );


  or
  g1386
  (
    n1618,
    n1314,
    n700,
    n682,
    n669
  );


  nor
  g1387
  (
    n1656,
    n768,
    n808,
    n1352,
    n1343
  );


  or
  g1388
  (
    n1397,
    n738,
    n1259,
    n658,
    n777
  );


  nor
  g1389
  (
    n1623,
    n656,
    n788,
    n800,
    n781
  );


  xor
  g1390
  (
    n1654,
    n840,
    n824,
    n723,
    n843
  );


  or
  g1391
  (
    n1719,
    n841,
    n712,
    n835,
    n1238
  );


  nor
  g1392
  (
    n1467,
    n766,
    n1230,
    n1228,
    n1212
  );


  or
  g1393
  (
    n1643,
    n752,
    n785,
    n666,
    n1329
  );


  and
  g1394
  (
    n1723,
    n686,
    n1198,
    n1328,
    n1215
  );


  nand
  g1395
  (
    n1405,
    n1339,
    n693,
    n1233,
    n783
  );


  or
  g1396
  (
    n1648,
    n825,
    n1304,
    n1300,
    n732
  );


  or
  g1397
  (
    n1594,
    n800,
    n1215,
    n791,
    n1210
  );


  xnor
  g1398
  (
    n1588,
    n789,
    n661,
    n1188,
    n1272
  );


  and
  g1399
  (
    n1398,
    n1265,
    n1335,
    n1250,
    n697
  );


  or
  g1400
  (
    n1378,
    n663,
    n711,
    n817,
    n1190
  );


  and
  g1401
  (
    n1721,
    n784,
    n748,
    n1228,
    n1015
  );


  xor
  g1402
  (
    n1614,
    n1247,
    n754,
    n752,
    n787
  );


  nor
  g1403
  (
    n1536,
    n820,
    n785,
    n698,
    n702
  );


  nor
  g1404
  (
    n1679,
    n705,
    n1345,
    n841,
    n1210
  );


  or
  g1405
  (
    n1619,
    n1239,
    n765,
    n489,
    n784
  );


  or
  g1406
  (
    n1470,
    n1313,
    n688,
    n810,
    n1321
  );


  nand
  g1407
  (
    n1627,
    n1326,
    n713,
    n687,
    n830
  );


  xor
  g1408
  (
    n1472,
    n1246,
    n684,
    n823,
    n820
  );


  or
  g1409
  (
    n1576,
    n811,
    n722,
    n784,
    n740
  );


  xnor
  g1410
  (
    n1542,
    n726,
    n1271,
    n829,
    n1356
  );


  xnor
  g1411
  (
    n1483,
    n1333,
    n675,
    n1225,
    n1275
  );


  or
  g1412
  (
    n1551,
    n802,
    n1261,
    n1298,
    n754
  );


  xnor
  g1413
  (
    n1587,
    n1205,
    n665,
    n682,
    n1288
  );


  xnor
  g1414
  (
    n1544,
    n1212,
    n1189,
    n1304,
    n700
  );


  xnor
  g1415
  (
    n1701,
    n488,
    n769,
    n1218,
    n1246
  );


  xnor
  g1416
  (
    n1543,
    n721,
    n734,
    n722,
    n688
  );


  xor
  g1417
  (
    n1605,
    n756,
    n1340,
    n757,
    n1195
  );


  xnor
  g1418
  (
    n1687,
    n767,
    n1330,
    n1259,
    n828
  );


  nor
  g1419
  (
    n1675,
    n1291,
    n786,
    n1359,
    n838
  );


  nor
  g1420
  (
    n1658,
    n668,
    n777,
    n1347,
    n797
  );


  and
  g1421
  (
    n1370,
    n1222,
    n684,
    n693,
    n718
  );


  xnor
  g1422
  (
    n1686,
    n1244,
    n827,
    n1230,
    n661
  );


  or
  g1423
  (
    n1638,
    n1246,
    n1328,
    n690,
    n1292
  );


  xor
  g1424
  (
    n1548,
    n1336,
    n1206,
    n657,
    n1352
  );


  xnor
  g1425
  (
    n1499,
    n1310,
    n1284,
    n774,
    n1290
  );


  xor
  g1426
  (
    n1577,
    n1268,
    n1247,
    n808,
    n1319
  );


  or
  g1427
  (
    n1570,
    n1342,
    n1261,
    n827,
    n725
  );


  or
  g1428
  (
    n1511,
    n764,
    n831,
    n694,
    n984
  );


  nand
  g1429
  (
    n1416,
    n666,
    n1276,
    n831,
    n1309
  );


  nand
  g1430
  (
    n1452,
    n1212,
    n794,
    n737,
    n1331
  );


  nor
  g1431
  (
    n1598,
    n817,
    n786,
    n698,
    n1234
  );


  nand
  g1432
  (
    n1404,
    n761,
    n703,
    n1238,
    n693
  );


  nor
  g1433
  (
    n1364,
    n675,
    n829,
    n984,
    n1349
  );


  nand
  g1434
  (
    n1437,
    n803,
    n1332,
    n1233,
    n1301
  );


  xor
  g1435
  (
    n1522,
    n1272,
    n1278,
    n719,
    n816
  );


  xnor
  g1436
  (
    n1698,
    n1189,
    n1225,
    n663,
    n743
  );


  xnor
  g1437
  (
    n1620,
    n694,
    n824,
    n1359,
    n829
  );


  and
  g1438
  (
    n1418,
    n759,
    n666,
    n821,
    n766
  );


  xor
  g1439
  (
    n1597,
    n1262,
    n1269,
    n746,
    n833
  );


  xnor
  g1440
  (
    n1479,
    n744,
    n734,
    n671,
    n790
  );


  nand
  g1441
  (
    n1586,
    n1322,
    n738,
    n1355,
    n670
  );


  nor
  g1442
  (
    n1705,
    n660,
    n1288,
    n793,
    n1293
  );


  and
  g1443
  (
    n1509,
    n785,
    n683,
    n723,
    n1345
  );


  nand
  g1444
  (
    n1412,
    n784,
    n775,
    n1353,
    n701
  );


  nor
  g1445
  (
    n1569,
    n760,
    n1188,
    n1189,
    n732
  );


  nor
  g1446
  (
    n1534,
    n1326,
    n1264,
    n487,
    n1245
  );


  nand
  g1447
  (
    n1440,
    n705,
    n679,
    n1341,
    n737
  );


  and
  g1448
  (
    n1402,
    n488,
    n1346,
    n805,
    n757
  );


  nand
  g1449
  (
    n1447,
    n653,
    n724,
    n1280,
    n1318
  );


  xor
  g1450
  (
    n1660,
    n1295,
    n1353,
    n813,
    n669
  );


  xnor
  g1451
  (
    n1446,
    n1324,
    n1265,
    n744,
    n755
  );


  nor
  g1452
  (
    n1510,
    n793,
    n1348,
    n1259,
    n1263
  );


  nor
  g1453
  (
    n1545,
    n1268,
    n1357,
    n779,
    n1348
  );


  nor
  g1454
  (
    n1393,
    n728,
    n730,
    n1192,
    n720
  );


  and
  g1455
  (
    n1451,
    n695,
    n1357,
    n805,
    n781
  );


  nor
  g1456
  (
    n1575,
    n748,
    n772,
    n832,
    n823
  );


  or
  g1457
  (
    n1517,
    n1291,
    n1280,
    n1279,
    n1338
  );


  and
  g1458
  (
    n1601,
    n1323,
    n1324,
    n1215,
    n1286
  );


  nor
  g1459
  (
    n1417,
    n680,
    n1341,
    n655,
    n1317
  );


  nand
  g1460
  (
    n1729,
    n654,
    n711,
    n751,
    n817
  );


  nor
  g1461
  (
    n1672,
    n1260,
    n1337,
    n745,
    n1319
  );


  or
  g1462
  (
    n1367,
    n800,
    n896,
    n1300,
    n1282
  );


  or
  g1463
  (
    n1603,
    n1270,
    n682,
    n1320,
    n757
  );


  xnor
  g1464
  (
    n1450,
    n1313,
    n683,
    n767,
    n1273
  );


  nand
  g1465
  (
    n1631,
    n1278,
    n1320,
    n1318,
    n708
  );


  xnor
  g1466
  (
    n1647,
    n1313,
    n833,
    n842,
    n1202
  );


  nand
  g1467
  (
    n1464,
    n1316,
    n1301,
    n1312,
    n733
  );


  or
  g1468
  (
    n1527,
    n779,
    n751,
    n790,
    n1206
  );


  and
  g1469
  (
    n1507,
    n741,
    n1193,
    n831,
    n730
  );


  nor
  g1470
  (
    n1371,
    n679,
    n1255,
    n1196,
    n658
  );


  nor
  g1471
  (
    n1730,
    n1306,
    n1334,
    n1200,
    n798
  );


  nand
  g1472
  (
    n1461,
    n1197,
    n690,
    n1258,
    n704
  );


  xor
  g1473
  (
    n1414,
    n794,
    n1337,
    n778,
    n834
  );


  nand
  g1474
  (
    n1408,
    n1322,
    n668,
    n1273,
    n755
  );


  and
  g1475
  (
    n1506,
    n487,
    n838,
    n737,
    n1245
  );


  or
  g1476
  (
    n1366,
    n1189,
    n731,
    n1219,
    n1355
  );


  nand
  g1477
  (
    n1425,
    n685,
    n729,
    n1253,
    n1267
  );


  nor
  g1478
  (
    n1681,
    n1309,
    n701,
    n731,
    n1228
  );


  xor
  g1479
  (
    n1637,
    n1264,
    n692,
    n748,
    n767
  );


  or
  g1480
  (
    n1693,
    n1346,
    n684,
    n707,
    n1249
  );


  xor
  g1481
  (
    n1494,
    n1204,
    n684,
    n1226,
    n1208
  );


  xnor
  g1482
  (
    n1428,
    n760,
    n659,
    n1211,
    n713
  );


  xnor
  g1483
  (
    n1573,
    n779,
    n1274,
    n683,
    n1333
  );


  xnor
  g1484
  (
    n1682,
    n673,
    n1257,
    n1213,
    n1305
  );


  and
  g1485
  (
    n1615,
    n762,
    n1354,
    n1269,
    n1200
  );


  or
  g1486
  (
    n1571,
    n1249,
    n735,
    n721,
    n716
  );


  or
  g1487
  (
    n1700,
    n656,
    n700,
    n1321,
    n1344
  );


  nor
  g1488
  (
    n1652,
    n1266,
    n1290,
    n809,
    n713
  );


  xor
  g1489
  (
    n1728,
    n1300,
    n782,
    n803,
    n796
  );


  or
  g1490
  (
    n1487,
    n1015,
    n1266,
    n1358,
    n1279
  );


  xnor
  g1491
  (
    n1668,
    n1342,
    n764,
    n1209,
    n1273
  );


  nand
  g1492
  (
    n1369,
    n679,
    n687,
    n1301,
    n790
  );


  xnor
  g1493
  (
    n1385,
    n763,
    n1250,
    n830,
    n490
  );


  nand
  g1494
  (
    n1726,
    n1187,
    n796,
    n1326,
    n724
  );


  or
  g1495
  (
    n1430,
    n731,
    n702,
    n1224,
    n1306
  );


  xnor
  g1496
  (
    n1733,
    n1257,
    n1351,
    n688,
    n1251
  );


  and
  g1497
  (
    n1667,
    n765,
    n1349,
    n1186,
    n1341
  );


  xor
  g1498
  (
    n1635,
    n487,
    n803,
    n1336,
    n701
  );


  and
  g1499
  (
    n1365,
    n768,
    n1345,
    n667,
    n1361
  );


  and
  g1500
  (
    n1566,
    n724,
    n766,
    n1262,
    n754
  );


  nand
  g1501
  (
    n1690,
    n1281,
    n733,
    n1214,
    n739
  );


  nand
  g1502
  (
    n1535,
    n1227,
    n664,
    n1336,
    n1190
  );


  nor
  g1503
  (
    n1531,
    n1240,
    n840,
    n796,
    n1354
  );


  xor
  g1504
  (
    n1489,
    n661,
    n1229,
    n821,
    n760
  );


  nand
  g1505
  (
    n1439,
    n1015,
    n671,
    n805,
    n1197
  );


  and
  g1506
  (
    n1478,
    n823,
    n1239,
    n1207,
    n768
  );


  xnor
  g1507
  (
    n1426,
    n1279,
    n1245,
    n1327,
    n1305
  );


  xnor
  g1508
  (
    n1607,
    n717,
    n662,
    n1197,
    n1254
  );


  or
  g1509
  (
    n1593,
    n764,
    n1316,
    n1284,
    n781
  );


  nand
  g1510
  (
    n1639,
    n1188,
    n1337,
    n691,
    n1232
  );


  nor
  g1511
  (
    n1659,
    n1295,
    n1252,
    n772,
    n686
  );


  xor
  g1512
  (
    n1488,
    n816,
    n714,
    n1200,
    n806
  );


  nor
  g1513
  (
    n1578,
    n812,
    n1266,
    n1303,
    n783
  );


  nand
  g1514
  (
    n1717,
    n691,
    n656,
    n487,
    n1271
  );


  nor
  g1515
  (
    n1703,
    n667,
    n1267,
    n775,
    n1359
  );


  xor
  g1516
  (
    n1716,
    n788,
    n1254,
    n798,
    n1355
  );


  xor
  g1517
  (
    n1554,
    n842,
    n1204,
    n1237,
    n1235
  );


  xnor
  g1518
  (
    n1589,
    n1324,
    n795,
    n820,
    n815
  );


  or
  g1519
  (
    n1604,
    n1344,
    n1351,
    n696,
    n804
  );


  or
  g1520
  (
    n1626,
    n680,
    n1200,
    n1190,
    n1214
  );


  and
  g1521
  (
    n1560,
    n1283,
    n678,
    n813,
    n1250
  );


  xnor
  g1522
  (
    n1676,
    n1273,
    n704,
    n819,
    n1340
  );


  xnor
  g1523
  (
    n1581,
    n697,
    n814,
    n1211,
    n1303
  );


  xor
  g1524
  (
    n1713,
    n1279,
    n1354,
    n676,
    n1233
  );


  nor
  g1525
  (
    n1410,
    n1334,
    n1341,
    n1207,
    n1221
  );


  nand
  g1526
  (
    n1584,
    n1223,
    n787,
    n1298,
    n1340
  );


  nand
  g1527
  (
    n1383,
    n1204,
    n1283,
    n1311,
    n1336
  );


  xnor
  g1528
  (
    n1495,
    n704,
    n667,
    n1242,
    n791
  );


  nand
  g1529
  (
    n1558,
    n1275,
    n712,
    n1284,
    n722
  );


  nand
  g1530
  (
    n1486,
    n802,
    n1206,
    n773,
    n775
  );


  nor
  g1531
  (
    n1424,
    n681,
    n743,
    n696,
    n1263
  );


  or
  g1532
  (
    n1420,
    n734,
    n719,
    n1217,
    n1357
  );


  nand
  g1533
  (
    n1629,
    n830,
    n1344,
    n747,
    n820
  );


  nand
  g1534
  (
    n1471,
    n1201,
    n1270,
    n723,
    n668
  );


  nor
  g1535
  (
    n1664,
    n674,
    n704,
    n756,
    n1251
  );


  nor
  g1536
  (
    n1436,
    n681,
    n1231,
    n1307,
    n736
  );


  nand
  g1537
  (
    n1691,
    n1350,
    n1248,
    n672,
    n1278
  );


  and
  g1538
  (
    n1688,
    n1358,
    n1229,
    n1203,
    n1343
  );


  xor
  g1539
  (
    n1621,
    n1307,
    n1218,
    n818,
    n799
  );


  nor
  g1540
  (
    n1583,
    n680,
    n1260,
    n725,
    n747
  );


  nor
  g1541
  (
    n1710,
    n1330,
    n1240,
    n1309,
    n828
  );


  xnor
  g1542
  (
    n1657,
    n1216,
    n1227,
    n840,
    n665
  );


  nand
  g1543
  (
    n1438,
    n810,
    n692,
    n1335,
    n1277
  );


  xor
  g1544
  (
    n1375,
    n1220,
    n778,
    n706,
    n745
  );


  or
  g1545
  (
    n1415,
    n1256,
    n1316,
    n1339,
    n675
  );


  xor
  g1546
  (
    n1482,
    n1194,
    n741,
    n674,
    n1246
  );


  and
  g1547
  (
    n1711,
    n1358,
    n1014,
    n1352,
    n489
  );


  xnor
  g1548
  (
    n1546,
    n1343,
    n827,
    n1335,
    n751
  );


  and
  g1549
  (
    n1674,
    n685,
    n804,
    n670,
    n1257
  );


  nand
  g1550
  (
    n1476,
    n814,
    n676,
    n669,
    n1281
  );


  or
  g1551
  (
    n1555,
    n766,
    n1206,
    n692,
    n1315
  );


  nor
  g1552
  (
    n1539,
    n1210,
    n1190,
    n1290,
    n753
  );


  or
  g1553
  (
    n1409,
    n1297,
    n1293,
    n759,
    n1347
  );


  xor
  g1554
  (
    n1666,
    n1216,
    n749,
    n792,
    n1220
  );


  nor
  g1555
  (
    n1411,
    n776,
    n758,
    n797,
    n843
  );


  xor
  g1556
  (
    n1481,
    n673,
    n772,
    n1198,
    n1238
  );


  nand
  g1557
  (
    n1538,
    n1251,
    n1216,
    n1338,
    n1287
  );


  xnor
  g1558
  (
    n1616,
    n801,
    n824,
    n655,
    n1310
  );


  and
  g1559
  (
    n1395,
    n1249,
    n1238,
    n1265,
    n663
  );


  xor
  g1560
  (
    n1724,
    n1235,
    n1291,
    n752,
    n836
  );


  xor
  g1561
  (
    n1683,
    n1353,
    n842,
    n714,
    n1191
  );


  nor
  g1562
  (
    n1463,
    n716,
    n787,
    n1207,
    n1296
  );


  or
  g1563
  (
    n1491,
    n1262,
    n703,
    n1296,
    n802
  );


  and
  g1564
  (
    n1649,
    n1229,
    n709,
    n809,
    n813
  );


  xor
  g1565
  (
    n1697,
    n1258,
    n777,
    n1244,
    n733
  );


  xor
  g1566
  (
    n1500,
    n664,
    n1285,
    n1318,
    n1210
  );


  xor
  g1567
  (
    n1427,
    n706,
    n789,
    n1353,
    n777
  );


  nor
  g1568
  (
    n1718,
    n708,
    n1361,
    n1241,
    n687
  );


  or
  g1569
  (
    n1445,
    n765,
    n821,
    n1289,
    n710
  );


  or
  g1570
  (
    n1610,
    n802,
    n742,
    n1264,
    n1234
  );


  or
  g1571
  (
    n1492,
    n1270,
    n1202,
    n735,
    n773
  );


  nand
  g1572
  (
    n1609,
    n703,
    n1269,
    n1264,
    n695
  );


  xnor
  g1573
  (
    n1595,
    n726,
    n657,
    n793,
    n1195
  );


  or
  g1574
  (
    n1612,
    n1302,
    n774,
    n792,
    n1339
  );


  nand
  g1575
  (
    n1391,
    n661,
    n1268,
    n1360,
    n665
  );


  or
  g1576
  (
    n1526,
    n1281,
    n1317,
    n756,
    n720
  );


  and
  g1577
  (
    n1377,
    n740,
    n818,
    n769,
    n1232
  );


  nand
  g1578
  (
    n1562,
    n1234,
    n668,
    n712,
    n672
  );


  nand
  g1579
  (
    n1421,
    n689,
    n1222,
    n1358,
    n815
  );


  xnor
  g1580
  (
    n1530,
    n683,
    n654,
    n678,
    n1327
  );


  and
  g1581
  (
    n1455,
    n1325,
    n1299,
    n776,
    n652
  );


  nor
  g1582
  (
    n1665,
    n698,
    n1218,
    n701,
    n1306
  );


  xor
  g1583
  (
    n1696,
    n842,
    n1356,
    n1319,
    n1354
  );


  and
  g1584
  (
    n1640,
    n676,
    n717,
    n800,
    n1348
  );


  nand
  g1585
  (
    n1663,
    n804,
    n776,
    n720,
    n664
  );


  and
  g1586
  (
    n1565,
    n809,
    n688,
    n1243,
    n1271
  );


  nor
  g1587
  (
    n1399,
    n681,
    n680,
    n738,
    n798
  );


  xnor
  g1588
  (
    n1448,
    n1274,
    n689,
    n745,
    n657
  );


  xor
  g1589
  (
    n1532,
    n1256,
    n1227,
    n797,
    n664
  );


  and
  g1590
  (
    n1473,
    n1227,
    n825,
    n488,
    n782
  );


  and
  g1591
  (
    n1707,
    n736,
    n843,
    n779,
    n1292
  );


  xnor
  g1592
  (
    n1559,
    n1221,
    n788,
    n1195,
    n1202
  );


  xnor
  g1593
  (
    n1734,
    n1280,
    n1289,
    n1216,
    n806
  );


  and
  g1594
  (
    n1422,
    n1274,
    n1293,
    n806,
    n1326
  );


  nor
  g1595
  (
    n1680,
    n1194,
    n490,
    n770
  );


  and
  g1596
  (
    n1722,
    n809,
    n1187,
    n1272,
    n769
  );


  xor
  g1597
  (
    n1591,
    n1290,
    n1237,
    n1292,
    n1320
  );


  and
  g1598
  (
    n1574,
    n1218,
    n1258,
    n660,
    n1360
  );


  xnor
  g1599
  (
    n1714,
    n717,
    n1230,
    n801,
    n658
  );


  xor
  g1600
  (
    n1561,
    n709,
    n686,
    n1355,
    n1208
  );


  xor
  g1601
  (
    n1466,
    n781,
    n686,
    n813,
    n1304
  );


  or
  g1602
  (
    n1403,
    n727,
    n765,
    n1331,
    n1330
  );


  nor
  g1603
  (
    n1547,
    n1209,
    n829,
    n1356,
    n1207
  );


  and
  g1604
  (
    n1596,
    n1323,
    n1317,
    n1242,
    n1307
  );


  and
  g1605
  (
    n1502,
    n1247,
    n692,
    n1235,
    n815
  );


  xnor
  g1606
  (
    n1564,
    n831,
    n671,
    n1225,
    n1198
  );


  or
  g1607
  (
    n1431,
    n1213,
    n834,
    n736,
    n1242
  );


  nand
  g1608
  (
    n1501,
    n1331,
    n739,
    n699,
    n797
  );


  nor
  g1609
  (
    n1661,
    n750,
    n806,
    n678,
    n1221
  );


  xor
  g1610
  (
    n1396,
    n796,
    n1303,
    n1219,
    n780
  );


  or
  g1611
  (
    n1376,
    n1302,
    n1342,
    n1308,
    n1255
  );


  xnor
  g1612
  (
    n1512,
    n1338,
    n1220,
    n742,
    n1361
  );


  xor
  g1613
  (
    n1394,
    n1233,
    n1226,
    n794,
    n1299
  );


  xnor
  g1614
  (
    n1362,
    n1299,
    n758,
    n761,
    n702
  );


  xor
  g1615
  (
    n1456,
    n677,
    n1308,
    n799,
    n1333
  );


  and
  g1616
  (
    n1613,
    n741,
    n1241,
    n1192,
    n794
  );


  xnor
  g1617
  (
    n1379,
    n750,
    n783,
    n1209,
    n1320
  );


  xnor
  g1618
  (
    n1720,
    n753,
    n1308,
    n743,
    n1254
  );


  or
  g1619
  (
    n1384,
    n1319,
    n728,
    n708,
    n1303
  );


  xor
  g1620
  (
    n1572,
    n698,
    n1277,
    n823,
    n709
  );


  xor
  g1621
  (
    n1386,
    n659,
    n1276,
    n706,
    n1327
  );


  or
  g1622
  (
    n1523,
    n1211,
    n747,
    n1261,
    n1240
  );


  xnor
  g1623
  (
    n1625,
    n1311,
    n1195,
    n1334,
    n763
  );


  xor
  g1624
  (
    n1557,
    n1307,
    n761,
    n1289,
    n677
  );


  nand
  g1625
  (
    n1580,
    n699,
    n718,
    n801,
    n1247
  );


  xor
  g1626
  (
    n1628,
    n750,
    n1208,
    n789,
    n1285
  );


  or
  g1627
  (
    n1490,
    n662,
    n1260,
    n760,
    n706
  );


  nand
  g1628
  (
    n1480,
    n812,
    n828,
    n1197,
    n780
  );


  and
  g1629
  (
    n1636,
    n1196,
    n726,
    n759,
    n837
  );


  or
  g1630
  (
    n1537,
    n1296,
    n984,
    n792,
    n763
  );


  xnor
  g1631
  (
    n1725,
    n716,
    n1283,
    n1328,
    n804
  );


  xor
  g1632
  (
    n1515,
    n741,
    n1332,
    n720,
    n1359
  );


  or
  g1633
  (
    n1454,
    n836,
    n763,
    n835,
    n670
  );


  xnor
  g1634
  (
    n1433,
    n655,
    n1192,
    n772,
    n1231
  );


  xor
  g1635
  (
    n1715,
    n732,
    n696,
    n1252
  );


  and
  g1636
  (
    n1541,
    n679,
    n749,
    n1349,
    n1278
  );


  xor
  g1637
  (
    n1390,
    n837,
    n771,
    n749,
    n488
  );


  nor
  g1638
  (
    n1453,
    n799,
    n1249,
    n1350,
    n1281
  );


  xor
  g1639
  (
    n1441,
    n1229,
    n778,
    n1324,
    n1203
  );


  or
  g1640
  (
    n1401,
    n773,
    n1241,
    n791,
    n1191
  );


  nand
  g1641
  (
    n1374,
    n1301,
    n1255,
    n1236,
    n814
  );


  or
  g1642
  (
    n1400,
    n776,
    n657,
    n1351,
    n1255
  );


  nand
  g1643
  (
    n1468,
    n755,
    n773,
    n1269,
    n729
  );


  nor
  g1644
  (
    n1600,
    n818,
    n1282,
    n762,
    n1201
  );


  nand
  g1645
  (
    n1732,
    n740,
    n826,
    n1302,
    n707
  );


  xnor
  g1646
  (
    n1465,
    n1325,
    n731,
    n834,
    n822
  );


  nor
  g1647
  (
    n1692,
    n687,
    n1228,
    n783,
    n1268
  );


  or
  g1648
  (
    n1550,
    n1275,
    n1327,
    n836,
    n1232
  );


  nand
  g1649
  (
    n1443,
    n762,
    n1333,
    n1196,
    n818
  );


  xnor
  g1650
  (
    n1653,
    n1193,
    n1315,
    n1267,
    n1295
  );


  nor
  g1651
  (
    n1624,
    n656,
    n1256,
    n834,
    n780
  );


  or
  g1652
  (
    n1516,
    n799,
    n1311,
    n1334,
    n727
  );


  or
  g1653
  (
    n1552,
    n702,
    n755,
    n703,
    n1286
  );


  xor
  g1654
  (
    n1671,
    n725,
    n833,
    n1205,
    n711
  );


  xnor
  g1655
  (
    n1380,
    n1323,
    n1344,
    n1263,
    n1350
  );


  nand
  g1656
  (
    n1504,
    n774,
    n739,
    n1315,
    n1328
  );


  xnor
  g1657
  (
    n1449,
    n748,
    n1224,
    n1220,
    n1287
  );


  nand
  g1658
  (
    n1513,
    n710,
    n1325,
    n1347,
    n816
  );


  xnor
  g1659
  (
    n1432,
    n1340,
    n665,
    n1314,
    n770
  );


  nor
  g1660
  (
    n1419,
    n1231,
    n795,
    n489,
    n807
  );


  xor
  g1661
  (
    n1622,
    n1280,
    n839,
    n744,
    n659
  );


  nand
  g1662
  (
    n1368,
    n693,
    n1205,
    n815,
    n826
  );


  xor
  g1663
  (
    n1388,
    n1244,
    n798,
    n715,
    n691
  );


  xor
  g1664
  (
    n1524,
    n1203,
    n709,
    n1248,
    n1297
  );


  xnor
  g1665
  (
    n1372,
    n1346,
    n1294,
    n1235,
    n673
  );


  nand
  g1666
  (
    n1709,
    n737,
    n730,
    n1321,
    n654
  );


  and
  g1667
  (
    n1706,
    n839,
    n659,
    n1349,
    n723
  );


  or
  g1668
  (
    n1678,
    n1284,
    n1199,
    n1203,
    n1286
  );


  nand
  g1669
  (
    n1632,
    n718,
    n1285,
    n1287,
    n1244
  );


  nand
  g1670
  (
    n1673,
    n1224,
    n678,
    n830,
    n1282
  );


  xor
  g1671
  (
    n1563,
    n1286,
    n660,
    n1186,
    n1321
  );


  or
  g1672
  (
    n1505,
    n791,
    n1287,
    n1338,
    n1305
  );


  xnor
  g1673
  (
    n1423,
    n1329,
    n835,
    n1258,
    n771
  );


  xnor
  g1674
  (
    n1642,
    n1325,
    n653,
    n824,
    n1248
  );


  or
  g1675
  (
    n1387,
    n835,
    n1191,
    n1288,
    n690
  );


  xor
  g1676
  (
    n1442,
    n1224,
    n1332,
    n744,
    n785
  );


  and
  g1677
  (
    n1498,
    n1188,
    n1294,
    n710,
    n807
  );


  xnor
  g1678
  (
    n1381,
    n795,
    n1240,
    n677,
    n1231
  );


  and
  g1679
  (
    n1582,
    n778,
    n1196,
    n1217
  );


  nor
  g1680
  (
    n1497,
    n730,
    n1310,
    n805,
    n768
  );


  or
  g1681
  (
    n1477,
    n695,
    n674,
    n489,
    n711
  );


  xnor
  g1682
  (
    n1702,
    n1187,
    n833,
    n752,
    n1357
  );


  xor
  g1683
  (
    n1549,
    n663,
    n660,
    n1236,
    n1277
  );


  xnor
  g1684
  (
    n1712,
    n714,
    n1201,
    n810,
    n786
  );


  xnor
  g1685
  (
    n1459,
    n1212,
    n721,
    n1332,
    n808
  );


  nand
  g1686
  (
    n1567,
    n1201,
    n735,
    n721,
    n1311
  );


  or
  g1687
  (
    n1508,
    n838,
    n707,
    n675,
    n705
  );


  xor
  g1688
  (
    n1611,
    n759,
    n1337,
    n654,
    n722
  );


  nand
  g1689
  (
    n1685,
    n1213,
    n1199,
    n696,
    n1282
  );


  or
  g1690
  (
    n1363,
    n733,
    n1274,
    n819,
    n1266
  );


  nor
  g1691
  (
    n1434,
    n1215,
    n1239,
    n1302,
    n672
  );


  xnor
  g1692
  (
    n1662,
    n708,
    n1304,
    n826,
    n1294
  );


  nor
  g1693
  (
    n1373,
    n667,
    n1225,
    n787,
    n803
  );


  xnor
  g1694
  (
    n1518,
    n1219,
    n810,
    n724,
    n754
  );


  xnor
  g1695
  (
    n1641,
    n738,
    n1193,
    n1348,
    n1312
  );


  xor
  g1696
  (
    n1651,
    n1254,
    n1312,
    n690,
    n746
  );


  nor
  g1697
  (
    n1457,
    n1308,
    n735,
    n1222,
    n1248
  );


  or
  g1698
  (
    n1617,
    n1199,
    n732,
    n822,
    n672
  );


  and
  g1699
  (
    n1462,
    n1193,
    n1350,
    n1260,
    n1297
  );


  nor
  g1700
  (
    n1469,
    n727,
    n1186,
    n1232,
    n713
  );


  or
  g1701
  (
    n1599,
    n841,
    n1234,
    n1275,
    n807
  );


  xnor
  g1702
  (
    n1901,
    n1721,
    n1545,
    n1553,
    n1717
  );


  nand
  g1703
  (
    n1891,
    n1638,
    n1501,
    n1632,
    n1424
  );


  nand
  g1704
  (
    n1831,
    n1394,
    n1660,
    n1435,
    n1649
  );


  nand
  g1705
  (
    n1922,
    n1630,
    n1664,
    n1556,
    n1384
  );


  xor
  g1706
  (
    n1929,
    n1730,
    n1622,
    n1665,
    n1643
  );


  nand
  g1707
  (
    n1907,
    n1674,
    n1632,
    n1424,
    n1543
  );


  nor
  g1708
  (
    n1939,
    n1633,
    n1451,
    n1453,
    n1720
  );


  xor
  g1709
  (
    n1777,
    n1492,
    n1416,
    n1641,
    n1387
  );


  nand
  g1710
  (
    n1743,
    n1418,
    n1579,
    n1440,
    n1386
  );


  xnor
  g1711
  (
    n1747,
    n1500,
    n1619,
    n148,
    n1493
  );


  and
  g1712
  (
    n1857,
    n1515,
    n1410,
    n1507,
    n1477
  );


  nand
  g1713
  (
    n1832,
    n1487,
    n1460,
    n1596,
    n1591
  );


  or
  g1714
  (
    n1790,
    n1636,
    n1372,
    n1590,
    n1415
  );


  or
  g1715
  (
    n1821,
    n1698,
    n1418,
    n1400,
    n1438
  );


  or
  g1716
  (
    n1896,
    n1557,
    n1587,
    n1699,
    n1459
  );


  xnor
  g1717
  (
    n1823,
    n1550,
    n1584,
    n1512,
    n1399
  );


  xor
  g1718
  (
    n1859,
    n1386,
    n1598,
    n1649,
    n1609
  );


  xor
  g1719
  (
    n1841,
    n1643,
    n1366,
    n1499,
    n1635
  );


  nand
  g1720
  (
    n1925,
    n1458,
    n1396,
    n1522,
    n1619
  );


  nor
  g1721
  (
    n1858,
    n1678,
    n1701,
    n1415,
    n1516
  );


  nor
  g1722
  (
    n1885,
    n1363,
    n1669,
    n1454,
    n1492
  );


  or
  g1723
  (
    n1931,
    n1373,
    n1392,
    n1696,
    n1442
  );


  or
  g1724
  (
    n1883,
    n1677,
    n1365,
    n1595,
    n1490
  );


  or
  g1725
  (
    n1869,
    n1711,
    n1661,
    n1589,
    n1726
  );


  nor
  g1726
  (
    n1873,
    n1468,
    n1497,
    n1607,
    n1517
  );


  nor
  g1727
  (
    n1765,
    n1568,
    n1731,
    n1684,
    n1608
  );


  and
  g1728
  (
    n1872,
    n1700,
    n1476,
    n1363,
    n1527
  );


  nand
  g1729
  (
    n1795,
    n1687,
    n1521,
    n1395,
    n1462
  );


  nand
  g1730
  (
    n1906,
    n1378,
    n1484,
    n1623,
    n1503
  );


  or
  g1731
  (
    n1825,
    n1715,
    n1392,
    n1618,
    n1641
  );


  and
  g1732
  (
    n1888,
    n1729,
    n1449,
    n1557,
    n1486
  );


  xor
  g1733
  (
    n1882,
    n1441,
    n1388,
    n1685,
    n1372
  );


  xor
  g1734
  (
    n1877,
    n1729,
    n1601,
    n1597,
    n1697
  );


  xnor
  g1735
  (
    n1932,
    n1672,
    n1465,
    n1376,
    n1658
  );


  and
  g1736
  (
    n1820,
    n1611,
    n1429,
    n1455,
    n1644
  );


  xnor
  g1737
  (
    n1785,
    n1514,
    n1651,
    n1606,
    n1555
  );


  nand
  g1738
  (
    n1921,
    n1369,
    n1627,
    n1658,
    n1642
  );


  xor
  g1739
  (
    n1833,
    n1437,
    n1634,
    n1534,
    n1652
  );


  and
  g1740
  (
    n1917,
    n1645,
    n1670,
    n1380,
    n1639
  );


  or
  g1741
  (
    n1770,
    n1620,
    n1434,
    n1382,
    n1423
  );


  or
  g1742
  (
    n1934,
    n1460,
    n1605,
    n1681,
    n1524
  );


  xnor
  g1743
  (
    n1937,
    n1693,
    n1399,
    n1649,
    n1527
  );


  and
  g1744
  (
    n1861,
    n1693,
    n1576,
    n1701,
    n1385
  );


  or
  g1745
  (
    n1766,
    n1447,
    n1463,
    n1488,
    n1600
  );


  nor
  g1746
  (
    n1864,
    n1519,
    n1398,
    n1544,
    n1564
  );


  nand
  g1747
  (
    n1830,
    n1474,
    n1521,
    n1431,
    n1432
  );


  xor
  g1748
  (
    n1868,
    n1540,
    n1725,
    n1549,
    n1525
  );


  xor
  g1749
  (
    n1920,
    n1433,
    n1570,
    n1412,
    n1502
  );


  or
  g1750
  (
    n1912,
    n1439,
    n1713,
    n1539,
    n1663
  );


  or
  g1751
  (
    n1769,
    n1678,
    n1377,
    n1592,
    n1468
  );


  nor
  g1752
  (
    n1783,
    n1593,
    n1715,
    n1532,
    n1498
  );


  xnor
  g1753
  (
    n1893,
    n1510,
    n1518,
    n1708,
    n1678
  );


  xnor
  g1754
  (
    n1835,
    n1421,
    n1669,
    n1504,
    n1637
  );


  or
  g1755
  (
    n1918,
    n1600,
    n1438,
    n1572,
    n1554
  );


  and
  g1756
  (
    n1749,
    n1490,
    n1587,
    n1531,
    n1564
  );


  and
  g1757
  (
    n1737,
    n1469,
    n1730,
    n1461,
    n1725
  );


  or
  g1758
  (
    n1863,
    n1670,
    n1730,
    n1709,
    n1429
  );


  xor
  g1759
  (
    n1940,
    n1463,
    n1441,
    n1653,
    n1425
  );


  nor
  g1760
  (
    n1881,
    n1481,
    n1727,
    n1596,
    n1419
  );


  or
  g1761
  (
    n1806,
    n1406,
    n1411,
    n1627,
    n1696
  );


  nand
  g1762
  (
    n1875,
    n1494,
    n1543,
    n1544,
    n1698
  );


  xor
  g1763
  (
    n1776,
    n1548,
    n1456,
    n1417,
    n1554
  );


  xor
  g1764
  (
    n1812,
    n1546,
    n1653,
    n1471,
    n1639
  );


  xor
  g1765
  (
    n1780,
    n1542,
    n1512,
    n1686,
    n1690
  );


  nand
  g1766
  (
    n1816,
    n1571,
    n1484,
    n1476,
    n1560
  );


  xnor
  g1767
  (
    n1928,
    n1452,
    n1407,
    n1640,
    n1657
  );


  or
  g1768
  (
    n1764,
    n1691,
    n1598,
    n1647,
    n1398
  );


  or
  g1769
  (
    n1930,
    n1673,
    n1660,
    n1653,
    n1644
  );


  xnor
  g1770
  (
    n1786,
    n1538,
    n1668,
    n1594,
    n1676
  );


  and
  g1771
  (
    n1935,
    n1505,
    n1532,
    n1546,
    n1537
  );


  xor
  g1772
  (
    n1916,
    n1690,
    n1621,
    n1614,
    n1535
  );


  nor
  g1773
  (
    n1754,
    n1648,
    n1426,
    n1697,
    n1671
  );


  xor
  g1774
  (
    n1814,
    n1613,
    n1378,
    n1430,
    n1731
  );


  nand
  g1775
  (
    n1760,
    n1699,
    n1401,
    n1466,
    n1505
  );


  or
  g1776
  (
    n1767,
    n1573,
    n1622,
    n1663,
    n1448
  );


  nand
  g1777
  (
    n1839,
    n1394,
    n1533,
    n1615,
    n1497
  );


  xor
  g1778
  (
    n1779,
    n1475,
    n1461,
    n1584,
    n1482
  );


  xor
  g1779
  (
    n1902,
    n1666,
    n1448,
    n1602,
    n1705
  );


  or
  g1780
  (
    n1889,
    n1721,
    n1561,
    n1666,
    n1665
  );


  nor
  g1781
  (
    n1746,
    n1577,
    n1430,
    n1595,
    n1605
  );


  and
  g1782
  (
    n1851,
    n1530,
    n1582,
    n1370,
    n1520
  );


  or
  g1783
  (
    n1813,
    n1526,
    n1703,
    n1674,
    n1523
  );


  xor
  g1784
  (
    n1761,
    n1650,
    n1624,
    n1694,
    n1464
  );


  xnor
  g1785
  (
    n1897,
    n1691,
    n1621,
    n1562,
    n1609
  );


  and
  g1786
  (
    n1850,
    n1513,
    n1422,
    n1580,
    n1453
  );


  nand
  g1787
  (
    n1910,
    n1528,
    n1408,
    n1610,
    n1680
  );


  xor
  g1788
  (
    n1755,
    n1370,
    n1716,
    n1379
  );


  xnor
  g1789
  (
    n1871,
    n1633,
    n1411,
    n1642,
    n1625
  );


  and
  g1790
  (
    n1890,
    n1570,
    n1679,
    n1626,
    n1648
  );


  xnor
  g1791
  (
    n1810,
    n1723,
    n1433,
    n1722,
    n1443
  );


  xnor
  g1792
  (
    n1900,
    n1599,
    n1593,
    n1470,
    n1629
  );


  xnor
  g1793
  (
    n1750,
    n1671,
    n1390,
    n1432,
    n1391
  );


  nand
  g1794
  (
    n1852,
    n1726,
    n1585,
    n1385,
    n1685
  );


  nand
  g1795
  (
    n1738,
    n1393,
    n1673,
    n1575,
    n1531
  );


  or
  g1796
  (
    n1751,
    n1727,
    n1686,
    n1585,
    n1575
  );


  nor
  g1797
  (
    n1775,
    n1533,
    n1455,
    n1501,
    n1526
  );


  nand
  g1798
  (
    n1778,
    n1374,
    n1643,
    n1634,
    n1608
  );


  or
  g1799
  (
    n1845,
    n1603,
    n1637,
    n1467,
    n1402
  );


  nor
  g1800
  (
    n1919,
    n1661,
    n1620,
    n1555,
    n1566
  );


  nand
  g1801
  (
    n1848,
    n1508,
    n1683,
    n1402,
    n1631
  );


  or
  g1802
  (
    n1745,
    n1556,
    n1642,
    n1450,
    n1569
  );


  and
  g1803
  (
    n1854,
    n1458,
    n1442,
    n1732,
    n1590
  );


  nand
  g1804
  (
    n1809,
    n1478,
    n1657,
    n1517,
    n1494
  );


  xnor
  g1805
  (
    n1791,
    n1695,
    n1375,
    n1405,
    n1439
  );


  nand
  g1806
  (
    n1773,
    n1698,
    n1446,
    n1478,
    n1450
  );


  and
  g1807
  (
    n1846,
    n1654,
    n1679,
    n1423,
    n1387
  );


  nor
  g1808
  (
    n1826,
    n1686,
    n1616,
    n1567,
    n1664
  );


  xnor
  g1809
  (
    n1894,
    n1718,
    n1537,
    n1528,
    n1367
  );


  nand
  g1810
  (
    n1739,
    n1727,
    n1507,
    n1456,
    n1731
  );


  xor
  g1811
  (
    n1899,
    n1647,
    n1539,
    n1547,
    n1617
  );


  xor
  g1812
  (
    n1753,
    n1656,
    n1702,
    n1565,
    n1722
  );


  nor
  g1813
  (
    n1886,
    n1706,
    n1662,
    n1612,
    n1444
  );


  nor
  g1814
  (
    n1815,
    n1413,
    n1583,
    n1700,
    n1524
  );


  xor
  g1815
  (
    n1879,
    n1541,
    n1445,
    n1364,
    n1707
  );


  xor
  g1816
  (
    n1756,
    n1371,
    n1683,
    n1519,
    n1389
  );


  or
  g1817
  (
    n1774,
    n1631,
    n1676,
    n1691,
    n1396
  );


  nand
  g1818
  (
    n1834,
    n1467,
    n1509,
    n1733,
    n1431
  );


  or
  g1819
  (
    n1862,
    n1628,
    n1655,
    n1509,
    n1495
  );


  nor
  g1820
  (
    n1838,
    n1688,
    n1713,
    n1413,
    n1664
  );


  or
  g1821
  (
    n1926,
    n1578,
    n1707,
    n1724,
    n1733
  );


  or
  g1822
  (
    n1874,
    n1583,
    n1542,
    n1475,
    n1651
  );


  xnor
  g1823
  (
    n1741,
    n1452,
    n1669,
    n1503,
    n1723
  );


  and
  g1824
  (
    n1803,
    n1706,
    n1491,
    n1551,
    n1661
  );


  xor
  g1825
  (
    n1938,
    n1485,
    n1606,
    n1684,
    n1734
  );


  or
  g1826
  (
    n1849,
    n1639,
    n1474,
    n1709,
    n1529
  );


  xnor
  g1827
  (
    n1933,
    n1658,
    n1485,
    n1719,
    n1705
  );


  xnor
  g1828
  (
    n1805,
    n1690,
    n1558,
    n1692,
    n1728
  );


  xor
  g1829
  (
    n1837,
    n1733,
    n1373,
    n1689,
    n1688
  );


  nor
  g1830
  (
    n1911,
    n1426,
    n1561,
    n1487,
    n1685
  );


  xor
  g1831
  (
    n1811,
    n1479,
    n1362,
    n1414,
    n1705
  );


  xor
  g1832
  (
    n1742,
    n1592,
    n937,
    n1529,
    n1571
  );


  and
  g1833
  (
    n1772,
    n1435,
    n1672,
    n1550,
    n1563
  );


  nand
  g1834
  (
    n1793,
    n1405,
    n1629,
    n1486,
    n1628
  );


  nor
  g1835
  (
    n1818,
    n1607,
    n1420,
    n1572,
    n1688
  );


  or
  g1836
  (
    n1822,
    n1717,
    n1687,
    n1397,
    n1470
  );


  nand
  g1837
  (
    n1752,
    n1708,
    n1651,
    n1623,
    n1511
  );


  and
  g1838
  (
    n1909,
    n1383,
    n1672,
    n1696,
    n1367
  );


  and
  g1839
  (
    n1903,
    n1481,
    n1580,
    n1417,
    n1626
  );


  xnor
  g1840
  (
    n1799,
    n1680,
    n1675,
    n1559,
    n1654
  );


  xnor
  g1841
  (
    n1904,
    n1506,
    n1703,
    n1719,
    n1720
  );


  or
  g1842
  (
    n1927,
    n1601,
    n1428,
    n1650,
    n1454
  );


  xnor
  g1843
  (
    n1840,
    n1712,
    n1469,
    n1710,
    n1728
  );


  xor
  g1844
  (
    n1807,
    n1662,
    n1711,
    n1582,
    n1420
  );


  nand
  g1845
  (
    n1788,
    n1638,
    n1610,
    n1404,
    n1687
  );


  nor
  g1846
  (
    n1943,
    n1547,
    n1446,
    n1704,
    n1694
  );


  or
  g1847
  (
    n1853,
    n1641,
    n1617,
    n1545,
    n1440
  );


  xor
  g1848
  (
    n1876,
    n1701,
    n1520,
    n1702,
    n1562
  );


  xor
  g1849
  (
    n1923,
    n1668,
    n1573,
    n1489,
    n1436
  );


  xor
  g1850
  (
    n1844,
    n1732,
    n1675,
    n1574,
    n1551
  );


  xor
  g1851
  (
    n1787,
    n1568,
    n1714,
    n1578,
    n1389
  );


  or
  g1852
  (
    n1798,
    n1612,
    n1427,
    n1722,
    n1645
  );


  or
  g1853
  (
    n1794,
    n1491,
    n1714,
    n1436,
    n1449
  );


  and
  g1854
  (
    n1781,
    n1563,
    n1704,
    n1522,
    n1644
  );


  xnor
  g1855
  (
    n1792,
    n1381,
    n1383,
    n1646,
    n1483
  );


  xor
  g1856
  (
    n1836,
    n1496,
    n1660,
    n1703,
    n1376
  );


  and
  g1857
  (
    n1842,
    n1699,
    n1422,
    n1530,
    n1707
  );


  xor
  g1858
  (
    n1913,
    n1684,
    n1498,
    n1393,
    n1419
  );


  and
  g1859
  (
    n1796,
    n1591,
    n1566,
    n1719,
    n1510
  );


  nor
  g1860
  (
    n1887,
    n1677,
    n1645,
    n1680,
    n1514
  );


  xor
  g1861
  (
    n1736,
    n1710,
    n1427,
    n1683,
    n1681
  );


  xor
  g1862
  (
    n1915,
    n1525,
    n1368,
    n1364,
    n1715
  );


  xor
  g1863
  (
    n1941,
    n147,
    n1692,
    n1388,
    n1451
  );


  nor
  g1864
  (
    n1735,
    n1586,
    n1709,
    n1681,
    n1700
  );


  and
  g1865
  (
    n1829,
    n1716,
    n1473,
    n1695,
    n1708
  );


  and
  g1866
  (
    n1784,
    n1535,
    n1734,
    n1613,
    n1671
  );


  and
  g1867
  (
    n1768,
    n1506,
    n1380,
    n1630,
    n1362
  );


  xor
  g1868
  (
    n1936,
    n1720,
    n1552,
    n1646,
    n1724
  );


  and
  g1869
  (
    n1867,
    n1646,
    n1656,
    n1712,
    n1473
  );


  xnor
  g1870
  (
    n1797,
    n1553,
    n1508,
    n1636,
    n1504
  );


  nor
  g1871
  (
    n1771,
    n1513,
    n1523,
    n1710,
    n1511
  );


  nor
  g1872
  (
    n1945,
    n1594,
    n1689,
    n1447,
    n1377
  );


  xor
  g1873
  (
    n1880,
    n1652,
    n1403,
    n1589,
    n1410
  );


  nor
  g1874
  (
    n1740,
    n1647,
    n1697,
    n1721,
    n1657
  );


  xor
  g1875
  (
    n1944,
    n1640,
    n1462,
    n1464,
    n1725
  );


  nand
  g1876
  (
    n1748,
    n1637,
    n1611,
    n1712,
    n1635
  );


  nor
  g1877
  (
    n1924,
    n1650,
    n1665,
    n1471,
    n1540
  );


  xnor
  g1878
  (
    n1870,
    n1662,
    n1673,
    n1412,
    n1401
  );


  nor
  g1879
  (
    n1800,
    n1659,
    n1404,
    n1729,
    n1586
  );


  and
  g1880
  (
    n1801,
    n1604,
    n1579,
    n1444,
    n1655
  );


  xnor
  g1881
  (
    n1855,
    n1384,
    n1655,
    n1652,
    n1569
  );


  nor
  g1882
  (
    n1819,
    n1407,
    n1479,
    n1574,
    n1567
  );


  and
  g1883
  (
    n1824,
    n1483,
    n1616,
    n148,
    n1718
  );


  nor
  g1884
  (
    n1762,
    n1654,
    n1638,
    n1443,
    n1682
  );


  and
  g1885
  (
    n1757,
    n1603,
    n1472,
    n1576,
    n1552
  );


  and
  g1886
  (
    n1843,
    n1714,
    n1706,
    n1676,
    n1499
  );


  xor
  g1887
  (
    n1860,
    n1548,
    n1732,
    n1488,
    n1711
  );


  nor
  g1888
  (
    n1856,
    n1395,
    n1675,
    n1391,
    n1480
  );


  and
  g1889
  (
    n1942,
    n1482,
    n1472,
    n1400,
    n1693
  );


  or
  g1890
  (
    n1828,
    n1434,
    n1480,
    n1581
  );


  nand
  g1891
  (
    n1895,
    n1397,
    n1659,
    n1489,
    n1677
  );


  xnor
  g1892
  (
    n1865,
    n1445,
    n1718,
    n1602,
    n1694
  );


  xnor
  g1893
  (
    n1808,
    n1559,
    n1409,
    n1667,
    n1516
  );


  nor
  g1894
  (
    n1789,
    n1428,
    n1459,
    n1382,
    n1536
  );


  and
  g1895
  (
    n1905,
    n1663,
    n1541,
    n1577,
    n1495
  );


  nor
  g1896
  (
    n1763,
    n1375,
    n1534,
    n1403,
    n1648
  );


  and
  g1897
  (
    n1866,
    n1502,
    n1549,
    n1695,
    n1518
  );


  and
  g1898
  (
    n1892,
    n1437,
    n1659,
    n1416,
    n1724
  );


  nand
  g1899
  (
    n1946,
    n1682,
    n147,
    n1666,
    n1565
  );


  or
  g1900
  (
    n1744,
    n1366,
    n1728,
    n1515,
    n1618
  );


  nand
  g1901
  (
    n1759,
    n1682,
    n1624,
    n1406,
    n1702
  );


  xor
  g1902
  (
    n1908,
    n1667,
    n1692,
    n1689,
    n1538
  );


  and
  g1903
  (
    n1782,
    n1599,
    n1408,
    n1588,
    n1381
  );


  and
  g1904
  (
    n1847,
    n1558,
    n1704,
    n1425,
    n1604
  );


  xnor
  g1905
  (
    n1804,
    n1597,
    n1588,
    n1457,
    n1496
  );


  nand
  g1906
  (
    n1827,
    n1614,
    n1466,
    n1723,
    n1379
  );


  or
  g1907
  (
    n1914,
    n1368,
    n1560,
    n1500,
    n1409
  );


  nand
  g1908
  (
    n1758,
    n1625,
    n1726,
    n1713,
    n1457
  );


  xnor
  g1909
  (
    n1884,
    n1674,
    n1615,
    n1365,
    n1493
  );


  nand
  g1910
  (
    n1817,
    n1421,
    n1465,
    n1679,
    n1390
  );


  and
  g1911
  (
    n1802,
    n1656,
    n1374,
    n1668,
    n1670
  );


  xnor
  g1912
  (
    n1898,
    n1667,
    n1371,
    n1717,
    n1414
  );


  xnor
  g1913
  (
    n1878,
    n1369,
    n1536,
    n1477,
    n1640
  );


  nor
  g1914
  (
    n1962,
    n1774,
    n1736
  );


  nand
  g1915
  (
    n1952,
    n1765,
    n1773,
    n1748,
    n1789
  );


  and
  g1916
  (
    n1957,
    n1794,
    n1762,
    n1788,
    n1784
  );


  nand
  g1917
  (
    n1955,
    n1780,
    n1778,
    n1792,
    n1783
  );


  xnor
  g1918
  (
    n1958,
    n1777,
    n1735,
    n1745,
    n1766
  );


  nand
  g1919
  (
    n1953,
    n1739,
    n1767,
    n1781,
    n1772
  );


  xnor
  g1920
  (
    n1959,
    n1790,
    n1741,
    n1787,
    n1760
  );


  nand
  g1921
  (
    n1954,
    n1779,
    n1768,
    n1743,
    n1755
  );


  and
  g1922
  (
    n1947,
    n1749,
    n1763,
    n1756,
    n1795
  );


  nor
  g1923
  (
    n1956,
    n1737,
    n1770,
    n1751,
    n1791
  );


  xnor
  g1924
  (
    n1950,
    n1793,
    n1744,
    n1771,
    n1776
  );


  nand
  g1925
  (
    n1951,
    n1764,
    n1769,
    n1786,
    n1747
  );


  xor
  g1926
  (
    n1961,
    n1758,
    n1738,
    n1742,
    n1757
  );


  xnor
  g1927
  (
    n1960,
    n1759,
    n1746,
    n1752,
    n1754
  );


  xnor
  g1928
  (
    n1949,
    n1761,
    n1796,
    n1785,
    n1740
  );


  nor
  g1929
  (
    n1948,
    n1782,
    n1750,
    n1753,
    n1775
  );


  and
  g1930
  (
    n1971,
    n1894,
    n1812,
    n1961,
    n1841
  );


  xor
  g1931
  (
    n2008,
    n1959,
    n1958,
    n1940
  );


  and
  g1932
  (
    n1963,
    n1844,
    n1955,
    n1822,
    n1905
  );


  nand
  g1933
  (
    n1989,
    n1956,
    n1957,
    n1814,
    n32
  );


  nor
  g1934
  (
    n1997,
    n1874,
    n1823,
    n1956,
    n1961
  );


  nor
  g1935
  (
    n2000,
    n1926,
    n1940,
    n1939,
    n1924
  );


  nor
  g1936
  (
    n1984,
    n1886,
    n1847,
    n1951,
    n1911
  );


  nand
  g1937
  (
    n1992,
    n1956,
    n1831,
    n1888,
    n1959
  );


  xnor
  g1938
  (
    n1968,
    n1914,
    n1806,
    n1908,
    n1933
  );


  xor
  g1939
  (
    n1973,
    n1931,
    n1798,
    n1856,
    n1862
  );


  nor
  g1940
  (
    n1974,
    n1954,
    n1938,
    n1951,
    n1960
  );


  or
  g1941
  (
    n1996,
    n1945,
    n1827,
    n1901,
    n1937
  );


  and
  g1942
  (
    n1980,
    n1870,
    n1896,
    n1839,
    n32
  );


  nand
  g1943
  (
    n1981,
    n1849,
    n1953,
    n1734,
    n1958
  );


  or
  g1944
  (
    n2013,
    n1962,
    n1957,
    n1951,
    n148
  );


  xnor
  g1945
  (
    n2002,
    n1880,
    n1962,
    n1939,
    n1868
  );


  nand
  g1946
  (
    n1977,
    n1900,
    n1799,
    n1819,
    n1854
  );


  or
  g1947
  (
    n2007,
    n1941,
    n1800,
    n1953,
    n1928
  );


  or
  g1948
  (
    n1969,
    n31,
    n1950,
    n1804,
    n1955
  );


  nor
  g1949
  (
    n1976,
    n1865,
    n1957,
    n1930,
    n1892
  );


  xnor
  g1950
  (
    n2018,
    n1863,
    n31,
    n1871,
    n1867
  );


  or
  g1951
  (
    n2017,
    n1866,
    n1912,
    n1801,
    n1835
  );


  or
  g1952
  (
    n2012,
    n1815,
    n1920,
    n1813,
    n1953
  );


  xnor
  g1953
  (
    n1965,
    n1932,
    n1950,
    n1942,
    n1952
  );


  nand
  g1954
  (
    n1988,
    n1898,
    n1845,
    n1927,
    n1837
  );


  or
  g1955
  (
    n1986,
    n1954,
    n1936,
    n1913,
    n1891
  );


  xor
  g1956
  (
    n2001,
    n1873,
    n1949,
    n1848,
    n1842
  );


  xnor
  g1957
  (
    n1998,
    n32,
    n1959,
    n1952,
    n1948
  );


  xnor
  g1958
  (
    n2006,
    n1950,
    n1910,
    n1917,
    n1810
  );


  or
  g1959
  (
    n1987,
    n1805,
    n1923,
    n1859,
    n32
  );


  xor
  g1960
  (
    n2004,
    n1944,
    n1952,
    n1828,
    n1878
  );


  nor
  g1961
  (
    n1970,
    n1961,
    n1958,
    n1904,
    n1885
  );


  xor
  g1962
  (
    n2009,
    n1941,
    n1889,
    n1851,
    n1949
  );


  nor
  g1963
  (
    n1979,
    n1960,
    n1809,
    n1834,
    n1943
  );


  xor
  g1964
  (
    n1978,
    n1949,
    n1853,
    n1893,
    n1852
  );


  xor
  g1965
  (
    n2010,
    n148,
    n1947,
    n31,
    n1820
  );


  nor
  g1966
  (
    n1985,
    n1925,
    n1816,
    n1959,
    n1869
  );


  nand
  g1967
  (
    n1983,
    n1843,
    n1846,
    n1922,
    n1811
  );


  nor
  g1968
  (
    n2003,
    n1947,
    n1855,
    n1955,
    n1879
  );


  xor
  g1969
  (
    n1975,
    n1946,
    n1954,
    n1919
  );


  xor
  g1970
  (
    n1972,
    n1961,
    n1836,
    n1887,
    n1877
  );


  xor
  g1971
  (
    n2005,
    n1860,
    n1817,
    n1829,
    n1909
  );


  xor
  g1972
  (
    n1991,
    n1872,
    n1882,
    n1883,
    n1915
  );


  xor
  g1973
  (
    n1982,
    n1861,
    n1962,
    n1832,
    n1956
  );


  and
  g1974
  (
    n1990,
    n1942,
    n1876,
    n1934,
    n1826
  );


  and
  g1975
  (
    n2011,
    n1962,
    n1825,
    n1821,
    n1857
  );


  or
  g1976
  (
    n2014,
    n1875,
    n1858,
    n1921,
    n1797
  );


  or
  g1977
  (
    n2016,
    n1960,
    n1895,
    n1808,
    n1902
  );


  nand
  g1978
  (
    n1964,
    n1803,
    n1944,
    n1864,
    n1903
  );


  or
  g1979
  (
    n1993,
    n1906,
    n1929,
    n1918,
    n1960
  );


  or
  g1980
  (
    n1966,
    n1884,
    n1943,
    n1840,
    n1890
  );


  and
  g1981
  (
    n2015,
    n1907,
    n1850,
    n1802,
    n1838
  );


  nor
  g1982
  (
    n1967,
    n1948,
    n1833,
    n1946,
    n1935
  );


  and
  g1983
  (
    n1994,
    n1916,
    n1945,
    n1948,
    n1957
  );


  xnor
  g1984
  (
    n1999,
    n1807,
    n1955,
    n1830,
    n1897
  );


  xor
  g1985
  (
    n1995,
    n1824,
    n1881,
    n1899,
    n1818
  );


  xnor
  g1986
  (
    n2032,
    n1996,
    n2004,
    n2017,
    n1973
  );


  xor
  g1987
  (
    n2019,
    n2007,
    n2008,
    n1989,
    n1991
  );


  nand
  g1988
  (
    n2029,
    n1966,
    n1987,
    n1975,
    n1985
  );


  nor
  g1989
  (
    n2025,
    n1971,
    n2012,
    n2003,
    n1992
  );


  xor
  g1990
  (
    n2027,
    n2000,
    n1969,
    n2016,
    n2002
  );


  nor
  g1991
  (
    n2020,
    n2013,
    n1983,
    n1986,
    n2005
  );


  or
  g1992
  (
    n2030,
    n1984,
    n1974,
    n1978,
    n2001
  );


  nand
  g1993
  (
    n2021,
    n2009,
    n1993,
    n1964,
    n1970
  );


  nor
  g1994
  (
    n2022,
    n1980,
    n1994,
    n1995,
    n2011
  );


  xnor
  g1995
  (
    n2028,
    n1967,
    n1972,
    n2014,
    n2015
  );


  nor
  g1996
  (
    n2026,
    n1968,
    n1997,
    n1981,
    n1965
  );


  nor
  g1997
  (
    n2023,
    n1979,
    n1998,
    n1976,
    n1977
  );


  or
  g1998
  (
    n2024,
    n2010,
    n1990,
    n1988,
    n2018
  );


  nand
  g1999
  (
    n2031,
    n2006,
    n1982,
    n1963,
    n1999
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n882,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

