

module Stat_1000_103
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1024,
  n1017,
  n1020,
  n1012,
  n1008,
  n1005,
  n1025,
  n1016,
  n1007,
  n1027,
  n1011,
  n1026,
  n1031,
  n1023,
  n1003,
  n1014,
  n1021,
  n1019,
  n1009,
  n1028,
  n1013,
  n1006,
  n1001,
  n1002,
  n1015,
  n1022,
  n1032,
  n1018,
  n1004,
  n1029,
  n1010,
  n1030,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n1024;
  output n1017;
  output n1020;
  output n1012;
  output n1008;
  output n1005;
  output n1025;
  output n1016;
  output n1007;
  output n1027;
  output n1011;
  output n1026;
  output n1031;
  output n1023;
  output n1003;
  output n1014;
  output n1021;
  output n1019;
  output n1009;
  output n1028;
  output n1013;
  output n1006;
  output n1001;
  output n1002;
  output n1015;
  output n1022;
  output n1032;
  output n1018;
  output n1004;
  output n1029;
  output n1010;
  output n1030;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyNOTWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    n145,
    n6
  );


  not
  g1
  (
    n34,
    n16
  );


  not
  g2
  (
    n160,
    n23
  );


  not
  g3
  (
    n157,
    n24
  );


  buf
  g4
  (
    n131,
    n10
  );


  not
  g5
  (
    n147,
    n17
  );


  not
  g6
  (
    n45,
    n22
  );


  not
  g7
  (
    n59,
    n6
  );


  not
  g8
  (
    n117,
    n11
  );


  buf
  g9
  (
    n62,
    n4
  );


  not
  g10
  (
    n115,
    n4
  );


  not
  g11
  (
    n119,
    n26
  );


  buf
  g12
  (
    n77,
    n9
  );


  buf
  g13
  (
    n42,
    n32
  );


  not
  g14
  (
    n100,
    n32
  );


  buf
  g15
  (
    n54,
    n3
  );


  not
  g16
  (
    n101,
    n27
  );


  buf
  g17
  (
    n57,
    n13
  );


  not
  g18
  (
    n134,
    n31
  );


  not
  g19
  (
    n116,
    n1
  );


  buf
  g20
  (
    n123,
    n8
  );


  buf
  g21
  (
    n105,
    n26
  );


  buf
  g22
  (
    n152,
    n6
  );


  not
  g23
  (
    n83,
    n9
  );


  buf
  g24
  (
    n149,
    n3
  );


  not
  g25
  (
    n60,
    n15
  );


  buf
  g26
  (
    n78,
    n18
  );


  buf
  g27
  (
    n108,
    n2
  );


  buf
  g28
  (
    n88,
    n4
  );


  buf
  g29
  (
    n70,
    n3
  );


  buf
  g30
  (
    n144,
    n14
  );


  buf
  g31
  (
    n67,
    n28
  );


  buf
  g32
  (
    n53,
    n11
  );


  buf
  g33
  (
    n76,
    n2
  );


  not
  g34
  (
    n107,
    n12
  );


  not
  g35
  (
    n95,
    n25
  );


  buf
  g36
  (
    n151,
    n28
  );


  not
  g37
  (
    n73,
    n15
  );


  not
  g38
  (
    n143,
    n2
  );


  not
  g39
  (
    n137,
    n31
  );


  buf
  g40
  (
    n75,
    n8
  );


  buf
  g41
  (
    n159,
    n16
  );


  not
  g42
  (
    n154,
    n5
  );


  not
  g43
  (
    n85,
    n7
  );


  not
  g44
  (
    n113,
    n30
  );


  buf
  g45
  (
    n132,
    n26
  );


  not
  g46
  (
    n71,
    n8
  );


  buf
  g47
  (
    n94,
    n23
  );


  not
  g48
  (
    KeyWire_0_20,
    n6
  );


  buf
  g49
  (
    n99,
    n30
  );


  buf
  g50
  (
    n40,
    n21
  );


  buf
  g51
  (
    n148,
    n29
  );


  not
  g52
  (
    n66,
    n27
  );


  buf
  g53
  (
    n140,
    n30
  );


  buf
  g54
  (
    n47,
    n22
  );


  not
  g55
  (
    n96,
    n20
  );


  buf
  g56
  (
    n43,
    n21
  );


  not
  g57
  (
    n102,
    n9
  );


  not
  g58
  (
    n86,
    n32
  );


  buf
  g59
  (
    n139,
    n16
  );


  buf
  g60
  (
    n61,
    n22
  );


  not
  g61
  (
    n52,
    n22
  );


  buf
  g62
  (
    KeyWire_0_59,
    n5
  );


  not
  g63
  (
    n93,
    n5
  );


  not
  g64
  (
    n121,
    n31
  );


  not
  g65
  (
    n36,
    n28
  );


  buf
  g66
  (
    n135,
    n25
  );


  buf
  g67
  (
    n138,
    n24
  );


  not
  g68
  (
    n82,
    n20
  );


  not
  g69
  (
    n87,
    n12
  );


  buf
  g70
  (
    n124,
    n5
  );


  buf
  g71
  (
    n63,
    n21
  );


  not
  g72
  (
    n158,
    n14
  );


  not
  g73
  (
    n58,
    n19
  );


  not
  g74
  (
    KeyWire_0_16,
    n15
  );


  buf
  g75
  (
    n103,
    n13
  );


  buf
  g76
  (
    n110,
    n27
  );


  buf
  g77
  (
    n129,
    n11
  );


  not
  g78
  (
    n79,
    n17
  );


  not
  g79
  (
    n56,
    n19
  );


  not
  g80
  (
    n48,
    n17
  );


  not
  g81
  (
    n127,
    n13
  );


  buf
  g82
  (
    n114,
    n2
  );


  buf
  g83
  (
    KeyWire_0_34,
    n25
  );


  buf
  g84
  (
    n89,
    n8
  );


  not
  g85
  (
    n128,
    n1
  );


  not
  g86
  (
    n133,
    n15
  );


  not
  g87
  (
    n122,
    n13
  );


  not
  g88
  (
    n141,
    n9
  );


  not
  g89
  (
    n118,
    n12
  );


  buf
  g90
  (
    n55,
    n19
  );


  buf
  g91
  (
    n37,
    n10
  );


  buf
  g92
  (
    KeyWire_0_19,
    n31
  );


  buf
  g93
  (
    n156,
    n28
  );


  buf
  g94
  (
    n92,
    n1
  );


  not
  g95
  (
    n64,
    n23
  );


  not
  g96
  (
    n65,
    n16
  );


  buf
  g97
  (
    n84,
    n24
  );


  buf
  g98
  (
    n130,
    n27
  );


  buf
  g99
  (
    n142,
    n12
  );


  buf
  g100
  (
    n146,
    n18
  );


  not
  g101
  (
    KeyWire_0_18,
    n14
  );


  buf
  g102
  (
    n72,
    n18
  );


  buf
  g103
  (
    n90,
    n7
  );


  buf
  g104
  (
    n91,
    n7
  );


  not
  g105
  (
    n126,
    n29
  );


  buf
  g106
  (
    n150,
    n26
  );


  not
  g107
  (
    n112,
    n1
  );


  buf
  g108
  (
    n68,
    n23
  );


  buf
  g109
  (
    n33,
    n21
  );


  not
  g110
  (
    n120,
    n18
  );


  not
  g111
  (
    n74,
    n20
  );


  buf
  g112
  (
    n51,
    n19
  );


  buf
  g113
  (
    n97,
    n20
  );


  buf
  g114
  (
    n46,
    n11
  );


  not
  g115
  (
    n98,
    n30
  );


  not
  g116
  (
    n111,
    n4
  );


  not
  g117
  (
    n109,
    n10
  );


  not
  g118
  (
    n69,
    n25
  );


  buf
  g119
  (
    n80,
    n29
  );


  buf
  g120
  (
    n125,
    n17
  );


  buf
  g121
  (
    n41,
    n32
  );


  not
  g122
  (
    KeyWire_0_21,
    n7
  );


  not
  g123
  (
    n153,
    n10
  );


  not
  g124
  (
    n104,
    n14
  );


  buf
  g125
  (
    n49,
    n3
  );


  buf
  g126
  (
    KeyWire_0_49,
    n29
  );


  not
  g127
  (
    KeyWire_0_30,
    n24
  );


  not
  g128
  (
    n294,
    n69
  );


  buf
  g129
  (
    n394,
    n75
  );


  not
  g130
  (
    n419,
    n112
  );


  buf
  g131
  (
    n300,
    n86
  );


  buf
  g132
  (
    n386,
    n125
  );


  buf
  g133
  (
    KeyWire_0_38,
    n112
  );


  buf
  g134
  (
    n485,
    n54
  );


  buf
  g135
  (
    n420,
    n78
  );


  not
  g136
  (
    KeyWire_0_53,
    n120
  );


  not
  g137
  (
    n208,
    n55
  );


  buf
  g138
  (
    KeyWire_0_37,
    n44
  );


  buf
  g139
  (
    n436,
    n85
  );


  not
  g140
  (
    n296,
    n85
  );


  buf
  g141
  (
    n343,
    n118
  );


  buf
  g142
  (
    n185,
    n54
  );


  buf
  g143
  (
    n166,
    n77
  );


  buf
  g144
  (
    n198,
    n123
  );


  not
  g145
  (
    n334,
    n70
  );


  not
  g146
  (
    n355,
    n69
  );


  not
  g147
  (
    n243,
    n74
  );


  buf
  g148
  (
    n517,
    n50
  );


  buf
  g149
  (
    n191,
    n60
  );


  not
  g150
  (
    n525,
    n60
  );


  buf
  g151
  (
    n324,
    n81
  );


  not
  g152
  (
    n384,
    n105
  );


  buf
  g153
  (
    n400,
    n52
  );


  buf
  g154
  (
    n427,
    n40
  );


  buf
  g155
  (
    n459,
    n93
  );


  not
  g156
  (
    n426,
    n105
  );


  buf
  g157
  (
    n197,
    n71
  );


  buf
  g158
  (
    n399,
    n112
  );


  buf
  g159
  (
    n402,
    n35
  );


  buf
  g160
  (
    n524,
    n34
  );


  buf
  g161
  (
    n377,
    n74
  );


  not
  g162
  (
    n266,
    n126
  );


  buf
  g163
  (
    n206,
    n51
  );


  buf
  g164
  (
    n240,
    n104
  );


  buf
  g165
  (
    n454,
    n44
  );


  buf
  g166
  (
    KeyWire_0_0,
    n83
  );


  not
  g167
  (
    n409,
    n88
  );


  not
  g168
  (
    n477,
    n39
  );


  not
  g169
  (
    n467,
    n80
  );


  not
  g170
  (
    n456,
    n94
  );


  not
  g171
  (
    n278,
    n83
  );


  not
  g172
  (
    KeyWire_0_32,
    n64
  );


  buf
  g173
  (
    n232,
    n80
  );


  not
  g174
  (
    n313,
    n73
  );


  not
  g175
  (
    KeyWire_0_24,
    n68
  );


  buf
  g176
  (
    n530,
    n102
  );


  not
  g177
  (
    n230,
    n90
  );


  not
  g178
  (
    n496,
    n39
  );


  not
  g179
  (
    n482,
    n68
  );


  not
  g180
  (
    n203,
    n108
  );


  buf
  g181
  (
    n209,
    n109
  );


  not
  g182
  (
    n455,
    n45
  );


  not
  g183
  (
    n210,
    n53
  );


  buf
  g184
  (
    n255,
    n86
  );


  buf
  g185
  (
    n319,
    n47
  );


  not
  g186
  (
    n219,
    n120
  );


  not
  g187
  (
    n483,
    n50
  );


  not
  g188
  (
    n336,
    n86
  );


  not
  g189
  (
    n171,
    n88
  );


  not
  g190
  (
    n441,
    n79
  );


  buf
  g191
  (
    n533,
    n51
  );


  buf
  g192
  (
    n186,
    n88
  );


  buf
  g193
  (
    n487,
    n37
  );


  not
  g194
  (
    n228,
    n82
  );


  not
  g195
  (
    n292,
    n87
  );


  not
  g196
  (
    n174,
    n103
  );


  not
  g197
  (
    n451,
    n81
  );


  not
  g198
  (
    n452,
    n107
  );


  buf
  g199
  (
    n453,
    n66
  );


  not
  g200
  (
    n225,
    n63
  );


  not
  g201
  (
    n463,
    n118
  );


  buf
  g202
  (
    n307,
    n51
  );


  buf
  g203
  (
    n254,
    n76
  );


  buf
  g204
  (
    n505,
    n117
  );


  buf
  g205
  (
    n393,
    n47
  );


  buf
  g206
  (
    n162,
    n56
  );


  not
  g207
  (
    n489,
    n114
  );


  not
  g208
  (
    KeyWire_0_46,
    n116
  );


  not
  g209
  (
    n207,
    n111
  );


  buf
  g210
  (
    n433,
    n54
  );


  buf
  g211
  (
    n305,
    n107
  );


  not
  g212
  (
    n301,
    n43
  );


  buf
  g213
  (
    n202,
    n115
  );


  not
  g214
  (
    n424,
    n52
  );


  not
  g215
  (
    n273,
    n95
  );


  buf
  g216
  (
    n371,
    n71
  );


  not
  g217
  (
    n217,
    n87
  );


  not
  g218
  (
    n309,
    n75
  );


  buf
  g219
  (
    n416,
    n121
  );


  buf
  g220
  (
    n182,
    n91
  );


  buf
  g221
  (
    n249,
    n103
  );


  buf
  g222
  (
    n381,
    n96
  );


  buf
  g223
  (
    n318,
    n50
  );


  not
  g224
  (
    n513,
    n111
  );


  not
  g225
  (
    KeyWire_0_60,
    n34
  );


  buf
  g226
  (
    n281,
    n58
  );


  buf
  g227
  (
    n368,
    n110
  );


  not
  g228
  (
    n448,
    n55
  );


  buf
  g229
  (
    n346,
    n97
  );


  not
  g230
  (
    n479,
    n104
  );


  buf
  g231
  (
    KeyWire_0_61,
    n105
  );


  buf
  g232
  (
    n231,
    n55
  );


  buf
  g233
  (
    n508,
    n47
  );


  not
  g234
  (
    n260,
    n36
  );


  buf
  g235
  (
    n366,
    n114
  );


  not
  g236
  (
    n196,
    n49
  );


  buf
  g237
  (
    n442,
    n48
  );


  buf
  g238
  (
    n507,
    n46
  );


  buf
  g239
  (
    n434,
    n110
  );


  buf
  g240
  (
    n311,
    n108
  );


  buf
  g241
  (
    n261,
    n59
  );


  not
  g242
  (
    n302,
    n71
  );


  not
  g243
  (
    n241,
    n50
  );


  buf
  g244
  (
    n474,
    n92
  );


  buf
  g245
  (
    n491,
    n38
  );


  buf
  g246
  (
    n326,
    n73
  );


  not
  g247
  (
    n445,
    n61
  );


  not
  g248
  (
    n526,
    n38
  );


  buf
  g249
  (
    KeyWire_0_2,
    n54
  );


  not
  g250
  (
    n520,
    n105
  );


  not
  g251
  (
    n527,
    n106
  );


  buf
  g252
  (
    KeyWire_0_22,
    n62
  );


  buf
  g253
  (
    n329,
    n120
  );


  not
  g254
  (
    n389,
    n123
  );


  not
  g255
  (
    n361,
    n120
  );


  buf
  g256
  (
    n413,
    n41
  );


  buf
  g257
  (
    n415,
    n70
  );


  buf
  g258
  (
    n330,
    n97
  );


  buf
  g259
  (
    n365,
    n95
  );


  buf
  g260
  (
    n164,
    n121
  );


  not
  g261
  (
    n481,
    n124
  );


  not
  g262
  (
    n170,
    n34
  );


  buf
  g263
  (
    n169,
    n41
  );


  not
  g264
  (
    n447,
    n63
  );


  buf
  g265
  (
    n475,
    n40
  );


  buf
  g266
  (
    n519,
    n77
  );


  buf
  g267
  (
    n175,
    n108
  );


  buf
  g268
  (
    n308,
    n84
  );


  not
  g269
  (
    n165,
    n61
  );


  not
  g270
  (
    n180,
    n119
  );


  buf
  g271
  (
    n177,
    n68
  );


  buf
  g272
  (
    n529,
    n89
  );


  buf
  g273
  (
    n504,
    n96
  );


  not
  g274
  (
    n316,
    n113
  );


  buf
  g275
  (
    n204,
    n84
  );


  not
  g276
  (
    n473,
    n35
  );


  buf
  g277
  (
    n417,
    n72
  );


  not
  g278
  (
    n512,
    n36
  );


  not
  g279
  (
    n471,
    n64
  );


  not
  g280
  (
    n468,
    n117
  );


  not
  g281
  (
    n276,
    n65
  );


  buf
  g282
  (
    n268,
    n35
  );


  not
  g283
  (
    n431,
    n75
  );


  not
  g284
  (
    n235,
    n98
  );


  buf
  g285
  (
    n347,
    n69
  );


  buf
  g286
  (
    n429,
    n103
  );


  buf
  g287
  (
    n299,
    n42
  );


  buf
  g288
  (
    n214,
    n125
  );


  buf
  g289
  (
    n398,
    n56
  );


  not
  g290
  (
    n488,
    n109
  );


  not
  g291
  (
    n353,
    n107
  );


  buf
  g292
  (
    n248,
    n80
  );


  buf
  g293
  (
    n161,
    n71
  );


  not
  g294
  (
    KeyWire_0_47,
    n125
  );


  buf
  g295
  (
    n221,
    n80
  );


  buf
  g296
  (
    n360,
    n91
  );


  buf
  g297
  (
    n211,
    n40
  );


  buf
  g298
  (
    n279,
    n59
  );


  buf
  g299
  (
    n460,
    n95
  );


  not
  g300
  (
    n335,
    n33
  );


  buf
  g301
  (
    n457,
    n94
  );


  buf
  g302
  (
    n163,
    n100
  );


  not
  g303
  (
    n262,
    n63
  );


  not
  g304
  (
    n523,
    n122
  );


  not
  g305
  (
    n500,
    n45
  );


  not
  g306
  (
    KeyWire_0_8,
    n96
  );


  not
  g307
  (
    n184,
    n124
  );


  not
  g308
  (
    n531,
    n83
  );


  not
  g309
  (
    n291,
    n92
  );


  buf
  g310
  (
    n282,
    n97
  );


  buf
  g311
  (
    n341,
    n113
  );


  not
  g312
  (
    n224,
    n123
  );


  buf
  g313
  (
    n369,
    n42
  );


  buf
  g314
  (
    n303,
    n53
  );


  not
  g315
  (
    n408,
    n62
  );


  buf
  g316
  (
    n338,
    n58
  );


  buf
  g317
  (
    n325,
    n42
  );


  buf
  g318
  (
    n256,
    n106
  );


  not
  g319
  (
    n193,
    n61
  );


  buf
  g320
  (
    n277,
    n35
  );


  not
  g321
  (
    n321,
    n81
  );


  buf
  g322
  (
    n480,
    n116
  );


  not
  g323
  (
    n484,
    n78
  );


  buf
  g324
  (
    n342,
    n58
  );


  not
  g325
  (
    n345,
    n39
  );


  not
  g326
  (
    n317,
    n45
  );


  buf
  g327
  (
    n287,
    n73
  );


  not
  g328
  (
    n444,
    n49
  );


  not
  g329
  (
    n357,
    n109
  );


  buf
  g330
  (
    n465,
    n116
  );


  not
  g331
  (
    n229,
    n74
  );


  buf
  g332
  (
    n476,
    n99
  );


  buf
  g333
  (
    n242,
    n51
  );


  buf
  g334
  (
    n337,
    n45
  );


  buf
  g335
  (
    n446,
    n79
  );


  not
  g336
  (
    n437,
    n76
  );


  buf
  g337
  (
    n315,
    n37
  );


  buf
  g338
  (
    n364,
    n91
  );


  not
  g339
  (
    n327,
    n101
  );


  not
  g340
  (
    n497,
    n101
  );


  not
  g341
  (
    n449,
    n56
  );


  buf
  g342
  (
    n323,
    n100
  );


  buf
  g343
  (
    n173,
    n46
  );


  not
  g344
  (
    n201,
    n84
  );


  buf
  g345
  (
    n199,
    n81
  );


  buf
  g346
  (
    KeyWire_0_48,
    n76
  );


  buf
  g347
  (
    n397,
    n44
  );


  buf
  g348
  (
    n227,
    n94
  );


  not
  g349
  (
    n438,
    n92
  );


  buf
  g350
  (
    n322,
    n79
  );


  buf
  g351
  (
    n295,
    n62
  );


  not
  g352
  (
    n352,
    n48
  );


  not
  g353
  (
    n430,
    n66
  );


  buf
  g354
  (
    n470,
    n59
  );


  buf
  g355
  (
    n403,
    n70
  );


  buf
  g356
  (
    n216,
    n98
  );


  not
  g357
  (
    n274,
    n75
  );


  buf
  g358
  (
    n469,
    n118
  );


  not
  g359
  (
    n250,
    n85
  );


  not
  g360
  (
    n267,
    n92
  );


  not
  g361
  (
    n306,
    n119
  );


  not
  g362
  (
    n220,
    n82
  );


  buf
  g363
  (
    n414,
    n83
  );


  not
  g364
  (
    n379,
    n43
  );


  not
  g365
  (
    n226,
    n115
  );


  buf
  g366
  (
    KeyWire_0_3,
    n62
  );


  not
  g367
  (
    n239,
    n72
  );


  not
  g368
  (
    n466,
    n111
  );


  buf
  g369
  (
    n298,
    n73
  );


  buf
  g370
  (
    n392,
    n104
  );


  buf
  g371
  (
    n189,
    n78
  );


  buf
  g372
  (
    n516,
    n47
  );


  not
  g373
  (
    n461,
    n67
  );


  not
  g374
  (
    n501,
    n112
  );


  buf
  g375
  (
    n304,
    n41
  );


  buf
  g376
  (
    n290,
    n122
  );


  buf
  g377
  (
    n506,
    n102
  );


  not
  g378
  (
    n511,
    n123
  );


  not
  g379
  (
    n222,
    n43
  );


  not
  g380
  (
    n258,
    n98
  );


  buf
  g381
  (
    n494,
    n91
  );


  buf
  g382
  (
    n532,
    n39
  );


  buf
  g383
  (
    n200,
    n90
  );


  not
  g384
  (
    n422,
    n61
  );


  not
  g385
  (
    n331,
    n33
  );


  not
  g386
  (
    n167,
    n38
  );


  not
  g387
  (
    n358,
    n57
  );


  not
  g388
  (
    n339,
    n113
  );


  buf
  g389
  (
    n406,
    n84
  );


  not
  g390
  (
    n236,
    n121
  );


  not
  g391
  (
    n458,
    n102
  );


  not
  g392
  (
    n275,
    n100
  );


  not
  g393
  (
    n411,
    n89
  );


  not
  g394
  (
    n396,
    n49
  );


  buf
  g395
  (
    n432,
    n57
  );


  not
  g396
  (
    n362,
    n89
  );


  buf
  g397
  (
    n499,
    n85
  );


  not
  g398
  (
    n401,
    n98
  );


  not
  g399
  (
    KeyWire_0_44,
    n41
  );


  not
  g400
  (
    n518,
    n57
  );


  buf
  g401
  (
    KeyWire_0_33,
    n34
  );


  buf
  g402
  (
    KeyWire_0_40,
    n33
  );


  not
  g403
  (
    n348,
    n65
  );


  buf
  g404
  (
    n359,
    n117
  );


  buf
  g405
  (
    n374,
    n82
  );


  not
  g406
  (
    n350,
    n101
  );


  not
  g407
  (
    KeyWire_0_4,
    n53
  );


  buf
  g408
  (
    n450,
    n67
  );


  not
  g409
  (
    n522,
    n63
  );


  buf
  g410
  (
    n195,
    n104
  );


  buf
  g411
  (
    KeyWire_0_27,
    n64
  );


  buf
  g412
  (
    n314,
    n72
  );


  not
  g413
  (
    n503,
    n36
  );


  not
  g414
  (
    n367,
    n90
  );


  buf
  g415
  (
    n247,
    n118
  );


  buf
  g416
  (
    n344,
    n76
  );


  buf
  g417
  (
    n190,
    n37
  );


  buf
  g418
  (
    n269,
    n67
  );


  not
  g419
  (
    n382,
    n113
  );


  not
  g420
  (
    n509,
    n124
  );


  buf
  g421
  (
    n237,
    n43
  );


  not
  g422
  (
    n478,
    n52
  );


  not
  g423
  (
    n443,
    n89
  );


  buf
  g424
  (
    n349,
    n88
  );


  not
  g425
  (
    n213,
    n114
  );


  not
  g426
  (
    n263,
    n101
  );


  buf
  g427
  (
    n312,
    n102
  );


  not
  g428
  (
    n390,
    n111
  );


  buf
  g429
  (
    n244,
    n56
  );


  not
  g430
  (
    n515,
    n79
  );


  not
  g431
  (
    n223,
    n59
  );


  buf
  g432
  (
    n259,
    n49
  );


  buf
  g433
  (
    n245,
    n36
  );


  buf
  g434
  (
    n412,
    n93
  );


  not
  g435
  (
    n383,
    n93
  );


  buf
  g436
  (
    n428,
    n97
  );


  not
  g437
  (
    n387,
    n99
  );


  not
  g438
  (
    n351,
    n38
  );


  buf
  g439
  (
    n404,
    n106
  );


  not
  g440
  (
    n283,
    n99
  );


  buf
  g441
  (
    n514,
    n107
  );


  buf
  g442
  (
    n238,
    n60
  );


  buf
  g443
  (
    n425,
    n86
  );


  buf
  g444
  (
    n297,
    n60
  );


  not
  g445
  (
    n320,
    n55
  );


  not
  g446
  (
    n192,
    n33
  );


  buf
  g447
  (
    n421,
    n53
  );


  buf
  g448
  (
    n233,
    n65
  );


  buf
  g449
  (
    KeyWire_0_9,
    n66
  );


  buf
  g450
  (
    n418,
    n70
  );


  buf
  g451
  (
    n179,
    n67
  );


  buf
  g452
  (
    n264,
    n69
  );


  buf
  g453
  (
    n176,
    n46
  );


  not
  g454
  (
    n521,
    n100
  );


  buf
  g455
  (
    n378,
    n64
  );


  not
  g456
  (
    n251,
    n65
  );


  buf
  g457
  (
    n486,
    n99
  );


  not
  g458
  (
    KeyWire_0_31,
    n77
  );


  not
  g459
  (
    n373,
    n124
  );


  buf
  g460
  (
    n272,
    n48
  );


  not
  g461
  (
    n385,
    n58
  );


  buf
  g462
  (
    n286,
    n93
  );


  not
  g463
  (
    n310,
    n74
  );


  not
  g464
  (
    n188,
    n37
  );


  not
  g465
  (
    n375,
    n96
  );


  buf
  g466
  (
    n372,
    n78
  );


  not
  g467
  (
    n356,
    n115
  );


  buf
  g468
  (
    n332,
    n122
  );


  not
  g469
  (
    n212,
    n77
  );


  not
  g470
  (
    n183,
    n109
  );


  not
  g471
  (
    n328,
    n82
  );


  buf
  g472
  (
    n462,
    n103
  );


  not
  g473
  (
    KeyWire_0_43,
    n72
  );


  not
  g474
  (
    n423,
    n119
  );


  buf
  g475
  (
    n495,
    n90
  );


  buf
  g476
  (
    n363,
    n42
  );


  buf
  g477
  (
    KeyWire_0_52,
    n115
  );


  buf
  g478
  (
    n498,
    n108
  );


  not
  g479
  (
    n388,
    n48
  );


  buf
  g480
  (
    n370,
    n95
  );


  buf
  g481
  (
    n246,
    n52
  );


  not
  g482
  (
    n253,
    n46
  );


  not
  g483
  (
    n178,
    n68
  );


  buf
  g484
  (
    n215,
    n121
  );


  not
  g485
  (
    n395,
    n40
  );


  not
  g486
  (
    n270,
    n114
  );


  not
  g487
  (
    n380,
    n119
  );


  buf
  g488
  (
    n280,
    n94
  );


  not
  g489
  (
    n293,
    n117
  );


  buf
  g490
  (
    KeyWire_0_55,
    n110
  );


  buf
  g491
  (
    n288,
    n106
  );


  buf
  g492
  (
    n234,
    n125
  );


  not
  g493
  (
    n492,
    n44
  );


  not
  g494
  (
    n289,
    n110
  );


  not
  g495
  (
    n528,
    n87
  );


  not
  g496
  (
    n194,
    n87
  );


  not
  g497
  (
    n435,
    n57
  );


  buf
  g498
  (
    n285,
    n116
  );


  buf
  g499
  (
    KeyWire_0_15,
    n122
  );


  not
  g500
  (
    n284,
    n66
  );


  not
  g501
  (
    n541,
    n164
  );


  buf
  g502
  (
    n540,
    n167
  );


  not
  g503
  (
    n537,
    n168
  );


  buf
  g504
  (
    n538,
    n166
  );


  not
  g505
  (
    n539,
    n163
  );


  buf
  g506
  (
    n543,
    n161
  );


  buf
  g507
  (
    n546,
    n161
  );


  not
  g508
  (
    n535,
    n162
  );


  buf
  g509
  (
    n542,
    n165
  );


  not
  g510
  (
    n544,
    n164
  );


  buf
  g511
  (
    n547,
    n162
  );


  not
  g512
  (
    n536,
    n167
  );


  not
  g513
  (
    n545,
    n163
  );


  not
  g514
  (
    KeyWire_0_13,
    n165
  );


  buf
  g515
  (
    KeyWire_0_6,
    n166
  );


  buf
  g516
  (
    n567,
    n538
  );


  not
  g517
  (
    n556,
    n174
  );


  buf
  g518
  (
    n580,
    n548
  );


  not
  g519
  (
    KeyWire_0_41,
    n182
  );


  not
  g520
  (
    n557,
    n169
  );


  not
  g521
  (
    n563,
    n179
  );


  not
  g522
  (
    n569,
    n176
  );


  buf
  g523
  (
    n553,
    n175
  );


  not
  g524
  (
    n559,
    n172
  );


  buf
  g525
  (
    n554,
    n180
  );


  not
  g526
  (
    n555,
    n547
  );


  not
  g527
  (
    n571,
    n537
  );


  not
  g528
  (
    n570,
    n548
  );


  not
  g529
  (
    n565,
    n534
  );


  not
  g530
  (
    n562,
    n540
  );


  not
  g531
  (
    n578,
    n543
  );


  buf
  g532
  (
    n551,
    n178
  );


  buf
  g533
  (
    n568,
    n539
  );


  buf
  g534
  (
    n566,
    n176
  );


  not
  g535
  (
    n579,
    n539
  );


  nor
  g536
  (
    n573,
    n538,
    n544
  );


  xnor
  g537
  (
    n576,
    n177,
    n171
  );


  nor
  g538
  (
    n577,
    n179,
    n548,
    n182,
    n541
  );


  nand
  g539
  (
    n549,
    n536,
    n543,
    n546,
    n169
  );


  and
  g540
  (
    n572,
    n168,
    n535,
    n546,
    n183
  );


  xnor
  g541
  (
    n564,
    n545,
    n175,
    n180,
    n542
  );


  nand
  g542
  (
    n550,
    n540,
    n171,
    n184,
    n534
  );


  xor
  g543
  (
    n558,
    n173,
    n542,
    n181,
    n537
  );


  and
  g544
  (
    n574,
    n170,
    n544,
    n545,
    n173
  );


  nor
  g545
  (
    n560,
    n178,
    n174,
    n172,
    n177
  );


  xnor
  g546
  (
    n552,
    n183,
    n170,
    n541,
    n547
  );


  xor
  g547
  (
    n575,
    n535,
    n181,
    n547,
    n536
  );


  not
  g548
  (
    n581,
    n159
  );


  xnor
  g549
  (
    n617,
    n552,
    n129,
    n155
  );


  or
  g550
  (
    n599,
    n550,
    n142,
    n137,
    n575
  );


  nand
  g551
  (
    n628,
    n566,
    n158,
    n141
  );


  nand
  g552
  (
    n586,
    n556,
    n128,
    n155,
    n159
  );


  and
  g553
  (
    n615,
    n566,
    n577,
    n155,
    n130
  );


  xnor
  g554
  (
    n601,
    n131,
    n156,
    n569,
    n149
  );


  or
  g555
  (
    n610,
    n127,
    n144,
    n568,
    n135
  );


  and
  g556
  (
    n627,
    n571,
    n159,
    n134,
    n140
  );


  or
  g557
  (
    n597,
    n576,
    n137,
    n160,
    n141
  );


  xor
  g558
  (
    n611,
    n148,
    n145,
    n144,
    n132
  );


  nor
  g559
  (
    n593,
    n553,
    n145,
    n160,
    n127
  );


  nand
  g560
  (
    n607,
    n568,
    n138,
    n145,
    n126
  );


  and
  g561
  (
    n620,
    n148,
    n147,
    n570,
    n150
  );


  xor
  g562
  (
    n624,
    n156,
    n128,
    n126,
    n555
  );


  or
  g563
  (
    n591,
    n154,
    n157,
    n142,
    n143
  );


  nand
  g564
  (
    n588,
    n129,
    n153,
    n133,
    n132
  );


  xor
  g565
  (
    n613,
    n146,
    n561,
    n152,
    n136
  );


  xnor
  g566
  (
    n606,
    n142,
    n133,
    n129,
    n562
  );


  xnor
  g567
  (
    n623,
    n151,
    n141,
    n549,
    n564
  );


  xor
  g568
  (
    n585,
    n133,
    n560,
    n134,
    n137
  );


  xnor
  g569
  (
    n582,
    n572,
    n158,
    n580,
    n154
  );


  xor
  g570
  (
    n618,
    n574,
    n138,
    n139,
    n145
  );


  and
  g571
  (
    n603,
    n141,
    n140,
    n142,
    n557
  );


  nor
  g572
  (
    n609,
    n136,
    n134,
    n135,
    n578
  );


  xnor
  g573
  (
    n600,
    n577,
    n148,
    n132,
    n147
  );


  xnor
  g574
  (
    n592,
    n149,
    n127,
    n152,
    n130
  );


  and
  g575
  (
    n604,
    n128,
    n576,
    n151,
    n156
  );


  nor
  g576
  (
    n583,
    n150,
    n155,
    n580,
    n579
  );


  xnor
  g577
  (
    n608,
    n135,
    n565,
    n156,
    n184
  );


  xor
  g578
  (
    n621,
    n154,
    n157,
    n132,
    n128
  );


  nand
  g579
  (
    n612,
    n143,
    n554,
    n579,
    n152
  );


  or
  g580
  (
    n622,
    n149,
    n139,
    n151,
    n129
  );


  xnor
  g581
  (
    n614,
    n127,
    n147,
    n572,
    n139
  );


  xnor
  g582
  (
    n598,
    n570,
    n131,
    n159,
    n573
  );


  nor
  g583
  (
    n596,
    n138,
    n146,
    n126,
    n143
  );


  or
  g584
  (
    n626,
    n569,
    n144,
    n150,
    n130
  );


  nand
  g585
  (
    n594,
    n136,
    n157,
    n151,
    n160
  );


  and
  g586
  (
    n616,
    n563,
    n130,
    n551,
    n131
  );


  nand
  g587
  (
    n590,
    n148,
    n137,
    n135,
    n147
  );


  nand
  g588
  (
    n625,
    n140,
    n157,
    n153,
    n138
  );


  xor
  g589
  (
    n602,
    n160,
    n149,
    n131,
    n559
  );


  or
  g590
  (
    n584,
    n152,
    n140,
    n578,
    n136
  );


  or
  g591
  (
    n605,
    n139,
    n158,
    n571,
    n146
  );


  xnor
  g592
  (
    n589,
    n153,
    n134,
    n150,
    n567
  );


  xnor
  g593
  (
    n595,
    n153,
    n133,
    n573,
    n558
  );


  nand
  g594
  (
    n587,
    n567,
    n574,
    n143,
    n575
  );


  xor
  g595
  (
    n619,
    n144,
    n146,
    n154,
    n565
  );


  xnor
  g596
  (
    n769,
    n246,
    n428,
    n285,
    n279
  );


  or
  g597
  (
    n807,
    n249,
    n304,
    n417,
    n289
  );


  nand
  g598
  (
    n638,
    n618,
    n430,
    n582,
    n213
  );


  xnor
  g599
  (
    KeyWire_0_28,
    n584,
    n315,
    n330,
    n269
  );


  xnor
  g600
  (
    n675,
    n380,
    n276,
    n364,
    n351
  );


  and
  g601
  (
    n810,
    n235,
    n411,
    n372,
    n207
  );


  nand
  g602
  (
    n713,
    n607,
    n367,
    n281,
    n604
  );


  xnor
  g603
  (
    n781,
    n602,
    n616,
    n322,
    n598
  );


  nor
  g604
  (
    n652,
    n432,
    n325,
    n233,
    n625
  );


  xor
  g605
  (
    n804,
    n311,
    n605,
    n410,
    n398
  );


  xnor
  g606
  (
    n635,
    n384,
    n241,
    n599,
    n219
  );


  xor
  g607
  (
    n703,
    n366,
    n308,
    n397,
    n215
  );


  and
  g608
  (
    n637,
    n365,
    n396,
    n298,
    n336
  );


  nand
  g609
  (
    KeyWire_0_42,
    n286,
    n323,
    n599,
    n400
  );


  xor
  g610
  (
    KeyWire_0_14,
    n185,
    n599,
    n387,
    n275
  );


  xor
  g611
  (
    n733,
    n618,
    n276,
    n262,
    n408
  );


  and
  g612
  (
    n661,
    n369,
    n423,
    n601,
    n387
  );


  nand
  g613
  (
    n654,
    n370,
    n583,
    n622,
    n595
  );


  or
  g614
  (
    n741,
    n194,
    n215,
    n195,
    n427
  );


  xor
  g615
  (
    n672,
    n399,
    n396,
    n258,
    n381
  );


  nand
  g616
  (
    n650,
    n360,
    n626,
    n384,
    n590
  );


  nand
  g617
  (
    n789,
    n366,
    n610,
    n585,
    n321
  );


  nor
  g618
  (
    n792,
    n415,
    n204,
    n342,
    n594
  );


  nor
  g619
  (
    n712,
    n244,
    n353,
    n200,
    n434
  );


  nand
  g620
  (
    n772,
    n191,
    n597,
    n598,
    n217
  );


  or
  g621
  (
    n734,
    n279,
    n299,
    n600,
    n388
  );


  and
  g622
  (
    n724,
    n375,
    n585,
    n384,
    n425
  );


  xor
  g623
  (
    n719,
    n257,
    n186,
    n342,
    n359
  );


  nand
  g624
  (
    n693,
    n374,
    n592,
    n431,
    n195
  );


  or
  g625
  (
    n641,
    n381,
    n583,
    n267,
    n404
  );


  and
  g626
  (
    KeyWire_0_17,
    n592,
    n240,
    n190,
    n365
  );


  and
  g627
  (
    n697,
    n604,
    n373,
    n418,
    n627
  );


  and
  g628
  (
    n629,
    n412,
    n613,
    n312,
    n232
  );


  and
  g629
  (
    n707,
    n263,
    n229,
    n372,
    n391
  );


  and
  g630
  (
    n680,
    n583,
    n305,
    n319,
    n626
  );


  nand
  g631
  (
    n720,
    n619,
    n264,
    n205,
    n227
  );


  and
  g632
  (
    n791,
    n380,
    n308,
    n406,
    n203
  );


  nand
  g633
  (
    n717,
    n303,
    n602,
    n407,
    n283
  );


  nand
  g634
  (
    n784,
    n258,
    n600,
    n259,
    n589
  );


  nand
  g635
  (
    n808,
    n313,
    n188,
    n289,
    n285
  );


  nand
  g636
  (
    n761,
    n290,
    n298,
    n251,
    n382
  );


  xnor
  g637
  (
    n766,
    n593,
    n619,
    n340,
    n364
  );


  or
  g638
  (
    n640,
    n601,
    n352,
    n241,
    n323
  );


  xor
  g639
  (
    n630,
    n286,
    n620,
    n347,
    n189
  );


  nor
  g640
  (
    n705,
    n331,
    n593,
    n261,
    n390
  );


  xor
  g641
  (
    n658,
    n603,
    n261,
    n226,
    n628
  );


  or
  g642
  (
    n753,
    n204,
    n584,
    n231,
    n617
  );


  xnor
  g643
  (
    KeyWire_0_7,
    n604,
    n292,
    n376,
    n277
  );


  xnor
  g644
  (
    n685,
    n387,
    n350,
    n347,
    n222
  );


  nand
  g645
  (
    n806,
    n581,
    n628,
    n357,
    n615
  );


  xor
  g646
  (
    KeyWire_0_12,
    n344,
    n349,
    n332,
    n328
  );


  nor
  g647
  (
    n696,
    n220,
    n314,
    n300,
    n252
  );


  or
  g648
  (
    n775,
    n586,
    n595,
    n296,
    n307
  );


  nand
  g649
  (
    n732,
    n605,
    n398,
    n217,
    n371
  );


  xor
  g650
  (
    n748,
    n197,
    n612,
    n594,
    n221
  );


  nor
  g651
  (
    n760,
    n366,
    n362,
    n211,
    n301
  );


  or
  g652
  (
    n715,
    n233,
    n268,
    n248,
    n198
  );


  and
  g653
  (
    KeyWire_0_25,
    n250,
    n414,
    n325,
    n318
  );


  nor
  g654
  (
    n723,
    n212,
    n346,
    n419,
    n402
  );


  and
  g655
  (
    n657,
    n412,
    n196,
    n343,
    n424
  );


  or
  g656
  (
    n721,
    n304,
    n327,
    n382,
    n256
  );


  or
  g657
  (
    n643,
    n311,
    n202,
    n406,
    n234
  );


  nor
  g658
  (
    n710,
    n411,
    n297,
    n612,
    n310
  );


  nand
  g659
  (
    n659,
    n592,
    n377,
    n238,
    n405
  );


  nor
  g660
  (
    n754,
    n395,
    n380,
    n605,
    n581
  );


  nor
  g661
  (
    n815,
    n602,
    n627,
    n225,
    n592
  );


  xnor
  g662
  (
    n737,
    n385,
    n274,
    n346,
    n378
  );


  and
  g663
  (
    n729,
    n374,
    n389,
    n350,
    n257
  );


  nor
  g664
  (
    n633,
    n255,
    n609,
    n269,
    n359
  );


  nor
  g665
  (
    n662,
    n400,
    n209,
    n392,
    n388
  );


  xor
  g666
  (
    n704,
    n418,
    n191,
    n622,
    n400
  );


  nor
  g667
  (
    n681,
    n406,
    n272,
    n337,
    n609
  );


  nand
  g668
  (
    n780,
    n596,
    n369,
    n589,
    n317
  );


  nor
  g669
  (
    n726,
    n193,
    n405,
    n208,
    n293
  );


  xnor
  g670
  (
    n798,
    n256,
    n377,
    n619,
    n620
  );


  and
  g671
  (
    n758,
    n421,
    n322,
    n231,
    n288
  );


  nand
  g672
  (
    n634,
    n588,
    n420,
    n303,
    n423
  );


  xnor
  g673
  (
    n777,
    n266,
    n333,
    n409,
    n582
  );


  nor
  g674
  (
    n788,
    n615,
    n302,
    n608,
    n382
  );


  xnor
  g675
  (
    n639,
    n392,
    n416,
    n225,
    n355
  );


  or
  g676
  (
    n631,
    n420,
    n594,
    n338,
    n324
  );


  nor
  g677
  (
    n664,
    n607,
    n265,
    n414,
    n356
  );


  and
  g678
  (
    n799,
    n287,
    n616,
    n393,
    n606
  );


  xor
  g679
  (
    n674,
    n343,
    n432,
    n429,
    n365
  );


  and
  g680
  (
    n790,
    n388,
    n613,
    n394,
    n620
  );


  or
  g681
  (
    n725,
    n430,
    n309,
    n591,
    n194
  );


  xnor
  g682
  (
    n689,
    n584,
    n598,
    n372,
    n317
  );


  nor
  g683
  (
    n809,
    n604,
    n273,
    n216,
    n211
  );


  or
  g684
  (
    n677,
    n422,
    n236,
    n377,
    n265
  );


  nand
  g685
  (
    n679,
    n198,
    n358,
    n433,
    n383
  );


  nand
  g686
  (
    n711,
    n368,
    n610,
    n586,
    n402
  );


  nor
  g687
  (
    n779,
    n354,
    n618,
    n282,
    n208
  );


  and
  g688
  (
    n814,
    n209,
    n623,
    n610,
    n606
  );


  or
  g689
  (
    n805,
    n207,
    n294,
    n245,
    n266
  );


  or
  g690
  (
    n671,
    n228,
    n214,
    n426,
    n353
  );


  and
  g691
  (
    n682,
    n363,
    n316,
    n603,
    n282
  );


  nor
  g692
  (
    n651,
    n415,
    n627,
    n288,
    n407
  );


  xor
  g693
  (
    n813,
    n583,
    n228,
    n597,
    n186
  );


  xnor
  g694
  (
    n770,
    n232,
    n330,
    n428,
    n414
  );


  xnor
  g695
  (
    n797,
    n433,
    n200,
    n278,
    n367
  );


  nand
  g696
  (
    n655,
    n223,
    n354,
    n416,
    n375
  );


  and
  g697
  (
    n660,
    n373,
    n326,
    n584,
    n293
  );


  and
  g698
  (
    n776,
    n267,
    n609,
    n251,
    n332
  );


  or
  g699
  (
    n708,
    n335,
    n612,
    n352,
    n296
  );


  nand
  g700
  (
    n714,
    n242,
    n421,
    n596,
    n606
  );


  or
  g701
  (
    n632,
    n320,
    n320,
    n334,
    n329
  );


  nor
  g702
  (
    n668,
    n611,
    n341,
    n614,
    n393
  );


  xor
  g703
  (
    n676,
    n386,
    n397,
    n588,
    n624
  );


  nand
  g704
  (
    n745,
    n621,
    n626,
    n284,
    n402
  );


  nor
  g705
  (
    n653,
    n278,
    n187,
    n290,
    n299
  );


  nor
  g706
  (
    n678,
    n240,
    n237,
    n202,
    n341
  );


  nand
  g707
  (
    n752,
    n610,
    n585,
    n606,
    n259
  );


  and
  g708
  (
    n730,
    n219,
    n218,
    n328,
    n415
  );


  nor
  g709
  (
    KeyWire_0_5,
    n254,
    n313,
    n431,
    n335
  );


  xnor
  g710
  (
    n787,
    n339,
    n295,
    n268,
    n427
  );


  xor
  g711
  (
    n667,
    n595,
    n603,
    n427,
    n401
  );


  and
  g712
  (
    n706,
    n395,
    n601,
    n401,
    n591
  );


  nor
  g713
  (
    n656,
    n331,
    n622,
    n260,
    n394
  );


  xor
  g714
  (
    n716,
    n242,
    n221,
    n581,
    n397
  );


  nor
  g715
  (
    n783,
    n621,
    n376,
    n389,
    n197
  );


  xor
  g716
  (
    n767,
    n609,
    n375,
    n587,
    n403
  );


  nor
  g717
  (
    n666,
    n612,
    n611,
    n422,
    n613
  );


  nor
  g718
  (
    n701,
    n420,
    n588,
    n607,
    n625
  );


  or
  g719
  (
    KeyWire_0_1,
    n199,
    n424,
    n274,
    n615
  );


  and
  g720
  (
    n751,
    n410,
    n391,
    n411,
    n602
  );


  nor
  g721
  (
    n687,
    n409,
    n199,
    n196,
    n315
  );


  and
  g722
  (
    n749,
    n409,
    n374,
    n404,
    n306
  );


  xor
  g723
  (
    n768,
    n300,
    n270,
    n364,
    n206
  );


  nand
  g724
  (
    n816,
    n255,
    n595,
    n403,
    n370
  );


  xor
  g725
  (
    n794,
    n248,
    n359,
    n246,
    n422
  );


  nor
  g726
  (
    n759,
    n203,
    n367,
    n608,
    n403
  );


  nand
  g727
  (
    n718,
    n386,
    n318,
    n433,
    n614
  );


  xor
  g728
  (
    n819,
    n376,
    n430,
    n625,
    n390
  );


  xnor
  g729
  (
    n699,
    n624,
    n357,
    n312,
    n192
  );


  and
  g730
  (
    n728,
    n361,
    n247,
    n249,
    n244
  );


  and
  g731
  (
    n636,
    n291,
    n434,
    n586,
    n316
  );


  or
  g732
  (
    n691,
    n396,
    n226,
    n611,
    n287
  );


  xnor
  g733
  (
    n818,
    n368,
    n608,
    n336,
    n213
  );


  xnor
  g734
  (
    n688,
    n424,
    n253,
    n413,
    n306
  );


  nor
  g735
  (
    n756,
    n363,
    n271,
    n264,
    n398
  );


  nor
  g736
  (
    n695,
    n239,
    n192,
    n385,
    n338
  );


  and
  g737
  (
    n742,
    n210,
    n379,
    n227,
    n371
  );


  nand
  g738
  (
    n743,
    n250,
    n408,
    n597,
    n613
  );


  xor
  g739
  (
    KeyWire_0_10,
    n628,
    n624,
    n247,
    n205
  );


  nand
  g740
  (
    n771,
    n294,
    n302,
    n324,
    n627
  );


  xnor
  g741
  (
    n642,
    n238,
    n301,
    n356,
    n587
  );


  nand
  g742
  (
    n665,
    n389,
    n607,
    n224,
    n235
  );


  xnor
  g743
  (
    n801,
    n337,
    n399,
    n410,
    n412
  );


  xnor
  g744
  (
    n750,
    n307,
    n230,
    n617,
    n297
  );


  nand
  g745
  (
    n663,
    n596,
    n582,
    n429,
    n349
  );


  nor
  g746
  (
    n786,
    n426,
    n362,
    n358,
    n621
  );


  and
  g747
  (
    n692,
    n236,
    n345,
    n419,
    n416
  );


  nand
  g748
  (
    n647,
    n405,
    n587,
    n362,
    n378
  );


  xnor
  g749
  (
    n709,
    n624,
    n622,
    n214,
    n587
  );


  xnor
  g750
  (
    KeyWire_0_26,
    n329,
    n421,
    n189,
    n237
  );


  and
  g751
  (
    n735,
    n425,
    n590,
    n361,
    n355
  );


  or
  g752
  (
    n785,
    n601,
    n585,
    n253,
    n210
  );


  xor
  g753
  (
    n736,
    n586,
    n385,
    n188,
    n399
  );


  xnor
  g754
  (
    n702,
    n611,
    n270,
    n190,
    n383
  );


  or
  g755
  (
    n796,
    n185,
    n392,
    n426,
    n321
  );


  nand
  g756
  (
    KeyWire_0_63,
    n419,
    n619,
    n348,
    n394
  );


  nor
  g757
  (
    n802,
    n272,
    n277,
    n594,
    n361
  );


  xnor
  g758
  (
    n757,
    n623,
    n327,
    n284,
    n617
  );


  xor
  g759
  (
    n765,
    n326,
    n234,
    n360,
    n589
  );


  or
  g760
  (
    n811,
    n423,
    n391,
    n281,
    n222
  );


  nand
  g761
  (
    n694,
    n379,
    n310,
    n344,
    n616
  );


  nor
  g762
  (
    n773,
    n589,
    n223,
    n368,
    n252
  );


  xor
  g763
  (
    KeyWire_0_51,
    n407,
    n254,
    n360,
    n401
  );


  nand
  g764
  (
    n739,
    n614,
    n220,
    n620,
    n370
  );


  xnor
  g765
  (
    n755,
    n418,
    n597,
    n334,
    n340
  );


  xor
  g766
  (
    n686,
    n600,
    n305,
    n617,
    n603
  );


  nor
  g767
  (
    n700,
    n333,
    n596,
    n363,
    n588
  );


  nand
  g768
  (
    n763,
    n206,
    n230,
    n605,
    n386
  );


  xnor
  g769
  (
    n803,
    n431,
    n623,
    n591,
    n593
  );


  and
  g770
  (
    n684,
    n383,
    n201,
    n291,
    n273
  );


  nor
  g771
  (
    KeyWire_0_35,
    n309,
    n615,
    n351,
    n339
  );


  nand
  g772
  (
    n820,
    n600,
    n239,
    n187,
    n413
  );


  or
  g773
  (
    n648,
    n369,
    n280,
    n582,
    n621
  );


  nor
  g774
  (
    n762,
    n245,
    n590,
    n432,
    n358
  );


  or
  g775
  (
    n778,
    n314,
    n243,
    n260,
    n425
  );


  nor
  g776
  (
    n690,
    n608,
    n591,
    n614,
    n628
  );


  and
  g777
  (
    n812,
    n345,
    n373,
    n283,
    n381
  );


  xnor
  g778
  (
    n747,
    n417,
    n201,
    n395,
    n616
  );


  nor
  g779
  (
    KeyWire_0_56,
    n393,
    n229,
    n428,
    n275
  );


  xnor
  g780
  (
    n645,
    n271,
    n348,
    n599,
    n408
  );


  or
  g781
  (
    n774,
    n263,
    n593,
    n598,
    n378
  );


  and
  g782
  (
    n764,
    n404,
    n623,
    n371,
    n581
  );


  or
  g783
  (
    n793,
    n379,
    n417,
    n413,
    n390
  );


  nor
  g784
  (
    n746,
    n280,
    n216,
    n590,
    n224
  );


  and
  g785
  (
    n683,
    n429,
    n212,
    n292,
    n625
  );


  nand
  g786
  (
    n740,
    n243,
    n295,
    n218,
    n618
  );


  nand
  g787
  (
    n722,
    n626,
    n262,
    n319,
    n193
  );


  nor
  g788
  (
    n889,
    n450,
    n446,
    n680
  );


  xnor
  g789
  (
    n896,
    n751,
    n694,
    n723,
    n481
  );


  and
  g790
  (
    n870,
    n479,
    n631,
    n688,
    n441
  );


  nand
  g791
  (
    n895,
    n482,
    n443,
    n752,
    n731
  );


  xor
  g792
  (
    n869,
    n746,
    n466,
    n739,
    n747
  );


  and
  g793
  (
    n863,
    n658,
    n467,
    n719,
    n718
  );


  xnor
  g794
  (
    n891,
    n482,
    n459,
    n455,
    n726
  );


  xnor
  g795
  (
    n829,
    n676,
    n467,
    n719,
    n705
  );


  xnor
  g796
  (
    n872,
    n703,
    n634,
    n444,
    n708
  );


  and
  g797
  (
    n883,
    n475,
    n737,
    n705,
    n460
  );


  or
  g798
  (
    n834,
    n749,
    n752,
    n739,
    n717
  );


  xor
  g799
  (
    n821,
    n468,
    n730,
    n448,
    n669
  );


  nor
  g800
  (
    n842,
    n469,
    n648,
    n735,
    n477
  );


  nor
  g801
  (
    KeyWire_0_62,
    n724,
    n629,
    n445,
    n704
  );


  xnor
  g802
  (
    n901,
    n753,
    n654,
    n438,
    n732
  );


  nand
  g803
  (
    n904,
    n464,
    n722,
    n652,
    n483
  );


  nand
  g804
  (
    n899,
    n714,
    n468,
    n734,
    n445
  );


  nand
  g805
  (
    n850,
    n711,
    n650,
    n447,
    n693
  );


  xor
  g806
  (
    n890,
    n734,
    n730,
    n703,
    n738
  );


  nand
  g807
  (
    n897,
    n720,
    n461,
    n463,
    n671
  );


  nor
  g808
  (
    n825,
    n720,
    n436,
    n651,
    n449
  );


  nand
  g809
  (
    n846,
    n732,
    n691,
    n684,
    n456
  );


  xnor
  g810
  (
    n868,
    n642,
    n667,
    n710,
    n466
  );


  nand
  g811
  (
    n884,
    n443,
    n449,
    n715,
    n462
  );


  nor
  g812
  (
    n903,
    n481,
    n461,
    n701,
    n483
  );


  or
  g813
  (
    n855,
    n662,
    n750,
    n475,
    n471
  );


  nand
  g814
  (
    n854,
    n630,
    n451,
    n440,
    n458
  );


  nand
  g815
  (
    n865,
    n702,
    n485,
    n456,
    n447
  );


  xnor
  g816
  (
    n885,
    n673,
    n687,
    n458,
    n663
  );


  or
  g817
  (
    n822,
    n641,
    n744,
    n476,
    n735
  );


  xnor
  g818
  (
    n827,
    n450,
    n701,
    n467,
    n440
  );


  nor
  g819
  (
    n849,
    n710,
    n683,
    n745,
    n460
  );


  xor
  g820
  (
    n881,
    n713,
    n475,
    n738,
    n472
  );


  and
  g821
  (
    n877,
    n485,
    n736,
    n465,
    n453
  );


  nor
  g822
  (
    n898,
    n706,
    n477,
    n714,
    n677
  );


  nand
  g823
  (
    n873,
    n440,
    n480,
    n674,
    n449
  );


  and
  g824
  (
    n862,
    n453,
    n653,
    n479,
    n438
  );


  xnor
  g825
  (
    n864,
    n468,
    n640,
    n482,
    n462
  );


  nor
  g826
  (
    n875,
    n457,
    n479,
    n435,
    n713
  );


  nand
  g827
  (
    n857,
    n721,
    n476,
    n463,
    n692
  );


  nor
  g828
  (
    n847,
    n478,
    n733,
    n698,
    n633
  );


  xnor
  g829
  (
    n838,
    n726,
    n477,
    n462,
    n459
  );


  and
  g830
  (
    n878,
    n457,
    n478,
    n473,
    n731
  );


  xor
  g831
  (
    n826,
    n472,
    n454,
    n727,
    n723
  );


  and
  g832
  (
    n893,
    n465,
    n753,
    n736,
    n439
  );


  xor
  g833
  (
    KeyWire_0_57,
    n451,
    n724,
    n708,
    n452
  );


  xnor
  g834
  (
    n880,
    n712,
    n469,
    n484,
    n747
  );


  and
  g835
  (
    n882,
    n469,
    n750,
    n727,
    n442
  );


  and
  g836
  (
    n874,
    n670,
    n453,
    n452,
    n743
  );


  nand
  g837
  (
    n839,
    n434,
    n473,
    n446,
    n741
  );


  xnor
  g838
  (
    n900,
    n480,
    n438,
    n442,
    n660
  );


  xnor
  g839
  (
    n871,
    n442,
    n483,
    n685,
    n718
  );


  nor
  g840
  (
    n886,
    n455,
    n444,
    n644,
    n668
  );


  nor
  g841
  (
    n894,
    n435,
    n729,
    n452,
    n679
  );


  nand
  g842
  (
    n833,
    n649,
    n743,
    n472,
    n484
  );


  xor
  g843
  (
    n841,
    n655,
    n721,
    n446,
    n742
  );


  xnor
  g844
  (
    n844,
    n725,
    n740,
    n733,
    n456
  );


  xnor
  g845
  (
    n830,
    n672,
    n437,
    n457
  );


  xor
  g846
  (
    n858,
    n441,
    n448,
    n635
  );


  or
  g847
  (
    n848,
    n450,
    n439,
    n666,
    n711
  );


  nand
  g848
  (
    n860,
    n741,
    n725,
    n704,
    n455
  );


  xor
  g849
  (
    n832,
    n436,
    n484,
    n678,
    n461
  );


  xor
  g850
  (
    n879,
    n745,
    n435,
    n746,
    n458
  );


  and
  g851
  (
    n835,
    n700,
    n695,
    n699,
    n643
  );


  nand
  g852
  (
    n866,
    n696,
    n751,
    n485,
    n445
  );


  and
  g853
  (
    KeyWire_0_45,
    n645,
    n690,
    n709,
    n451
  );


  nor
  g854
  (
    n853,
    n647,
    n748,
    n636,
    n664
  );


  or
  g855
  (
    n824,
    n470,
    n480,
    n682,
    n689
  );


  nand
  g856
  (
    n861,
    n742,
    n439,
    n748,
    n728
  );


  nand
  g857
  (
    n840,
    n675,
    n471,
    n459,
    n470
  );


  xor
  g858
  (
    n888,
    n481,
    n637,
    n646,
    n717
  );


  and
  g859
  (
    n836,
    n436,
    n656,
    n447,
    n702
  );


  xnor
  g860
  (
    n828,
    n737,
    n698,
    n638,
    n639
  );


  nor
  g861
  (
    n823,
    n709,
    n686,
    n470,
    n454
  );


  xnor
  g862
  (
    KeyWire_0_29,
    n699,
    n749,
    n478,
    n632
  );


  or
  g863
  (
    KeyWire_0_11,
    n707,
    n716,
    n657
  );


  xor
  g864
  (
    n859,
    n661,
    n715,
    n441,
    n722
  );


  nor
  g865
  (
    n831,
    n444,
    n463,
    n465,
    n460
  );


  xnor
  g866
  (
    n867,
    n476,
    n473,
    n740,
    n474
  );


  nand
  g867
  (
    n851,
    n700,
    n437,
    n454,
    n659
  );


  xor
  g868
  (
    n856,
    n471,
    n706,
    n474,
    n665
  );


  or
  g869
  (
    n852,
    n707,
    n466,
    n697,
    n474
  );


  and
  g870
  (
    n887,
    n728,
    n712,
    n729,
    n681
  );


  nor
  g871
  (
    n902,
    n744,
    n464,
    n443
  );


  nand
  g872
  (
    n928,
    n767,
    n755,
    n889,
    n757
  );


  and
  g873
  (
    n930,
    n842,
    n761,
    n859,
    n825
  );


  nor
  g874
  (
    n927,
    n757,
    n759,
    n892,
    n832
  );


  or
  g875
  (
    n920,
    n755,
    n847,
    n831,
    n769
  );


  and
  g876
  (
    KeyWire_0_58,
    n871,
    n764,
    n767,
    n844
  );


  nor
  g877
  (
    n919,
    n770,
    n861,
    n766,
    n875
  );


  nor
  g878
  (
    n931,
    n874,
    n860,
    n835,
    n754
  );


  xnor
  g879
  (
    n915,
    n756,
    n821,
    n771,
    n853
  );


  nand
  g880
  (
    n916,
    n758,
    n893,
    n837,
    n888
  );


  xnor
  g881
  (
    n911,
    n851,
    n858,
    n823,
    n824
  );


  and
  g882
  (
    n932,
    n879,
    n840,
    n882,
    n761
  );


  nor
  g883
  (
    n908,
    n893,
    n770,
    n829,
    n890
  );


  or
  g884
  (
    n914,
    n870,
    n872,
    n856,
    n852
  );


  xnor
  g885
  (
    n912,
    n830,
    n892,
    n839,
    n854
  );


  nor
  g886
  (
    n922,
    n841,
    n869,
    n876,
    n765
  );


  nand
  g887
  (
    n923,
    n862,
    n887,
    n891,
    n769
  );


  nor
  g888
  (
    n921,
    n754,
    n891,
    n836,
    n762
  );


  or
  g889
  (
    n909,
    n765,
    n877,
    n885,
    n886
  );


  xnor
  g890
  (
    n910,
    n846,
    n771,
    n822,
    n867
  );


  xnor
  g891
  (
    n925,
    n855,
    n766,
    n880,
    n884
  );


  and
  g892
  (
    n918,
    n843,
    n760,
    n865,
    n763
  );


  or
  g893
  (
    n905,
    n826,
    n764,
    n827,
    n834
  );


  or
  g894
  (
    n906,
    n863,
    n828,
    n768,
    n838
  );


  xnor
  g895
  (
    n913,
    n878,
    n848,
    n868,
    n759
  );


  nand
  g896
  (
    n917,
    n756,
    n763,
    n768,
    n864
  );


  nor
  g897
  (
    n929,
    n849,
    n845,
    n760,
    n833
  );


  xor
  g898
  (
    n926,
    n873,
    n883,
    n850,
    n758
  );


  xor
  g899
  (
    n924,
    n881,
    n866,
    n762,
    n857
  );


  or
  g900
  (
    n959,
    n908,
    n526,
    n900,
    n508
  );


  and
  g901
  (
    n980,
    n490,
    n507,
    n906,
    n504
  );


  or
  g902
  (
    n952,
    n913,
    n533,
    n490,
    n512
  );


  and
  g903
  (
    n943,
    n898,
    n488,
    n503,
    n904
  );


  xnor
  g904
  (
    n937,
    n487,
    n498,
    n497
  );


  and
  g905
  (
    n957,
    n785,
    n531,
    n528,
    n506
  );


  xor
  g906
  (
    n999,
    n530,
    n488,
    n912,
    n780
  );


  or
  g907
  (
    n1000,
    n905,
    n511,
    n489,
    n932
  );


  nor
  g908
  (
    n998,
    n775,
    n932,
    n505,
    n780
  );


  or
  g909
  (
    n987,
    n517,
    n486,
    n903,
    n495
  );


  and
  g910
  (
    n949,
    n921,
    n492,
    n923
  );


  nor
  g911
  (
    n939,
    n782,
    n516,
    n925,
    n928
  );


  nand
  g912
  (
    n990,
    n521,
    n513,
    n508,
    n533
  );


  or
  g913
  (
    n965,
    n899,
    n924,
    n919,
    n529
  );


  xor
  g914
  (
    KeyWire_0_36,
    n500,
    n514,
    n789,
    n907
  );


  nand
  g915
  (
    n981,
    n509,
    n533,
    n492,
    n503
  );


  nand
  g916
  (
    n935,
    n510,
    n906,
    n777,
    n496
  );


  nor
  g917
  (
    n984,
    n914,
    n529,
    n526,
    n496
  );


  and
  g918
  (
    KeyWire_0_54,
    n532,
    n530,
    n510,
    n494
  );


  nand
  g919
  (
    n960,
    n929,
    n923,
    n527,
    n517
  );


  or
  g920
  (
    n955,
    n911,
    n529,
    n774,
    n511
  );


  or
  g921
  (
    n977,
    n500,
    n501,
    n927,
    n907
  );


  nand
  g922
  (
    n988,
    n521,
    n912,
    n896,
    n498
  );


  xnor
  g923
  (
    n974,
    n897,
    n782,
    n909,
    n775
  );


  xnor
  g924
  (
    n972,
    n510,
    n491,
    n928,
    n895
  );


  nand
  g925
  (
    n953,
    n506,
    n788,
    n524,
    n523
  );


  and
  g926
  (
    n950,
    n489,
    n486,
    n505,
    n904
  );


  xnor
  g927
  (
    n954,
    n911,
    n908,
    n515,
    n790
  );


  xor
  g928
  (
    n975,
    n518,
    n897,
    n773,
    n772
  );


  nand
  g929
  (
    n970,
    n926,
    n504,
    n919,
    n520
  );


  and
  g930
  (
    n986,
    n895,
    n777,
    n493,
    n931
  );


  or
  g931
  (
    n961,
    n930,
    n527,
    n913,
    n524
  );


  xnor
  g932
  (
    n942,
    n503,
    n926,
    n514,
    n778
  );


  and
  g933
  (
    n940,
    n516,
    n917,
    n920,
    n929
  );


  and
  g934
  (
    n936,
    n920,
    n531,
    n916,
    n491
  );


  nand
  g935
  (
    n951,
    n776,
    n786,
    n523
  );


  nor
  g936
  (
    n946,
    n921,
    n488,
    n525
  );


  and
  g937
  (
    n976,
    n783,
    n512,
    n894,
    n778
  );


  nor
  g938
  (
    n982,
    n495,
    n511,
    n521,
    n513
  );


  nor
  g939
  (
    KeyWire_0_23,
    n784,
    n910,
    n520,
    n519
  );


  xor
  g940
  (
    n947,
    n502,
    n519,
    n513,
    n495
  );


  and
  g941
  (
    n978,
    n528,
    n517,
    n507,
    n518
  );


  xor
  g942
  (
    n962,
    n499,
    n499,
    n494,
    n903
  );


  nor
  g943
  (
    n979,
    n506,
    n779,
    n531,
    n923
  );


  or
  g944
  (
    n983,
    n505,
    n902,
    n523,
    n772
  );


  or
  g945
  (
    n969,
    n925,
    n931,
    n501,
    n526
  );


  nor
  g946
  (
    n985,
    n779,
    n783,
    n929,
    n532
  );


  xor
  g947
  (
    n996,
    n930,
    n785,
    n901,
    n902
  );


  xor
  g948
  (
    n948,
    n915,
    n916,
    n930,
    n918
  );


  or
  g949
  (
    n989,
    n784,
    n905,
    n787,
    n781
  );


  and
  g950
  (
    KeyWire_0_50,
    n900,
    n932,
    n776,
    n787
  );


  or
  g951
  (
    n964,
    n774,
    n924,
    n490,
    n527
  );


  or
  g952
  (
    n994,
    n493,
    n520,
    n512,
    n927
  );


  nor
  g953
  (
    n973,
    n910,
    n922,
    n491,
    n516
  );


  or
  g954
  (
    n967,
    n508,
    n493,
    n486,
    n918
  );


  and
  g955
  (
    n971,
    n926,
    n494,
    n928,
    n922
  );


  or
  g956
  (
    n956,
    n530,
    n509,
    n524,
    n489
  );


  nand
  g957
  (
    n968,
    n525,
    n502,
    n915,
    n522
  );


  xnor
  g958
  (
    n933,
    n497,
    n788,
    n515,
    n773
  );


  nand
  g959
  (
    n938,
    n790,
    n924,
    n500,
    n921
  );


  and
  g960
  (
    n945,
    n497,
    n899,
    n528,
    n532
  );


  nor
  g961
  (
    n963,
    n931,
    n894,
    n917,
    n927
  );


  and
  g962
  (
    n966,
    n914,
    n518,
    n507,
    n909
  );


  and
  g963
  (
    n991,
    n781,
    n509,
    n499,
    n901
  );


  or
  g964
  (
    n958,
    n487,
    n487,
    n496,
    n898
  );


  nand
  g965
  (
    n941,
    n925,
    n922,
    n502,
    n789
  );


  xor
  g966
  (
    n944,
    n522,
    n896,
    n504,
    n515
  );


  nor
  g967
  (
    n993,
    n514,
    n522,
    n501,
    n519
  );


  nor
  g968
  (
    n1001,
    n958,
    n808,
    n977,
    n798
  );


  xor
  g969
  (
    n1020,
    n991,
    n986,
    n818,
    n972
  );


  and
  g970
  (
    n1017,
    n955,
    n808,
    n959,
    n935
  );


  xor
  g971
  (
    n1021,
    n957,
    n966,
    n814,
    n968
  );


  xnor
  g972
  (
    KeyWire_0_39,
    n794,
    n797,
    n796,
    n814
  );


  or
  g973
  (
    n1004,
    n953,
    n817,
    n940,
    n795
  );


  and
  g974
  (
    n1008,
    n799,
    n795,
    n811,
    n796
  );


  and
  g975
  (
    n1002,
    n792,
    n815,
    n818,
    n987
  );


  or
  g976
  (
    n1030,
    n800,
    n807,
    n819,
    n944
  );


  xnor
  g977
  (
    n1019,
    n943,
    n812,
    n952,
    n817
  );


  or
  g978
  (
    n1024,
    n996,
    n806,
    n976,
    n961
  );


  xor
  g979
  (
    n1032,
    n1000,
    n819,
    n992,
    n820
  );


  and
  g980
  (
    n1011,
    n933,
    n791,
    n816,
    n970
  );


  or
  g981
  (
    n1003,
    n979,
    n969,
    n975,
    n806
  );


  and
  g982
  (
    n1016,
    n960,
    n948,
    n815,
    n978
  );


  nand
  g983
  (
    n1023,
    n994,
    n988,
    n809,
    n813
  );


  xor
  g984
  (
    n1014,
    n956,
    n934,
    n983,
    n985
  );


  and
  g985
  (
    n1025,
    n981,
    n938,
    n945,
    n995
  );


  nand
  g986
  (
    n1007,
    n941,
    n816,
    n980,
    n802
  );


  or
  g987
  (
    n1029,
    n813,
    n947,
    n982,
    n792
  );


  and
  g988
  (
    n1027,
    n964,
    n974,
    n967,
    n807
  );


  and
  g989
  (
    n1015,
    n803,
    n793,
    n794
  );


  or
  g990
  (
    n1026,
    n800,
    n803,
    n950,
    n999
  );


  xor
  g991
  (
    n1009,
    n809,
    n939,
    n810,
    n984
  );


  xor
  g992
  (
    n1018,
    n954,
    n804,
    n942,
    n812
  );


  or
  g993
  (
    n1022,
    n998,
    n805,
    n971,
    n997
  );


  or
  g994
  (
    n1006,
    n965,
    n799,
    n949,
    n990
  );


  or
  g995
  (
    n1012,
    n937,
    n820,
    n804,
    n798
  );


  or
  g996
  (
    n1031,
    n802,
    n811,
    n801,
    n791
  );


  and
  g997
  (
    n1013,
    n797,
    n951,
    n989,
    n962
  );


  and
  g998
  (
    n1005,
    n993,
    n963,
    n801,
    n946
  );


  xnor
  g999
  (
    n1028,
    n805,
    n973,
    n810,
    n936
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n391,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n649,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n187,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n354,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n510,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n644,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n548,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n800,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n181,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n464,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n744,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n892,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n731,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n534,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n646,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n333,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n39,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n817,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n44,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n35,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n81,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n106,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n439,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n997,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n257,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n673,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n782,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n407,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n698,
    KeyNOTWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n845,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n50,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n172,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n265,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n376,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    KeyNOTWire_0_34,
    keyIn_0_34,
    KeyWire_0_34
  );


  not
  KeyNOTGate_0_34
  (
    n155,
    KeyNOTWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n670,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n934,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n472,
    KeyNOTWire_0_37
  );


  xnor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n440,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n1010,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n493,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n561,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n738,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n340,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n218,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n837,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n405,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n205,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n502,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n136,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n992,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n727,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n252,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    n410,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n995,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n271,
    KeyNOTWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n795,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n876,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n907,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n38,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n490,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n168,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n843,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n669,
    KeyNOTWire_0_63
  );


endmodule

