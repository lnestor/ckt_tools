

module Stat_3000_321
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2121,
  n2106,
  n2084,
  n2093,
  n2088,
  n2107,
  n2092,
  n2091,
  n2099,
  n2116,
  n2109,
  n2101,
  n2083,
  n2081,
  n2709,
  n2710,
  n2713,
  n2705,
  n2704,
  n2714,
  n2712,
  n2707,
  n2715,
  n2706,
  n2711,
  n2754,
  n2749,
  n3030,
  n3029,
  n3028,
  n3032,
  n3031
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n2121;output n2106;output n2084;output n2093;output n2088;output n2107;output n2092;output n2091;output n2099;output n2116;output n2109;output n2101;output n2083;output n2081;output n2709;output n2710;output n2713;output n2705;output n2704;output n2714;output n2712;output n2707;output n2715;output n2706;output n2711;output n2754;output n2749;output n3030;output n3029;output n3028;output n3032;output n3031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2082;wire n2085;wire n2086;wire n2087;wire n2089;wire n2090;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2100;wire n2102;wire n2103;wire n2104;wire n2105;wire n2108;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2117;wire n2118;wire n2119;wire n2120;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2708;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2750;wire n2751;wire n2752;wire n2753;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire n3010;wire n3011;wire n3012;wire n3013;wire n3014;wire n3015;wire n3016;wire n3017;wire n3018;wire n3019;wire n3020;wire n3021;wire n3022;wire n3023;wire n3024;wire n3025;wire n3026;wire n3027;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  buf
  g0
  (
    n58,
    n14
  );


  not
  g1
  (
    n55,
    n6
  );


  buf
  g2
  (
    n64,
    n18
  );


  not
  g3
  (
    n75,
    n25
  );


  buf
  g4
  (
    n59,
    n5
  );


  not
  g5
  (
    n68,
    n13
  );


  buf
  g6
  (
    n54,
    n9
  );


  not
  g7
  (
    n85,
    n16
  );


  buf
  g8
  (
    n110,
    n7
  );


  not
  g9
  (
    n79,
    n12
  );


  buf
  g10
  (
    n33,
    n21
  );


  buf
  g11
  (
    n116,
    n15
  );


  not
  g12
  (
    n52,
    n18
  );


  buf
  g13
  (
    n86,
    n1
  );


  not
  g14
  (
    n95,
    n22
  );


  buf
  g15
  (
    n60,
    n27
  );


  not
  g16
  (
    n129,
    n31
  );


  buf
  g17
  (
    n132,
    n2
  );


  buf
  g18
  (
    n121,
    n11
  );


  buf
  g19
  (
    n158,
    n10
  );


  buf
  g20
  (
    n35,
    n25
  );


  buf
  g21
  (
    n100,
    n11
  );


  buf
  g22
  (
    n126,
    n6
  );


  not
  g23
  (
    n71,
    n1
  );


  buf
  g24
  (
    n154,
    n20
  );


  not
  g25
  (
    n144,
    n4
  );


  not
  g26
  (
    n36,
    n3
  );


  buf
  g27
  (
    n50,
    n26
  );


  buf
  g28
  (
    n136,
    n18
  );


  buf
  g29
  (
    n115,
    n2
  );


  buf
  g30
  (
    n112,
    n19
  );


  buf
  g31
  (
    n76,
    n16
  );


  not
  g32
  (
    n145,
    n20
  );


  buf
  g33
  (
    n133,
    n12
  );


  buf
  g34
  (
    n149,
    n23
  );


  not
  g35
  (
    n135,
    n4
  );


  buf
  g36
  (
    n97,
    n15
  );


  buf
  g37
  (
    n34,
    n25
  );


  not
  g38
  (
    n93,
    n24
  );


  not
  g39
  (
    n140,
    n22
  );


  buf
  g40
  (
    n99,
    n14
  );


  not
  g41
  (
    n104,
    n1
  );


  not
  g42
  (
    n118,
    n26
  );


  buf
  g43
  (
    n57,
    n8
  );


  buf
  g44
  (
    n125,
    n21
  );


  not
  g45
  (
    n137,
    n15
  );


  buf
  g46
  (
    n160,
    n24
  );


  buf
  g47
  (
    n130,
    n8
  );


  buf
  g48
  (
    n88,
    n16
  );


  buf
  g49
  (
    n41,
    n15
  );


  not
  g50
  (
    n152,
    n19
  );


  not
  g51
  (
    n123,
    n10
  );


  buf
  g52
  (
    n142,
    n4
  );


  buf
  g53
  (
    n157,
    n12
  );


  buf
  g54
  (
    n107,
    n13
  );


  not
  g55
  (
    n138,
    n32
  );


  not
  g56
  (
    n156,
    n30
  );


  not
  g57
  (
    n141,
    n17
  );


  buf
  g58
  (
    n44,
    n8
  );


  buf
  g59
  (
    n70,
    n13
  );


  not
  g60
  (
    n83,
    n27
  );


  buf
  g61
  (
    n62,
    n28
  );


  buf
  g62
  (
    n113,
    n9
  );


  not
  g63
  (
    n150,
    n32
  );


  buf
  g64
  (
    n39,
    n16
  );


  not
  g65
  (
    n131,
    n7
  );


  buf
  g66
  (
    n127,
    n6
  );


  not
  g67
  (
    n81,
    n24
  );


  buf
  g68
  (
    n146,
    n6
  );


  buf
  g69
  (
    n98,
    n5
  );


  buf
  g70
  (
    n147,
    n25
  );


  not
  g71
  (
    n91,
    n17
  );


  not
  g72
  (
    n90,
    n30
  );


  not
  g73
  (
    n74,
    n18
  );


  buf
  g74
  (
    n61,
    n29
  );


  buf
  g75
  (
    KeyWire_0_5,
    n23
  );


  not
  g76
  (
    n42,
    n22
  );


  not
  g77
  (
    n72,
    n28
  );


  not
  g78
  (
    n49,
    n11
  );


  not
  g79
  (
    n92,
    n29
  );


  buf
  g80
  (
    n69,
    n4
  );


  not
  g81
  (
    n46,
    n30
  );


  buf
  g82
  (
    n96,
    n19
  );


  buf
  g83
  (
    n124,
    n12
  );


  buf
  g84
  (
    n120,
    n3
  );


  buf
  g85
  (
    n43,
    n29
  );


  buf
  g86
  (
    n159,
    n24
  );


  not
  g87
  (
    n122,
    n31
  );


  not
  g88
  (
    n111,
    n5
  );


  not
  g89
  (
    n51,
    n9
  );


  buf
  g90
  (
    n134,
    n9
  );


  buf
  g91
  (
    n47,
    n7
  );


  buf
  g92
  (
    n87,
    n19
  );


  not
  g93
  (
    n38,
    n8
  );


  not
  g94
  (
    n109,
    n32
  );


  not
  g95
  (
    n155,
    n14
  );


  not
  g96
  (
    n77,
    n28
  );


  buf
  g97
  (
    n80,
    n30
  );


  not
  g98
  (
    n139,
    n21
  );


  not
  g99
  (
    n65,
    n20
  );


  not
  g100
  (
    n73,
    n21
  );


  not
  g101
  (
    n78,
    n2
  );


  buf
  g102
  (
    n102,
    n32
  );


  buf
  g103
  (
    n48,
    n10
  );


  buf
  g104
  (
    n148,
    n17
  );


  buf
  g105
  (
    n56,
    n5
  );


  not
  g106
  (
    n82,
    n10
  );


  not
  g107
  (
    n119,
    n14
  );


  not
  g108
  (
    n143,
    n20
  );


  buf
  g109
  (
    n37,
    n23
  );


  not
  g110
  (
    n101,
    n2
  );


  buf
  g111
  (
    n128,
    n29
  );


  not
  g112
  (
    n66,
    n31
  );


  not
  g113
  (
    n108,
    n31
  );


  buf
  g114
  (
    n53,
    n13
  );


  not
  g115
  (
    n89,
    n22
  );


  not
  g116
  (
    n103,
    n7
  );


  not
  g117
  (
    n67,
    n23
  );


  buf
  g118
  (
    n40,
    n3
  );


  buf
  g119
  (
    n63,
    n28
  );


  buf
  g120
  (
    n114,
    n1
  );


  buf
  g121
  (
    n117,
    n3
  );


  buf
  g122
  (
    n153,
    n11
  );


  not
  g123
  (
    n45,
    n27
  );


  not
  g124
  (
    n106,
    n26
  );


  buf
  g125
  (
    n94,
    n17
  );


  buf
  g126
  (
    n151,
    n26
  );


  not
  g127
  (
    n84,
    n27
  );


  buf
  g128
  (
    n251,
    n103
  );


  buf
  g129
  (
    n439,
    n127
  );


  not
  g130
  (
    n248,
    n38
  );


  buf
  g131
  (
    n459,
    n140
  );


  not
  g132
  (
    n493,
    n39
  );


  buf
  g133
  (
    n175,
    n110
  );


  not
  g134
  (
    n256,
    n134
  );


  buf
  g135
  (
    n216,
    n65
  );


  not
  g136
  (
    n243,
    n85
  );


  not
  g137
  (
    n408,
    n61
  );


  not
  g138
  (
    n524,
    n108
  );


  not
  g139
  (
    n537,
    n50
  );


  buf
  g140
  (
    n491,
    n104
  );


  not
  g141
  (
    n205,
    n151
  );


  not
  g142
  (
    n601,
    n106
  );


  buf
  g143
  (
    n183,
    n108
  );


  buf
  g144
  (
    n286,
    n145
  );


  not
  g145
  (
    n220,
    n50
  );


  buf
  g146
  (
    n283,
    n72
  );


  not
  g147
  (
    n237,
    n50
  );


  not
  g148
  (
    n435,
    n110
  );


  buf
  g149
  (
    n277,
    n130
  );


  not
  g150
  (
    n377,
    n123
  );


  not
  g151
  (
    n416,
    n156
  );


  buf
  g152
  (
    n249,
    n108
  );


  buf
  g153
  (
    n461,
    n48
  );


  not
  g154
  (
    n521,
    n69
  );


  buf
  g155
  (
    n638,
    n158
  );


  buf
  g156
  (
    n653,
    n153
  );


  not
  g157
  (
    n492,
    n91
  );


  buf
  g158
  (
    n647,
    n41
  );


  not
  g159
  (
    n621,
    n131
  );


  buf
  g160
  (
    n213,
    n132
  );


  not
  g161
  (
    n543,
    n142
  );


  buf
  g162
  (
    n557,
    n105
  );


  buf
  g163
  (
    n629,
    n84
  );


  buf
  g164
  (
    n460,
    n79
  );


  not
  g165
  (
    n566,
    n154
  );


  buf
  g166
  (
    n184,
    n84
  );


  buf
  g167
  (
    n645,
    n85
  );


  not
  g168
  (
    n354,
    n45
  );


  not
  g169
  (
    n480,
    n97
  );


  buf
  g170
  (
    n507,
    n99
  );


  not
  g171
  (
    n185,
    n72
  );


  buf
  g172
  (
    n455,
    n155
  );


  not
  g173
  (
    n196,
    n48
  );


  not
  g174
  (
    n208,
    n116
  );


  not
  g175
  (
    n431,
    n143
  );


  buf
  g176
  (
    n533,
    n104
  );


  buf
  g177
  (
    n371,
    n123
  );


  not
  g178
  (
    n167,
    n91
  );


  buf
  g179
  (
    n226,
    n121
  );


  not
  g180
  (
    n475,
    n78
  );


  buf
  g181
  (
    n336,
    n138
  );


  not
  g182
  (
    n280,
    n82
  );


  not
  g183
  (
    n578,
    n74
  );


  buf
  g184
  (
    n378,
    n49
  );


  buf
  g185
  (
    n463,
    n64
  );


  not
  g186
  (
    n197,
    n66
  );


  buf
  g187
  (
    n209,
    n98
  );


  not
  g188
  (
    n514,
    n144
  );


  not
  g189
  (
    n267,
    n116
  );


  buf
  g190
  (
    n652,
    n70
  );


  not
  g191
  (
    n258,
    n100
  );


  not
  g192
  (
    n562,
    n139
  );


  buf
  g193
  (
    n485,
    n46
  );


  not
  g194
  (
    n328,
    n74
  );


  not
  g195
  (
    n487,
    n148
  );


  not
  g196
  (
    n335,
    n76
  );


  buf
  g197
  (
    n546,
    n139
  );


  not
  g198
  (
    n319,
    n108
  );


  not
  g199
  (
    n164,
    n35
  );


  buf
  g200
  (
    n229,
    n130
  );


  not
  g201
  (
    n607,
    n120
  );


  not
  g202
  (
    n173,
    n145
  );


  not
  g203
  (
    n632,
    n89
  );


  not
  g204
  (
    n482,
    n41
  );


  buf
  g205
  (
    n238,
    n102
  );


  not
  g206
  (
    n574,
    n142
  );


  buf
  g207
  (
    n577,
    n73
  );


  buf
  g208
  (
    n585,
    n128
  );


  buf
  g209
  (
    n279,
    n92
  );


  buf
  g210
  (
    KeyWire_0_12,
    n46
  );


  not
  g211
  (
    n409,
    n61
  );


  not
  g212
  (
    n307,
    n127
  );


  buf
  g213
  (
    n413,
    n142
  );


  buf
  g214
  (
    n497,
    n75
  );


  buf
  g215
  (
    n594,
    n125
  );


  buf
  g216
  (
    n490,
    n114
  );


  not
  g217
  (
    n344,
    n43
  );


  not
  g218
  (
    n270,
    n111
  );


  not
  g219
  (
    n468,
    n150
  );


  buf
  g220
  (
    n644,
    n150
  );


  not
  g221
  (
    n244,
    n131
  );


  buf
  g222
  (
    n452,
    n132
  );


  buf
  g223
  (
    n355,
    n59
  );


  buf
  g224
  (
    n275,
    n74
  );


  not
  g225
  (
    n473,
    n148
  );


  not
  g226
  (
    n253,
    n84
  );


  not
  g227
  (
    n457,
    n57
  );


  buf
  g228
  (
    n387,
    n106
  );


  buf
  g229
  (
    n373,
    n100
  );


  buf
  g230
  (
    n260,
    n89
  );


  buf
  g231
  (
    n611,
    n141
  );


  not
  g232
  (
    n414,
    n113
  );


  buf
  g233
  (
    n215,
    n44
  );


  not
  g234
  (
    n222,
    n82
  );


  not
  g235
  (
    n450,
    n68
  );


  not
  g236
  (
    n659,
    n88
  );


  buf
  g237
  (
    n360,
    n36
  );


  not
  g238
  (
    n615,
    n99
  );


  not
  g239
  (
    n194,
    n62
  );


  not
  g240
  (
    n412,
    n35
  );


  buf
  g241
  (
    n227,
    n112
  );


  not
  g242
  (
    n564,
    n63
  );


  not
  g243
  (
    n470,
    n67
  );


  not
  g244
  (
    n458,
    n123
  );


  buf
  g245
  (
    n626,
    n34
  );


  not
  g246
  (
    n247,
    n134
  );


  not
  g247
  (
    n516,
    n55
  );


  buf
  g248
  (
    n329,
    n35
  );


  not
  g249
  (
    n366,
    n95
  );


  buf
  g250
  (
    n231,
    n93
  );


  buf
  g251
  (
    n365,
    n99
  );


  not
  g252
  (
    n558,
    n115
  );


  not
  g253
  (
    n643,
    n58
  );


  not
  g254
  (
    n177,
    n42
  );


  buf
  g255
  (
    n271,
    n39
  );


  not
  g256
  (
    KeyWire_0_1,
    n40
  );


  buf
  g257
  (
    n515,
    n147
  );


  buf
  g258
  (
    n437,
    n72
  );


  not
  g259
  (
    n424,
    n117
  );


  not
  g260
  (
    n363,
    n46
  );


  buf
  g261
  (
    n265,
    n49
  );


  not
  g262
  (
    n320,
    n151
  );


  buf
  g263
  (
    n269,
    n144
  );


  not
  g264
  (
    n372,
    n48
  );


  not
  g265
  (
    n657,
    n119
  );


  buf
  g266
  (
    n297,
    n56
  );


  not
  g267
  (
    n565,
    n81
  );


  buf
  g268
  (
    n405,
    n145
  );


  not
  g269
  (
    n655,
    n102
  );


  not
  g270
  (
    n534,
    n113
  );


  not
  g271
  (
    n625,
    n52
  );


  not
  g272
  (
    n614,
    n116
  );


  buf
  g273
  (
    n567,
    n53
  );


  buf
  g274
  (
    n547,
    n110
  );


  not
  g275
  (
    n342,
    n112
  );


  not
  g276
  (
    n636,
    n113
  );


  not
  g277
  (
    n464,
    n101
  );


  not
  g278
  (
    n593,
    n55
  );


  not
  g279
  (
    n230,
    n68
  );


  not
  g280
  (
    n207,
    n141
  );


  not
  g281
  (
    n592,
    n103
  );


  not
  g282
  (
    n358,
    n107
  );


  buf
  g283
  (
    n392,
    n118
  );


  not
  g284
  (
    n648,
    n95
  );


  buf
  g285
  (
    n660,
    n71
  );


  not
  g286
  (
    n390,
    n152
  );


  not
  g287
  (
    n428,
    n86
  );


  not
  g288
  (
    n300,
    n71
  );


  not
  g289
  (
    n393,
    n54
  );


  not
  g290
  (
    n356,
    n61
  );


  buf
  g291
  (
    n471,
    n158
  );


  not
  g292
  (
    n600,
    n137
  );


  buf
  g293
  (
    n606,
    n49
  );


  buf
  g294
  (
    n406,
    n54
  );


  not
  g295
  (
    n523,
    n129
  );


  buf
  g296
  (
    n654,
    n146
  );


  buf
  g297
  (
    n536,
    n107
  );


  not
  g298
  (
    n576,
    n51
  );


  not
  g299
  (
    n500,
    n149
  );


  buf
  g300
  (
    n224,
    n149
  );


  buf
  g301
  (
    n206,
    n79
  );


  buf
  g302
  (
    n287,
    n143
  );


  not
  g303
  (
    n189,
    n152
  );


  buf
  g304
  (
    n379,
    n41
  );


  not
  g305
  (
    n642,
    n119
  );


  buf
  g306
  (
    n338,
    n80
  );


  not
  g307
  (
    n649,
    n123
  );


  not
  g308
  (
    n272,
    n85
  );


  not
  g309
  (
    n282,
    n60
  );


  not
  g310
  (
    n199,
    n107
  );


  buf
  g311
  (
    n318,
    n90
  );


  not
  g312
  (
    n404,
    n64
  );


  not
  g313
  (
    n651,
    n86
  );


  not
  g314
  (
    n326,
    n44
  );


  not
  g315
  (
    n628,
    n125
  );


  buf
  g316
  (
    n563,
    n144
  );


  not
  g317
  (
    n496,
    n130
  );


  not
  g318
  (
    n637,
    n55
  );


  buf
  g319
  (
    n560,
    n125
  );


  not
  g320
  (
    n165,
    n65
  );


  not
  g321
  (
    n257,
    n76
  );


  buf
  g322
  (
    n433,
    n33
  );


  buf
  g323
  (
    n436,
    n34
  );


  buf
  g324
  (
    n420,
    n91
  );


  not
  g325
  (
    n223,
    n62
  );


  buf
  g326
  (
    n448,
    n81
  );


  buf
  g327
  (
    n417,
    n112
  );


  buf
  g328
  (
    n346,
    n124
  );


  not
  g329
  (
    n617,
    n62
  );


  not
  g330
  (
    n597,
    n88
  );


  not
  g331
  (
    n332,
    n124
  );


  buf
  g332
  (
    n411,
    n105
  );


  buf
  g333
  (
    n242,
    n63
  );


  buf
  g334
  (
    n246,
    n69
  );


  not
  g335
  (
    n402,
    n133
  );


  buf
  g336
  (
    n664,
    n42
  );


  buf
  g337
  (
    n398,
    n134
  );


  buf
  g338
  (
    n559,
    n37
  );


  buf
  g339
  (
    n488,
    n107
  );


  not
  g340
  (
    n353,
    n109
  );


  not
  g341
  (
    n364,
    n88
  );


  not
  g342
  (
    n303,
    n127
  );


  buf
  g343
  (
    n174,
    n45
  );


  buf
  g344
  (
    n449,
    n117
  );


  not
  g345
  (
    n650,
    n97
  );


  not
  g346
  (
    n631,
    n56
  );


  buf
  g347
  (
    n445,
    n105
  );


  buf
  g348
  (
    n661,
    n82
  );


  buf
  g349
  (
    n550,
    n67
  );


  buf
  g350
  (
    n212,
    n44
  );


  buf
  g351
  (
    n423,
    n117
  );


  not
  g352
  (
    n292,
    n87
  );


  buf
  g353
  (
    n598,
    n72
  );


  not
  g354
  (
    n376,
    n133
  );


  buf
  g355
  (
    n484,
    n146
  );


  buf
  g356
  (
    n389,
    n128
  );


  buf
  g357
  (
    n234,
    n151
  );


  buf
  g358
  (
    n603,
    n59
  );


  not
  g359
  (
    n453,
    n57
  );


  buf
  g360
  (
    n434,
    n141
  );


  buf
  g361
  (
    n314,
    n93
  );


  buf
  g362
  (
    n370,
    n132
  );


  buf
  g363
  (
    n587,
    n129
  );


  not
  g364
  (
    n368,
    n98
  );


  buf
  g365
  (
    n568,
    n53
  );


  not
  g366
  (
    n232,
    n144
  );


  not
  g367
  (
    n278,
    n69
  );


  buf
  g368
  (
    n362,
    n100
  );


  not
  g369
  (
    n465,
    n54
  );


  not
  g370
  (
    n306,
    n36
  );


  not
  g371
  (
    n214,
    n66
  );


  not
  g372
  (
    n217,
    n46
  );


  not
  g373
  (
    n211,
    n38
  );


  buf
  g374
  (
    n361,
    n74
  );


  buf
  g375
  (
    n489,
    n79
  );


  not
  g376
  (
    n410,
    n111
  );


  buf
  g377
  (
    n202,
    n76
  );


  not
  g378
  (
    n438,
    n77
  );


  not
  g379
  (
    n178,
    n52
  );


  not
  g380
  (
    n323,
    n120
  );


  buf
  g381
  (
    n443,
    n153
  );


  not
  g382
  (
    n384,
    n115
  );


  buf
  g383
  (
    n513,
    n44
  );


  buf
  g384
  (
    n570,
    n68
  );


  buf
  g385
  (
    n252,
    n146
  );


  not
  g386
  (
    n508,
    n100
  );


  not
  g387
  (
    n401,
    n52
  );


  not
  g388
  (
    n193,
    n109
  );


  buf
  g389
  (
    n343,
    n89
  );


  buf
  g390
  (
    n274,
    n99
  );


  buf
  g391
  (
    n289,
    n94
  );


  buf
  g392
  (
    n198,
    n67
  );


  buf
  g393
  (
    n381,
    n43
  );


  buf
  g394
  (
    n203,
    n70
  );


  not
  g395
  (
    n495,
    n40
  );


  buf
  g396
  (
    n419,
    n39
  );


  buf
  g397
  (
    n191,
    n114
  );


  buf
  g398
  (
    n351,
    n36
  );


  not
  g399
  (
    n308,
    n86
  );


  buf
  g400
  (
    n309,
    n135
  );


  not
  g401
  (
    n575,
    n60
  );


  not
  g402
  (
    n315,
    n149
  );


  not
  g403
  (
    n172,
    n114
  );


  buf
  g404
  (
    n472,
    n152
  );


  buf
  g405
  (
    n474,
    n121
  );


  not
  g406
  (
    n456,
    n92
  );


  not
  g407
  (
    n168,
    n45
  );


  buf
  g408
  (
    n656,
    n122
  );


  not
  g409
  (
    n608,
    n70
  );


  buf
  g410
  (
    n561,
    n150
  );


  buf
  g411
  (
    n188,
    n38
  );


  buf
  g412
  (
    n469,
    n156
  );


  buf
  g413
  (
    n569,
    n71
  );


  not
  g414
  (
    n181,
    n42
  );


  buf
  g415
  (
    n486,
    n62
  );


  buf
  g416
  (
    KeyWire_0_8,
    n148
  );


  not
  g417
  (
    n334,
    n154
  );


  not
  g418
  (
    n333,
    n122
  );


  buf
  g419
  (
    n293,
    n120
  );


  buf
  g420
  (
    n294,
    n157
  );


  buf
  g421
  (
    n432,
    n94
  );


  buf
  g422
  (
    n499,
    n78
  );


  buf
  g423
  (
    n602,
    n136
  );


  buf
  g424
  (
    n582,
    n111
  );


  not
  g425
  (
    n646,
    n70
  );


  buf
  g426
  (
    n618,
    n88
  );


  not
  g427
  (
    n446,
    n65
  );


  not
  g428
  (
    n298,
    n55
  );


  not
  g429
  (
    n310,
    n90
  );


  buf
  g430
  (
    n324,
    n124
  );


  not
  g431
  (
    n240,
    n78
  );


  buf
  g432
  (
    n662,
    n119
  );


  not
  g433
  (
    n261,
    n92
  );


  not
  g434
  (
    n161,
    n47
  );


  not
  g435
  (
    n476,
    n38
  );


  buf
  g436
  (
    n520,
    n90
  );


  not
  g437
  (
    n532,
    n36
  );


  buf
  g438
  (
    n612,
    n131
  );


  buf
  g439
  (
    n375,
    n63
  );


  buf
  g440
  (
    n162,
    n138
  );


  not
  g441
  (
    n540,
    n126
  );


  buf
  g442
  (
    n504,
    n43
  );


  buf
  g443
  (
    n425,
    n140
  );


  buf
  g444
  (
    n284,
    n96
  );


  buf
  g445
  (
    n589,
    n135
  );


  buf
  g446
  (
    n407,
    n125
  );


  buf
  g447
  (
    n583,
    n139
  );


  not
  g448
  (
    n531,
    n105
  );


  buf
  g449
  (
    n388,
    n89
  );


  not
  g450
  (
    n259,
    n80
  );


  buf
  g451
  (
    n290,
    n45
  );


  buf
  g452
  (
    n322,
    n90
  );


  buf
  g453
  (
    n221,
    n158
  );


  buf
  g454
  (
    n610,
    n138
  );


  buf
  g455
  (
    n352,
    n136
  );


  not
  g456
  (
    n421,
    n41
  );


  buf
  g457
  (
    n201,
    n51
  );


  buf
  g458
  (
    n192,
    n40
  );


  buf
  g459
  (
    n517,
    n102
  );


  not
  g460
  (
    n288,
    n83
  );


  not
  g461
  (
    n228,
    n117
  );


  buf
  g462
  (
    n399,
    n34
  );


  buf
  g463
  (
    n317,
    n87
  );


  not
  g464
  (
    n316,
    n86
  );


  buf
  g465
  (
    n444,
    n59
  );


  buf
  g466
  (
    n605,
    n136
  );


  buf
  g467
  (
    n325,
    n47
  );


  buf
  g468
  (
    n299,
    n80
  );


  buf
  g469
  (
    n302,
    n146
  );


  buf
  g470
  (
    n529,
    n133
  );


  not
  g471
  (
    n553,
    n155
  );


  buf
  g472
  (
    n179,
    n135
  );


  not
  g473
  (
    n180,
    n94
  );


  buf
  g474
  (
    n170,
    n142
  );


  not
  g475
  (
    n327,
    n104
  );


  not
  g476
  (
    n541,
    n119
  );


  not
  g477
  (
    n619,
    n126
  );


  not
  g478
  (
    n281,
    n52
  );


  buf
  g479
  (
    n639,
    n96
  );


  buf
  g480
  (
    n386,
    n143
  );


  not
  g481
  (
    n586,
    n118
  );


  buf
  g482
  (
    n255,
    n128
  );


  buf
  g483
  (
    n385,
    n153
  );


  not
  g484
  (
    n163,
    n147
  );


  not
  g485
  (
    n451,
    n75
  );


  not
  g486
  (
    n341,
    n134
  );


  not
  g487
  (
    n658,
    n121
  );


  not
  g488
  (
    n512,
    n140
  );


  buf
  g489
  (
    n518,
    n77
  );


  buf
  g490
  (
    n219,
    n154
  );


  not
  g491
  (
    n528,
    n106
  );


  buf
  g492
  (
    n519,
    n114
  );


  not
  g493
  (
    n494,
    n57
  );


  buf
  g494
  (
    n573,
    n60
  );


  not
  g495
  (
    n526,
    n96
  );


  buf
  g496
  (
    n525,
    n56
  );


  buf
  g497
  (
    n542,
    n33
  );


  not
  g498
  (
    n285,
    n106
  );


  not
  g499
  (
    n171,
    n118
  );


  buf
  g500
  (
    n266,
    n113
  );


  not
  g501
  (
    n331,
    n101
  );


  not
  g502
  (
    n581,
    n104
  );


  buf
  g503
  (
    n596,
    n122
  );


  buf
  g504
  (
    n441,
    n98
  );


  buf
  g505
  (
    n166,
    n121
  );


  buf
  g506
  (
    n295,
    n95
  );


  not
  g507
  (
    n218,
    n73
  );


  buf
  g508
  (
    n511,
    n51
  );


  not
  g509
  (
    n454,
    n157
  );


  not
  g510
  (
    n572,
    n79
  );


  buf
  g511
  (
    n502,
    n84
  );


  not
  g512
  (
    n627,
    n75
  );


  not
  g513
  (
    n383,
    n87
  );


  buf
  g514
  (
    n640,
    n129
  );


  buf
  g515
  (
    n613,
    n67
  );


  not
  g516
  (
    n225,
    n54
  );


  not
  g517
  (
    n241,
    n137
  );


  not
  g518
  (
    n584,
    n50
  );


  buf
  g519
  (
    n305,
    n33
  );


  buf
  g520
  (
    n169,
    n68
  );


  buf
  g521
  (
    n239,
    n58
  );


  not
  g522
  (
    n478,
    n60
  );


  not
  g523
  (
    n429,
    n103
  );


  not
  g524
  (
    n620,
    n102
  );


  not
  g525
  (
    n609,
    n140
  );


  buf
  g526
  (
    n467,
    n103
  );


  not
  g527
  (
    n622,
    n58
  );


  not
  g528
  (
    n254,
    n157
  );


  not
  g529
  (
    n591,
    n37
  );


  not
  g530
  (
    n397,
    n92
  );


  buf
  g531
  (
    n250,
    n98
  );


  buf
  g532
  (
    n348,
    n111
  );


  not
  g533
  (
    n588,
    n122
  );


  not
  g534
  (
    n479,
    n116
  );


  buf
  g535
  (
    n347,
    n153
  );


  not
  g536
  (
    n527,
    n63
  );


  not
  g537
  (
    n330,
    n132
  );


  buf
  g538
  (
    n590,
    n97
  );


  buf
  g539
  (
    n466,
    n101
  );


  buf
  g540
  (
    n580,
    n58
  );


  buf
  g541
  (
    n291,
    n97
  );


  buf
  g542
  (
    n522,
    n131
  );


  not
  g543
  (
    n235,
    n82
  );


  not
  g544
  (
    n633,
    n81
  );


  buf
  g545
  (
    n195,
    n137
  );


  buf
  g546
  (
    n395,
    n37
  );


  not
  g547
  (
    n311,
    n126
  );


  not
  g548
  (
    n634,
    n115
  );


  not
  g549
  (
    n663,
    n33
  );


  not
  g550
  (
    n503,
    n95
  );


  not
  g551
  (
    n604,
    n83
  );


  not
  g552
  (
    n262,
    n96
  );


  not
  g553
  (
    n263,
    n73
  );


  not
  g554
  (
    n276,
    n147
  );


  not
  g555
  (
    n340,
    n156
  );


  not
  g556
  (
    n369,
    n56
  );


  buf
  g557
  (
    n304,
    n93
  );


  not
  g558
  (
    n396,
    n48
  );


  buf
  g559
  (
    n483,
    n149
  );


  not
  g560
  (
    n264,
    n81
  );


  not
  g561
  (
    n204,
    n37
  );


  buf
  g562
  (
    n176,
    n109
  );


  not
  g563
  (
    n312,
    n66
  );


  not
  g564
  (
    n374,
    n135
  );


  not
  g565
  (
    n641,
    n35
  );


  buf
  g566
  (
    n481,
    n42
  );


  buf
  g567
  (
    n391,
    n109
  );


  buf
  g568
  (
    n539,
    n78
  );


  not
  g569
  (
    n555,
    n83
  );


  buf
  g570
  (
    n415,
    n150
  );


  not
  g571
  (
    n418,
    n75
  );


  buf
  g572
  (
    n296,
    n124
  );


  buf
  g573
  (
    n359,
    n83
  );


  not
  g574
  (
    n623,
    n133
  );


  buf
  g575
  (
    n616,
    n76
  );


  buf
  g576
  (
    n571,
    n77
  );


  not
  g577
  (
    n556,
    n154
  );


  not
  g578
  (
    n535,
    n112
  );


  not
  g579
  (
    n579,
    n64
  );


  not
  g580
  (
    n538,
    n69
  );


  buf
  g581
  (
    n422,
    n59
  );


  buf
  g582
  (
    n426,
    n65
  );


  not
  g583
  (
    n440,
    n129
  );


  buf
  g584
  (
    n545,
    n147
  );


  buf
  g585
  (
    n554,
    n115
  );


  buf
  g586
  (
    n544,
    n49
  );


  buf
  g587
  (
    n442,
    n110
  );


  not
  g588
  (
    n599,
    n43
  );


  not
  g589
  (
    n394,
    n39
  );


  not
  g590
  (
    n505,
    n128
  );


  buf
  g591
  (
    n548,
    n91
  );


  not
  g592
  (
    n350,
    n152
  );


  buf
  g593
  (
    n549,
    n47
  );


  buf
  g594
  (
    n268,
    n127
  );


  not
  g595
  (
    n301,
    n145
  );


  not
  g596
  (
    n382,
    n141
  );


  not
  g597
  (
    n635,
    n120
  );


  not
  g598
  (
    n551,
    n51
  );


  buf
  g599
  (
    n339,
    n118
  );


  not
  g600
  (
    n233,
    n53
  );


  buf
  g601
  (
    n403,
    n143
  );


  not
  g602
  (
    n349,
    n148
  );


  buf
  g603
  (
    n321,
    n155
  );


  buf
  g604
  (
    n530,
    n34
  );


  buf
  g605
  (
    n313,
    n126
  );


  buf
  g606
  (
    n357,
    n156
  );


  buf
  g607
  (
    n345,
    n101
  );


  buf
  g608
  (
    n501,
    n71
  );


  buf
  g609
  (
    n337,
    n77
  );


  not
  g610
  (
    n498,
    n53
  );


  not
  g611
  (
    n186,
    n73
  );


  not
  g612
  (
    n509,
    n47
  );


  not
  g613
  (
    n182,
    n94
  );


  not
  g614
  (
    KeyWire_0_7,
    n61
  );


  not
  g615
  (
    n624,
    n80
  );


  not
  g616
  (
    n477,
    n136
  );


  buf
  g617
  (
    n427,
    n158
  );


  not
  g618
  (
    n462,
    n66
  );


  buf
  g619
  (
    n430,
    n57
  );


  buf
  g620
  (
    n273,
    n40
  );


  buf
  g621
  (
    n245,
    n157
  );


  buf
  g622
  (
    n187,
    n85
  );


  buf
  g623
  (
    n552,
    n130
  );


  not
  g624
  (
    n595,
    n151
  );


  buf
  g625
  (
    n630,
    n93
  );


  not
  g626
  (
    n210,
    n139
  );


  buf
  g627
  (
    n400,
    n137
  );


  not
  g628
  (
    n506,
    n155
  );


  not
  g629
  (
    n447,
    n87
  );


  not
  g630
  (
    n367,
    n64
  );


  not
  g631
  (
    n236,
    n138
  );


  buf
  g632
  (
    n734,
    n243
  );


  buf
  g633
  (
    n717,
    n311
  );


  buf
  g634
  (
    n1074,
    n310
  );


  buf
  g635
  (
    n942,
    n538
  );


  not
  g636
  (
    n1087,
    n606
  );


  not
  g637
  (
    n1656,
    n231
  );


  not
  g638
  (
    n1834,
    n636
  );


  not
  g639
  (
    n1850,
    n652
  );


  not
  g640
  (
    n1530,
    n354
  );


  not
  g641
  (
    n887,
    n544
  );


  buf
  g642
  (
    n893,
    n474
  );


  not
  g643
  (
    n715,
    n508
  );


  not
  g644
  (
    n692,
    n169
  );


  buf
  g645
  (
    n1624,
    n617
  );


  buf
  g646
  (
    n1822,
    n457
  );


  not
  g647
  (
    n1302,
    n324
  );


  buf
  g648
  (
    n1386,
    n496
  );


  not
  g649
  (
    n1028,
    n608
  );


  buf
  g650
  (
    n1538,
    n580
  );


  buf
  g651
  (
    n1715,
    n313
  );


  not
  g652
  (
    n733,
    n167
  );


  not
  g653
  (
    n1470,
    n592
  );


  buf
  g654
  (
    n991,
    n542
  );


  not
  g655
  (
    n1472,
    n406
  );


  not
  g656
  (
    n995,
    n408
  );


  buf
  g657
  (
    n1291,
    n578
  );


  not
  g658
  (
    n1736,
    n624
  );


  not
  g659
  (
    n1553,
    n364
  );


  buf
  g660
  (
    n879,
    n413
  );


  buf
  g661
  (
    n1458,
    n206
  );


  buf
  g662
  (
    n1285,
    n373
  );


  not
  g663
  (
    n1403,
    n357
  );


  not
  g664
  (
    n1245,
    n179
  );


  not
  g665
  (
    n752,
    n547
  );


  not
  g666
  (
    n726,
    n619
  );


  not
  g667
  (
    n1443,
    n637
  );


  buf
  g668
  (
    n1801,
    n335
  );


  not
  g669
  (
    n874,
    n440
  );


  not
  g670
  (
    n1617,
    n175
  );


  not
  g671
  (
    n754,
    n649
  );


  not
  g672
  (
    n1208,
    n525
  );


  buf
  g673
  (
    n1852,
    n607
  );


  not
  g674
  (
    n957,
    n420
  );


  buf
  g675
  (
    n1788,
    n260
  );


  buf
  g676
  (
    n974,
    n553
  );


  not
  g677
  (
    n687,
    n222
  );


  not
  g678
  (
    n1740,
    n221
  );


  buf
  g679
  (
    n1427,
    n179
  );


  not
  g680
  (
    n825,
    n255
  );


  not
  g681
  (
    n978,
    n639
  );


  not
  g682
  (
    n1312,
    n251
  );


  not
  g683
  (
    n1535,
    n387
  );


  not
  g684
  (
    n1151,
    n571
  );


  buf
  g685
  (
    n1071,
    n493
  );


  not
  g686
  (
    n1693,
    n379
  );


  not
  g687
  (
    n1336,
    n333
  );


  buf
  g688
  (
    KeyWire_0_10,
    n165
  );


  not
  g689
  (
    n667,
    n230
  );


  not
  g690
  (
    n1186,
    n391
  );


  not
  g691
  (
    n1197,
    n202
  );


  not
  g692
  (
    n1388,
    n474
  );


  not
  g693
  (
    n1545,
    n443
  );


  not
  g694
  (
    n1728,
    n611
  );


  not
  g695
  (
    n965,
    n247
  );


  buf
  g696
  (
    n1340,
    n327
  );


  buf
  g697
  (
    n776,
    n273
  );


  not
  g698
  (
    n1253,
    n471
  );


  buf
  g699
  (
    n1582,
    n229
  );


  not
  g700
  (
    n761,
    n591
  );


  not
  g701
  (
    n1397,
    n535
  );


  buf
  g702
  (
    n712,
    n185
  );


  not
  g703
  (
    n1366,
    n654
  );


  not
  g704
  (
    n1325,
    n205
  );


  buf
  g705
  (
    n1131,
    n337
  );


  buf
  g706
  (
    n1556,
    n444
  );


  buf
  g707
  (
    n1601,
    n619
  );


  buf
  g708
  (
    n1464,
    n332
  );


  not
  g709
  (
    n1865,
    n207
  );


  not
  g710
  (
    n1434,
    n573
  );


  not
  g711
  (
    n1425,
    n262
  );


  not
  g712
  (
    n1328,
    n166
  );


  not
  g713
  (
    n1305,
    n336
  );


  not
  g714
  (
    n952,
    n162
  );


  not
  g715
  (
    n820,
    n604
  );


  buf
  g716
  (
    n1461,
    n181
  );


  buf
  g717
  (
    n1271,
    n373
  );


  buf
  g718
  (
    n1407,
    n464
  );


  not
  g719
  (
    n1255,
    n333
  );


  not
  g720
  (
    n759,
    n420
  );


  not
  g721
  (
    n1089,
    n410
  );


  buf
  g722
  (
    n1679,
    n603
  );


  buf
  g723
  (
    n972,
    n276
  );


  buf
  g724
  (
    n767,
    n295
  );


  not
  g725
  (
    n1172,
    n215
  );


  buf
  g726
  (
    n1207,
    n437
  );


  not
  g727
  (
    n1573,
    n445
  );


  buf
  g728
  (
    n1560,
    n473
  );


  buf
  g729
  (
    n773,
    n637
  );


  not
  g730
  (
    n1554,
    n458
  );


  buf
  g731
  (
    n852,
    n212
  );


  buf
  g732
  (
    n1571,
    n526
  );


  not
  g733
  (
    n827,
    n298
  );


  not
  g734
  (
    n1252,
    n429
  );


  buf
  g735
  (
    n1404,
    n557
  );


  buf
  g736
  (
    n1733,
    n522
  );


  not
  g737
  (
    n807,
    n271
  );


  not
  g738
  (
    n1048,
    n525
  );


  buf
  g739
  (
    n1501,
    n331
  );


  buf
  g740
  (
    n1024,
    n388
  );


  not
  g741
  (
    n1615,
    n584
  );


  buf
  g742
  (
    n675,
    n575
  );


  not
  g743
  (
    n815,
    n421
  );


  buf
  g744
  (
    n836,
    n528
  );


  not
  g745
  (
    n1797,
    n185
  );


  not
  g746
  (
    n1045,
    n360
  );


  buf
  g747
  (
    KeyWire_0_11,
    n180
  );


  buf
  g748
  (
    n1260,
    n171
  );


  not
  g749
  (
    n1754,
    n330
  );


  buf
  g750
  (
    n1382,
    n649
  );


  buf
  g751
  (
    n1787,
    n338
  );


  not
  g752
  (
    n1775,
    n189
  );


  not
  g753
  (
    n1198,
    n342
  );


  not
  g754
  (
    n1647,
    n451
  );


  not
  g755
  (
    n1332,
    n393
  );


  not
  g756
  (
    n876,
    n604
  );


  not
  g757
  (
    n732,
    n247
  );


  buf
  g758
  (
    n1796,
    n471
  );


  buf
  g759
  (
    n762,
    n293
  );


  not
  g760
  (
    n904,
    n536
  );


  buf
  g761
  (
    n912,
    n251
  );


  not
  g762
  (
    n889,
    n378
  );


  not
  g763
  (
    n1568,
    n224
  );


  not
  g764
  (
    n832,
    n532
  );


  buf
  g765
  (
    n1264,
    n481
  );


  not
  g766
  (
    n1581,
    n564
  );


  not
  g767
  (
    n951,
    n256
  );


  buf
  g768
  (
    n1256,
    n546
  );


  not
  g769
  (
    n1484,
    n503
  );


  buf
  g770
  (
    n826,
    n611
  );


  not
  g771
  (
    n1625,
    n621
  );


  buf
  g772
  (
    n672,
    n468
  );


  buf
  g773
  (
    n1149,
    n198
  );


  not
  g774
  (
    n1135,
    n390
  );


  not
  g775
  (
    n1194,
    n516
  );


  not
  g776
  (
    n1579,
    n386
  );


  not
  g777
  (
    n1043,
    n503
  );


  buf
  g778
  (
    n981,
    n268
  );


  buf
  g779
  (
    n1537,
    n395
  );


  buf
  g780
  (
    n741,
    n454
  );


  buf
  g781
  (
    n1534,
    n377
  );


  buf
  g782
  (
    n1130,
    n629
  );


  buf
  g783
  (
    n1278,
    n562
  );


  buf
  g784
  (
    n1844,
    n241
  );


  buf
  g785
  (
    n1126,
    n462
  );


  not
  g786
  (
    n897,
    n442
  );


  not
  g787
  (
    n1379,
    n222
  );


  not
  g788
  (
    n1666,
    n441
  );


  buf
  g789
  (
    n1631,
    n634
  );


  not
  g790
  (
    n794,
    n321
  );


  buf
  g791
  (
    n1743,
    n464
  );


  not
  g792
  (
    n1313,
    n602
  );


  not
  g793
  (
    n1677,
    n187
  );


  buf
  g794
  (
    n1712,
    n382
  );


  not
  g795
  (
    n786,
    n588
  );


  not
  g796
  (
    n1858,
    n402
  );


  buf
  g797
  (
    n731,
    n614
  );


  not
  g798
  (
    n756,
    n635
  );


  not
  g799
  (
    n1008,
    n408
  );


  buf
  g800
  (
    n757,
    n354
  );


  buf
  g801
  (
    n1494,
    n200
  );


  buf
  g802
  (
    n923,
    n444
  );


  not
  g803
  (
    n1828,
    n286
  );


  buf
  g804
  (
    n1117,
    n422
  );


  not
  g805
  (
    n903,
    n235
  );


  not
  g806
  (
    n682,
    n454
  );


  not
  g807
  (
    n1523,
    n227
  );


  not
  g808
  (
    n1184,
    n472
  );


  buf
  g809
  (
    n1497,
    n599
  );


  not
  g810
  (
    n1299,
    n388
  );


  not
  g811
  (
    n783,
    n632
  );


  buf
  g812
  (
    n683,
    n624
  );


  not
  g813
  (
    n1350,
    n271
  );


  buf
  g814
  (
    n1761,
    n503
  );


  not
  g815
  (
    n746,
    n570
  );


  not
  g816
  (
    n1006,
    n510
  );


  buf
  g817
  (
    n1481,
    n534
  );


  buf
  g818
  (
    n1767,
    n261
  );


  buf
  g819
  (
    n1279,
    n556
  );


  buf
  g820
  (
    n1516,
    n315
  );


  buf
  g821
  (
    n1393,
    n433
  );


  buf
  g822
  (
    n1794,
    n415
  );


  buf
  g823
  (
    n1069,
    n418
  );


  buf
  g824
  (
    n1244,
    n331
  );


  buf
  g825
  (
    n907,
    n529
  );


  not
  g826
  (
    n1499,
    n191
  );


  buf
  g827
  (
    n1540,
    n250
  );


  buf
  g828
  (
    n1163,
    n249
  );


  not
  g829
  (
    n830,
    n256
  );


  buf
  g830
  (
    n1511,
    n295
  );


  buf
  g831
  (
    n968,
    n199
  );


  buf
  g832
  (
    n1696,
    n280
  );


  not
  g833
  (
    n1300,
    n298
  );


  not
  g834
  (
    n1463,
    n224
  );


  buf
  g835
  (
    n1093,
    n653
  );


  buf
  g836
  (
    n1584,
    n596
  );


  not
  g837
  (
    n1334,
    n436
  );


  buf
  g838
  (
    n1210,
    n430
  );


  not
  g839
  (
    n1588,
    n568
  );


  not
  g840
  (
    n1751,
    n317
  );


  not
  g841
  (
    n1552,
    n359
  );


  buf
  g842
  (
    n1124,
    n268
  );


  buf
  g843
  (
    n1395,
    n593
  );


  not
  g844
  (
    n701,
    n628
  );


  not
  g845
  (
    n1506,
    n531
  );


  not
  g846
  (
    n1112,
    n286
  );


  not
  g847
  (
    n1837,
    n533
  );


  buf
  g848
  (
    n841,
    n639
  );


  buf
  g849
  (
    n774,
    n645
  );


  buf
  g850
  (
    n1756,
    n337
  );


  buf
  g851
  (
    n950,
    n555
  );


  not
  g852
  (
    n1842,
    n302
  );


  buf
  g853
  (
    n750,
    n201
  );


  not
  g854
  (
    n1092,
    n285
  );


  not
  g855
  (
    n1373,
    n372
  );


  buf
  g856
  (
    n778,
    n568
  );


  buf
  g857
  (
    n899,
    n325
  );


  not
  g858
  (
    n1031,
    n426
  );


  not
  g859
  (
    n1578,
    n600
  );


  not
  g860
  (
    n865,
    n205
  );


  not
  g861
  (
    n697,
    n202
  );


  not
  g862
  (
    n670,
    n451
  );


  not
  g863
  (
    n816,
    n242
  );


  not
  g864
  (
    n1555,
    n564
  );


  not
  g865
  (
    n1103,
    n285
  );


  not
  g866
  (
    n798,
    n339
  );


  not
  g867
  (
    n1166,
    n367
  );


  not
  g868
  (
    n1070,
    n268
  );


  buf
  g869
  (
    n1349,
    n639
  );


  not
  g870
  (
    n1303,
    n222
  );


  buf
  g871
  (
    n673,
    n616
  );


  not
  g872
  (
    n686,
    n527
  );


  not
  g873
  (
    n1058,
    n580
  );


  buf
  g874
  (
    n1222,
    n197
  );


  buf
  g875
  (
    n1680,
    n560
  );


  not
  g876
  (
    n1780,
    n395
  );


  buf
  g877
  (
    n1372,
    n372
  );


  not
  g878
  (
    n735,
    n339
  );


  not
  g879
  (
    n1577,
    n577
  );


  buf
  g880
  (
    n1655,
    n190
  );


  not
  g881
  (
    n1121,
    n647
  );


  not
  g882
  (
    n1747,
    n359
  );


  buf
  g883
  (
    n1218,
    n541
  );


  buf
  g884
  (
    n1468,
    n163
  );


  not
  g885
  (
    n785,
    n365
  );


  not
  g886
  (
    n846,
    n162
  );


  not
  g887
  (
    n1485,
    n487
  );


  not
  g888
  (
    n1737,
    n439
  );


  buf
  g889
  (
    n1778,
    n296
  );


  not
  g890
  (
    n743,
    n240
  );


  not
  g891
  (
    n1167,
    n412
  );


  not
  g892
  (
    n1115,
    n166
  );


  not
  g893
  (
    n1384,
    n264
  );


  not
  g894
  (
    n1640,
    n488
  );


  not
  g895
  (
    n1620,
    n299
  );


  not
  g896
  (
    n1802,
    n227
  );


  buf
  g897
  (
    n1800,
    n426
  );


  buf
  g898
  (
    n1100,
    n466
  );


  not
  g899
  (
    n1380,
    n241
  );


  not
  g900
  (
    n890,
    n193
  );


  buf
  g901
  (
    n881,
    n329
  );


  buf
  g902
  (
    n1091,
    n200
  );


  not
  g903
  (
    n1745,
    n552
  );


  not
  g904
  (
    n1290,
    n493
  );


  buf
  g905
  (
    n1385,
    n583
  );


  buf
  g906
  (
    n997,
    n254
  );


  not
  g907
  (
    n1663,
    n258
  );


  not
  g908
  (
    n986,
    n447
  );


  not
  g909
  (
    n1645,
    n220
  );


  not
  g910
  (
    n884,
    n256
  );


  buf
  g911
  (
    n1205,
    n586
  );


  buf
  g912
  (
    n1433,
    n525
  );


  buf
  g913
  (
    n1575,
    n561
  );


  not
  g914
  (
    n848,
    n418
  );


  buf
  g915
  (
    n745,
    n272
  );


  not
  g916
  (
    n822,
    n206
  );


  buf
  g917
  (
    n1414,
    n504
  );


  buf
  g918
  (
    n850,
    n537
  );


  buf
  g919
  (
    n1360,
    n475
  );


  buf
  g920
  (
    n961,
    n526
  );


  buf
  g921
  (
    n1862,
    n462
  );


  not
  g922
  (
    n1227,
    n574
  );


  not
  g923
  (
    n791,
    n276
  );


  buf
  g924
  (
    n1232,
    n530
  );


  not
  g925
  (
    n674,
    n274
  );


  not
  g926
  (
    n722,
    n575
  );


  not
  g927
  (
    n1042,
    n258
  );


  not
  g928
  (
    n1758,
    n557
  );


  not
  g929
  (
    n1243,
    n561
  );


  not
  g930
  (
    n1280,
    n437
  );


  buf
  g931
  (
    n1032,
    n245
  );


  not
  g932
  (
    n1014,
    n618
  );


  not
  g933
  (
    n1532,
    n464
  );


  buf
  g934
  (
    n1790,
    n576
  );


  not
  g935
  (
    n924,
    n225
  );


  not
  g936
  (
    n1719,
    n180
  );


  not
  g937
  (
    n1002,
    n404
  );


  buf
  g938
  (
    KeyWire_0_15,
    n218
  );


  buf
  g939
  (
    n1399,
    n516
  );


  buf
  g940
  (
    n1864,
    n228
  );


  not
  g941
  (
    n1049,
    n393
  );


  not
  g942
  (
    n1847,
    n523
  );


  buf
  g943
  (
    n931,
    n574
  );


  buf
  g944
  (
    n999,
    n465
  );


  not
  g945
  (
    n1426,
    n602
  );


  not
  g946
  (
    n1576,
    n329
  );


  buf
  g947
  (
    n1216,
    n293
  );


  buf
  g948
  (
    n1835,
    n330
  );


  not
  g949
  (
    n1085,
    n386
  );


  not
  g950
  (
    n1519,
    n465
  );


  not
  g951
  (
    n1439,
    n520
  );


  buf
  g952
  (
    n1611,
    n304
  );


  not
  g953
  (
    n703,
    n226
  );


  not
  g954
  (
    n956,
    n233
  );


  buf
  g955
  (
    n925,
    n435
  );


  not
  g956
  (
    n1122,
    n553
  );


  not
  g957
  (
    n1750,
    n357
  );


  buf
  g958
  (
    n1202,
    n634
  );


  buf
  g959
  (
    n1355,
    n299
  );


  not
  g960
  (
    n1410,
    n304
  );


  not
  g961
  (
    n1354,
    n651
  );


  buf
  g962
  (
    n806,
    n300
  );


  not
  g963
  (
    n679,
    n343
  );


  not
  g964
  (
    n1717,
    n277
  );


  not
  g965
  (
    n1396,
    n416
  );


  buf
  g966
  (
    n1642,
    n457
  );


  not
  g967
  (
    n1479,
    n165
  );


  buf
  g968
  (
    n1812,
    n653
  );


  buf
  g969
  (
    n724,
    n165
  );


  buf
  g970
  (
    n869,
    n609
  );


  buf
  g971
  (
    n892,
    n302
  );


  buf
  g972
  (
    n1466,
    n561
  );


  buf
  g973
  (
    n811,
    n269
  );


  buf
  g974
  (
    n813,
    n301
  );


  buf
  g975
  (
    n1176,
    n462
  );


  buf
  g976
  (
    n1709,
    n278
  );


  buf
  g977
  (
    n760,
    n282
  );


  not
  g978
  (
    n1816,
    n173
  );


  buf
  g979
  (
    n1318,
    n528
  );


  not
  g980
  (
    n1213,
    n450
  );


  buf
  g981
  (
    n1016,
    n476
  );


  not
  g982
  (
    n1254,
    n628
  );


  buf
  g983
  (
    n1586,
    n196
  );


  not
  g984
  (
    n1589,
    n199
  );


  not
  g985
  (
    n1192,
    n338
  );


  buf
  g986
  (
    n1664,
    n266
  );


  buf
  g987
  (
    n1001,
    n443
  );


  buf
  g988
  (
    n849,
    n451
  );


  not
  g989
  (
    n1561,
    n377
  );


  not
  g990
  (
    n1017,
    n442
  );


  buf
  g991
  (
    n1729,
    n653
  );


  buf
  g992
  (
    n1572,
    n595
  );


  not
  g993
  (
    n720,
    n367
  );


  not
  g994
  (
    n1627,
    n258
  );


  not
  g995
  (
    n983,
    n581
  );


  buf
  g996
  (
    n1452,
    n420
  );


  buf
  g997
  (
    n839,
    n620
  );


  not
  g998
  (
    n1162,
    n438
  );


  buf
  g999
  (
    n1595,
    n632
  );


  buf
  g1000
  (
    n1261,
    n233
  );


  buf
  g1001
  (
    n1798,
    n448
  );


  buf
  g1002
  (
    n740,
    n474
  );


  not
  g1003
  (
    n1766,
    n599
  );


  not
  g1004
  (
    n862,
    n624
  );


  not
  g1005
  (
    n1480,
    n528
  );


  buf
  g1006
  (
    n1843,
    n240
  );


  not
  g1007
  (
    n902,
    n477
  );


  buf
  g1008
  (
    n1310,
    n590
  );


  buf
  g1009
  (
    n769,
    n352
  );


  not
  g1010
  (
    n1212,
    n172
  );


  not
  g1011
  (
    n1409,
    n550
  );


  not
  g1012
  (
    n1609,
    n300
  );


  buf
  g1013
  (
    n1214,
    n332
  );


  buf
  g1014
  (
    n955,
    n440
  );


  buf
  g1015
  (
    n1308,
    n351
  );


  not
  g1016
  (
    n1619,
    n507
  );


  buf
  g1017
  (
    n1814,
    n582
  );


  not
  g1018
  (
    n1341,
    n450
  );


  not
  g1019
  (
    n1453,
    n603
  );


  buf
  g1020
  (
    n1339,
    n381
  );


  not
  g1021
  (
    n963,
    n648
  );


  buf
  g1022
  (
    n962,
    n442
  );


  buf
  g1023
  (
    n1653,
    n221
  );


  not
  g1024
  (
    n1451,
    n243
  );


  not
  g1025
  (
    n1171,
    n325
  );


  buf
  g1026
  (
    n1287,
    n567
  );


  buf
  g1027
  (
    n1518,
    n252
  );


  buf
  g1028
  (
    n1174,
    n420
  );


  buf
  g1029
  (
    n1752,
    n320
  );


  buf
  g1030
  (
    n1598,
    n170
  );


  buf
  g1031
  (
    n926,
    n504
  );


  buf
  g1032
  (
    n1825,
    n309
  );


  not
  g1033
  (
    n855,
    n257
  );


  not
  g1034
  (
    n840,
    n213
  );


  not
  g1035
  (
    n1551,
    n423
  );


  not
  g1036
  (
    n1226,
    n409
  );


  buf
  g1037
  (
    n1265,
    n340
  );


  not
  g1038
  (
    n1759,
    n412
  );


  buf
  g1039
  (
    n1514,
    n405
  );


  buf
  g1040
  (
    n1053,
    n572
  );


  buf
  g1041
  (
    n1533,
    n427
  );


  not
  g1042
  (
    n1228,
    n537
  );


  not
  g1043
  (
    n964,
    n320
  );


  buf
  g1044
  (
    n1169,
    n284
  );


  not
  g1045
  (
    n1829,
    n311
  );


  buf
  g1046
  (
    n937,
    n551
  );


  buf
  g1047
  (
    n1527,
    n322
  );


  not
  g1048
  (
    n1830,
    n534
  );


  buf
  g1049
  (
    n797,
    n406
  );


  buf
  g1050
  (
    n1134,
    n335
  );


  buf
  g1051
  (
    n1723,
    n502
  );


  not
  g1052
  (
    n1512,
    n162
  );


  buf
  g1053
  (
    n975,
    n437
  );


  not
  g1054
  (
    n960,
    n320
  );


  buf
  g1055
  (
    n1605,
    n366
  );


  not
  g1056
  (
    n1565,
    n430
  );


  not
  g1057
  (
    n1587,
    n221
  );


  buf
  g1058
  (
    n875,
    n217
  );


  buf
  g1059
  (
    n843,
    n304
  );


  buf
  g1060
  (
    n977,
    n369
  );


  buf
  g1061
  (
    n969,
    n479
  );


  buf
  g1062
  (
    n1809,
    n625
  );


  buf
  g1063
  (
    n725,
    n632
  );


  buf
  g1064
  (
    n1805,
    n489
  );


  buf
  g1065
  (
    n1522,
    n413
  );


  not
  g1066
  (
    n1495,
    n357
  );


  buf
  g1067
  (
    n1082,
    n341
  );


  buf
  g1068
  (
    n1724,
    n339
  );


  buf
  g1069
  (
    n666,
    n239
  );


  not
  g1070
  (
    n1607,
    n436
  );


  buf
  g1071
  (
    n1636,
    n204
  );


  not
  g1072
  (
    n1604,
    n448
  );


  buf
  g1073
  (
    n1118,
    n498
  );


  buf
  g1074
  (
    n1764,
    n206
  );


  buf
  g1075
  (
    n707,
    n246
  );


  not
  g1076
  (
    n1866,
    n288
  );


  not
  g1077
  (
    n1297,
    n360
  );


  not
  g1078
  (
    n1155,
    n216
  );


  buf
  g1079
  (
    n1060,
    n497
  );


  buf
  g1080
  (
    n1274,
    n591
  );


  buf
  g1081
  (
    n1020,
    n429
  );


  not
  g1082
  (
    n787,
    n611
  );


  not
  g1083
  (
    n919,
    n524
  );


  not
  g1084
  (
    n1282,
    n522
  );


  buf
  g1085
  (
    n1068,
    n397
  );


  not
  g1086
  (
    n1023,
    n225
  );


  buf
  g1087
  (
    n1133,
    n586
  );


  buf
  g1088
  (
    n1187,
    n569
  );


  buf
  g1089
  (
    n1346,
    n623
  );


  buf
  g1090
  (
    n1301,
    n360
  );


  not
  g1091
  (
    n915,
    n348
  );


  buf
  g1092
  (
    n1786,
    n478
  );


  buf
  g1093
  (
    n1784,
    n161
  );


  not
  g1094
  (
    n1036,
    n330
  );


  not
  g1095
  (
    n910,
    n515
  );


  not
  g1096
  (
    n1030,
    n400
  );


  not
  g1097
  (
    n1566,
    n642
  );


  not
  g1098
  (
    n1544,
    n267
  );


  not
  g1099
  (
    n859,
    n497
  );


  buf
  g1100
  (
    n1281,
    n369
  );


  buf
  g1101
  (
    n788,
    n260
  );


  not
  g1102
  (
    n771,
    n253
  );


  buf
  g1103
  (
    n1503,
    n549
  );


  not
  g1104
  (
    n976,
    n645
  );


  buf
  g1105
  (
    n1026,
    n169
  );


  buf
  g1106
  (
    n810,
    n161
  );


  buf
  g1107
  (
    n1543,
    n453
  );


  not
  g1108
  (
    n1189,
    n287
  );


  buf
  g1109
  (
    n1513,
    n546
  );


  not
  g1110
  (
    n1277,
    n178
  );


  not
  g1111
  (
    n1455,
    n551
  );


  not
  g1112
  (
    n1034,
    n205
  );


  buf
  g1113
  (
    n1447,
    n610
  );


  buf
  g1114
  (
    n1056,
    n268
  );


  not
  g1115
  (
    n958,
    n392
  );


  not
  g1116
  (
    n1580,
    n344
  );


  not
  g1117
  (
    n1086,
    n582
  );


  not
  g1118
  (
    n980,
    n469
  );


  not
  g1119
  (
    n1137,
    n517
  );


  not
  g1120
  (
    n1773,
    n558
  );


  buf
  g1121
  (
    n684,
    n278
  );


  buf
  g1122
  (
    n1259,
    n270
  );


  buf
  g1123
  (
    n1483,
    n513
  );


  buf
  g1124
  (
    n706,
    n243
  );


  not
  g1125
  (
    n1700,
    n412
  );


  buf
  g1126
  (
    n1487,
    n443
  );


  buf
  g1127
  (
    n1361,
    n469
  );


  not
  g1128
  (
    n1153,
    n480
  );


  buf
  g1129
  (
    n1033,
    n207
  );


  not
  g1130
  (
    n1055,
    n350
  );


  not
  g1131
  (
    n1105,
    n633
  );


  not
  g1132
  (
    n1690,
    n521
  );


  buf
  g1133
  (
    n863,
    n411
  );


  buf
  g1134
  (
    n765,
    n338
  );


  not
  g1135
  (
    n700,
    n167
  );


  buf
  g1136
  (
    n1613,
    n650
  );


  buf
  g1137
  (
    n1567,
    n308
  );


  not
  g1138
  (
    n954,
    n270
  );


  not
  g1139
  (
    n1708,
    n188
  );


  buf
  g1140
  (
    n1757,
    n345
  );


  not
  g1141
  (
    n1658,
    n254
  );


  buf
  g1142
  (
    n934,
    n650
  );


  not
  g1143
  (
    n1368,
    n316
  );


  buf
  g1144
  (
    n990,
    n500
  );


  buf
  g1145
  (
    n1141,
    n262
  );


  buf
  g1146
  (
    n1622,
    n592
  );


  buf
  g1147
  (
    n1389,
    n592
  );


  buf
  g1148
  (
    n1027,
    n584
  );


  not
  g1149
  (
    n1375,
    n568
  );


  not
  g1150
  (
    n883,
    n587
  );


  buf
  g1151
  (
    n1818,
    n424
  );


  buf
  g1152
  (
    n766,
    n215
  );


  buf
  g1153
  (
    n1789,
    n565
  );


  not
  g1154
  (
    n1722,
    n432
  );


  buf
  g1155
  (
    n1691,
    n394
  );


  buf
  g1156
  (
    n970,
    n305
  );


  not
  g1157
  (
    n1639,
    n211
  );


  not
  g1158
  (
    n1116,
    n372
  );


  buf
  g1159
  (
    n709,
    n283
  );


  buf
  g1160
  (
    n1687,
    n589
  );


  not
  g1161
  (
    n1734,
    n544
  );


  not
  g1162
  (
    n940,
    n456
  );


  buf
  g1163
  (
    n1569,
    n370
  );


  buf
  g1164
  (
    n819,
    n534
  );


  not
  g1165
  (
    n1777,
    n164
  );


  buf
  g1166
  (
    n1128,
    n576
  );


  buf
  g1167
  (
    n1306,
    n520
  );


  not
  g1168
  (
    n719,
    n404
  );


  not
  g1169
  (
    n1046,
    n643
  );


  buf
  g1170
  (
    n1857,
    n518
  );


  buf
  g1171
  (
    n671,
    n489
  );


  not
  g1172
  (
    n861,
    n242
  );


  not
  g1173
  (
    n1840,
    n411
  );


  not
  g1174
  (
    n1462,
    n512
  );


  not
  g1175
  (
    n1436,
    n642
  );


  buf
  g1176
  (
    n1596,
    n169
  );


  buf
  g1177
  (
    n1526,
    n261
  );


  not
  g1178
  (
    n1183,
    n410
  );


  not
  g1179
  (
    n1348,
    n342
  );


  not
  g1180
  (
    KeyWire_0_2,
    n491
  );


  buf
  g1181
  (
    n1698,
    n191
  );


  buf
  g1182
  (
    n1353,
    n509
  );


  not
  g1183
  (
    n1154,
    n503
  );


  not
  g1184
  (
    n1637,
    n485
  );


  buf
  g1185
  (
    n1145,
    n167
  );


  not
  g1186
  (
    n1839,
    n577
  );


  not
  g1187
  (
    n1242,
    n606
  );


  buf
  g1188
  (
    n1635,
    n449
  );


  buf
  g1189
  (
    n779,
    n523
  );


  not
  g1190
  (
    n1249,
    n449
  );


  not
  g1191
  (
    n920,
    n589
  );


  not
  g1192
  (
    n1614,
    n549
  );


  not
  g1193
  (
    n1633,
    n445
  );


  buf
  g1194
  (
    n665,
    n216
  );


  not
  g1195
  (
    n784,
    n417
  );


  buf
  g1196
  (
    n1422,
    n397
  );


  buf
  g1197
  (
    n1109,
    n622
  );


  buf
  g1198
  (
    n1748,
    n611
  );


  buf
  g1199
  (
    n871,
    n264
  );


  buf
  g1200
  (
    n1623,
    n228
  );


  buf
  g1201
  (
    n694,
    n529
  );


  not
  g1202
  (
    n1224,
    n385
  );


  buf
  g1203
  (
    n1168,
    n607
  );


  not
  g1204
  (
    n1536,
    n355
  );


  buf
  g1205
  (
    n748,
    n225
  );


  not
  g1206
  (
    n1490,
    n482
  );


  not
  g1207
  (
    n699,
    n249
  );


  not
  g1208
  (
    n1165,
    n569
  );


  not
  g1209
  (
    n1358,
    n612
  );


  buf
  g1210
  (
    n1482,
    n626
  );


  not
  g1211
  (
    n930,
    n394
  );


  not
  g1212
  (
    n1474,
    n492
  );


  buf
  g1213
  (
    n1321,
    n498
  );


  buf
  g1214
  (
    n872,
    n524
  );


  not
  g1215
  (
    n1402,
    n281
  );


  not
  g1216
  (
    n1446,
    n427
  );


  buf
  g1217
  (
    n1492,
    n406
  );


  not
  g1218
  (
    n1782,
    n189
  );


  buf
  g1219
  (
    n1159,
    n316
  );


  buf
  g1220
  (
    n831,
    n328
  );


  buf
  g1221
  (
    n1442,
    n326
  );


  buf
  g1222
  (
    n1196,
    n355
  );


  buf
  g1223
  (
    n1559,
    n417
  );


  not
  g1224
  (
    n677,
    n274
  );


  buf
  g1225
  (
    n1599,
    n495
  );


  not
  g1226
  (
    n1003,
    n651
  );


  buf
  g1227
  (
    n1469,
    n425
  );


  buf
  g1228
  (
    n1689,
    n222
  );


  buf
  g1229
  (
    n906,
    n407
  );


  buf
  g1230
  (
    n1201,
    n466
  );


  not
  g1231
  (
    n1018,
    n314
  );


  not
  g1232
  (
    n1846,
    n560
  );


  not
  g1233
  (
    n781,
    n358
  );


  buf
  g1234
  (
    n1072,
    n601
  );


  buf
  g1235
  (
    n1667,
    n570
  );


  buf
  g1236
  (
    n1090,
    n334
  );


  buf
  g1237
  (
    n1147,
    n183
  );


  buf
  g1238
  (
    n1792,
    n612
  );


  buf
  g1239
  (
    n1190,
    n643
  );


  buf
  g1240
  (
    n1275,
    n506
  );


  buf
  g1241
  (
    n1294,
    n627
  );


  not
  g1242
  (
    n808,
    n334
  );


  buf
  g1243
  (
    n1225,
    n508
  );


  buf
  g1244
  (
    n1525,
    n494
  );


  buf
  g1245
  (
    n1721,
    n493
  );


  buf
  g1246
  (
    n1419,
    n599
  );


  buf
  g1247
  (
    n932,
    n325
  );


  not
  g1248
  (
    n1127,
    n646
  );


  buf
  g1249
  (
    n1477,
    n482
  );


  not
  g1250
  (
    n1838,
    n169
  );


  buf
  g1251
  (
    n790,
    n317
  );


  not
  g1252
  (
    n1638,
    n187
  );


  not
  g1253
  (
    n1570,
    n600
  );


  buf
  g1254
  (
    n1673,
    n376
  );


  not
  g1255
  (
    n1239,
    n638
  );


  buf
  g1256
  (
    n1316,
    n553
  );


  not
  g1257
  (
    n1517,
    n458
  );


  buf
  g1258
  (
    n1738,
    n530
  );


  not
  g1259
  (
    n993,
    n460
  );


  buf
  g1260
  (
    n1597,
    n190
  );


  not
  g1261
  (
    n864,
    n459
  );


  buf
  g1262
  (
    n695,
    n523
  );


  buf
  g1263
  (
    n1819,
    n285
  );


  not
  g1264
  (
    n1420,
    n227
  );


  buf
  g1265
  (
    n918,
    n251
  );


  not
  g1266
  (
    n775,
    n389
  );


  not
  g1267
  (
    n1320,
    n399
  );


  not
  g1268
  (
    n1111,
    n291
  );


  buf
  g1269
  (
    n891,
    n542
  );


  not
  g1270
  (
    n1803,
    n414
  );


  not
  g1271
  (
    n1558,
    n511
  );


  buf
  g1272
  (
    n1125,
    n585
  );


  not
  g1273
  (
    n1094,
    n231
  );


  buf
  g1274
  (
    n1753,
    n249
  );


  buf
  g1275
  (
    n1370,
    n230
  );


  not
  g1276
  (
    n845,
    n384
  );


  not
  g1277
  (
    n1000,
    n613
  );


  not
  g1278
  (
    n1441,
    n341
  );


  not
  g1279
  (
    n1714,
    n312
  );


  not
  g1280
  (
    n1185,
    n435
  );


  not
  g1281
  (
    n1013,
    n323
  );


  buf
  g1282
  (
    n1528,
    n501
  );


  not
  g1283
  (
    n959,
    n342
  );


  not
  g1284
  (
    n1749,
    n566
  );


  not
  g1285
  (
    n1025,
    n453
  );


  buf
  g1286
  (
    n1705,
    n387
  );


  buf
  g1287
  (
    n1272,
    n621
  );


  buf
  g1288
  (
    n796,
    n252
  );


  buf
  g1289
  (
    n768,
    n324
  );


  buf
  g1290
  (
    n1779,
    n254
  );


  buf
  g1291
  (
    n1374,
    n194
  );


  buf
  g1292
  (
    n1289,
    n647
  );


  buf
  g1293
  (
    n838,
    n239
  );


  not
  g1294
  (
    n1266,
    n516
  );


  buf
  g1295
  (
    n1457,
    n487
  );


  buf
  g1296
  (
    n1686,
    n581
  );


  not
  g1297
  (
    n966,
    n237
  );


  not
  g1298
  (
    n1697,
    n310
  );


  buf
  g1299
  (
    n888,
    n585
  );


  buf
  g1300
  (
    n1548,
    n510
  );


  buf
  g1301
  (
    n1132,
    n481
  );


  not
  g1302
  (
    n1010,
    n227
  );


  buf
  g1303
  (
    n1233,
    n275
  );


  buf
  g1304
  (
    n1634,
    n388
  );


  not
  g1305
  (
    n1195,
    n383
  );


  not
  g1306
  (
    n823,
    n192
  );


  not
  g1307
  (
    n1701,
    n293
  );


  buf
  g1308
  (
    n728,
    n648
  );


  not
  g1309
  (
    n1012,
    n210
  );


  buf
  g1310
  (
    n1539,
    n472
  );


  buf
  g1311
  (
    n973,
    n419
  );


  buf
  g1312
  (
    n789,
    n416
  );


  not
  g1313
  (
    n1238,
    n438
  );


  not
  g1314
  (
    n1342,
    n588
  );


  buf
  g1315
  (
    n1344,
    n535
  );


  not
  g1316
  (
    n929,
    n344
  );


  buf
  g1317
  (
    n947,
    n347
  );


  buf
  g1318
  (
    n994,
    n377
  );


  buf
  g1319
  (
    n758,
    n585
  );


  buf
  g1320
  (
    n867,
    n518
  );


  buf
  g1321
  (
    n1220,
    n455
  );


  not
  g1322
  (
    n1813,
    n201
  );


  buf
  g1323
  (
    n837,
    n439
  );


  buf
  g1324
  (
    n1524,
    n402
  );


  buf
  g1325
  (
    n1508,
    n640
  );


  not
  g1326
  (
    n1448,
    n429
  );


  buf
  g1327
  (
    n1630,
    n501
  );


  buf
  g1328
  (
    n805,
    n234
  );


  buf
  g1329
  (
    n943,
    n248
  );


  not
  g1330
  (
    n835,
    n486
  );


  not
  g1331
  (
    n1073,
    n164
  );


  buf
  g1332
  (
    n1098,
    n499
  );


  buf
  g1333
  (
    n1345,
    n353
  );


  not
  g1334
  (
    n1454,
    n476
  );


  buf
  g1335
  (
    n1083,
    n409
  );


  not
  g1336
  (
    n1707,
    n626
  );


  buf
  g1337
  (
    n1610,
    n223
  );


  not
  g1338
  (
    n693,
    n299
  );


  buf
  g1339
  (
    n1182,
    n264
  );


  not
  g1340
  (
    n1199,
    n468
  );


  not
  g1341
  (
    n928,
    n501
  );


  not
  g1342
  (
    n1730,
    n511
  );


  not
  g1343
  (
    n1178,
    n515
  );


  buf
  g1344
  (
    n1270,
    n237
  );


  not
  g1345
  (
    n669,
    n592
  );


  buf
  g1346
  (
    n1641,
    n549
  );


  buf
  g1347
  (
    n744,
    n537
  );


  buf
  g1348
  (
    n1815,
    n248
  );


  buf
  g1349
  (
    n917,
    n323
  );


  buf
  g1350
  (
    n1237,
    n447
  );


  buf
  g1351
  (
    n1080,
    n188
  );


  not
  g1352
  (
    n1104,
    n433
  );


  not
  g1353
  (
    n1646,
    n403
  );


  buf
  g1354
  (
    n1651,
    n476
  );


  not
  g1355
  (
    n1699,
    n467
  );


  not
  g1356
  (
    n1337,
    n533
  );


  not
  g1357
  (
    n1273,
    n321
  );


  not
  g1358
  (
    n1095,
    n375
  );


  buf
  g1359
  (
    n1381,
    n575
  );


  not
  g1360
  (
    n1826,
    n466
  );


  not
  g1361
  (
    n885,
    n393
  );


  buf
  g1362
  (
    n1283,
    n253
  );


  not
  g1363
  (
    n1250,
    n534
  );


  not
  g1364
  (
    n939,
    n623
  );


  not
  g1365
  (
    n702,
    n476
  );


  not
  g1366
  (
    n873,
    n176
  );


  not
  g1367
  (
    n1047,
    n263
  );


  buf
  g1368
  (
    n1262,
    n626
  );


  not
  g1369
  (
    n1488,
    n363
  );


  buf
  g1370
  (
    n1428,
    n492
  );


  buf
  g1371
  (
    n833,
    n204
  );


  not
  g1372
  (
    n913,
    n307
  );


  not
  g1373
  (
    n1175,
    n349
  );


  not
  g1374
  (
    n1665,
    n620
  );


  not
  g1375
  (
    n1096,
    n584
  );


  not
  g1376
  (
    n933,
    n319
  );


  buf
  g1377
  (
    n1621,
    n509
  );


  not
  g1378
  (
    n1241,
    n638
  );


  not
  g1379
  (
    n792,
    n196
  );


  buf
  g1380
  (
    n1181,
    n241
  );


  buf
  g1381
  (
    n1574,
    n219
  );


  buf
  g1382
  (
    n1052,
    n610
  );


  buf
  g1383
  (
    n1504,
    n234
  );


  not
  g1384
  (
    n753,
    n184
  );


  buf
  g1385
  (
    n1076,
    n355
  );


  not
  g1386
  (
    n1438,
    n205
  );


  buf
  g1387
  (
    n1593,
    n507
  );


  not
  g1388
  (
    n1859,
    n382
  );


  buf
  g1389
  (
    n1437,
    n375
  );


  not
  g1390
  (
    n1845,
    n272
  );


  not
  g1391
  (
    n1661,
    n613
  );


  not
  g1392
  (
    n1236,
    n349
  );


  not
  g1393
  (
    n1746,
    n604
  );


  not
  g1394
  (
    n1231,
    n326
  );


  not
  g1395
  (
    n1343,
    n620
  );


  buf
  g1396
  (
    n1288,
    n631
  );


  buf
  g1397
  (
    n985,
    n269
  );


  buf
  g1398
  (
    n1505,
    n570
  );


  buf
  g1399
  (
    n1520,
    n400
  );


  buf
  g1400
  (
    n1333,
    n401
  );


  buf
  g1401
  (
    n770,
    n549
  );


  buf
  g1402
  (
    n1836,
    n164
  );


  not
  g1403
  (
    n1742,
    n492
  );


  buf
  g1404
  (
    n1824,
    n548
  );


  not
  g1405
  (
    n834,
    n230
  );


  not
  g1406
  (
    n858,
    n210
  );


  buf
  g1407
  (
    n1867,
    n267
  );


  not
  g1408
  (
    n842,
    n170
  );


  not
  g1409
  (
    n1510,
    n446
  );


  not
  g1410
  (
    n1762,
    n239
  );


  not
  g1411
  (
    n1107,
    n299
  );


  not
  g1412
  (
    n1716,
    n439
  );


  buf
  g1413
  (
    n1772,
    n607
  );


  not
  g1414
  (
    n1449,
    n536
  );


  buf
  g1415
  (
    n1413,
    n526
  );


  not
  g1416
  (
    n1247,
    n378
  );


  buf
  g1417
  (
    n1223,
    n488
  );


  not
  g1418
  (
    n1869,
    n486
  );


  buf
  g1419
  (
    n1440,
    n396
  );


  not
  g1420
  (
    n1157,
    n500
  );


  not
  g1421
  (
    n705,
    n226
  );


  buf
  g1422
  (
    n801,
    n182
  );


  not
  g1423
  (
    n1390,
    n376
  );


  not
  g1424
  (
    n1177,
    n575
  );


  buf
  g1425
  (
    n1507,
    n272
  );


  buf
  g1426
  (
    n1136,
    n269
  );


  buf
  g1427
  (
    n1486,
    n392
  );


  buf
  g1428
  (
    n1685,
    n514
  );


  buf
  g1429
  (
    n895,
    n347
  );


  not
  g1430
  (
    n860,
    n180
  );


  buf
  g1431
  (
    n1652,
    n599
  );


  not
  g1432
  (
    n1097,
    n382
  );


  not
  g1433
  (
    n1327,
    n290
  );


  not
  g1434
  (
    n945,
    n305
  );


  buf
  g1435
  (
    n847,
    n243
  );


  not
  g1436
  (
    n668,
    n480
  );


  not
  g1437
  (
    n1063,
    n364
  );


  buf
  g1438
  (
    n1331,
    n395
  );


  buf
  g1439
  (
    n866,
    n493
  );


  buf
  g1440
  (
    n987,
    n537
  );


  not
  g1441
  (
    n911,
    n168
  );


  buf
  g1442
  (
    n1084,
    n458
  );


  not
  g1443
  (
    n812,
    n443
  );


  buf
  g1444
  (
    n1459,
    n427
  );


  buf
  g1445
  (
    n922,
    n404
  );


  not
  g1446
  (
    n1806,
    n444
  );


  not
  g1447
  (
    n1602,
    n472
  );


  buf
  g1448
  (
    n1811,
    n649
  );


  buf
  g1449
  (
    n1005,
    n491
  );


  buf
  g1450
  (
    n1315,
    n527
  );


  buf
  g1451
  (
    n1654,
    n220
  );


  buf
  g1452
  (
    n854,
    n494
  );


  not
  g1453
  (
    n886,
    n229
  );


  not
  g1454
  (
    n927,
    n310
  );


  not
  g1455
  (
    n1832,
    n216
  );


  not
  g1456
  (
    n1180,
    n210
  );


  not
  g1457
  (
    n680,
    n595
  );


  buf
  g1458
  (
    n1509,
    n577
  );


  buf
  g1459
  (
    n898,
    n550
  );


  buf
  g1460
  (
    n1079,
    n616
  );


  not
  g1461
  (
    n1521,
    n539
  );


  not
  g1462
  (
    n1755,
    n504
  );


  buf
  g1463
  (
    n1744,
    n378
  );


  buf
  g1464
  (
    n908,
    n593
  );


  buf
  g1465
  (
    n708,
    n346
  );


  buf
  g1466
  (
    n1557,
    n365
  );


  not
  g1467
  (
    n1234,
    n363
  );


  buf
  g1468
  (
    n1804,
    n434
  );


  buf
  g1469
  (
    n880,
    n475
  );


  not
  g1470
  (
    n1276,
    n462
  );


  buf
  g1471
  (
    n1323,
    n535
  );


  not
  g1472
  (
    n1412,
    n312
  );


  not
  g1473
  (
    n1774,
    n531
  );


  buf
  g1474
  (
    n1550,
    n255
  );


  not
  g1475
  (
    n1763,
    n297
  );


  not
  g1476
  (
    n1720,
    n608
  );


  buf
  g1477
  (
    n1161,
    n397
  );


  buf
  g1478
  (
    n1099,
    n391
  );


  not
  g1479
  (
    n1668,
    n246
  );


  not
  g1480
  (
    n1541,
    n168
  );


  not
  g1481
  (
    n1211,
    n518
  );


  buf
  g1482
  (
    n688,
    n380
  );


  not
  g1483
  (
    n909,
    n538
  );


  buf
  g1484
  (
    n992,
    n415
  );


  buf
  g1485
  (
    n1430,
    n303
  );


  not
  g1486
  (
    n1606,
    n640
  );


  buf
  g1487
  (
    n1785,
    n361
  );


  not
  g1488
  (
    n1703,
    n366
  );


  buf
  g1489
  (
    n710,
    n447
  );


  buf
  g1490
  (
    n870,
    n448
  );


  not
  g1491
  (
    n691,
    n444
  );


  buf
  g1492
  (
    n1383,
    n479
  );


  not
  g1493
  (
    n730,
    n307
  );


  buf
  g1494
  (
    n1317,
    n309
  );


  buf
  g1495
  (
    n1657,
    n330
  );


  not
  g1496
  (
    n1860,
    n286
  );


  buf
  g1497
  (
    n751,
    n403
  );


  not
  g1498
  (
    n821,
    n593
  );


  not
  g1499
  (
    n896,
    n405
  );


  buf
  g1500
  (
    n1841,
    n204
  );


  not
  g1501
  (
    n1088,
    n632
  );


  buf
  g1502
  (
    n1776,
    n453
  );


  buf
  g1503
  (
    n996,
    n321
  );


  buf
  g1504
  (
    n1515,
    n348
  );


  buf
  g1505
  (
    n1191,
    n398
  );


  not
  g1506
  (
    n1081,
    n486
  );


  buf
  g1507
  (
    n1319,
    n257
  );


  not
  g1508
  (
    n1411,
    n391
  );


  not
  g1509
  (
    n1681,
    n468
  );


  not
  g1510
  (
    n1037,
    n387
  );


  buf
  g1511
  (
    n795,
    n573
  );


  buf
  g1512
  (
    n989,
    n500
  );


  not
  g1513
  (
    n772,
    n217
  );


  buf
  g1514
  (
    n723,
    n456
  );


  not
  g1515
  (
    n844,
    n541
  );


  not
  g1516
  (
    n878,
    n591
  );


  buf
  g1517
  (
    n1377,
    n296
  );


  not
  g1518
  (
    n1102,
    n617
  );


  not
  g1519
  (
    n1146,
    n598
  );


  buf
  g1520
  (
    n1007,
    n540
  );


  buf
  g1521
  (
    n1467,
    n574
  );


  buf
  g1522
  (
    n1678,
    n325
  );


  not
  g1523
  (
    n1240,
    n259
  );


  not
  g1524
  (
    n690,
    n454
  );


  not
  g1525
  (
    n1591,
    n441
  );


  not
  g1526
  (
    n1029,
    n433
  );


  not
  g1527
  (
    n1676,
    n192
  );


  buf
  g1528
  (
    n1435,
    n530
  );


  not
  g1529
  (
    n1365,
    n200
  );


  not
  g1530
  (
    n737,
    n641
  );


  buf
  g1531
  (
    n1156,
    n409
  );


  not
  g1532
  (
    n1502,
    n362
  );


  not
  g1533
  (
    n1418,
    n551
  );


  not
  g1534
  (
    n824,
    n400
  );


  buf
  g1535
  (
    n729,
    n554
  );


  buf
  g1536
  (
    n742,
    n385
  );


  buf
  g1537
  (
    n1429,
    n361
  );


  not
  g1538
  (
    n1741,
    n499
  );


  not
  g1539
  (
    n1406,
    n543
  );


  not
  g1540
  (
    n1648,
    n203
  );


  not
  g1541
  (
    n1330,
    n630
  );


  buf
  g1542
  (
    n1626,
    n239
  );


  not
  g1543
  (
    n678,
    n479
  );


  not
  g1544
  (
    n1129,
    n419
  );


  buf
  g1545
  (
    n1362,
    n258
  );


  not
  g1546
  (
    n948,
    n589
  );


  buf
  g1547
  (
    n946,
    n395
  );


  not
  g1548
  (
    n1590,
    n292
  );


  buf
  g1549
  (
    n1051,
    n491
  );


  buf
  g1550
  (
    n802,
    n636
  );


  not
  g1551
  (
    n851,
    n220
  );


  not
  g1552
  (
    n1322,
    n428
  );


  buf
  g1553
  (
    n1771,
    n277
  );


  buf
  g1554
  (
    n1478,
    n212
  );


  buf
  g1555
  (
    n1347,
    n635
  );


  not
  g1556
  (
    n877,
    n556
  );


  not
  g1557
  (
    n967,
    n275
  );


  not
  g1558
  (
    n1284,
    n284
  );


  buf
  g1559
  (
    n1387,
    n332
  );


  buf
  g1560
  (
    n739,
    n280
  );


  buf
  g1561
  (
    n1608,
    n586
  );


  not
  g1562
  (
    n782,
    n422
  );


  not
  g1563
  (
    n1307,
    n182
  );


  not
  g1564
  (
    n941,
    n209
  );


  not
  g1565
  (
    n681,
    n473
  );


  not
  g1566
  (
    n1143,
    n301
  );


  buf
  g1567
  (
    n1173,
    n563
  );


  buf
  g1568
  (
    n1148,
    n350
  );


  not
  g1569
  (
    n1713,
    n162
  );


  buf
  g1570
  (
    n1861,
    n351
  );


  buf
  g1571
  (
    n777,
    n331
  );


  not
  g1572
  (
    n1731,
    n638
  );


  buf
  g1573
  (
    n1204,
    n459
  );


  buf
  g1574
  (
    n1400,
    n335
  );


  buf
  g1575
  (
    n905,
    n247
  );


  not
  g1576
  (
    n1618,
    n362
  );


  buf
  g1577
  (
    n1391,
    n583
  );


  not
  g1578
  (
    n809,
    n485
  );


  not
  g1579
  (
    n1491,
    n572
  );


  buf
  g1580
  (
    n764,
    n195
  );


  nor
  g1581
  (
    n1041,
    n263,
    n382,
    n448,
    n521
  );


  and
  g1582
  (
    n1113,
    n166,
    n583,
    n540,
    n636
  );


  and
  g1583
  (
    n1314,
    n356,
    n519,
    n481,
    n470
  );


  xor
  g1584
  (
    n1363,
    n590,
    n328,
    n215,
    n235
  );


  nand
  g1585
  (
    n1781,
    n197,
    n482,
    n425,
    n273
  );


  nand
  g1586
  (
    n1823,
    n438,
    n594,
    n371,
    n275
  );


  nor
  g1587
  (
    n1674,
    n279,
    n484,
    n204,
    n321
  );


  or
  g1588
  (
    n1768,
    n389,
    n289,
    n343,
    n541
  );


  xnor
  g1589
  (
    n1765,
    n338,
    n371,
    n579,
    n224
  );


  nor
  g1590
  (
    n1263,
    n428,
    n300,
    n542,
    n177
  );


  xnor
  g1591
  (
    n982,
    n605,
    n492,
    n246,
    n490
  );


  nand
  g1592
  (
    n1295,
    n345,
    n175,
    n389,
    n327
  );


  xnor
  g1593
  (
    n1039,
    n449,
    n231,
    n623,
    n228
  );


  nor
  g1594
  (
    n829,
    n609,
    n434,
    n629,
    n618
  );


  xor
  g1595
  (
    n900,
    n414,
    n539,
    n218,
    n232
  );


  and
  g1596
  (
    n1695,
    n624,
    n615,
    n312,
    n489
  );


  or
  g1597
  (
    n1398,
    n625,
    n279,
    n306,
    n225
  );


  xnor
  g1598
  (
    n1015,
    n471,
    n340,
    n260,
    n428
  );


  xnor
  g1599
  (
    n1529,
    n525,
    n288,
    n254,
    n533
  );


  and
  g1600
  (
    n1547,
    n625,
    n297,
    n219,
    n431
  );


  and
  g1601
  (
    n1367,
    n229,
    n375,
    n426,
    n524
  );


  and
  g1602
  (
    n828,
    n601,
    n570,
    n405,
    n415
  );


  nor
  g1603
  (
    n1471,
    n407,
    n631,
    n376,
    n373
  );


  xor
  g1604
  (
    n817,
    n226,
    n560,
    n423,
    n479
  );


  nor
  g1605
  (
    n1795,
    n265,
    n545,
    n452,
    n587
  );


  nor
  g1606
  (
    n1329,
    n270,
    n242,
    n419,
    n647
  );


  nor
  g1607
  (
    n1267,
    n654,
    n463,
    n641,
    n460
  );


  nor
  g1608
  (
    n1603,
    n244,
    n489,
    n215,
    n379
  );


  nor
  g1609
  (
    n921,
    n517,
    n430,
    n612,
    n441
  );


  xor
  g1610
  (
    n1203,
    n374,
    n198,
    n253,
    n250
  );


  xor
  g1611
  (
    n704,
    n274,
    n285,
    n370,
    n235
  );


  xnor
  g1612
  (
    n1357,
    n571,
    n356,
    n618,
    n625
  );


  xor
  g1613
  (
    n1235,
    n557,
    n277,
    n576,
    n559
  );


  xor
  g1614
  (
    n747,
    n326,
    n391,
    n651,
    n334
  );


  nand
  g1615
  (
    n944,
    n352,
    n652,
    n304,
    n167
  );


  or
  g1616
  (
    n1465,
    n578,
    n333,
    n642,
    n194
  );


  xor
  g1617
  (
    n1500,
    n463,
    n483,
    n348,
    n636
  );


  nor
  g1618
  (
    n1160,
    n560,
    n548,
    n581,
    n633
  );


  nor
  g1619
  (
    n1292,
    n424,
    n564,
    n384,
    n360
  );


  nand
  g1620
  (
    n1009,
    n281,
    n174,
    n343,
    n520
  );


  nand
  g1621
  (
    n1810,
    n441,
    n552,
    n455,
    n486
  );


  and
  g1622
  (
    n721,
    n484,
    n530,
    n535,
    n362
  );


  nor
  g1623
  (
    n711,
    n454,
    n189,
    n381,
    n252
  );


  xnor
  g1624
  (
    n1549,
    n315,
    n384,
    n318,
    n540
  );


  nand
  g1625
  (
    n1335,
    n195,
    n318,
    n273,
    n554
  );


  and
  g1626
  (
    n1140,
    n328,
    n517,
    n562,
    n640
  );


  nand
  g1627
  (
    n1616,
    n177,
    n341,
    n257,
    n170
  );


  or
  g1628
  (
    n1044,
    n173,
    n545,
    n507,
    n519
  );


  xor
  g1629
  (
    n868,
    n371,
    n213,
    n319,
    n287
  );


  nor
  g1630
  (
    n1683,
    n597,
    n202,
    n265,
    n450
  );


  xnor
  g1631
  (
    n1632,
    n237,
    n652,
    n502,
    n432
  );


  xnor
  g1632
  (
    n1493,
    n520,
    n439,
    n378,
    n198
  );


  and
  g1633
  (
    n1531,
    n627,
    n214,
    n219,
    n346
  );


  nor
  g1634
  (
    n1445,
    n292,
    n354,
    n544,
    n234
  );


  xor
  g1635
  (
    n1706,
    n186,
    n329,
    n336,
    n358
  );


  and
  g1636
  (
    n1123,
    n349,
    n248,
    n293,
    n475
  );


  nand
  g1637
  (
    n1120,
    n461,
    n457,
    n380,
    n414
  );


  and
  g1638
  (
    n716,
    n437,
    n459,
    n452,
    n429
  );


  nor
  g1639
  (
    n1612,
    n366,
    n470,
    n212,
    n233
  );


  nor
  g1640
  (
    n1268,
    n176,
    n240,
    n644,
    n505
  );


  nand
  g1641
  (
    n1688,
    n237,
    n282,
    n261,
    n463
  );


  xnor
  g1642
  (
    n696,
    n176,
    n445,
    n244,
    n584
  );


  xor
  g1643
  (
    n1732,
    n166,
    n344,
    n245,
    n402
  );


  and
  g1644
  (
    n1421,
    n600,
    n543,
    n361,
    n649
  );


  xnor
  g1645
  (
    n1692,
    n440,
    n366,
    n445,
    n571
  );


  and
  g1646
  (
    n1251,
    n365,
    n597,
    n226,
    n234
  );


  and
  g1647
  (
    n1643,
    n432,
    n416,
    n333,
    n244
  );


  nor
  g1648
  (
    n1416,
    n547,
    n418,
    n586,
    n291
  );


  xor
  g1649
  (
    n1496,
    n296,
    n627,
    n641,
    n498
  );


  nand
  g1650
  (
    n1863,
    n308,
    n490,
    n351,
    n256
  );


  and
  g1651
  (
    n856,
    n353,
    n384,
    n456,
    n643
  );


  nand
  g1652
  (
    n1338,
    n390,
    n436,
    n267,
    n347
  );


  nand
  g1653
  (
    n1417,
    n515,
    n316,
    n641,
    n352
  );


  xnor
  g1654
  (
    n1065,
    n244,
    n519,
    n580,
    n334
  );


  xor
  g1655
  (
    n1546,
    n442,
    n650,
    n191,
    n288
  );


  xor
  g1656
  (
    n998,
    n513,
    n546,
    n340,
    n569
  );


  nand
  g1657
  (
    n1670,
    n474,
    n301,
    n522,
    n238
  );


  nand
  g1658
  (
    n1456,
    n388,
    n213,
    n634,
    n468
  );


  or
  g1659
  (
    n713,
    n529,
    n172,
    n294,
    n262
  );


  xnor
  g1660
  (
    n718,
    n371,
    n403,
    n194,
    n543
  );


  xnor
  g1661
  (
    n1498,
    n435,
    n208,
    n380,
    n579
  );


  nor
  g1662
  (
    n1671,
    n543,
    n352,
    n253,
    n187
  );


  and
  g1663
  (
    n1628,
    n446,
    n368,
    n422,
    n359
  );


  xor
  g1664
  (
    n1769,
    n323,
    n412,
    n513,
    n606
  );


  nor
  g1665
  (
    n1078,
    n558,
    n411,
    n587,
    n495
  );


  nand
  g1666
  (
    n1054,
    n556,
    n202,
    n572,
    n531
  );


  and
  g1667
  (
    n1711,
    n590,
    n470,
    n340,
    n579
  );


  nand
  g1668
  (
    n914,
    n601,
    n421,
    n414,
    n571
  );


  nand
  g1669
  (
    n1672,
    n320,
    n413,
    n386,
    n614
  );


  nor
  g1670
  (
    n1760,
    n559,
    n481,
    n326,
    n255
  );


  xor
  g1671
  (
    n1444,
    n259,
    n275,
    n650,
    n508
  );


  nand
  g1672
  (
    n1820,
    n316,
    n282,
    n175,
    n350
  );


  and
  g1673
  (
    n1660,
    n303,
    n495,
    n283,
    n502
  );


  xnor
  g1674
  (
    n1248,
    n562,
    n280,
    n536,
    n313
  );


  xnor
  g1675
  (
    n1423,
    n613,
    n609,
    n183,
    n417
  );


  xnor
  g1676
  (
    n1564,
    n183,
    n423,
    n287,
    n531
  );


  xnor
  g1677
  (
    n1827,
    n339,
    n396,
    n399,
    n514
  );


  xnor
  g1678
  (
    n1062,
    n618,
    n452,
    n446,
    n516
  );


  and
  g1679
  (
    n1684,
    n174,
    n403,
    n431,
    n473
  );


  nor
  g1680
  (
    n1269,
    n177,
    n168,
    n458,
    n289
  );


  xor
  g1681
  (
    n857,
    n273,
    n218,
    n375,
    n367
  );


  xor
  g1682
  (
    n1791,
    n182,
    n483,
    n562,
    n400
  );


  nor
  g1683
  (
    n1359,
    n259,
    n615,
    n298,
    n302
  );


  or
  g1684
  (
    n1718,
    n466,
    n203,
    n348,
    n594
  );


  xor
  g1685
  (
    n953,
    n223,
    n236,
    n628,
    n231
  );


  xnor
  g1686
  (
    n1075,
    n432,
    n629,
    n544,
    n506
  );


  and
  g1687
  (
    n1258,
    n383,
    n309,
    n567,
    n356
  );


  nand
  g1688
  (
    n727,
    n620,
    n524,
    n175,
    n478
  );


  nor
  g1689
  (
    n1179,
    n606,
    n396,
    n346,
    n538
  );


  or
  g1690
  (
    n979,
    n582,
    n242,
    n424,
    n472
  );


  nor
  g1691
  (
    n1415,
    n461,
    n434,
    n511,
    n532
  );


  or
  g1692
  (
    n1309,
    n617,
    n217,
    n596,
    n417
  );


  and
  g1693
  (
    n1110,
    n173,
    n627,
    n464,
    n566
  );


  nand
  g1694
  (
    n1324,
    n367,
    n278,
    n588,
    n556
  );


  or
  g1695
  (
    n1585,
    n346,
    n499,
    n480,
    n461
  );


  or
  g1696
  (
    n1600,
    n208,
    n259,
    n488,
    n281
  );


  xnor
  g1697
  (
    n1649,
    n265,
    n644,
    n192
  );


  xor
  g1698
  (
    n1592,
    n596,
    n447,
    n283,
    n327
  );


  and
  g1699
  (
    n1035,
    n460,
    n643,
    n475,
    n598
  );


  nor
  g1700
  (
    n1022,
    n623,
    n374,
    n179,
    n170
  );


  or
  g1701
  (
    n1057,
    n190,
    n510,
    n477,
    n401
  );


  or
  g1702
  (
    n1401,
    n171,
    n637,
    n648,
    n482
  );


  xnor
  g1703
  (
    n1378,
    n212,
    n188,
    n568,
    n344
  );


  or
  g1704
  (
    n1217,
    n186,
    n555,
    n196,
    n354
  );


  xnor
  g1705
  (
    n971,
    n221,
    n207,
    n430,
    n590
  );


  xnor
  g1706
  (
    n988,
    n329,
    n469,
    n548,
    n494
  );


  nand
  g1707
  (
    n1286,
    n196,
    n467,
    n416,
    n297
  );


  nand
  g1708
  (
    n1142,
    n223,
    n457,
    n621,
    n295
  );


  nand
  g1709
  (
    n1298,
    n602,
    n203,
    n264,
    n490
  );


  nor
  g1710
  (
    n1004,
    n369,
    n436,
    n399,
    n463
  );


  or
  g1711
  (
    n1326,
    n305,
    n609,
    n383,
    n314
  );


  and
  g1712
  (
    n763,
    n640,
    n291,
    n385,
    n512
  );


  and
  g1713
  (
    n780,
    n402,
    n161,
    n597,
    n616
  );


  and
  g1714
  (
    n1629,
    n653,
    n633,
    n461,
    n201
  );


  or
  g1715
  (
    n1215,
    n342,
    n601,
    n306,
    n637
  );


  xnor
  g1716
  (
    n1011,
    n502,
    n351,
    n539,
    n613
  );


  and
  g1717
  (
    n1562,
    n290,
    n517,
    n418,
    n477
  );


  xnor
  g1718
  (
    n1119,
    n255,
    n283,
    n305,
    n389
  );


  xnor
  g1719
  (
    n736,
    n290,
    n246,
    n452,
    n349
  );


  and
  g1720
  (
    n1476,
    n605,
    n280,
    n232,
    n455
  );


  nand
  g1721
  (
    n1392,
    n327,
    n614,
    n595,
    n449
  );


  and
  g1722
  (
    n1101,
    n455,
    n262,
    n614,
    n547
  );


  xor
  g1723
  (
    n1702,
    n642,
    n583,
    n201,
    n178
  );


  xor
  g1724
  (
    n1848,
    n287,
    n487,
    n183,
    n427
  );


  nor
  g1725
  (
    n804,
    n197,
    n313,
    n240,
    n163
  );


  nor
  g1726
  (
    n1594,
    n545,
    n605,
    n648,
    n453
  );


  nor
  g1727
  (
    n1304,
    n195,
    n211,
    n440,
    n610
  );


  xnor
  g1728
  (
    n803,
    n485,
    n318,
    n379,
    n184
  );


  xnor
  g1729
  (
    n1352,
    n421,
    n306,
    n228
  );


  or
  g1730
  (
    n1019,
    n282,
    n577,
    n182,
    n421
  );


  or
  g1731
  (
    n1739,
    n343,
    n594,
    n199,
    n279
  );


  nand
  g1732
  (
    n1489,
    n451,
    n257,
    n260,
    n358
  );


  nand
  g1733
  (
    n1144,
    n646,
    n397,
    n465,
    n210
  );


  xnor
  g1734
  (
    n1221,
    n174,
    n487,
    n359,
    n565
  );


  nor
  g1735
  (
    n1219,
    n428,
    n284,
    n450,
    n235
  );


  nand
  g1736
  (
    n1682,
    n298,
    n184,
    n552,
    n631
  );


  and
  g1737
  (
    n894,
    n634,
    n506,
    n322,
    n401
  );


  or
  g1738
  (
    n1870,
    n365,
    n526,
    n187,
    n274
  );


  and
  g1739
  (
    n1293,
    n341,
    n281,
    n423,
    n410
  );


  nand
  g1740
  (
    n1077,
    n622,
    n361,
    n434,
    n401
  );


  nor
  g1741
  (
    n1431,
    n550,
    n377,
    n300,
    n303
  );


  xnor
  g1742
  (
    n1209,
    n200,
    n380,
    n297,
    n245
  );


  nand
  g1743
  (
    n1807,
    n336,
    n557,
    n408,
    n179
  );


  and
  g1744
  (
    n676,
    n496,
    n459,
    n185,
    n460
  );


  xor
  g1745
  (
    n1114,
    n368,
    n207,
    n467,
    n631
  );


  nand
  g1746
  (
    n1164,
    n501,
    n188,
    n272,
    n587
  );


  nand
  g1747
  (
    n935,
    n394,
    n379,
    n633,
    n184
  );


  nor
  g1748
  (
    KeyWire_0_9,
    n473,
    n353,
    n267,
    n399
  );


  nand
  g1749
  (
    n793,
    n390,
    n638,
    n197,
    n392
  );


  nor
  g1750
  (
    n1849,
    n317,
    n383,
    n567,
    n394
  );


  nand
  g1751
  (
    n1563,
    n532,
    n527,
    n573,
    n546
  );


  and
  g1752
  (
    n1170,
    n252,
    n602,
    n193,
    n607
  );


  or
  g1753
  (
    n1855,
    n596,
    n355,
    n236,
    n251
  );


  and
  g1754
  (
    n1475,
    n600,
    n521,
    n480,
    n194
  );


  nor
  g1755
  (
    n1460,
    n630,
    n186,
    n622,
    n249
  );


  nand
  g1756
  (
    n1364,
    n393,
    n435,
    n313,
    n617
  );


  nand
  g1757
  (
    n1257,
    n646,
    n324,
    n276,
    n363
  );


  and
  g1758
  (
    n1735,
    n236,
    n619,
    n589,
    n192
  );


  nand
  g1759
  (
    n1152,
    n515,
    n604,
    n644,
    n309
  );


  nor
  g1760
  (
    n1200,
    n566,
    n478,
    n217,
    n193
  );


  nand
  g1761
  (
    n1246,
    n191,
    n506,
    n337,
    n195
  );


  or
  g1762
  (
    n1727,
    n446,
    n178,
    n209,
    n370
  );


  or
  g1763
  (
    n1356,
    n161,
    n554,
    n213,
    n483
  );


  nand
  g1764
  (
    n1659,
    n598,
    n433,
    n233,
    n301
  );


  or
  g1765
  (
    n853,
    n595,
    n621,
    n579,
    n172
  );


  or
  g1766
  (
    n1583,
    n211,
    n319,
    n630,
    n406
  );


  nor
  g1767
  (
    n1206,
    n290,
    n467,
    n364,
    n172
  );


  or
  g1768
  (
    n1040,
    n209,
    n574,
    n496,
    n409
  );


  and
  g1769
  (
    n1821,
    n263,
    n390,
    n563,
    n295
  );


  xor
  g1770
  (
    n1831,
    n314,
    n419,
    n241,
    n171
  );


  and
  g1771
  (
    n1394,
    n539,
    n323,
    n218,
    n294
  );


  nand
  g1772
  (
    n1675,
    n512,
    n647,
    n491,
    n294
  );


  or
  g1773
  (
    n800,
    n630,
    n456,
    n163,
    n542
  );


  and
  g1774
  (
    n1817,
    n425,
    n559,
    n315,
    n519
  );


  nand
  g1775
  (
    n799,
    n407,
    n307,
    n431,
    n386
  );


  nor
  g1776
  (
    n1662,
    n193,
    n608,
    n362,
    n507
  );


  nor
  g1777
  (
    n1351,
    n372,
    n347,
    n622,
    n585
  );


  xnor
  g1778
  (
    n1229,
    n211,
    n163,
    n478,
    n573
  );


  or
  g1779
  (
    n1704,
    n425,
    n353,
    n219,
    n165
  );


  xor
  g1780
  (
    n1405,
    n490,
    n363,
    n654,
    n610
  );


  and
  g1781
  (
    n1473,
    n407,
    n186,
    n578,
    n496
  );


  and
  g1782
  (
    n1432,
    n181,
    n465,
    n426,
    n296
  );


  or
  g1783
  (
    n1158,
    n471,
    n424,
    n266,
    n550
  );


  or
  g1784
  (
    n1694,
    n398,
    n522,
    n356,
    n178
  );


  nand
  g1785
  (
    n1064,
    n385,
    n396,
    n214,
    n229
  );


  nor
  g1786
  (
    n1854,
    n312,
    n619,
    n499,
    n358
  );


  xnor
  g1787
  (
    n1856,
    n250,
    n569,
    n404,
    n488
  );


  nand
  g1788
  (
    n1851,
    n278,
    n580,
    n336,
    n248
  );


  nand
  g1789
  (
    n1371,
    n497,
    n654,
    n368,
    n216
  );


  and
  g1790
  (
    n1106,
    n565,
    n308,
    n357,
    n223
  );


  or
  g1791
  (
    n1067,
    n286,
    n608,
    n639,
    n572
  );


  nor
  g1792
  (
    n1296,
    n368,
    n505,
    n284,
    n581
  );


  xnor
  g1793
  (
    n1770,
    n238,
    n269,
    n232,
    n504
  );


  xor
  g1794
  (
    n1061,
    n289,
    n513,
    n345,
    n224
  );


  and
  g1795
  (
    n1369,
    n265,
    n209,
    n250,
    n483
  );


  and
  g1796
  (
    n1799,
    n387,
    n315,
    n603,
    n276
  );


  nor
  g1797
  (
    n1050,
    n245,
    n214,
    n616,
    n494
  );


  nand
  g1798
  (
    n698,
    n552,
    n203,
    n337,
    n232
  );


  nand
  g1799
  (
    n1066,
    n370,
    n405,
    n392,
    n553
  );


  or
  g1800
  (
    n1650,
    n561,
    n477,
    n398,
    n238
  );


  or
  g1801
  (
    n949,
    n220,
    n311,
    n547,
    n605
  );


  or
  g1802
  (
    n916,
    n176,
    n545,
    n576,
    n518
  );


  or
  g1803
  (
    n1669,
    n261,
    n291,
    n266,
    n431
  );


  or
  g1804
  (
    n938,
    n415,
    n185,
    n532,
    n206
  );


  nor
  g1805
  (
    n1408,
    n551,
    n318,
    n512,
    n413
  );


  nand
  g1806
  (
    n818,
    n646,
    n190,
    n555,
    n374
  );


  nor
  g1807
  (
    n1833,
    n350,
    n376,
    n495,
    n514
  );


  or
  g1808
  (
    n1150,
    n369,
    n266,
    n538,
    n307
  );


  nor
  g1809
  (
    n1376,
    n626,
    n555,
    n527,
    n508
  );


  xnor
  g1810
  (
    n1193,
    n529,
    n485,
    n208,
    n615
  );


  nand
  g1811
  (
    n1138,
    n509,
    n655,
    n422,
    n308
  );


  xnor
  g1812
  (
    n1726,
    n279,
    n594,
    n180,
    n198
  );


  and
  g1813
  (
    n1542,
    n469,
    n398,
    n498,
    n470
  );


  nor
  g1814
  (
    n1311,
    n497,
    n603,
    n271,
    n381
  );


  xor
  g1815
  (
    n1059,
    n635,
    n303,
    n364,
    n500
  );


  nand
  g1816
  (
    n1424,
    n505,
    n270,
    n289,
    n593
  );


  nand
  g1817
  (
    n1853,
    n635,
    n345,
    n311,
    n177
  );


  nor
  g1818
  (
    n901,
    n558,
    n324,
    n174,
    n374
  );


  or
  g1819
  (
    n738,
    n288,
    n588,
    n317,
    n292
  );


  xnor
  g1820
  (
    n1783,
    n373,
    n238,
    n181,
    n319
  );


  nor
  g1821
  (
    n814,
    n168,
    n578,
    n263,
    n189
  );


  and
  g1822
  (
    n1450,
    n214,
    n563,
    n484,
    n615
  );


  nor
  g1823
  (
    n1108,
    n328,
    n511,
    n505,
    n302
  );


  nand
  g1824
  (
    n1021,
    n523,
    n528,
    n564,
    n559
  );


  xnor
  g1825
  (
    n1644,
    n510,
    n310,
    n236,
    n271
  );


  xor
  g1826
  (
    n714,
    n199,
    n208,
    n598,
    n566
  );


  xnor
  g1827
  (
    n1230,
    n173,
    n410,
    n652,
    n181
  );


  and
  g1828
  (
    n984,
    n331,
    n438,
    n645,
    n230
  );


  and
  g1829
  (
    n1868,
    n645,
    n514,
    n247,
    n314
  );


  xnor
  g1830
  (
    n1710,
    n533,
    n521,
    n277,
    n628
  );


  and
  g1831
  (
    n1793,
    n171,
    n558,
    n408,
    n567
  );


  xor
  g1832
  (
    n1725,
    n381,
    n563,
    n582,
    n509
  );


  xor
  g1833
  (
    n936,
    n292,
    n536,
    n565,
    n335
  );


  nor
  g1834
  (
    n1808,
    n541,
    n484,
    n591,
    n411
  );


  nor
  g1835
  (
    n1038,
    n294,
    n554,
    n322,
    n612
  );


  xor
  g1836
  (
    n749,
    n164,
    n548,
    n322,
    n332
  );


  and
  g1837
  (
    n685,
    n597,
    n629,
    n651,
    n540
  );


  and
  g1838
  (
    n1886,
    n1035,
    n755,
    n1467,
    n1053
  );


  and
  g1839
  (
    n1997,
    n1311,
    n1294,
    n1172,
    n1232
  );


  nor
  g1840
  (
    n1925,
    n857,
    n975,
    n1335,
    n1039
  );


  xnor
  g1841
  (
    n1882,
    n876,
    n1427,
    n1176,
    n767
  );


  xor
  g1842
  (
    n1878,
    n672,
    n955,
    n1451,
    n1491
  );


  xnor
  g1843
  (
    n1981,
    n1403,
    n800,
    n757,
    n1309
  );


  or
  g1844
  (
    n2002,
    n692,
    n895,
    n1436,
    n1296
  );


  or
  g1845
  (
    n1892,
    n827,
    n1002,
    n1069,
    n718
  );


  nand
  g1846
  (
    n1988,
    n978,
    n690,
    n1394,
    n1047
  );


  nand
  g1847
  (
    n1896,
    n1236,
    n1262,
    n1355,
    n1315
  );


  and
  g1848
  (
    n2067,
    n1033,
    n1182,
    n1192,
    n1246
  );


  and
  g1849
  (
    n2001,
    n779,
    n1054,
    n925,
    n860
  );


  nand
  g1850
  (
    n2044,
    n1361,
    n1185,
    n1010,
    n1241
  );


  nand
  g1851
  (
    n2063,
    n1282,
    n1046,
    n1444,
    n1215
  );


  xnor
  g1852
  (
    n1999,
    n1257,
    n818,
    n709,
    n1050
  );


  xor
  g1853
  (
    n1962,
    n1199,
    n959,
    n1382,
    n1051
  );


  or
  g1854
  (
    n1969,
    n1169,
    n1098,
    n970,
    n765
  );


  nand
  g1855
  (
    n1924,
    n795,
    n778,
    n770,
    n1374
  );


  xnor
  g1856
  (
    n1996,
    n986,
    n930,
    n1300,
    n904
  );


  nand
  g1857
  (
    n1898,
    n826,
    n989,
    n1020,
    n1022
  );


  xor
  g1858
  (
    n2054,
    n1235,
    n1250,
    n813,
    n674
  );


  nand
  g1859
  (
    n1971,
    n1493,
    n802,
    n1214,
    n1011
  );


  or
  g1860
  (
    n2017,
    n1462,
    n845,
    n1177,
    n931
  );


  and
  g1861
  (
    n1985,
    n784,
    n1299,
    n1005,
    n1408
  );


  nor
  g1862
  (
    n1923,
    n710,
    n744,
    n803,
    n1225
  );


  nand
  g1863
  (
    n1955,
    n1256,
    n1433,
    n1230,
    n712
  );


  xor
  g1864
  (
    n1880,
    n878,
    n753,
    n1237,
    n886
  );


  and
  g1865
  (
    n1940,
    n1305,
    n1026,
    n764,
    n748
  );


  nor
  g1866
  (
    n2018,
    n797,
    n864,
    n677,
    n1063
  );


  nor
  g1867
  (
    n1909,
    n1340,
    n916,
    n1395,
    n965
  );


  or
  g1868
  (
    n1871,
    n1324,
    n841,
    n920,
    n1146
  );


  xor
  g1869
  (
    n1968,
    n1401,
    n1188,
    n1306,
    n1056
  );


  or
  g1870
  (
    n2015,
    n1000,
    n1397,
    n990,
    n790
  );


  and
  g1871
  (
    n2010,
    n1065,
    n840,
    n1226,
    n1435
  );


  nor
  g1872
  (
    n2039,
    n1460,
    n811,
    n1084,
    n882
  );


  nand
  g1873
  (
    n2007,
    n819,
    n880,
    n734,
    n1052
  );


  and
  g1874
  (
    n2020,
    n1371,
    n1121,
    n906,
    n694
  );


  xor
  g1875
  (
    n1876,
    n1287,
    n736,
    n1245,
    n936
  );


  and
  g1876
  (
    n2013,
    n786,
    n1399,
    n1476,
    n834
  );


  nor
  g1877
  (
    n1984,
    n1320,
    n820,
    n1437,
    n1152
  );


  nand
  g1878
  (
    n1980,
    n1113,
    n666,
    n785,
    n1348
  );


  and
  g1879
  (
    n2040,
    n948,
    n1271,
    n1273,
    n768
  );


  and
  g1880
  (
    n1914,
    n1148,
    n681,
    n1466,
    n1071
  );


  nand
  g1881
  (
    n2027,
    n1195,
    n1290,
    n1074,
    n1420
  );


  xor
  g1882
  (
    n1961,
    n836,
    n749,
    n838,
    n972
  );


  and
  g1883
  (
    n2076,
    n964,
    n1464,
    n829,
    n750
  );


  xor
  g1884
  (
    n2045,
    n1203,
    n730,
    n1304,
    n943
  );


  and
  g1885
  (
    n2071,
    n1062,
    n1267,
    n809,
    n1406
  );


  nand
  g1886
  (
    n2077,
    n998,
    n898,
    n954,
    n1380
  );


  or
  g1887
  (
    n2078,
    n1345,
    n1298,
    n1030,
    n725
  );


  and
  g1888
  (
    n1992,
    n837,
    n810,
    n1123,
    n1137
  );


  xnor
  g1889
  (
    n1901,
    n1354,
    n1258,
    n1356,
    n1372
  );


  nand
  g1890
  (
    KeyWire_0_3,
    n740,
    n950,
    n947,
    n1446
  );


  nor
  g1891
  (
    n2038,
    n1163,
    n977,
    n1249,
    n1313
  );


  nand
  g1892
  (
    n1904,
    n1244,
    n957,
    n1014,
    n1102
  );


  xor
  g1893
  (
    n2056,
    n721,
    n1207,
    n1331,
    n889
  );


  xnor
  g1894
  (
    n1894,
    n1119,
    n1392,
    n706,
    n900
  );


  xnor
  g1895
  (
    n1946,
    n1106,
    n969,
    n1027,
    n1202
  );


  or
  g1896
  (
    n2024,
    n1162,
    n828,
    n974,
    n1293
  );


  and
  g1897
  (
    n1908,
    n1254,
    n1131,
    n1066,
    n1301
  );


  nor
  g1898
  (
    n2026,
    n967,
    n912,
    n1314,
    n722
  );


  nand
  g1899
  (
    n2036,
    n1150,
    n1068,
    n933,
    n891
  );


  xnor
  g1900
  (
    n2011,
    n1191,
    n1283,
    n1440,
    n1449
  );


  nand
  g1901
  (
    n2022,
    n669,
    n997,
    n804,
    n1253
  );


  nand
  g1902
  (
    n1976,
    n942,
    n1402,
    n919,
    n1339
  );


  xnor
  g1903
  (
    n1929,
    n714,
    n1292,
    n1180,
    n1090
  );


  xor
  g1904
  (
    n1982,
    n1155,
    n1019,
    n910,
    n1473
  );


  nand
  g1905
  (
    n1891,
    n1139,
    n793,
    n1379,
    n1307
  );


  nor
  g1906
  (
    n1972,
    n962,
    n1417,
    n1222,
    n1455
  );


  or
  g1907
  (
    n1884,
    n869,
    n745,
    n1461,
    n1213
  );


  nor
  g1908
  (
    n1915,
    n874,
    n679,
    n1398,
    n1431
  );


  xor
  g1909
  (
    n1998,
    n862,
    n1322,
    n1468,
    n752
  );


  and
  g1910
  (
    n2041,
    n1198,
    n1388,
    n1099,
    n1092
  );


  xor
  g1911
  (
    n1935,
    n1492,
    n759,
    n1409,
    n1040
  );


  and
  g1912
  (
    n2014,
    n897,
    n1057,
    n1110,
    n1284
  );


  nor
  g1913
  (
    n2050,
    n1209,
    n1327,
    n1434,
    n1197
  );


  nor
  g1914
  (
    n1907,
    n853,
    n817,
    n1329,
    n846
  );


  nand
  g1915
  (
    n1989,
    n1089,
    n956,
    n1489,
    n830
  );


  or
  g1916
  (
    n1913,
    n871,
    n1488,
    n1079,
    n1456
  );


  xnor
  g1917
  (
    n1975,
    n807,
    n1370,
    n901,
    n1481
  );


  xnor
  g1918
  (
    n1918,
    n1366,
    n852,
    n1483,
    n999
  );


  xnor
  g1919
  (
    n2061,
    n856,
    n703,
    n1142,
    n913
  );


  and
  g1920
  (
    n1943,
    n831,
    n1404,
    n934,
    n918
  );


  xnor
  g1921
  (
    n1895,
    n1042,
    n1414,
    n1485,
    n713
  );


  xor
  g1922
  (
    n1952,
    n756,
    n704,
    n1423,
    n1413
  );


  and
  g1923
  (
    n1977,
    n1337,
    n1268,
    n842,
    n991
  );


  or
  g1924
  (
    n1939,
    n1269,
    n1297,
    n775,
    n1109
  );


  xnor
  g1925
  (
    n2051,
    n1077,
    n1187,
    n1239,
    n984
  );


  or
  g1926
  (
    n1920,
    n1091,
    n1428,
    n1333,
    n890
  );


  xor
  g1927
  (
    n1900,
    n1012,
    n915,
    n1334,
    n1031
  );


  xnor
  g1928
  (
    n2030,
    n1487,
    n1234,
    n1183,
    n1007
  );


  and
  g1929
  (
    n2042,
    n760,
    n774,
    n1075,
    n708
  );


  nand
  g1930
  (
    n2025,
    n1160,
    n855,
    n1044,
    n911
  );


  nand
  g1931
  (
    n1957,
    n1164,
    n1144,
    n1438,
    n958
  );


  and
  g1932
  (
    n2021,
    n1286,
    n1318,
    n1263,
    n1096
  );


  xnor
  g1933
  (
    n1890,
    n1450,
    n1251,
    n1278,
    n1132
  );


  nand
  g1934
  (
    n1995,
    n1006,
    n1114,
    n1439,
    n682
  );


  nand
  g1935
  (
    n2057,
    n766,
    n700,
    n926,
    n1359
  );


  xnor
  g1936
  (
    n1916,
    n1126,
    n973,
    n1470,
    n732
  );


  nand
  g1937
  (
    n1948,
    n963,
    n798,
    n1458,
    n1325
  );


  or
  g1938
  (
    n1937,
    n742,
    n769,
    n1454,
    n1127
  );


  xnor
  g1939
  (
    n1917,
    n1117,
    n1343,
    n994,
    n667
  );


  nor
  g1940
  (
    n1942,
    n858,
    n726,
    n1393,
    n1463
  );


  nor
  g1941
  (
    n2059,
    n678,
    n1120,
    n686,
    n717
  );


  xnor
  g1942
  (
    n1994,
    n1432,
    n938,
    n787,
    n1149
  );


  nor
  g1943
  (
    n1899,
    n822,
    n1145,
    n1342,
    n1457
  );


  xnor
  g1944
  (
    n1978,
    n1328,
    n1274,
    n727,
    n935
  );


  and
  g1945
  (
    n1965,
    n1336,
    n1264,
    n1415,
    n1422
  );


  nand
  g1946
  (
    n2005,
    n747,
    n1344,
    n1083,
    n731
  );


  nor
  g1947
  (
    n2074,
    n1025,
    n739,
    n1326,
    n908
  );


  and
  g1948
  (
    n2029,
    n940,
    n1216,
    n903,
    n691
  );


  xor
  g1949
  (
    n1979,
    n1484,
    n1049,
    n684,
    n1303
  );


  nor
  g1950
  (
    n2028,
    n1276,
    n1338,
    n1008,
    n1261
  );


  xnor
  g1951
  (
    n1902,
    n1101,
    n697,
    n1368,
    n1078
  );


  xor
  g1952
  (
    n1954,
    n1255,
    n1472,
    n881,
    n1194
  );


  and
  g1953
  (
    n1963,
    n1229,
    n1351,
    n1217,
    n676
  );


  nor
  g1954
  (
    n1888,
    n872,
    n1087,
    n952,
    n1064
  );


  or
  g1955
  (
    n1881,
    n1242,
    n1107,
    n1469,
    n723
  );


  nor
  g1956
  (
    n1910,
    n1243,
    n814,
    n701,
    n1224
  );


  nand
  g1957
  (
    n1986,
    n1167,
    n1181,
    n833,
    n1363
  );


  nand
  g1958
  (
    n2047,
    n1453,
    n914,
    n961,
    n894
  );


  and
  g1959
  (
    n1974,
    n1174,
    n1032,
    n1289,
    n823
  );


  xnor
  g1960
  (
    n1987,
    n1111,
    n929,
    n1426,
    n1412
  );


  xnor
  g1961
  (
    n2004,
    n763,
    n1475,
    n854,
    n680
  );


  nor
  g1962
  (
    n1958,
    n980,
    n932,
    n945,
    n1265
  );


  nand
  g1963
  (
    n1945,
    n1391,
    n1159,
    n1352,
    n1266
  );


  or
  g1964
  (
    n1947,
    n1178,
    n687,
    n981,
    n780
  );


  and
  g1965
  (
    n2052,
    n1059,
    n1387,
    n1386,
    n861
  );


  xor
  g1966
  (
    n2072,
    n1248,
    n1093,
    n1227,
    n1165
  );


  and
  g1967
  (
    n1905,
    n728,
    n796,
    n976,
    n698
  );


  nand
  g1968
  (
    n1873,
    n937,
    n685,
    n673,
    n782
  );


  nor
  g1969
  (
    n2012,
    n1041,
    n905,
    n988,
    n693
  );


  nand
  g1970
  (
    n2035,
    n777,
    n859,
    n1317,
    n699
  );


  xor
  g1971
  (
    n1936,
    n1003,
    n1474,
    n1103,
    n983
  );


  xor
  g1972
  (
    n1887,
    n1017,
    n1373,
    n815,
    n1158
  );


  nor
  g1973
  (
    n2043,
    n866,
    n996,
    n1240,
    n1024
  );


  and
  g1974
  (
    n2066,
    n1443,
    n1009,
    n773,
    n702
  );


  nand
  g1975
  (
    KeyWire_0_0,
    n1105,
    n875,
    n1396,
    n1061
  );


  and
  g1976
  (
    n1949,
    n792,
    n689,
    n1424,
    n1316
  );


  and
  g1977
  (
    n1911,
    n1347,
    n1441,
    n1085,
    n1094
  );


  xnor
  g1978
  (
    n2068,
    n1048,
    n1425,
    n743,
    n1411
  );


  and
  g1979
  (
    n1912,
    n1319,
    n1125,
    n1482,
    n1410
  );


  or
  g1980
  (
    n1879,
    n1259,
    n995,
    n1072,
    n849
  );


  and
  g1981
  (
    n1956,
    n953,
    n668,
    n868,
    n1252
  );


  xnor
  g1982
  (
    n2000,
    n1465,
    n1369,
    n1153,
    n1358
  );


  and
  g1983
  (
    n2009,
    n761,
    n949,
    n848,
    n1362
  );


  nor
  g1984
  (
    n1877,
    n839,
    n789,
    n907,
    n1405
  );


  nor
  g1985
  (
    n2008,
    n1034,
    n772,
    n939,
    n1349
  );


  or
  g1986
  (
    n1928,
    n899,
    n808,
    n873,
    n1004
  );


  xnor
  g1987
  (
    n2019,
    n1218,
    n1452,
    n1134,
    n843
  );


  xnor
  g1988
  (
    n2034,
    n821,
    n1384,
    n979,
    n917
  );


  and
  g1989
  (
    n2060,
    n1070,
    n1055,
    n987,
    n799
  );


  xnor
  g1990
  (
    n1990,
    n879,
    n1201,
    n720,
    n951
  );


  nor
  g1991
  (
    n1919,
    n982,
    n1043,
    n1280,
    n781
  );


  or
  g1992
  (
    n2046,
    n1140,
    n865,
    n1021,
    n960
  );


  and
  g1993
  (
    n1960,
    n1193,
    n1357,
    n1383,
    n707
  );


  nand
  g1994
  (
    n1964,
    n1365,
    n1036,
    n902,
    n1001
  );


  nor
  g1995
  (
    n1933,
    n1175,
    n1295,
    n1170,
    n1166
  );


  nand
  g1996
  (
    n1950,
    n665,
    n1168,
    n887,
    n1205
  );


  xnor
  g1997
  (
    n1983,
    n1407,
    n1233,
    n791,
    n1184
  );


  xor
  g1998
  (
    n2049,
    n893,
    n1138,
    n1442,
    n1122
  );


  nand
  g1999
  (
    n1872,
    n1260,
    n1228,
    n1416,
    n1073
  );


  xor
  g2000
  (
    n1885,
    n883,
    n1486,
    n776,
    n922
  );


  xnor
  g2001
  (
    n2058,
    n1038,
    n1141,
    n1088,
    n1129
  );


  and
  g2002
  (
    n1893,
    n1151,
    n1367,
    n1028,
    n1419
  );


  xor
  g2003
  (
    n1934,
    n1496,
    n1018,
    n675,
    n794
  );


  xor
  g2004
  (
    n1993,
    n1128,
    n1156,
    n705,
    n941
  );


  nor
  g2005
  (
    n2031,
    n719,
    n1029,
    n1448,
    n1157
  );


  or
  g2006
  (
    n1973,
    n1058,
    n1323,
    n1060,
    n968
  );


  and
  g2007
  (
    n1959,
    n1196,
    n1275,
    n1381,
    n1223
  );


  nor
  g2008
  (
    n2037,
    n1389,
    n746,
    n806,
    n1480
  );


  nor
  g2009
  (
    n2023,
    n923,
    n695,
    n1346,
    n724
  );


  xor
  g2010
  (
    n1951,
    n1376,
    n683,
    n1238,
    n1067
  );


  and
  g2011
  (
    n1966,
    n847,
    n754,
    n1112,
    n788
  );


  nor
  g2012
  (
    n2073,
    n1211,
    n715,
    n1179,
    n870
  );


  and
  g2013
  (
    n2033,
    n885,
    n1459,
    n1378,
    n1321
  );


  or
  g2014
  (
    n1927,
    n1291,
    n1400,
    n1350,
    n1288
  );


  xor
  g2015
  (
    n1889,
    n1173,
    n1277,
    n1360,
    n758
  );


  and
  g2016
  (
    n2055,
    n1108,
    n1076,
    n1186,
    n1015
  );


  nor
  g2017
  (
    n2053,
    n1221,
    n1478,
    n1281,
    n877
  );


  nand
  g2018
  (
    n1874,
    n1082,
    n1097,
    n844,
    n1135
  );


  xor
  g2019
  (
    n1944,
    n892,
    n1429,
    n1390,
    n716
  );


  and
  g2020
  (
    n1903,
    n801,
    n741,
    n1341,
    n771
  );


  xnor
  g2021
  (
    n2064,
    n1308,
    n867,
    n921,
    n1136
  );


  nor
  g2022
  (
    n2065,
    n1118,
    n1045,
    n1143,
    n1385
  );


  nor
  g2023
  (
    n2006,
    n1247,
    n1204,
    n1086,
    n1115
  );


  and
  g2024
  (
    n2032,
    n738,
    n1285,
    n1206,
    n729
  );


  or
  g2025
  (
    n1875,
    n1364,
    n762,
    n909,
    n850
  );


  and
  g2026
  (
    n1991,
    n711,
    n966,
    n1430,
    n1130
  );


  and
  g2027
  (
    n1938,
    n832,
    n884,
    n1471,
    n993
  );


  or
  g2028
  (
    n1953,
    n1220,
    n1154,
    n737,
    n1124
  );


  or
  g2029
  (
    n2048,
    n733,
    n1023,
    n1494,
    n696
  );


  and
  g2030
  (
    n2003,
    n670,
    n1210,
    n1016,
    n928
  );


  nor
  g2031
  (
    n1897,
    n1104,
    n985,
    n688,
    n1171
  );


  and
  g2032
  (
    n1932,
    n1302,
    n1147,
    n944,
    n1272
  );


  or
  g2033
  (
    n2069,
    n805,
    n1037,
    n1100,
    n896
  );


  and
  g2034
  (
    n1941,
    n1189,
    n835,
    n1161,
    n924
  );


  and
  g2035
  (
    n1921,
    n1080,
    n1445,
    n1490,
    n1312
  );


  xnor
  g2036
  (
    n1926,
    n1116,
    n1353,
    n1310,
    n863
  );


  nand
  g2037
  (
    n2016,
    n816,
    n751,
    n1208,
    n888
  );


  nand
  g2038
  (
    n2075,
    n946,
    n971,
    n1279,
    n824
  );


  or
  g2039
  (
    n1970,
    n1212,
    n1095,
    n1421,
    n783
  );


  xnor
  g2040
  (
    n2062,
    n1219,
    n992,
    n1479,
    n812
  );


  and
  g2041
  (
    n1883,
    n1133,
    n825,
    n1377,
    n1013
  );


  and
  g2042
  (
    n1906,
    n1231,
    n1330,
    n1200,
    n1418
  );


  or
  g2043
  (
    n1930,
    n1270,
    n1495,
    n1477,
    n927
  );


  xor
  g2044
  (
    n1922,
    n851,
    n1332,
    n671,
    n1081
  );


  and
  g2045
  (
    n2070,
    n1190,
    n1447,
    n1375,
    n735
  );


  nor
  g2046
  (
    n2112,
    n1523,
    n1987
  );


  xnor
  g2047
  (
    n2101,
    n1970,
    n1930,
    n1906,
    n1947
  );


  or
  g2048
  (
    n2113,
    n1916,
    n1914,
    n1886,
    n1997
  );


  nand
  g2049
  (
    n2097,
    n1907,
    n1932,
    n2002,
    n1893
  );


  nor
  g2050
  (
    n2121,
    n1931,
    n1954,
    n1961,
    n1502
  );


  or
  g2051
  (
    n2088,
    n1887,
    n1876,
    n1875,
    n1955
  );


  or
  g2052
  (
    n2082,
    n1927,
    n1950,
    n1964,
    n1873
  );


  xnor
  g2053
  (
    n2109,
    n1943,
    n1968,
    n1963,
    n1958
  );


  xnor
  g2054
  (
    n2079,
    n1911,
    n2011,
    n1908,
    n1497
  );


  or
  g2055
  (
    n2110,
    n1872,
    n2008,
    n1976,
    n2009
  );


  nor
  g2056
  (
    n2083,
    n1915,
    n1500,
    n1939,
    n1888
  );


  nand
  g2057
  (
    n2080,
    n1903,
    n1882,
    n1501,
    n1510
  );


  nand
  g2058
  (
    n2111,
    n1509,
    n2012,
    n1919,
    n1986
  );


  xor
  g2059
  (
    n2085,
    n1877,
    n1994,
    n1996,
    n2006
  );


  xor
  g2060
  (
    n2103,
    n1965,
    n1973,
    n1953,
    n1917
  );


  and
  g2061
  (
    n2084,
    n1979,
    n1514,
    n1940,
    n1505
  );


  xnor
  g2062
  (
    n2086,
    n1522,
    n1900,
    n1972,
    n1896
  );


  xor
  g2063
  (
    n2118,
    n1913,
    n1895,
    n1946,
    n1974
  );


  and
  g2064
  (
    n2096,
    n1881,
    n1934,
    n1993,
    n1982
  );


  xor
  g2065
  (
    n2120,
    n1520,
    n1515,
    n1519,
    n1948
  );


  nor
  g2066
  (
    n2104,
    n2000,
    n1909,
    n1524,
    n1902
  );


  xor
  g2067
  (
    n2081,
    n1905,
    n1945,
    n1518,
    n1525
  );


  or
  g2068
  (
    n2108,
    n1526,
    n1962,
    n1508,
    n1923
  );


  and
  g2069
  (
    n2122,
    n1960,
    n1999,
    n1504,
    n1924
  );


  xor
  g2070
  (
    n2099,
    n1527,
    n1951,
    n1897,
    n1922
  );


  xnor
  g2071
  (
    n2095,
    n1984,
    n1498,
    n1894,
    n1891
  );


  and
  g2072
  (
    n2115,
    n1991,
    n1938,
    n1884,
    n1899
  );


  xor
  g2073
  (
    n2119,
    n1977,
    n1998,
    n1507,
    n1921
  );


  and
  g2074
  (
    n2114,
    n1918,
    n1517,
    n1995,
    n1901
  );


  and
  g2075
  (
    n2100,
    n1942,
    n1949,
    n1925,
    n1521
  );


  and
  g2076
  (
    n2106,
    n1983,
    n1499,
    n1898,
    n1966
  );


  and
  g2077
  (
    n2116,
    n1883,
    n2005,
    n2004,
    n1513
  );


  nor
  g2078
  (
    n2093,
    n1885,
    n1969,
    n1989,
    n1910
  );


  or
  g2079
  (
    n2090,
    n1516,
    n1959,
    n1912,
    n1952
  );


  or
  g2080
  (
    n2117,
    n1511,
    n1957,
    n1920,
    n1941
  );


  and
  g2081
  (
    n2107,
    n1512,
    n1904,
    n1937,
    n1506
  );


  xnor
  g2082
  (
    n2091,
    n1936,
    n1878,
    n1944,
    n1929
  );


  or
  g2083
  (
    n2098,
    n1928,
    n1503,
    n2013,
    n1935
  );


  nand
  g2084
  (
    n2089,
    n1992,
    n2001,
    n1889,
    n1880
  );


  nor
  g2085
  (
    n2102,
    n1874,
    n1879,
    n2007,
    n1871
  );


  xnor
  g2086
  (
    n2094,
    n2010,
    n1892,
    n1967,
    n1988
  );


  and
  g2087
  (
    n2092,
    n1981,
    n1980,
    n1978,
    n1956
  );


  xor
  g2088
  (
    n2087,
    n1933,
    n1971,
    n1890,
    n1990
  );


  or
  g2089
  (
    n2105,
    n2003,
    n1985,
    n1975,
    n1926
  );


  buf
  g2090
  (
    n2129,
    n2119
  );


  buf
  g2091
  (
    n2123,
    n2106
  );


  not
  g2092
  (
    n2147,
    n1550
  );


  not
  g2093
  (
    n2132,
    n2120
  );


  not
  g2094
  (
    n2135,
    n1541
  );


  not
  g2095
  (
    n2145,
    n1559
  );


  buf
  g2096
  (
    n2149,
    n1534
  );


  not
  g2097
  (
    n2146,
    n1532
  );


  not
  g2098
  (
    n2140,
    n2107
  );


  buf
  g2099
  (
    n2152,
    n1564
  );


  not
  g2100
  (
    n2150,
    n1546
  );


  nor
  g2101
  (
    n2142,
    n1543,
    n2112,
    n1549
  );


  nand
  g2102
  (
    n2148,
    n1535,
    n1539,
    n2114
  );


  nand
  g2103
  (
    n2141,
    n1555,
    n1533,
    n1558
  );


  nor
  g2104
  (
    n2139,
    n2096,
    n2099,
    n2094
  );


  and
  g2105
  (
    n2136,
    n2122,
    n1529,
    n1547
  );


  xor
  g2106
  (
    n2138,
    n2105,
    n1553,
    n2115
  );


  xor
  g2107
  (
    n2127,
    n1562,
    n2116,
    n1566
  );


  or
  g2108
  (
    n2124,
    n2121,
    n1540,
    n1528
  );


  and
  g2109
  (
    n2131,
    n1561,
    n1537,
    n2102
  );


  nand
  g2110
  (
    n2134,
    n2097,
    n1544,
    n2093
  );


  or
  g2111
  (
    n2128,
    n2118,
    n2108,
    n2111
  );


  nor
  g2112
  (
    n2151,
    n2113,
    n2101,
    n2110
  );


  or
  g2113
  (
    n2130,
    n2100,
    n1552,
    n1530
  );


  nor
  g2114
  (
    n2137,
    n2103,
    n1560,
    n1565
  );


  or
  g2115
  (
    n2143,
    n1538,
    n2104,
    n1542
  );


  nor
  g2116
  (
    n2125,
    n1551,
    n2117,
    n1536
  );


  xor
  g2117
  (
    n2144,
    n1545,
    n1568,
    n1563,
    n1531
  );


  and
  g2118
  (
    n2126,
    n1557,
    n1556,
    n2098,
    n1567
  );


  or
  g2119
  (
    n2133,
    n1554,
    n2109,
    n2095,
    n1548
  );


  xor
  g2120
  (
    n2161,
    n1573,
    n2123,
    n1593
  );


  or
  g2121
  (
    n2156,
    n1585,
    n1576,
    n1589,
    n1598
  );


  xor
  g2122
  (
    n2155,
    n2123,
    n1587,
    n2125,
    n2124
  );


  and
  g2123
  (
    n2160,
    n1586,
    n2125,
    n1596,
    n1591
  );


  xnor
  g2124
  (
    n2157,
    n1570,
    n1569,
    n2123,
    n2124
  );


  nand
  g2125
  (
    n2159,
    n1584,
    n1580,
    n1595,
    n1572
  );


  or
  g2126
  (
    n2158,
    n1579,
    n1594,
    n1574,
    n1597
  );


  nand
  g2127
  (
    n2162,
    n1575,
    n1577,
    n1588,
    n2124
  );


  xnor
  g2128
  (
    n2154,
    n1582,
    n1590,
    n1581,
    n1578
  );


  and
  g2129
  (
    n2153,
    n1571,
    n1583,
    n1592,
    n2124
  );


  buf
  g2130
  (
    n2163,
    n2153
  );


  buf
  g2131
  (
    n2164,
    n2163
  );


  buf
  g2132
  (
    n2165,
    n2163
  );


  buf
  g2133
  (
    n2166,
    n2163
  );


  buf
  g2134
  (
    n2168,
    n2164
  );


  buf
  g2135
  (
    n2167,
    n2164
  );


  nand
  g2136
  (
    n2169,
    n1600,
    n1599,
    n1601,
    n2167
  );


  not
  g2137
  (
    n2170,
    n2169
  );


  buf
  g2138
  (
    n2171,
    n2169
  );


  xnor
  g2139
  (
    n2176,
    n1604,
    n2170
  );


  or
  g2140
  (
    n2172,
    n1612,
    n1603
  );


  or
  g2141
  (
    n2174,
    n2170,
    n1611,
    n1608,
    n1607
  );


  xnor
  g2142
  (
    n2175,
    n1606,
    n1602,
    n2170,
    n2171
  );


  xnor
  g2143
  (
    n2173,
    n1609,
    n1605,
    n1610,
    n2170
  );


  xnor
  g2144
  (
    n2178,
    n1645,
    n1642,
    n1636,
    n2172
  );


  xor
  g2145
  (
    n2188,
    n1620,
    n1616,
    n1637,
    n1622
  );


  xor
  g2146
  (
    n2190,
    n1630,
    n2174,
    n1633,
    n1657
  );


  nand
  g2147
  (
    n2186,
    n2175,
    n1631,
    n1656,
    n1648
  );


  xor
  g2148
  (
    n2180,
    n1640,
    n1627,
    n1613,
    n2173
  );


  nand
  g2149
  (
    n2187,
    n1652,
    n1650,
    n1632,
    n2173
  );


  and
  g2150
  (
    n2185,
    n2175,
    n2174,
    n1644,
    n1641
  );


  and
  g2151
  (
    n2189,
    n1653,
    n1639,
    n1647,
    n1619
  );


  xor
  g2152
  (
    n2182,
    n1618,
    n1643,
    n2173,
    n1614
  );


  nand
  g2153
  (
    n2179,
    n1649,
    n1628,
    n1638,
    n2174
  );


  xnor
  g2154
  (
    n2183,
    n2173,
    n1651,
    n1655,
    n1624
  );


  xnor
  g2155
  (
    n2181,
    n1629,
    n2172,
    n1634,
    n1625
  );


  or
  g2156
  (
    n2191,
    n1626,
    n1646,
    n2172,
    n1623
  );


  and
  g2157
  (
    n2177,
    n2172,
    n2175,
    n2174,
    n1617
  );


  or
  g2158
  (
    n2184,
    n1635,
    n1621,
    n1615,
    n1654
  );


  buf
  g2159
  (
    n2224,
    n2041
  );


  buf
  g2160
  (
    n2235,
    n2184
  );


  not
  g2161
  (
    n2217,
    n2038
  );


  not
  g2162
  (
    n2232,
    n2186
  );


  buf
  g2163
  (
    n2199,
    n2182
  );


  buf
  g2164
  (
    n2196,
    n2040
  );


  buf
  g2165
  (
    n2193,
    n2188
  );


  not
  g2166
  (
    n2212,
    n1660
  );


  buf
  g2167
  (
    n2205,
    n2191
  );


  not
  g2168
  (
    n2222,
    n1662
  );


  buf
  g2169
  (
    n2210,
    n2019
  );


  not
  g2170
  (
    n2238,
    n2033
  );


  buf
  g2171
  (
    n2214,
    n2186
  );


  buf
  g2172
  (
    n2227,
    n2188
  );


  not
  g2173
  (
    n2192,
    n2183
  );


  not
  g2174
  (
    n2202,
    n2021
  );


  not
  g2175
  (
    n2207,
    n2025
  );


  not
  g2176
  (
    n2213,
    n2184
  );


  buf
  g2177
  (
    n2230,
    n2187
  );


  buf
  g2178
  (
    n2206,
    n2185
  );


  not
  g2179
  (
    n2211,
    n2187
  );


  buf
  g2180
  (
    n2226,
    n2188
  );


  buf
  g2181
  (
    n2201,
    n2039
  );


  buf
  g2182
  (
    n2239,
    n2032
  );


  not
  g2183
  (
    n2218,
    n2185
  );


  not
  g2184
  (
    n2229,
    n2027
  );


  not
  g2185
  (
    n2216,
    n2178
  );


  not
  g2186
  (
    n2195,
    n2185
  );


  not
  g2187
  (
    n2209,
    n2182
  );


  not
  g2188
  (
    n2228,
    n2183
  );


  not
  g2189
  (
    n2204,
    n2183
  );


  not
  g2190
  (
    n2194,
    n1659
  );


  not
  g2191
  (
    n2236,
    n2020
  );


  not
  g2192
  (
    n2200,
    n2018
  );


  not
  g2193
  (
    n2225,
    n2037
  );


  buf
  g2194
  (
    n2198,
    n2177
  );


  or
  g2195
  (
    n2220,
    n2181,
    n2181,
    n2017,
    n2028
  );


  nand
  g2196
  (
    n2203,
    n2029,
    n2184,
    n2034,
    n2190
  );


  xor
  g2197
  (
    n2231,
    n2187,
    n2026,
    n1661,
    n2023
  );


  or
  g2198
  (
    n2208,
    n2189,
    n2044,
    n2190
  );


  and
  g2199
  (
    n2215,
    n2014,
    n2180,
    n2030,
    n2181
  );


  xor
  g2200
  (
    n2237,
    n2186,
    n2191,
    n2022,
    n2189
  );


  xor
  g2201
  (
    n2197,
    n2179,
    n2189,
    n2185,
    n2035
  );


  and
  g2202
  (
    n2223,
    n2186,
    n2188,
    n2031,
    n2015
  );


  or
  g2203
  (
    n2233,
    n2182,
    n2182,
    n2024,
    n2183
  );


  nand
  g2204
  (
    n2219,
    n2189,
    n2191,
    n2043,
    n2016
  );


  or
  g2205
  (
    n2234,
    n2042,
    n2191,
    n1658,
    n2036
  );


  or
  g2206
  (
    n2221,
    n2187,
    n2181,
    n2184,
    n2190
  );


  not
  g2207
  (
    n2378,
    n2214
  );


  not
  g2208
  (
    n2358,
    n2129
  );


  not
  g2209
  (
    n2262,
    n2200
  );


  not
  g2210
  (
    n2368,
    n2136
  );


  buf
  g2211
  (
    n2314,
    n2147
  );


  buf
  g2212
  (
    n2281,
    n2213
  );


  not
  g2213
  (
    n2252,
    n1670
  );


  not
  g2214
  (
    n2316,
    n2146
  );


  not
  g2215
  (
    n2332,
    n2209
  );


  buf
  g2216
  (
    n2406,
    n2224
  );


  not
  g2217
  (
    n2244,
    n2142
  );


  buf
  g2218
  (
    n2359,
    n2144
  );


  buf
  g2219
  (
    n2257,
    n2217
  );


  buf
  g2220
  (
    n2404,
    n2128
  );


  buf
  g2221
  (
    n2256,
    n2225
  );


  not
  g2222
  (
    n2301,
    n2200
  );


  not
  g2223
  (
    n2347,
    n2131
  );


  not
  g2224
  (
    n2280,
    n2151
  );


  buf
  g2225
  (
    n2289,
    n2234
  );


  buf
  g2226
  (
    n2299,
    n2132
  );


  buf
  g2227
  (
    n2381,
    n2222
  );


  buf
  g2228
  (
    n2421,
    n2232
  );


  buf
  g2229
  (
    n2428,
    n2215
  );


  buf
  g2230
  (
    n2330,
    n2149
  );


  not
  g2231
  (
    n2350,
    n1669
  );


  buf
  g2232
  (
    n2339,
    n2147
  );


  not
  g2233
  (
    n2279,
    n2223
  );


  not
  g2234
  (
    n2354,
    n2142
  );


  buf
  g2235
  (
    n2411,
    n2143
  );


  not
  g2236
  (
    n2352,
    n2236
  );


  buf
  g2237
  (
    n2310,
    n2210
  );


  buf
  g2238
  (
    n2304,
    n2144
  );


  not
  g2239
  (
    n2284,
    n2211
  );


  buf
  g2240
  (
    n2265,
    n2208
  );


  buf
  g2241
  (
    n2372,
    n2148
  );


  not
  g2242
  (
    n2349,
    n2216
  );


  not
  g2243
  (
    n2241,
    n2233
  );


  buf
  g2244
  (
    n2313,
    n2146
  );


  not
  g2245
  (
    n2306,
    n2221
  );


  not
  g2246
  (
    n2401,
    n2228
  );


  buf
  g2247
  (
    n2371,
    n2202
  );


  not
  g2248
  (
    n2373,
    n2131
  );


  buf
  g2249
  (
    n2375,
    n2229
  );


  not
  g2250
  (
    n2245,
    n2222
  );


  buf
  g2251
  (
    n2335,
    n2223
  );


  not
  g2252
  (
    n2282,
    n2136
  );


  not
  g2253
  (
    n2324,
    n2209
  );


  buf
  g2254
  (
    n2308,
    n2213
  );


  not
  g2255
  (
    n2278,
    n2149
  );


  not
  g2256
  (
    n2402,
    n2137
  );


  buf
  g2257
  (
    n2248,
    n2216
  );


  buf
  g2258
  (
    n2361,
    n2126
  );


  not
  g2259
  (
    n2420,
    n2233
  );


  buf
  g2260
  (
    n2276,
    n2136
  );


  not
  g2261
  (
    n2261,
    n2237
  );


  buf
  g2262
  (
    n2283,
    n2225
  );


  not
  g2263
  (
    n2394,
    n2203
  );


  buf
  g2264
  (
    n2321,
    n2237
  );


  buf
  g2265
  (
    n2254,
    n2231
  );


  not
  g2266
  (
    n2398,
    n2140
  );


  not
  g2267
  (
    n2247,
    n2150
  );


  buf
  g2268
  (
    n2318,
    n2230
  );


  not
  g2269
  (
    n2385,
    n2148
  );


  not
  g2270
  (
    n2382,
    n2195
  );


  not
  g2271
  (
    n2274,
    n1665
  );


  not
  g2272
  (
    n2386,
    n2203
  );


  buf
  g2273
  (
    n2425,
    n2138
  );


  not
  g2274
  (
    n2342,
    n2234
  );


  buf
  g2275
  (
    n2374,
    n2224
  );


  buf
  g2276
  (
    n2240,
    n2215
  );


  buf
  g2277
  (
    n2391,
    n2221
  );


  buf
  g2278
  (
    n2414,
    n2134
  );


  buf
  g2279
  (
    n2267,
    n2203
  );


  buf
  g2280
  (
    n2343,
    n2125
  );


  not
  g2281
  (
    n2333,
    n2206
  );


  not
  g2282
  (
    n2380,
    n2127
  );


  buf
  g2283
  (
    n2345,
    n2204
  );


  not
  g2284
  (
    n2360,
    n2138
  );


  buf
  g2285
  (
    n2426,
    n2141
  );


  not
  g2286
  (
    n2334,
    n2125
  );


  buf
  g2287
  (
    n2258,
    n2144
  );


  buf
  g2288
  (
    n2326,
    n2196
  );


  not
  g2289
  (
    n2251,
    n2128
  );


  not
  g2290
  (
    n2407,
    n2194
  );


  buf
  g2291
  (
    n2430,
    n2215
  );


  buf
  g2292
  (
    n2364,
    n1663
  );


  buf
  g2293
  (
    n2270,
    n2218
  );


  not
  g2294
  (
    n2341,
    n2239
  );


  buf
  g2295
  (
    n2396,
    n2218
  );


  buf
  g2296
  (
    n2250,
    n2197
  );


  not
  g2297
  (
    n2388,
    n2210
  );


  not
  g2298
  (
    n2295,
    n2150
  );


  not
  g2299
  (
    n2323,
    n2147
  );


  not
  g2300
  (
    n2246,
    n2212
  );


  buf
  g2301
  (
    n2379,
    n2192
  );


  not
  g2302
  (
    n2410,
    n2136
  );


  not
  g2303
  (
    n2331,
    n2201
  );


  buf
  g2304
  (
    n2336,
    n2225
  );


  not
  g2305
  (
    n2431,
    n2211
  );


  not
  g2306
  (
    n2303,
    n2207
  );


  not
  g2307
  (
    n2292,
    n2198
  );


  buf
  g2308
  (
    n2325,
    n2227
  );


  not
  g2309
  (
    n2285,
    n2233
  );


  buf
  g2310
  (
    n2312,
    n2140
  );


  buf
  g2311
  (
    n2287,
    n2198
  );


  buf
  g2312
  (
    n2348,
    n2209
  );


  not
  g2313
  (
    n2387,
    n2226
  );


  not
  g2314
  (
    n2424,
    n2206
  );


  not
  g2315
  (
    n2357,
    n2142
  );


  buf
  g2316
  (
    n2255,
    n1667
  );


  not
  g2317
  (
    n2400,
    n2195
  );


  not
  g2318
  (
    n2363,
    n2129
  );


  not
  g2319
  (
    n2418,
    n2230
  );


  not
  g2320
  (
    n2242,
    n2141
  );


  not
  g2321
  (
    n2302,
    n2230
  );


  not
  g2322
  (
    n2290,
    n2139
  );


  buf
  g2323
  (
    n2297,
    n2148
  );


  buf
  g2324
  (
    n2367,
    n2228
  );


  not
  g2325
  (
    n2293,
    n2221
  );


  not
  g2326
  (
    n2413,
    n2148
  );


  not
  g2327
  (
    n2416,
    n2194
  );


  not
  g2328
  (
    n2291,
    n2239
  );


  buf
  g2329
  (
    n2305,
    n2134
  );


  not
  g2330
  (
    n2403,
    n2204
  );


  buf
  g2331
  (
    n2307,
    n2146
  );


  buf
  g2332
  (
    n2337,
    n2132
  );


  not
  g2333
  (
    n2329,
    n2201
  );


  not
  g2334
  (
    n2275,
    n2201
  );


  not
  g2335
  (
    n2365,
    n2205
  );


  not
  g2336
  (
    n2429,
    n2227
  );


  not
  g2337
  (
    n2389,
    n2238
  );


  buf
  g2338
  (
    n2355,
    n2221
  );


  buf
  g2339
  (
    n2263,
    n2139
  );


  not
  g2340
  (
    n2405,
    n2194
  );


  buf
  g2341
  (
    n2393,
    n2231
  );


  not
  g2342
  (
    n2369,
    n2196
  );


  or
  g2343
  (
    n2259,
    n2130,
    n2213,
    n2126
  );


  nand
  g2344
  (
    n2409,
    n2149,
    n2138,
    n2234
  );


  nor
  g2345
  (
    n2427,
    n2228,
    n2139,
    n2212
  );


  xor
  g2346
  (
    n2408,
    n2145,
    n2217,
    n2146
  );


  xor
  g2347
  (
    n2351,
    n2235,
    n2213,
    n2236
  );


  xnor
  g2348
  (
    n2327,
    n2217,
    n2129,
    n1666
  );


  nor
  g2349
  (
    n2412,
    n2223,
    n2126,
    n2235
  );


  nand
  g2350
  (
    n2422,
    n2239,
    n2223,
    n2141
  );


  or
  g2351
  (
    n2286,
    n2216,
    n2197,
    n2209
  );


  xnor
  g2352
  (
    n2260,
    n2138,
    n2214,
    n2199
  );


  nor
  g2353
  (
    n2397,
    n2193,
    n2224,
    n2192
  );


  nand
  g2354
  (
    n2423,
    n2202,
    n2233,
    n2204
  );


  nand
  g2355
  (
    n2269,
    n2237,
    n2201,
    n2199
  );


  xor
  g2356
  (
    n2264,
    n2219,
    n2231,
    n2208
  );


  or
  g2357
  (
    n2315,
    n2200,
    n2210,
    n2199
  );


  xnor
  g2358
  (
    n2272,
    n2229,
    n2130,
    n2207
  );


  xnor
  g2359
  (
    n2288,
    n2214,
    n2228,
    n2198
  );


  xor
  g2360
  (
    n2419,
    n2128,
    n2229,
    n2226
  );


  xor
  g2361
  (
    n2384,
    n2211,
    n2218,
    n2150
  );


  xnor
  g2362
  (
    n2377,
    n2135,
    n2197,
    n2226
  );


  xor
  g2363
  (
    n2266,
    n2132,
    n1664,
    n2220
  );


  or
  g2364
  (
    n2338,
    n2232,
    n2226,
    n2140
  );


  xnor
  g2365
  (
    n2417,
    n2151,
    n2215,
    n2238
  );


  xor
  g2366
  (
    n2356,
    n2133,
    n2137,
    n2127
  );


  nor
  g2367
  (
    n2249,
    n2143,
    n2217,
    n2211
  );


  nor
  g2368
  (
    n2294,
    n2205,
    n2208,
    n2149
  );


  or
  g2369
  (
    n2340,
    n2225,
    n2230,
    n2132
  );


  or
  g2370
  (
    n2320,
    n2137,
    n2130,
    n2231
  );


  nand
  g2371
  (
    n2300,
    n2238,
    n2198,
    n2196
  );


  and
  g2372
  (
    n2395,
    n2145,
    n2133,
    n2207
  );


  xor
  g2373
  (
    n2243,
    n2238,
    n2195,
    n2236
  );


  xnor
  g2374
  (
    n2353,
    n2210,
    n2207,
    n2219
  );


  and
  g2375
  (
    n2399,
    n2143,
    n2212,
    n2144
  );


  or
  g2376
  (
    n2328,
    n2220,
    n2139,
    n2200
  );


  or
  g2377
  (
    n2311,
    n2239,
    n2199,
    n2137
  );


  nand
  g2378
  (
    n2309,
    n2220,
    n2129,
    n2206
  );


  nand
  g2379
  (
    n2362,
    n2135,
    n2232,
    n2206
  );


  or
  g2380
  (
    n2415,
    n2143,
    n2145,
    n2193
  );


  nand
  g2381
  (
    n2298,
    n2145,
    n2204,
    n2194
  );


  xnor
  g2382
  (
    n2296,
    n2140,
    n2212,
    n2147
  );


  nand
  g2383
  (
    n2392,
    n2236,
    n2192,
    n2235
  );


  or
  g2384
  (
    n2366,
    n2134,
    n2222,
    n2235
  );


  nor
  g2385
  (
    n2277,
    n2222,
    n2205,
    n2141
  );


  nor
  g2386
  (
    n2390,
    n2227,
    n2131,
    n2196
  );


  xnor
  g2387
  (
    n2273,
    n2220,
    n2192,
    n2150
  );


  nor
  g2388
  (
    n2383,
    n2232,
    n2219
  );


  and
  g2389
  (
    n2322,
    n2216,
    n2227,
    n2195
  );


  nand
  g2390
  (
    n2370,
    n2130,
    n2135,
    n2214
  );


  and
  g2391
  (
    n2317,
    n2218,
    n2237,
    n2127
  );


  or
  g2392
  (
    n2268,
    n1668,
    n2131,
    n2193
  );


  nor
  g2393
  (
    n2319,
    n2133,
    n2224,
    n2127
  );


  xor
  g2394
  (
    n2344,
    n2193,
    n2234,
    n2135
  );


  and
  g2395
  (
    n2346,
    n2197,
    n2142,
    n2202
  );


  and
  g2396
  (
    n2253,
    n2128,
    n2134,
    n2205
  );


  nand
  g2397
  (
    n2271,
    n2133,
    n2229,
    n2126
  );


  nand
  g2398
  (
    n2376,
    n2208,
    n2202,
    n2203
  );


  not
  g2399
  (
    n2691,
    n2271
  );


  not
  g2400
  (
    n2554,
    n2361
  );


  buf
  g2401
  (
    n2533,
    n1671
  );


  buf
  g2402
  (
    n2577,
    n2429
  );


  not
  g2403
  (
    n2612,
    n2329
  );


  buf
  g2404
  (
    n2499,
    n2326
  );


  buf
  g2405
  (
    n2607,
    n2364
  );


  buf
  g2406
  (
    n2483,
    n2395
  );


  buf
  g2407
  (
    n2681,
    n2243
  );


  not
  g2408
  (
    n2588,
    n2364
  );


  not
  g2409
  (
    n2509,
    n2302
  );


  buf
  g2410
  (
    n2506,
    n2410
  );


  not
  g2411
  (
    n2538,
    n2278
  );


  not
  g2412
  (
    n2504,
    n2337
  );


  buf
  g2413
  (
    n2470,
    n2295
  );


  buf
  g2414
  (
    n2647,
    n2257
  );


  not
  g2415
  (
    n2702,
    n2346
  );


  buf
  g2416
  (
    n2585,
    n2251
  );


  not
  g2417
  (
    n2675,
    n2322
  );


  buf
  g2418
  (
    n2646,
    n2360
  );


  buf
  g2419
  (
    n2477,
    n2376
  );


  buf
  g2420
  (
    n2476,
    n2317
  );


  not
  g2421
  (
    n2676,
    n2295
  );


  not
  g2422
  (
    n2443,
    n2276
  );


  not
  g2423
  (
    n2463,
    n2280
  );


  buf
  g2424
  (
    n2446,
    n2273
  );


  buf
  g2425
  (
    n2464,
    n2257
  );


  not
  g2426
  (
    n2497,
    n2424
  );


  not
  g2427
  (
    n2621,
    n2394
  );


  buf
  g2428
  (
    n2454,
    n2323
  );


  buf
  g2429
  (
    n2573,
    n2427
  );


  buf
  g2430
  (
    n2677,
    n2280
  );


  not
  g2431
  (
    n2540,
    n2405
  );


  not
  g2432
  (
    n2518,
    n2263
  );


  not
  g2433
  (
    n2479,
    n2422
  );


  buf
  g2434
  (
    n2461,
    n2416
  );


  buf
  g2435
  (
    n2694,
    n2297
  );


  buf
  g2436
  (
    n2629,
    n2404
  );


  not
  g2437
  (
    n2650,
    n2304
  );


  not
  g2438
  (
    n2609,
    n2343
  );


  buf
  g2439
  (
    n2468,
    n2253
  );


  buf
  g2440
  (
    n2571,
    n2289
  );


  buf
  g2441
  (
    n2553,
    n1682
  );


  buf
  g2442
  (
    n2486,
    n2276
  );


  not
  g2443
  (
    n2665,
    n2265
  );


  not
  g2444
  (
    n2433,
    n2389
  );


  buf
  g2445
  (
    n2542,
    n2322
  );


  not
  g2446
  (
    n2682,
    n2342
  );


  not
  g2447
  (
    n2439,
    n2303
  );


  buf
  g2448
  (
    n2654,
    n2373
  );


  buf
  g2449
  (
    n2556,
    n2268
  );


  not
  g2450
  (
    n2572,
    n2273
  );


  buf
  g2451
  (
    n2586,
    n2261
  );


  not
  g2452
  (
    n2482,
    n2301
  );


  not
  g2453
  (
    n2597,
    n2262
  );


  buf
  g2454
  (
    n2467,
    n2306
  );


  buf
  g2455
  (
    n2655,
    n2385
  );


  not
  g2456
  (
    n2643,
    n2341
  );


  not
  g2457
  (
    n2667,
    n2332
  );


  buf
  g2458
  (
    n2445,
    n2254
  );


  buf
  g2459
  (
    n2594,
    n2305
  );


  buf
  g2460
  (
    n2531,
    n2289
  );


  buf
  g2461
  (
    KeyWire_0_13,
    n2408
  );


  buf
  g2462
  (
    n2434,
    n2272
  );


  buf
  g2463
  (
    n2458,
    n2290
  );


  buf
  g2464
  (
    n2671,
    n2392
  );


  not
  g2465
  (
    n2641,
    n2412
  );


  not
  g2466
  (
    n2590,
    n2348
  );


  buf
  g2467
  (
    n2489,
    n2409
  );


  not
  g2468
  (
    n2537,
    n2255
  );


  not
  g2469
  (
    n2669,
    n2316
  );


  not
  g2470
  (
    n2508,
    n2242
  );


  not
  g2471
  (
    n2605,
    n2403
  );


  not
  g2472
  (
    n2640,
    n2391
  );


  buf
  g2473
  (
    n2440,
    n2267
  );


  buf
  g2474
  (
    n2633,
    n2393
  );


  buf
  g2475
  (
    n2644,
    n2384
  );


  not
  g2476
  (
    n2601,
    n2308
  );


  buf
  g2477
  (
    n2471,
    n2289
  );


  not
  g2478
  (
    n2432,
    n2242
  );


  not
  g2479
  (
    n2611,
    n2348
  );


  not
  g2480
  (
    n2545,
    n2329
  );


  not
  g2481
  (
    n2657,
    n2381
  );


  not
  g2482
  (
    n2539,
    n2297
  );


  buf
  g2483
  (
    n2604,
    n2412
  );


  not
  g2484
  (
    n2466,
    n2421
  );


  not
  g2485
  (
    n2630,
    n2339
  );


  not
  g2486
  (
    n2460,
    n2371
  );


  buf
  g2487
  (
    n2664,
    n2303
  );


  not
  g2488
  (
    n2560,
    n2385
  );


  buf
  g2489
  (
    n2700,
    n2397
  );


  not
  g2490
  (
    n2498,
    n2330
  );


  buf
  g2491
  (
    n2478,
    n2251
  );


  not
  g2492
  (
    n2645,
    n2362
  );


  buf
  g2493
  (
    n2634,
    n2283
  );


  buf
  g2494
  (
    n2503,
    n2429
  );


  not
  g2495
  (
    n2561,
    n2351
  );


  buf
  g2496
  (
    n2473,
    n2405
  );


  nor
  g2497
  (
    n2510,
    n2264,
    n2249,
    n655,
    n2418
  );


  xnor
  g2498
  (
    n2485,
    n2260,
    n2313,
    n2290,
    n2392
  );


  xnor
  g2499
  (
    n2666,
    n2382,
    n2429,
    n2256,
    n2344
  );


  nand
  g2500
  (
    n2622,
    n2285,
    n2298,
    n2262,
    n2331
  );


  nand
  g2501
  (
    n2493,
    n2390,
    n2255,
    n2360,
    n2329
  );


  and
  g2502
  (
    n2521,
    n2350,
    n2383,
    n2375,
    n2334
  );


  xnor
  g2503
  (
    n2557,
    n2373,
    n2384,
    n2254,
    n2319
  );


  or
  g2504
  (
    n2680,
    n2283,
    n2391,
    n2345,
    n2325
  );


  xor
  g2505
  (
    n2505,
    n2427,
    n2309,
    n2381,
    n2262
  );


  nand
  g2506
  (
    n2444,
    n2247,
    n2408,
    n2250,
    n2396
  );


  xor
  g2507
  (
    n2673,
    n2301,
    n2295,
    n2245,
    n2240
  );


  nand
  g2508
  (
    n2579,
    n2296,
    n2269,
    n2426,
    n2318
  );


  xor
  g2509
  (
    n2481,
    n2277,
    n2286,
    n2268,
    n2347
  );


  xnor
  g2510
  (
    n2547,
    n2318,
    n2268,
    n2328,
    n2305
  );


  and
  g2511
  (
    n2462,
    n2302,
    n2294,
    n2335,
    n2282
  );


  xnor
  g2512
  (
    n2626,
    n2328,
    n2341,
    n2420,
    n2271
  );


  xnor
  g2513
  (
    n2610,
    n2306,
    n2310,
    n2256,
    n2361
  );


  xnor
  g2514
  (
    n2490,
    n2395,
    n2257,
    n2423,
    n2258
  );


  or
  g2515
  (
    n2628,
    n2351,
    n2384,
    n2352,
    n2345
  );


  xor
  g2516
  (
    n2514,
    n2323,
    n2361,
    n2352,
    n2401
  );


  nand
  g2517
  (
    n2501,
    n2324,
    n2404,
    n2307,
    n2311
  );


  xor
  g2518
  (
    n2492,
    n2317,
    n2377,
    n2367,
    n2411
  );


  nor
  g2519
  (
    n2566,
    n2339,
    n2400,
    n2313,
    n2419
  );


  nand
  g2520
  (
    n2529,
    n2356,
    n2293,
    n2374,
    n2304
  );


  xor
  g2521
  (
    n2496,
    n2336,
    n2312,
    n2252,
    n2417
  );


  nor
  g2522
  (
    n2550,
    n655,
    n2354,
    n656,
    n2387
  );


  xor
  g2523
  (
    n2686,
    n657,
    n2375,
    n2290,
    n2427
  );


  and
  g2524
  (
    n2692,
    n2365,
    n2279,
    n2369,
    n2302
  );


  or
  g2525
  (
    n2652,
    n2377,
    n2376,
    n2399,
    n2420
  );


  xnor
  g2526
  (
    n2639,
    n2365,
    n2372,
    n2309,
    n2403
  );


  or
  g2527
  (
    n2638,
    n2426,
    n2353,
    n2247,
    n2367
  );


  or
  g2528
  (
    n2624,
    n2336,
    n2345,
    n2299,
    n2241
  );


  nand
  g2529
  (
    n2581,
    n2176,
    n2269,
    n2379,
    n2383
  );


  xor
  g2530
  (
    n2599,
    n2356,
    n2261,
    n2346,
    n2315
  );


  nor
  g2531
  (
    n2447,
    n2388,
    n2303,
    n2335,
    n2416
  );


  nor
  g2532
  (
    n2526,
    n656,
    n2332,
    n2331,
    n2257
  );


  nor
  g2533
  (
    n2578,
    n2369,
    n2279,
    n2326,
    n2410
  );


  xnor
  g2534
  (
    n2457,
    n2306,
    n2251,
    n2314,
    n2285
  );


  xor
  g2535
  (
    n2491,
    n2368,
    n2306,
    n2409,
    n2381
  );


  and
  g2536
  (
    n2649,
    n2390,
    n2270,
    n2294,
    n2176
  );


  xnor
  g2537
  (
    n2635,
    n2413,
    n2419,
    n2320,
    n2275
  );


  or
  g2538
  (
    n2475,
    n2278,
    n2422,
    n2358,
    n2248
  );


  xor
  g2539
  (
    n2683,
    n2259,
    n2412,
    n2328,
    n2418
  );


  xnor
  g2540
  (
    n2519,
    n2259,
    n2249,
    n2250,
    n2381
  );


  nor
  g2541
  (
    n2502,
    n2425,
    n2315,
    n2313,
    n2284
  );


  and
  g2542
  (
    n2661,
    n2351,
    n1681,
    n2415,
    n2247
  );


  and
  g2543
  (
    n2651,
    n2350,
    n2365,
    n2272,
    n2340
  );


  xnor
  g2544
  (
    n2688,
    n2388,
    n2407,
    n2273,
    n2309
  );


  or
  g2545
  (
    n2699,
    n2318,
    n2253,
    n2305,
    n2284
  );


  xnor
  g2546
  (
    n2484,
    n2314,
    n2406,
    n2401,
    n2291
  );


  xor
  g2547
  (
    n2695,
    n2330,
    n2398,
    n2360,
    n2349
  );


  xnor
  g2548
  (
    n2619,
    n2371,
    n2408,
    n2287,
    n2364
  );


  nor
  g2549
  (
    n2441,
    n2398,
    n2263,
    n2255,
    n2249
  );


  xor
  g2550
  (
    n2679,
    n2345,
    n2277,
    n2260,
    n2382
  );


  or
  g2551
  (
    n2528,
    n2343,
    n2363,
    n2273,
    n2400
  );


  nor
  g2552
  (
    n2552,
    n2382,
    n2349,
    n2317,
    n2368
  );


  nor
  g2553
  (
    n2564,
    n2332,
    n1679,
    n2372,
    n2414
  );


  xnor
  g2554
  (
    n2642,
    n2280,
    n2398,
    n2251,
    n2283
  );


  and
  g2555
  (
    n2690,
    n2357,
    n2312,
    n2396,
    n2418
  );


  xnor
  g2556
  (
    n2534,
    n2308,
    n2355,
    n2311,
    n2416
  );


  or
  g2557
  (
    n2555,
    n2335,
    n2240,
    n2367,
    n2322
  );


  and
  g2558
  (
    n2696,
    n2321,
    n2423,
    n2387,
    n2354
  );


  nand
  g2559
  (
    n2449,
    n2378,
    n2292,
    n2308,
    n2364
  );


  nor
  g2560
  (
    n2659,
    n2415,
    n2326,
    n2366,
    n2265
  );


  xor
  g2561
  (
    n2516,
    n2384,
    n2279,
    n2175,
    n2259
  );


  nor
  g2562
  (
    n2697,
    n2262,
    n2275,
    n2418,
    n2248
  );


  nand
  g2563
  (
    n2636,
    n2417,
    n2347,
    n2324,
    n2366
  );


  xor
  g2564
  (
    n2522,
    n656,
    n2366,
    n2327,
    n2417
  );


  xor
  g2565
  (
    n2631,
    n2245,
    n2344,
    n2243,
    n2320
  );


  or
  g2566
  (
    n2495,
    n2339,
    n656,
    n2430,
    n2420
  );


  xor
  g2567
  (
    n2563,
    n2299,
    n2410,
    n2281,
    n2375
  );


  nand
  g2568
  (
    n2625,
    n2380,
    n2285,
    n2265,
    n2370
  );


  xor
  g2569
  (
    n2544,
    n2407,
    n2281,
    n2356,
    n2403
  );


  and
  g2570
  (
    n2623,
    n2404,
    n2292,
    n2367,
    n2379
  );


  xor
  g2571
  (
    n2451,
    n2419,
    n2356,
    n2369,
    n2293
  );


  xor
  g2572
  (
    n2615,
    n2313,
    n2252,
    n2320,
    n2342
  );


  nand
  g2573
  (
    n2620,
    n2291,
    n2246,
    n2404,
    n2380
  );


  xor
  g2574
  (
    n2567,
    n2430,
    n2405,
    n2307,
    n2304
  );


  nand
  g2575
  (
    n2687,
    n2299,
    n2406,
    n2242,
    n2294
  );


  or
  g2576
  (
    n2465,
    n2296,
    n2346,
    n2390,
    n2263
  );


  nand
  g2577
  (
    n2435,
    n2421,
    n2274,
    n1672,
    n2424
  );


  or
  g2578
  (
    n2513,
    n2275,
    n2250,
    n2387,
    n2244
  );


  nor
  g2579
  (
    n2472,
    n2425,
    n2395,
    n2389,
    n657
  );


  and
  g2580
  (
    n2469,
    n2346,
    n2292,
    n2413,
    n2344
  );


  or
  g2581
  (
    n2523,
    n2286,
    n2358,
    n2390,
    n2340
  );


  or
  g2582
  (
    n2559,
    n2382,
    n2380,
    n2316,
    n2355
  );


  and
  g2583
  (
    n2576,
    n2288,
    n2321,
    n2378,
    n2373
  );


  nand
  g2584
  (
    n2515,
    n2282,
    n2298,
    n2386,
    n2403
  );


  or
  g2585
  (
    n2592,
    n2338,
    n2300,
    n2406,
    n2317
  );


  nor
  g2586
  (
    n2580,
    n2368,
    n2250,
    n2412,
    n2347
  );


  nand
  g2587
  (
    n2520,
    n2427,
    n2308,
    n2430,
    n2389
  );


  nand
  g2588
  (
    n2600,
    n2415,
    n2343,
    n2271,
    n2319
  );


  nor
  g2589
  (
    n2584,
    n2282,
    n2407,
    n2402,
    n2253
  );


  or
  g2590
  (
    n2674,
    n2336,
    n2296,
    n2241,
    n2270
  );


  and
  g2591
  (
    n2589,
    n2402,
    n2341,
    n2242,
    n2339
  );


  nor
  g2592
  (
    n2596,
    n2377,
    n2325,
    n2413,
    n2241
  );


  nor
  g2593
  (
    n2480,
    n2428,
    n2426,
    n2287,
    n2337
  );


  and
  g2594
  (
    n2525,
    n2304,
    n2293,
    n2373,
    n2254
  );


  nand
  g2595
  (
    n2570,
    n2342,
    n2376,
    n2297,
    n2325
  );


  nor
  g2596
  (
    n2512,
    n2423,
    n2295,
    n2411,
    n2399
  );


  nor
  g2597
  (
    n2587,
    n2374,
    n2248,
    n2342,
    n1677
  );


  xor
  g2598
  (
    n2653,
    n2334,
    n2386,
    n2315,
    n2359
  );


  nand
  g2599
  (
    n2494,
    n2337,
    n2350,
    n2422,
    n2335
  );


  or
  g2600
  (
    n2703,
    n2288,
    n2408,
    n2413,
    n2300
  );


  or
  g2601
  (
    n2453,
    n2371,
    n2396,
    n2301,
    n2269
  );


  xor
  g2602
  (
    n2618,
    n2284,
    n2425,
    n2329,
    n2288
  );


  and
  g2603
  (
    n2617,
    n2314,
    n2285,
    n2316,
    n2315
  );


  or
  g2604
  (
    n2698,
    n2275,
    n2428,
    n2300,
    n2328
  );


  nor
  g2605
  (
    n2575,
    n2286,
    n2246,
    n2385,
    n2376
  );


  nand
  g2606
  (
    n2684,
    n2414,
    n2348,
    n2318,
    n2391
  );


  and
  g2607
  (
    n2583,
    n2264,
    n2353,
    n2246,
    n2341
  );


  nor
  g2608
  (
    n2551,
    n2340,
    n2319,
    n2349,
    n2360
  );


  xnor
  g2609
  (
    n2685,
    n2281,
    n2379,
    n2401,
    n2338
  );


  or
  g2610
  (
    n2701,
    n2331,
    n2266,
    n2402,
    n2374
  );


  and
  g2611
  (
    n2437,
    n2398,
    n1678,
    n2176,
    n2321
  );


  or
  g2612
  (
    n2662,
    n2271,
    n2423,
    n2312,
    n2245
  );


  and
  g2613
  (
    n2658,
    n2378,
    n2266,
    n2368,
    n2290
  );


  xnor
  g2614
  (
    n2438,
    n2385,
    n2350,
    n2258,
    n2420
  );


  nand
  g2615
  (
    n2616,
    n2305,
    n2399,
    n2243,
    n2358
  );


  nand
  g2616
  (
    n2672,
    n2307,
    n2327,
    n2301,
    n2354
  );


  xor
  g2617
  (
    n2456,
    n1675,
    n2355,
    n2325,
    n2370
  );


  xor
  g2618
  (
    n2614,
    n2431,
    n2270,
    n2246,
    n1683
  );


  nor
  g2619
  (
    n2511,
    n2297,
    n2248,
    n2151,
    n2333
  );


  xnor
  g2620
  (
    n2648,
    n2354,
    n2407,
    n2425,
    n2293
  );


  xor
  g2621
  (
    n2530,
    n2326,
    n2362,
    n2399,
    n2299
  );


  xor
  g2622
  (
    n2569,
    n2245,
    n2348,
    n2421,
    n2298
  );


  xnor
  g2623
  (
    n2455,
    n2362,
    n2372,
    n2283,
    n2291
  );


  nor
  g2624
  (
    n2595,
    n2258,
    n2380,
    n2319,
    n2268
  );


  or
  g2625
  (
    n2668,
    n2400,
    n2288,
    n2252,
    n2260
  );


  nor
  g2626
  (
    n2474,
    n2274,
    n2388,
    n2337,
    n2414
  );


  xnor
  g2627
  (
    n2670,
    n2289,
    n2379,
    n2426,
    n2406
  );


  xor
  g2628
  (
    n2632,
    n2402,
    n2281,
    n2276,
    n2256
  );


  and
  g2629
  (
    n2693,
    n2411,
    n2363,
    n2298,
    n1684
  );


  and
  g2630
  (
    n2663,
    n2401,
    n2267,
    n2409,
    n2269
  );


  and
  g2631
  (
    n2452,
    n655,
    n2357,
    n2372,
    n2278
  );


  nand
  g2632
  (
    n2582,
    n2409,
    n2430,
    n2393,
    n2359
  );


  nand
  g2633
  (
    n2598,
    n2428,
    n2424,
    n2277,
    n2327
  );


  and
  g2634
  (
    n2543,
    n2397,
    n2333,
    n2370,
    n2296
  );


  or
  g2635
  (
    n2442,
    n1674,
    n2343,
    n2351,
    n2278
  );


  and
  g2636
  (
    n2507,
    n2387,
    n2357,
    n2276,
    n2265
  );


  nor
  g2637
  (
    n2603,
    n2240,
    n2307,
    n2310,
    n1680
  );


  xnor
  g2638
  (
    n2487,
    n2378,
    n2331,
    n2386,
    n2353
  );


  and
  g2639
  (
    n2593,
    n2415,
    n2272,
    n2332,
    n2397
  );


  and
  g2640
  (
    n2536,
    n2353,
    n2388,
    n2312,
    n2243
  );


  nand
  g2641
  (
    n2436,
    n1673,
    n2428,
    n2416,
    n2252
  );


  xnor
  g2642
  (
    n2548,
    n2322,
    n2424,
    n2310,
    n2272
  );


  xnor
  g2643
  (
    n2541,
    n2270,
    n2383,
    n2274,
    n2359
  );


  xnor
  g2644
  (
    n2591,
    n2261,
    n2261,
    n2303,
    n2247
  );


  xor
  g2645
  (
    n2500,
    n2371,
    n2340,
    n2392,
    n2300
  );


  xor
  g2646
  (
    n2558,
    n2258,
    n2417,
    n2311,
    n2347
  );


  nor
  g2647
  (
    n2535,
    n2405,
    n2421,
    n2333,
    n2267
  );


  xnor
  g2648
  (
    n2459,
    n2369,
    n2309,
    n2358,
    n2241
  );


  xor
  g2649
  (
    n2568,
    n2291,
    n2256,
    n2282,
    n2264
  );


  xnor
  g2650
  (
    n2602,
    n2310,
    n2311,
    n2254,
    n2287
  );


  or
  g2651
  (
    n2637,
    n2333,
    n2349,
    n2323,
    n2253
  );


  xor
  g2652
  (
    n2524,
    n2176,
    n2316,
    n2320,
    n2352
  );


  and
  g2653
  (
    n2546,
    n1676,
    n2374,
    n2394,
    n2344
  );


  nor
  g2654
  (
    n2678,
    n2414,
    n2294,
    n2327,
    n2393
  );


  xor
  g2655
  (
    n2608,
    n2263,
    n2244,
    n2330,
    n2264
  );


  nand
  g2656
  (
    n2574,
    n2277,
    n2361,
    n2287,
    n2284
  );


  xor
  g2657
  (
    n2660,
    n2324,
    n2274,
    n2338,
    n2362
  );


  and
  g2658
  (
    n2656,
    n2429,
    n2396,
    n2324,
    n2292
  );


  nor
  g2659
  (
    n2689,
    n2260,
    n2338,
    n2334,
    n2323
  );


  and
  g2660
  (
    n2565,
    n2410,
    n2383,
    n2400,
    n2244
  );


  nor
  g2661
  (
    n2627,
    n2370,
    n2355,
    n2394,
    n2321
  );


  nor
  g2662
  (
    n2532,
    n2334,
    n2259,
    n2366,
    n2266
  );


  and
  g2663
  (
    n2606,
    n2280,
    n2389,
    n2422,
    n2266
  );


  and
  g2664
  (
    n2562,
    n2352,
    n2386,
    n2395,
    n2244
  );


  and
  g2665
  (
    n2488,
    n2365,
    n2393,
    n2267,
    n2286
  );


  xnor
  g2666
  (
    n2450,
    n2375,
    n2377,
    n2419,
    n2255
  );


  nand
  g2667
  (
    n2448,
    n2359,
    n2397,
    n2302,
    n2314
  );


  or
  g2668
  (
    n2517,
    n2330,
    n2357,
    n2411,
    n2336
  );


  or
  g2669
  (
    n2527,
    n2249,
    n2279,
    n2392,
    n2391
  );


  nor
  g2670
  (
    n2549,
    n2363,
    n2363,
    n2394,
    n2240
  );


  or
  g2671
  (
    n2715,
    n2438,
    n2462,
    n2466,
    n2464
  );


  and
  g2672
  (
    n2711,
    n2479,
    n2448,
    n2440,
    n2434
  );


  xnor
  g2673
  (
    n2704,
    n2473,
    n2447,
    n2457,
    n2446
  );


  or
  g2674
  (
    n2709,
    n2432,
    n2441,
    n2437,
    n2444
  );


  xor
  g2675
  (
    n2710,
    n2471,
    n2454,
    n2474,
    n2472
  );


  nand
  g2676
  (
    KeyWire_0_14,
    n2433,
    n2456,
    n2451,
    n2435
  );


  xnor
  g2677
  (
    n2714,
    n2478,
    n2460,
    n2468,
    n2443
  );


  and
  g2678
  (
    n2707,
    n2458,
    n2477,
    n2453,
    n2465
  );


  xnor
  g2679
  (
    n2713,
    n2467,
    n2452,
    n2463,
    n2455
  );


  nor
  g2680
  (
    n2706,
    n2449,
    n2476,
    n2442,
    n2445
  );


  nand
  g2681
  (
    n2708,
    n2439,
    n2459,
    n2436,
    n2469
  );


  and
  g2682
  (
    n2705,
    n2475,
    n2461,
    n2470,
    n2450
  );


  and
  g2683
  (
    n2716,
    n1685,
    n2715
  );


  xnor
  g2684
  (
    n2719,
    n2168,
    n2716,
    n2166
  );


  xnor
  g2685
  (
    n2718,
    n2166,
    n2165
  );


  or
  g2686
  (
    n2720,
    n2164,
    n2165,
    n2166,
    n2716
  );


  xnor
  g2687
  (
    n2717,
    n2166,
    n1686,
    n2716,
    n2164
  );


  or
  g2688
  (
    n2722,
    n2488,
    n2502,
    n2489,
    n2494
  );


  nor
  g2689
  (
    n2725,
    n2497,
    n2485,
    n2501,
    n2481
  );


  nand
  g2690
  (
    n2727,
    n2482,
    n2720,
    n2719,
    n2500
  );


  xnor
  g2691
  (
    n2724,
    n2498,
    n2490,
    n2484,
    n2491
  );


  xor
  g2692
  (
    n2726,
    n2492,
    n2717,
    n2486,
    n2499
  );


  and
  g2693
  (
    n2723,
    n2503,
    n2496,
    n2720,
    n2483
  );


  or
  g2694
  (
    n2721,
    n2480,
    n2487,
    n2495,
    n2493
  );


  and
  g2695
  (
    n2728,
    n2720,
    n2719,
    n2718
  );


  nor
  g2696
  (
    n2730,
    n2723,
    n2158,
    n2057
  );


  nor
  g2697
  (
    n2734,
    n2171,
    n2061,
    n2506
  );


  nand
  g2698
  (
    n2739,
    n2728,
    n2724,
    n2054
  );


  xnor
  g2699
  (
    n2735,
    n2052,
    n2725,
    n2058
  );


  or
  g2700
  (
    n2745,
    n657,
    n2171,
    n2045
  );


  nand
  g2701
  (
    n2729,
    n658,
    n2726,
    n2060
  );


  xor
  g2702
  (
    n2737,
    n2431,
    n2727,
    n2728
  );


  and
  g2703
  (
    n2738,
    n2155,
    n2726
  );


  nor
  g2704
  (
    n2742,
    n2055,
    n2727
  );


  or
  g2705
  (
    n2736,
    n659,
    n2050,
    n2059
  );


  xor
  g2706
  (
    n2731,
    n2046,
    n2431,
    n2504
  );


  and
  g2707
  (
    n2741,
    n2721,
    n2156,
    n2505
  );


  xor
  g2708
  (
    n2740,
    n2726,
    n2154,
    n658
  );


  nand
  g2709
  (
    n2732,
    n2049,
    n2171,
    n2048
  );


  nor
  g2710
  (
    n2744,
    n2157,
    n2056,
    n2047,
    n2728
  );


  or
  g2711
  (
    n2733,
    n2431,
    n2725,
    n2051,
    n658
  );


  xnor
  g2712
  (
    n2743,
    n2728,
    n2053,
    n659,
    n2722
  );


  nor
  g2713
  (
    n2746,
    n2159,
    n657,
    n2727,
    n658
  );


  and
  g2714
  (
    n2748,
    n2731,
    n2733,
    n2734
  );


  xnor
  g2715
  (
    n2747,
    n2732,
    n2730,
    n2733,
    n2729
  );


  xnor
  g2716
  (
    n2753,
    n662,
    n662,
    n660,
    n661
  );


  or
  g2717
  (
    n2754,
    n2748,
    n2748,
    n2747,
    n660
  );


  and
  g2718
  (
    n2749,
    n661,
    n659,
    n2747,
    n2748
  );


  or
  g2719
  (
    n2751,
    n1688,
    n659,
    n2747,
    n662
  );


  nand
  g2720
  (
    n2752,
    n1689,
    n660,
    n1690,
    n1687
  );


  nand
  g2721
  (
    n2750,
    n660,
    n661,
    n662
  );


  nor
  g2722
  (
    n2755,
    n1693,
    n1691,
    n1692,
    n2751
  );


  not
  g2723
  (
    n2758,
    n2755
  );


  not
  g2724
  (
    n2756,
    n2755
  );


  buf
  g2725
  (
    n2759,
    n2755
  );


  buf
  g2726
  (
    n2757,
    n2755
  );


  nor
  g2727
  (
    n2771,
    n1700,
    n1708,
    n2527,
    n1698
  );


  nor
  g2728
  (
    n2774,
    n1709,
    n1703,
    n2523,
    n2756
  );


  nand
  g2729
  (
    n2763,
    n2524,
    n2510,
    n2759,
    n2520
  );


  xnor
  g2730
  (
    n2772,
    n2757,
    n2758,
    n2521,
    n2756
  );


  and
  g2731
  (
    n2764,
    n2512,
    n2519,
    n1697,
    n1699
  );


  or
  g2732
  (
    n2773,
    n2511,
    n2757,
    n2758,
    n2526
  );


  xnor
  g2733
  (
    n2769,
    n2756,
    n2535,
    n2525,
    n1705
  );


  or
  g2734
  (
    n2775,
    n2518,
    n2536,
    n2517,
    n1702
  );


  xnor
  g2735
  (
    n2765,
    n2759,
    n1706,
    n2513,
    n2516
  );


  and
  g2736
  (
    n2760,
    n1704,
    n2515,
    n2758,
    n2528
  );


  or
  g2737
  (
    n2767,
    n1696,
    n2507,
    n2532,
    n2514
  );


  nor
  g2738
  (
    n2762,
    n1694,
    n1695,
    n1710,
    n2759
  );


  xnor
  g2739
  (
    n2766,
    n2757,
    n2509,
    n2756,
    n2530
  );


  xnor
  g2740
  (
    n2768,
    n2537,
    n2534,
    n2508,
    n2758
  );


  xor
  g2741
  (
    n2761,
    n1707,
    n2533,
    n2757,
    n2522
  );


  xnor
  g2742
  (
    n2770,
    n1701,
    n2531,
    n2759,
    n2529
  );


  nor
  g2743
  (
    n2791,
    n2588,
    n2687,
    n2761,
    n2626
  );


  xor
  g2744
  (
    n2809,
    n2736,
    n2701,
    n2676,
    n2615
  );


  xnor
  g2745
  (
    n2784,
    n2735,
    n2663,
    n2702,
    n2654
  );


  and
  g2746
  (
    n2804,
    n2584,
    n2586,
    n2734,
    n2764
  );


  or
  g2747
  (
    n2796,
    n2762,
    n2567,
    n2631,
    n2774
  );


  xor
  g2748
  (
    n2832,
    n2700,
    n2598,
    n2601,
    n2703
  );


  nor
  g2749
  (
    n2837,
    n2738,
    n2760,
    n2590,
    n2648
  );


  xnor
  g2750
  (
    n2821,
    n2630,
    n2671,
    n2769,
    n2653
  );


  and
  g2751
  (
    n2806,
    n2565,
    n2766,
    n2612,
    n2682
  );


  nand
  g2752
  (
    n2786,
    n2675,
    n2763,
    n2664
  );


  and
  g2753
  (
    n2826,
    n2568,
    n2774,
    n2622,
    n2760
  );


  or
  g2754
  (
    n2816,
    n2634,
    n2636,
    n2608,
    n2555
  );


  xnor
  g2755
  (
    n2798,
    n2587,
    n2538,
    n2703,
    n2667
  );


  xor
  g2756
  (
    n2793,
    n2592,
    n2767,
    n2771,
    n2600
  );


  xor
  g2757
  (
    n2787,
    n2605,
    n2574,
    n2623,
    n2641
  );


  nand
  g2758
  (
    n2778,
    n2762,
    n2647,
    n2694,
    n2738
  );


  xor
  g2759
  (
    n2822,
    n2625,
    n2765,
    n2772,
    n2734
  );


  nand
  g2760
  (
    n2820,
    n2558,
    n2657,
    n2775,
    n2769
  );


  and
  g2761
  (
    n2810,
    n2770,
    n2646,
    n2661,
    n2580
  );


  and
  g2762
  (
    n2818,
    n2775,
    n2596,
    n2550,
    n2616
  );


  nand
  g2763
  (
    n2788,
    n2585,
    n2698,
    n2774,
    n2767
  );


  and
  g2764
  (
    n2780,
    n2762,
    n2763,
    n2603,
    n2611
  );


  or
  g2765
  (
    n2779,
    n2665,
    n2607,
    n2610,
    n2768
  );


  or
  g2766
  (
    n2785,
    n2668,
    n2547,
    n2770,
    n2570
  );


  nor
  g2767
  (
    n2789,
    n2695,
    n2613,
    n2540,
    n2666
  );


  nor
  g2768
  (
    n2802,
    n2650,
    n2738,
    n2633,
    n2674
  );


  xor
  g2769
  (
    n2819,
    n2737,
    n2770,
    n2573,
    n2539
  );


  xnor
  g2770
  (
    n2811,
    n2579,
    n2548,
    n2583,
    n2771
  );


  and
  g2771
  (
    n2834,
    n2762,
    n2761,
    n2639
  );


  nor
  g2772
  (
    n2792,
    n2774,
    n2702,
    n2699,
    n2770
  );


  xor
  g2773
  (
    n2783,
    n2768,
    n2752,
    n2739,
    n2649
  );


  or
  g2774
  (
    n2790,
    n2638,
    n2703,
    n2739,
    n2686
  );


  or
  g2775
  (
    n2812,
    n2754,
    n2673,
    n2589,
    n2618
  );


  xor
  g2776
  (
    n2813,
    n2651,
    n2609,
    n2542,
    n2652
  );


  xnor
  g2777
  (
    n2795,
    n2659,
    n2689,
    n2576,
    n2735
  );


  xor
  g2778
  (
    n2830,
    n2572,
    n2697,
    n2563,
    n2771
  );


  or
  g2779
  (
    n2825,
    n2760,
    n2645,
    n2703,
    n2696
  );


  nand
  g2780
  (
    n2815,
    n2684,
    n2629,
    n2594,
    n2593
  );


  or
  g2781
  (
    n2801,
    n2736,
    n2578,
    n2559,
    n2562
  );


  xor
  g2782
  (
    n2777,
    n2672,
    n2632,
    n2566,
    n2766
  );


  xnor
  g2783
  (
    n2814,
    n2602,
    n2761,
    n2736,
    n2753
  );


  xor
  g2784
  (
    n2839,
    n2771,
    n2677,
    n2678,
    n2561
  );


  nor
  g2785
  (
    n2829,
    n2617,
    n2560,
    n2693,
    n2557
  );


  and
  g2786
  (
    n2781,
    n2766,
    n2546,
    n2772,
    n2564
  );


  nor
  g2787
  (
    n2776,
    n2599,
    n2551,
    n2552,
    n2637
  );


  nand
  g2788
  (
    n2799,
    n2670,
    n2569,
    n2773,
    n2679
  );


  xnor
  g2789
  (
    n2817,
    n2549,
    n2614,
    n2642,
    n2553
  );


  xor
  g2790
  (
    n2803,
    n2773,
    n2760,
    n2620,
    n2739
  );


  xnor
  g2791
  (
    n2782,
    n2764,
    n2621,
    n2767,
    n2635
  );


  xor
  g2792
  (
    n2836,
    n2680,
    n2765,
    n2628,
    n2767
  );


  nor
  g2793
  (
    n2823,
    n2768,
    n2737,
    n2692,
    n2773
  );


  and
  g2794
  (
    n2807,
    n2702,
    n2683,
    n2571,
    n2606
  );


  xnor
  g2795
  (
    n2835,
    n2624,
    n2581,
    n2769,
    n2768
  );


  xor
  g2796
  (
    n2797,
    n2597,
    n2764,
    n2765
  );


  nand
  g2797
  (
    n2800,
    n2545,
    n2658,
    n2643,
    n2766
  );


  nand
  g2798
  (
    n2805,
    n2575,
    n2543,
    n2773,
    n2772
  );


  xnor
  g2799
  (
    n2794,
    n2619,
    n2556,
    n2769,
    n2656
  );


  xor
  g2800
  (
    n2824,
    n2681,
    n2775,
    n2604,
    n2737
  );


  nor
  g2801
  (
    n2828,
    n2765,
    n2627,
    n2595,
    n2685
  );


  xor
  g2802
  (
    n2833,
    n2690,
    n2541,
    n2669,
    n2662
  );


  or
  g2803
  (
    n2831,
    n2775,
    n2688,
    n2582,
    n2763
  );


  or
  g2804
  (
    n2808,
    n2554,
    n2644,
    n2655,
    n2544
  );


  or
  g2805
  (
    n2838,
    n2640,
    n2735,
    n2691,
    n2577
  );


  xor
  g2806
  (
    n2827,
    n2591,
    n2702,
    n2772,
    n2660
  );


  buf
  g2807
  (
    n2909,
    n2821
  );


  not
  g2808
  (
    n2854,
    n2833
  );


  not
  g2809
  (
    n2917,
    n2152
  );


  buf
  g2810
  (
    n2870,
    n2787
  );


  not
  g2811
  (
    n2879,
    n2071
  );


  not
  g2812
  (
    n2896,
    n2786
  );


  buf
  g2813
  (
    n2884,
    n2790
  );


  buf
  g2814
  (
    n2856,
    n2805
  );


  not
  g2815
  (
    n2888,
    n2778
  );


  buf
  g2816
  (
    n2895,
    n2831
  );


  buf
  g2817
  (
    n2867,
    n2069
  );


  buf
  g2818
  (
    n2920,
    n2836
  );


  buf
  g2819
  (
    n2868,
    n2776
  );


  buf
  g2820
  (
    n2864,
    n2795
  );


  nand
  g2821
  (
    n2858,
    n2817,
    n2777,
    n2795
  );


  nand
  g2822
  (
    n2902,
    n2829,
    n2066,
    n2834
  );


  nand
  g2823
  (
    n2878,
    n2160,
    n2812,
    n2789,
    n2835
  );


  xor
  g2824
  (
    n2911,
    n2838,
    n2802,
    n2742,
    n2784
  );


  xor
  g2825
  (
    n2872,
    n2786,
    n2828,
    n2788,
    n2799
  );


  or
  g2826
  (
    n2883,
    n2835,
    n2804,
    n2834,
    n2825
  );


  xor
  g2827
  (
    n2910,
    n2808,
    n2797,
    n2805
  );


  nor
  g2828
  (
    n2904,
    n2793,
    n2806,
    n2805,
    n2839
  );


  nand
  g2829
  (
    n2846,
    n2801,
    n2793,
    n2790,
    n2741
  );


  nand
  g2830
  (
    n2926,
    n2748,
    n2781,
    n2741,
    n2830
  );


  nor
  g2831
  (
    n2885,
    n2779,
    n2797,
    n2819,
    n2821
  );


  nand
  g2832
  (
    KeyWire_0_4,
    n2790,
    n2829,
    n2816,
    n2778
  );


  xnor
  g2833
  (
    n2924,
    n2831,
    n2785,
    n2784,
    n2827
  );


  nor
  g2834
  (
    n2892,
    n2809,
    n2744,
    n2161,
    n2806
  );


  xnor
  g2835
  (
    n2842,
    n2819,
    n2073,
    n2162,
    n2783
  );


  xor
  g2836
  (
    n2906,
    n2818,
    n2152,
    n2075,
    n2072
  );


  nand
  g2837
  (
    n2922,
    n2817,
    n2798,
    n2804,
    n2814
  );


  nand
  g2838
  (
    n2890,
    n2794,
    n2797,
    n2791,
    n2780
  );


  xnor
  g2839
  (
    n2899,
    n2744,
    n2743,
    n2780,
    n2806
  );


  nand
  g2840
  (
    n2871,
    n2813,
    n2833,
    n2791,
    n2151
  );


  xnor
  g2841
  (
    n2914,
    n664,
    n2816,
    n2776,
    n2783
  );


  and
  g2842
  (
    n2915,
    n2070,
    n2809,
    n2815,
    n2787
  );


  or
  g2843
  (
    n2865,
    n2807,
    n2818,
    n2800,
    n2779
  );


  xnor
  g2844
  (
    n2873,
    n2821,
    n2819,
    n2782,
    n2777
  );


  or
  g2845
  (
    n2841,
    n2836,
    n2829,
    n2810
  );


  or
  g2846
  (
    n2863,
    n2826,
    n2823,
    n2780,
    n2798
  );


  or
  g2847
  (
    n2894,
    n2067,
    n2798,
    n2810,
    n2782
  );


  xnor
  g2848
  (
    n2855,
    n2807,
    n2828,
    n2800,
    n2794
  );


  xnor
  g2849
  (
    n2848,
    n2815,
    n2802,
    n663,
    n2831
  );


  nor
  g2850
  (
    n2921,
    n2828,
    n2813,
    n2817,
    n2838
  );


  or
  g2851
  (
    n2887,
    n2832,
    n2800,
    n2824,
    n2792
  );


  or
  g2852
  (
    n2908,
    n2792,
    n2839,
    n2815,
    n2786
  );


  and
  g2853
  (
    n2925,
    n2785,
    n2828,
    n2792,
    n2818
  );


  and
  g2854
  (
    n2851,
    n2835,
    n2837,
    n2791,
    n2825
  );


  nand
  g2855
  (
    n2869,
    n2838,
    n2783,
    n2076,
    n2832
  );


  nand
  g2856
  (
    n2893,
    n2827,
    n2744,
    n2815,
    n2796
  );


  xnor
  g2857
  (
    n2903,
    n2830,
    n2832,
    n2793,
    n2822
  );


  nor
  g2858
  (
    n2875,
    n663,
    n2064,
    n2778,
    n2823
  );


  nor
  g2859
  (
    n2844,
    n2810,
    n2824,
    n2789,
    n2811
  );


  nand
  g2860
  (
    n2886,
    n2822,
    n2801,
    n2812,
    n2065
  );


  nand
  g2861
  (
    n2861,
    n2837,
    n2826,
    n2787,
    n2740
  );


  and
  g2862
  (
    n2847,
    n2063,
    n2793,
    n2068,
    n2810
  );


  nand
  g2863
  (
    n2891,
    n2796,
    n2807,
    n2812,
    n2789
  );


  nand
  g2864
  (
    n2859,
    n2794,
    n2152,
    n2742,
    n2832
  );


  or
  g2865
  (
    n2882,
    n2839,
    n2802,
    n2804,
    n2788
  );


  nand
  g2866
  (
    n2860,
    n2740,
    n2801,
    n2786,
    n2074
  );


  or
  g2867
  (
    n2843,
    n2823,
    n2789,
    n2797,
    n2803
  );


  xor
  g2868
  (
    n2877,
    n2742,
    n2780,
    n2821,
    n2787
  );


  or
  g2869
  (
    n2900,
    n2796,
    n2062,
    n2812,
    n2830
  );


  xnor
  g2870
  (
    n2850,
    n2781,
    n2811,
    n2839,
    n2794
  );


  or
  g2871
  (
    n2857,
    n159,
    n2824,
    n2778,
    n2152
  );


  and
  g2872
  (
    n2852,
    n2783,
    n2799,
    n2795,
    n2745
  );


  nand
  g2873
  (
    n2918,
    n2818,
    n2835,
    n664,
    n2814
  );


  xnor
  g2874
  (
    n2905,
    n2816,
    n664,
    n2830,
    n2798
  );


  nand
  g2875
  (
    n2862,
    n2788,
    n2792,
    n2784,
    n2811
  );


  xnor
  g2876
  (
    n2913,
    n2808,
    n2836,
    n2807,
    n663
  );


  nor
  g2877
  (
    n2876,
    n2809,
    n2825,
    n2813,
    n2820
  );


  nand
  g2878
  (
    n2912,
    n2800,
    n2833,
    n2804,
    n2809
  );


  or
  g2879
  (
    n2866,
    n2808,
    n2796,
    n663,
    n2777
  );


  xnor
  g2880
  (
    n2881,
    n1712,
    n2826,
    n1711,
    n2777
  );


  nor
  g2881
  (
    n2919,
    n2827,
    n2808,
    n2781,
    n2803
  );


  and
  g2882
  (
    n2907,
    n2785,
    n2802,
    n2790,
    n2799
  );


  xor
  g2883
  (
    n2898,
    n2831,
    n2781,
    n2803,
    n2784
  );


  nor
  g2884
  (
    n2840,
    n2799,
    n2814,
    n2782,
    n2827
  );


  nand
  g2885
  (
    n2897,
    n2820,
    n2078,
    n2823,
    n2838
  );


  or
  g2886
  (
    n2916,
    n2788,
    n2817,
    n2833,
    n2779
  );


  nand
  g2887
  (
    n2889,
    n2825,
    n2813,
    n2803,
    n2837
  );


  xnor
  g2888
  (
    n2901,
    n2785,
    n2791,
    n2740,
    n2820
  );


  nor
  g2889
  (
    n2853,
    n2819,
    n2779,
    n2077,
    n2741
  );


  xor
  g2890
  (
    n2880,
    n2782,
    n2826,
    n2834,
    n2822
  );


  xor
  g2891
  (
    n2849,
    n2795,
    n2801,
    n2776,
    n2743
  );


  or
  g2892
  (
    n2874,
    n2837,
    n2834,
    n2811,
    n2820
  );


  nor
  g2893
  (
    n2927,
    n2814,
    n2836,
    n2776,
    n2824
  );


  nor
  g2894
  (
    n2845,
    n2816,
    n2822,
    n2806,
    n2743
  );


  xor
  g2895
  (
    n2979,
    n1869,
    n2893,
    n1807,
    n1861
  );


  xnor
  g2896
  (
    n2942,
    n2884,
    n2856,
    n2910,
    n1776
  );


  or
  g2897
  (
    n2991,
    n1866,
    n1813,
    n2916,
    n1865
  );


  nand
  g2898
  (
    n2971,
    n2845,
    n1727,
    n2887,
    n1865
  );


  or
  g2899
  (
    n2988,
    n1815,
    n2915,
    n1792,
    n2863
  );


  nor
  g2900
  (
    n2953,
    n160,
    n1848,
    n1866,
    n1855
  );


  nor
  g2901
  (
    n2963,
    n1844,
    n1858,
    n1769,
    n1751
  );


  or
  g2902
  (
    n2978,
    n1836,
    n1863,
    n1851
  );


  xnor
  g2903
  (
    n2999,
    n2907,
    n1851,
    n1857,
    n664
  );


  and
  g2904
  (
    n2959,
    n2858,
    n1771,
    n1854,
    n1859
  );


  xnor
  g2905
  (
    n2954,
    n1862,
    n1828,
    n1820,
    n1869
  );


  xor
  g2906
  (
    n3003,
    n2889,
    n1808,
    n1765,
    n2859
  );


  or
  g2907
  (
    n2969,
    n1866,
    n2869,
    n1846,
    n2853
  );


  xor
  g2908
  (
    n2981,
    n1737,
    n1746,
    n1852,
    n2855
  );


  or
  g2909
  (
    n2935,
    n2849,
    n2852,
    n2908,
    n1859
  );


  or
  g2910
  (
    n2984,
    n2909,
    n1854,
    n1858,
    n2918
  );


  or
  g2911
  (
    n2929,
    n1809,
    n2898,
    n2857,
    n1806
  );


  xnor
  g2912
  (
    n2933,
    n1744,
    n1837,
    n1817,
    n1855
  );


  and
  g2913
  (
    n2985,
    n2904,
    n1719,
    n1868,
    n159
  );


  or
  g2914
  (
    n2974,
    n1790,
    n1849,
    n1735,
    n2850
  );


  and
  g2915
  (
    n3007,
    n1862,
    n1868,
    n2870,
    n1739
  );


  nand
  g2916
  (
    n2968,
    n2842,
    n1802,
    n2861,
    n1755
  );


  xnor
  g2917
  (
    n3004,
    n2905,
    n2906,
    n1731,
    n1754
  );


  nor
  g2918
  (
    n3005,
    n1821,
    n1866,
    n1716,
    n2872
  );


  or
  g2919
  (
    n2998,
    n1785,
    n1814,
    n2920,
    n1858
  );


  xnor
  g2920
  (
    n2943,
    n2883,
    n1779,
    n1732,
    n1852
  );


  nand
  g2921
  (
    n2931,
    n159,
    n1819,
    n1864,
    n2868
  );


  nand
  g2922
  (
    n2964,
    n1834,
    n2913,
    n1729,
    n2924
  );


  nor
  g2923
  (
    n2958,
    n2745,
    n1822,
    n1767,
    n2854
  );


  xnor
  g2924
  (
    n2962,
    n1870,
    n1800,
    n1838,
    n1862
  );


  nor
  g2925
  (
    n2966,
    n1781,
    n1845,
    n2886,
    n1870
  );


  nor
  g2926
  (
    n2994,
    n1825,
    n1853,
    n2874,
    n1856
  );


  xor
  g2927
  (
    n2945,
    n1860,
    n1859,
    n1753,
    n2919
  );


  or
  g2928
  (
    n2996,
    n2746,
    n1861,
    n2876,
    n2894
  );


  and
  g2929
  (
    n2970,
    n1823,
    n2925,
    n1730,
    n1832
  );


  xor
  g2930
  (
    n2987,
    n2921,
    n1861,
    n2903,
    n1852
  );


  nor
  g2931
  (
    n2976,
    n1782,
    n2891,
    n1840,
    n1750
  );


  xnor
  g2932
  (
    n2977,
    n160,
    n1714,
    n1853,
    n1775
  );


  and
  g2933
  (
    n3001,
    n1718,
    n1864,
    n2896,
    n1830
  );


  and
  g2934
  (
    n2975,
    n2864,
    n1827,
    n2846,
    n1851
  );


  nand
  g2935
  (
    KeyWire_0_6,
    n1855,
    n2892,
    n2871,
    n1867
  );


  xnor
  g2936
  (
    n2997,
    n1864,
    n1763,
    n1784,
    n1768
  );


  and
  g2937
  (
    n2993,
    n2746,
    n1804,
    n2911,
    n1868
  );


  and
  g2938
  (
    n2948,
    n1764,
    n2923,
    n1824,
    n1724
  );


  xnor
  g2939
  (
    n2952,
    n2897,
    n1863,
    n1852,
    n1810
  );


  and
  g2940
  (
    n2934,
    n1799,
    n1793,
    n1738,
    n1812
  );


  or
  g2941
  (
    n2946,
    n1795,
    n1788,
    n1783,
    n1854
  );


  xor
  g2942
  (
    n2967,
    n1869,
    n2878,
    n2888,
    n1756
  );


  nor
  g2943
  (
    n2972,
    n2865,
    n1863,
    n2917,
    n1777
  );


  nand
  g2944
  (
    n2951,
    n2745,
    n2746,
    n1722,
    n2862
  );


  and
  g2945
  (
    n2955,
    n1839,
    n2879,
    n1752,
    n1715
  );


  nor
  g2946
  (
    n2986,
    n1857,
    n1717,
    n1797,
    n1859
  );


  xnor
  g2947
  (
    n2932,
    n1831,
    n1794,
    n1721,
    n2900
  );


  nand
  g2948
  (
    n2982,
    n1860,
    n1726,
    n2844,
    n1857
  );


  xor
  g2949
  (
    n2956,
    n2877,
    n1851,
    n1842,
    n1816
  );


  nor
  g2950
  (
    n2950,
    n2847,
    n1780,
    n160,
    n1854
  );


  or
  g2951
  (
    n2980,
    n2848,
    n2901,
    n1833,
    n1855
  );


  nor
  g2952
  (
    n2990,
    n1742,
    n1869,
    n1868,
    n1856
  );


  nand
  g2953
  (
    n2992,
    n2843,
    n2890,
    n1749,
    n1748
  );


  nand
  g2954
  (
    n2938,
    n2902,
    n2841,
    n1857,
    n1772
  );


  xnor
  g2955
  (
    n2949,
    n2840,
    n1762,
    n2880,
    n1743
  );


  or
  g2956
  (
    n2995,
    n160,
    n1811,
    n1829,
    n1853
  );


  and
  g2957
  (
    n2965,
    n2866,
    n1757,
    n1734,
    n1801
  );


  nor
  g2958
  (
    n2937,
    n1761,
    n2895,
    n1865,
    n2860
  );


  xor
  g2959
  (
    n3006,
    n1741,
    n1728,
    n1870,
    n1745
  );


  xnor
  g2960
  (
    n2947,
    n2885,
    n1747,
    n1867,
    n2922
  );


  nand
  g2961
  (
    n2983,
    n2875,
    n1870,
    n1826,
    n1733
  );


  and
  g2962
  (
    n2936,
    n1865,
    n159,
    n1856,
    n1867
  );


  nor
  g2963
  (
    n3000,
    n1861,
    n2882,
    n1860,
    n1758
  );


  xor
  g2964
  (
    n2928,
    n1740,
    n2899,
    n2926,
    n1847
  );


  xor
  g2965
  (
    n2939,
    n2914,
    n1856,
    n1759,
    n1736
  );


  xnor
  g2966
  (
    n2944,
    n1770,
    n1713,
    n1789,
    n1760
  );


  xnor
  g2967
  (
    n2961,
    n2867,
    n1786,
    n1725,
    n1773
  );


  xnor
  g2968
  (
    n2957,
    n1818,
    n1864,
    n1860,
    n1805
  );


  or
  g2969
  (
    n2930,
    n1841,
    n1774,
    n1835,
    n1853
  );


  or
  g2970
  (
    n2940,
    n1803,
    n1720,
    n1850,
    n1766
  );


  xor
  g2971
  (
    n3002,
    n2881,
    n1796,
    n1843,
    n1867
  );


  xor
  g2972
  (
    n2973,
    n1787,
    n1791,
    n2851,
    n1862
  );


  xor
  g2973
  (
    n2941,
    n1858,
    n2912,
    n2927,
    n1778
  );


  xor
  g2974
  (
    n2989,
    n1850,
    n1798,
    n2873,
    n1723
  );


  and
  g2975
  (
    n3026,
    n3000,
    n2929,
    n2983,
    n2941
  );


  nand
  g2976
  (
    n3017,
    n2966,
    n2982,
    n2958,
    n2994
  );


  nand
  g2977
  (
    n3009,
    n2988,
    n2951,
    n2997,
    n2972
  );


  xor
  g2978
  (
    n3018,
    n2938,
    n2931,
    n2948,
    n2947
  );


  nor
  g2979
  (
    n3013,
    n2976,
    n3001,
    n2980,
    n2991
  );


  nor
  g2980
  (
    n3024,
    n2946,
    n2993,
    n3006,
    n2943
  );


  xnor
  g2981
  (
    n3015,
    n2928,
    n2952,
    n2978,
    n2975
  );


  nor
  g2982
  (
    n3014,
    n2995,
    n3002,
    n2945,
    n2998
  );


  xor
  g2983
  (
    n3011,
    n2942,
    n2956,
    n2973,
    n2930
  );


  xor
  g2984
  (
    n3019,
    n2974,
    n2970,
    n2962,
    n2944
  );


  nor
  g2985
  (
    n3025,
    n2981,
    n2939,
    n2969,
    n2977
  );


  xnor
  g2986
  (
    n3023,
    n2936,
    n2953,
    n2985,
    n2999
  );


  or
  g2987
  (
    n3027,
    n2984,
    n2955,
    n2933,
    n2940
  );


  nand
  g2988
  (
    n3008,
    n2971,
    n2963,
    n2996,
    n2937
  );


  xnor
  g2989
  (
    n3021,
    n2967,
    n2932,
    n3005,
    n2957
  );


  and
  g2990
  (
    n3020,
    n2934,
    n2960,
    n2986,
    n2954
  );


  nor
  g2991
  (
    n3012,
    n3003,
    n2968,
    n2989,
    n3007
  );


  nand
  g2992
  (
    n3016,
    n2950,
    n2961,
    n3004,
    n2959
  );


  or
  g2993
  (
    n3010,
    n2935,
    n2965,
    n2990,
    n2949
  );


  xor
  g2994
  (
    n3022,
    n2964,
    n2987,
    n2979,
    n2992
  );


  and
  g2995
  (
    n3028,
    n3008,
    n3012,
    n3026,
    n3021
  );


  xnor
  g2996
  (
    n3029,
    n3011,
    n3027,
    n3019,
    n3013
  );


  nor
  g2997
  (
    n3030,
    n3016,
    n3020,
    n3014,
    n3015
  );


  nand
  g2998
  (
    n3032,
    n3018,
    n3024,
    n3010,
    n3009
  );


  xnor
  g2999
  (
    n3031,
    n3017,
    n3023,
    n3022,
    n3025
  );


  xor
  KeyGate_0_0
  (
    n1967,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n200,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n1188,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1931,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n2923,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n105,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n2960,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n510,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n190,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n689,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n755,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1139,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n380,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n2613,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n2712,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n882,
    KeyNOTWire_0_15
  );


endmodule


