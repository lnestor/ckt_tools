

module Stat_1000_154
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n981,
  n976,
  n959,
  n969,
  n961,
  n978,
  n972,
  n974,
  n970,
  n973,
  n966,
  n971,
  n983,
  n965,
  n982,
  n963,
  n985,
  n977,
  n960,
  n968,
  n1022,
  n1030,
  n1032,
  n1021,
  n1024,
  n1031,
  n1025,
  n1029,
  n1027,
  n1028,
  n1026,
  n1023,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n981;
  output n976;
  output n959;
  output n969;
  output n961;
  output n978;
  output n972;
  output n974;
  output n970;
  output n973;
  output n966;
  output n971;
  output n983;
  output n965;
  output n982;
  output n963;
  output n985;
  output n977;
  output n960;
  output n968;
  output n1022;
  output n1030;
  output n1032;
  output n1021;
  output n1024;
  output n1031;
  output n1025;
  output n1029;
  output n1027;
  output n1028;
  output n1026;
  output n1023;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n962;
  wire n964;
  wire n967;
  wire n975;
  wire n979;
  wire n980;
  wire n984;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n62,
    n14
  );


  not
  g1
  (
    n59,
    n11
  );


  not
  g2
  (
    n112,
    n5
  );


  buf
  g3
  (
    n33,
    n26
  );


  buf
  g4
  (
    n94,
    n19
  );


  buf
  g5
  (
    n48,
    n20
  );


  not
  g6
  (
    n149,
    n2
  );


  buf
  g7
  (
    n63,
    n13
  );


  not
  g8
  (
    n86,
    n2
  );


  not
  g9
  (
    n46,
    n25
  );


  buf
  g10
  (
    n148,
    n22
  );


  not
  g11
  (
    n66,
    n7
  );


  buf
  g12
  (
    n41,
    n29
  );


  not
  g13
  (
    n141,
    n9
  );


  buf
  g14
  (
    n95,
    n17
  );


  not
  g15
  (
    n42,
    n10
  );


  buf
  g16
  (
    n151,
    n18
  );


  buf
  g17
  (
    n134,
    n26
  );


  buf
  g18
  (
    n113,
    n1
  );


  buf
  g19
  (
    n103,
    n4
  );


  not
  g20
  (
    n89,
    n15
  );


  buf
  g21
  (
    n64,
    n12
  );


  buf
  g22
  (
    n138,
    n32
  );


  buf
  g23
  (
    KeyWire_0_25,
    n1
  );


  not
  g24
  (
    n101,
    n28
  );


  not
  g25
  (
    n39,
    n24
  );


  buf
  g26
  (
    n58,
    n24
  );


  buf
  g27
  (
    n72,
    n19
  );


  not
  g28
  (
    n84,
    n30
  );


  buf
  g29
  (
    KeyWire_0_40,
    n20
  );


  buf
  g30
  (
    n73,
    n9
  );


  buf
  g31
  (
    KeyWire_0_30,
    n3
  );


  buf
  g32
  (
    n36,
    n8
  );


  not
  g33
  (
    n99,
    n11
  );


  not
  g34
  (
    n126,
    n31
  );


  not
  g35
  (
    n82,
    n5
  );


  not
  g36
  (
    n109,
    n28
  );


  buf
  g37
  (
    n37,
    n23
  );


  not
  g38
  (
    n106,
    n13
  );


  not
  g39
  (
    n156,
    n12
  );


  buf
  g40
  (
    n91,
    n20
  );


  buf
  g41
  (
    n52,
    n21
  );


  not
  g42
  (
    n108,
    n3
  );


  not
  g43
  (
    n107,
    n28
  );


  not
  g44
  (
    n60,
    n19
  );


  not
  g45
  (
    n140,
    n29
  );


  buf
  g46
  (
    n50,
    n4
  );


  not
  g47
  (
    n90,
    n30
  );


  not
  g48
  (
    n74,
    n10
  );


  buf
  g49
  (
    n133,
    n22
  );


  buf
  g50
  (
    KeyWire_0_22,
    n24
  );


  not
  g51
  (
    KeyWire_0_5,
    n27
  );


  not
  g52
  (
    n104,
    n16
  );


  buf
  g53
  (
    n155,
    n12
  );


  not
  g54
  (
    n81,
    n17
  );


  not
  g55
  (
    n157,
    n6
  );


  not
  g56
  (
    n145,
    n15
  );


  buf
  g57
  (
    n160,
    n9
  );


  not
  g58
  (
    n150,
    n12
  );


  buf
  g59
  (
    n122,
    n27
  );


  not
  g60
  (
    n100,
    n3
  );


  buf
  g61
  (
    n47,
    n4
  );


  buf
  g62
  (
    n142,
    n23
  );


  not
  g63
  (
    n130,
    n3
  );


  not
  g64
  (
    n132,
    n29
  );


  not
  g65
  (
    n131,
    n22
  );


  buf
  g66
  (
    n35,
    n15
  );


  not
  g67
  (
    n68,
    n19
  );


  buf
  g68
  (
    n143,
    n21
  );


  not
  g69
  (
    n111,
    n22
  );


  not
  g70
  (
    n61,
    n7
  );


  not
  g71
  (
    n96,
    n4
  );


  buf
  g72
  (
    n51,
    n9
  );


  buf
  g73
  (
    n98,
    n6
  );


  buf
  g74
  (
    KeyWire_0_38,
    n17
  );


  not
  g75
  (
    KeyWire_0_24,
    n1
  );


  buf
  g76
  (
    n57,
    n27
  );


  buf
  g77
  (
    n80,
    n6
  );


  buf
  g78
  (
    n158,
    n31
  );


  not
  g79
  (
    n144,
    n6
  );


  not
  g80
  (
    n45,
    n10
  );


  not
  g81
  (
    n127,
    n1
  );


  not
  g82
  (
    n117,
    n27
  );


  not
  g83
  (
    n67,
    n16
  );


  buf
  g84
  (
    n135,
    n10
  );


  buf
  g85
  (
    n136,
    n7
  );


  buf
  g86
  (
    n105,
    n30
  );


  buf
  g87
  (
    n124,
    n13
  );


  not
  g88
  (
    n76,
    n8
  );


  buf
  g89
  (
    n38,
    n29
  );


  not
  g90
  (
    n128,
    n25
  );


  buf
  g91
  (
    n85,
    n32
  );


  not
  g92
  (
    n116,
    n23
  );


  not
  g93
  (
    n137,
    n25
  );


  buf
  g94
  (
    n70,
    n8
  );


  not
  g95
  (
    n87,
    n28
  );


  buf
  g96
  (
    n88,
    n15
  );


  not
  g97
  (
    n102,
    n32
  );


  buf
  g98
  (
    n154,
    n18
  );


  buf
  g99
  (
    n93,
    n26
  );


  buf
  g100
  (
    n65,
    n21
  );


  buf
  g101
  (
    n53,
    n16
  );


  buf
  g102
  (
    n147,
    n21
  );


  not
  g103
  (
    n120,
    n16
  );


  not
  g104
  (
    n79,
    n26
  );


  not
  g105
  (
    n114,
    n30
  );


  buf
  g106
  (
    n153,
    n23
  );


  buf
  g107
  (
    KeyWire_0_0,
    n18
  );


  not
  g108
  (
    n123,
    n7
  );


  buf
  g109
  (
    n110,
    n18
  );


  buf
  g110
  (
    n40,
    n5
  );


  buf
  g111
  (
    n83,
    n17
  );


  buf
  g112
  (
    n129,
    n24
  );


  buf
  g113
  (
    n54,
    n25
  );


  not
  g114
  (
    n115,
    n5
  );


  buf
  g115
  (
    n34,
    n14
  );


  buf
  g116
  (
    n55,
    n11
  );


  not
  g117
  (
    n69,
    n14
  );


  not
  g118
  (
    n139,
    n2
  );


  buf
  g119
  (
    n75,
    n2
  );


  buf
  g120
  (
    n97,
    n20
  );


  not
  g121
  (
    n146,
    n11
  );


  buf
  g122
  (
    n78,
    n14
  );


  not
  g123
  (
    n152,
    n31
  );


  not
  g124
  (
    n121,
    n13
  );


  buf
  g125
  (
    n56,
    n32
  );


  buf
  g126
  (
    n159,
    n31
  );


  not
  g127
  (
    n119,
    n8
  );


  buf
  g128
  (
    n318,
    n40
  );


  buf
  g129
  (
    KeyWire_0_62,
    n51
  );


  not
  g130
  (
    n244,
    n84
  );


  not
  g131
  (
    n339,
    n61
  );


  not
  g132
  (
    n271,
    n93
  );


  buf
  g133
  (
    n192,
    n94
  );


  not
  g134
  (
    n463,
    n87
  );


  not
  g135
  (
    n414,
    n94
  );


  buf
  g136
  (
    n406,
    n98
  );


  not
  g137
  (
    n377,
    n80
  );


  buf
  g138
  (
    n447,
    n44
  );


  not
  g139
  (
    n472,
    n64
  );


  not
  g140
  (
    n188,
    n103
  );


  not
  g141
  (
    n213,
    n98
  );


  buf
  g142
  (
    n410,
    n45
  );


  not
  g143
  (
    KeyWire_0_20,
    n99
  );


  not
  g144
  (
    n415,
    n50
  );


  not
  g145
  (
    n223,
    n68
  );


  not
  g146
  (
    n400,
    n65
  );


  buf
  g147
  (
    n428,
    n76
  );


  not
  g148
  (
    n220,
    n92
  );


  not
  g149
  (
    n373,
    n39
  );


  not
  g150
  (
    n227,
    n73
  );


  not
  g151
  (
    n245,
    n87
  );


  buf
  g152
  (
    n198,
    n67
  );


  not
  g153
  (
    KeyWire_0_46,
    n39
  );


  buf
  g154
  (
    n385,
    n37
  );


  not
  g155
  (
    n430,
    n43
  );


  not
  g156
  (
    KeyWire_0_26,
    n48
  );


  not
  g157
  (
    KeyWire_0_50,
    n70
  );


  buf
  g158
  (
    n222,
    n103
  );


  not
  g159
  (
    n446,
    n108
  );


  buf
  g160
  (
    n181,
    n72
  );


  not
  g161
  (
    n405,
    n109
  );


  buf
  g162
  (
    n233,
    n60
  );


  not
  g163
  (
    n289,
    n35
  );


  not
  g164
  (
    n379,
    n80
  );


  not
  g165
  (
    n403,
    n110
  );


  buf
  g166
  (
    n243,
    n46
  );


  buf
  g167
  (
    n176,
    n60
  );


  buf
  g168
  (
    n298,
    n96
  );


  buf
  g169
  (
    n407,
    n78
  );


  buf
  g170
  (
    n388,
    n36
  );


  not
  g171
  (
    n255,
    n101
  );


  buf
  g172
  (
    KeyWire_0_39,
    n54
  );


  not
  g173
  (
    n445,
    n89
  );


  buf
  g174
  (
    n320,
    n86
  );


  buf
  g175
  (
    n349,
    n42
  );


  not
  g176
  (
    n288,
    n81
  );


  buf
  g177
  (
    n285,
    n47
  );


  not
  g178
  (
    KeyWire_0_19,
    n71
  );


  buf
  g179
  (
    n356,
    n88
  );


  not
  g180
  (
    n440,
    n105
  );


  not
  g181
  (
    n380,
    n58
  );


  not
  g182
  (
    n208,
    n41
  );


  not
  g183
  (
    n260,
    n99
  );


  not
  g184
  (
    n185,
    n45
  );


  not
  g185
  (
    n342,
    n58
  );


  not
  g186
  (
    n221,
    n87
  );


  not
  g187
  (
    n467,
    n102
  );


  buf
  g188
  (
    n392,
    n38
  );


  not
  g189
  (
    n319,
    n67
  );


  not
  g190
  (
    n471,
    n49
  );


  not
  g191
  (
    n376,
    n65
  );


  not
  g192
  (
    n393,
    n33
  );


  buf
  g193
  (
    n276,
    n90
  );


  not
  g194
  (
    n335,
    n34
  );


  buf
  g195
  (
    n402,
    n54
  );


  not
  g196
  (
    n351,
    n98
  );


  not
  g197
  (
    KeyWire_0_58,
    n40
  );


  buf
  g198
  (
    n206,
    n75
  );


  buf
  g199
  (
    n470,
    n93
  );


  not
  g200
  (
    n182,
    n105
  );


  not
  g201
  (
    n404,
    n40
  );


  buf
  g202
  (
    n168,
    n63
  );


  buf
  g203
  (
    n346,
    n79
  );


  not
  g204
  (
    n209,
    n61
  );


  buf
  g205
  (
    n417,
    n57
  );


  buf
  g206
  (
    n273,
    n96
  );


  not
  g207
  (
    n332,
    n53
  );


  buf
  g208
  (
    n418,
    n88
  );


  buf
  g209
  (
    n241,
    n74
  );


  buf
  g210
  (
    n237,
    n35
  );


  not
  g211
  (
    n193,
    n104
  );


  not
  g212
  (
    n432,
    n77
  );


  buf
  g213
  (
    n306,
    n68
  );


  buf
  g214
  (
    n341,
    n44
  );


  not
  g215
  (
    n210,
    n78
  );


  not
  g216
  (
    n161,
    n81
  );


  not
  g217
  (
    n473,
    n43
  );


  buf
  g218
  (
    KeyWire_0_54,
    n107
  );


  not
  g219
  (
    n300,
    n102
  );


  not
  g220
  (
    KeyWire_0_56,
    n80
  );


  not
  g221
  (
    n304,
    n46
  );


  not
  g222
  (
    n308,
    n109
  );


  buf
  g223
  (
    n202,
    n48
  );


  not
  g224
  (
    n256,
    n74
  );


  buf
  g225
  (
    n189,
    n73
  );


  not
  g226
  (
    n266,
    n100
  );


  buf
  g227
  (
    n448,
    n110
  );


  not
  g228
  (
    n167,
    n65
  );


  not
  g229
  (
    n216,
    n107
  );


  not
  g230
  (
    n283,
    n38
  );


  not
  g231
  (
    n230,
    n101
  );


  buf
  g232
  (
    n437,
    n74
  );


  not
  g233
  (
    n229,
    n89
  );


  buf
  g234
  (
    n282,
    n97
  );


  not
  g235
  (
    n372,
    n37
  );


  not
  g236
  (
    n426,
    n56
  );


  not
  g237
  (
    n184,
    n57
  );


  buf
  g238
  (
    n186,
    n53
  );


  not
  g239
  (
    KeyWire_0_57,
    n108
  );


  not
  g240
  (
    n169,
    n44
  );


  not
  g241
  (
    n452,
    n92
  );


  not
  g242
  (
    n324,
    n51
  );


  buf
  g243
  (
    n343,
    n103
  );


  buf
  g244
  (
    n360,
    n72
  );


  not
  g245
  (
    n171,
    n60
  );


  buf
  g246
  (
    n329,
    n96
  );


  not
  g247
  (
    n201,
    n41
  );


  buf
  g248
  (
    n228,
    n90
  );


  not
  g249
  (
    n424,
    n36
  );


  not
  g250
  (
    n162,
    n85
  );


  buf
  g251
  (
    n163,
    n102
  );


  not
  g252
  (
    KeyWire_0_6,
    n108
  );


  buf
  g253
  (
    n225,
    n71
  );


  not
  g254
  (
    n441,
    n37
  );


  buf
  g255
  (
    n179,
    n79
  );


  buf
  g256
  (
    n174,
    n82
  );


  buf
  g257
  (
    n173,
    n83
  );


  buf
  g258
  (
    n468,
    n83
  );


  not
  g259
  (
    n199,
    n104
  );


  not
  g260
  (
    n257,
    n66
  );


  buf
  g261
  (
    n338,
    n64
  );


  not
  g262
  (
    n164,
    n55
  );


  not
  g263
  (
    n365,
    n41
  );


  not
  g264
  (
    n313,
    n84
  );


  not
  g265
  (
    n390,
    n57
  );


  not
  g266
  (
    n270,
    n103
  );


  not
  g267
  (
    n328,
    n93
  );


  buf
  g268
  (
    n358,
    n34
  );


  not
  g269
  (
    n369,
    n33
  );


  buf
  g270
  (
    n262,
    n47
  );


  buf
  g271
  (
    n361,
    n100
  );


  buf
  g272
  (
    n327,
    n106
  );


  buf
  g273
  (
    n195,
    n100
  );


  buf
  g274
  (
    n226,
    n63
  );


  buf
  g275
  (
    n239,
    n38
  );


  buf
  g276
  (
    n170,
    n91
  );


  buf
  g277
  (
    n389,
    n58
  );


  buf
  g278
  (
    n333,
    n49
  );


  buf
  g279
  (
    n317,
    n55
  );


  buf
  g280
  (
    n409,
    n102
  );


  not
  g281
  (
    n190,
    n69
  );


  buf
  g282
  (
    n457,
    n62
  );


  not
  g283
  (
    n314,
    n76
  );


  not
  g284
  (
    n235,
    n83
  );


  not
  g285
  (
    n427,
    n50
  );


  not
  g286
  (
    n362,
    n110
  );


  buf
  g287
  (
    n382,
    n79
  );


  buf
  g288
  (
    n269,
    n54
  );


  not
  g289
  (
    n302,
    n99
  );


  buf
  g290
  (
    n419,
    n91
  );


  buf
  g291
  (
    n279,
    n42
  );


  buf
  g292
  (
    n316,
    n72
  );


  not
  g293
  (
    n453,
    n46
  );


  not
  g294
  (
    n197,
    n48
  );


  not
  g295
  (
    n178,
    n35
  );


  not
  g296
  (
    n461,
    n106
  );


  buf
  g297
  (
    n194,
    n66
  );


  not
  g298
  (
    n462,
    n86
  );


  buf
  g299
  (
    n175,
    n55
  );


  not
  g300
  (
    n251,
    n94
  );


  not
  g301
  (
    n310,
    n78
  );


  buf
  g302
  (
    n284,
    n106
  );


  not
  g303
  (
    n224,
    n45
  );


  buf
  g304
  (
    n207,
    n51
  );


  not
  g305
  (
    n305,
    n58
  );


  buf
  g306
  (
    n394,
    n43
  );


  buf
  g307
  (
    n259,
    n61
  );


  not
  g308
  (
    n177,
    n105
  );


  buf
  g309
  (
    n435,
    n109
  );


  not
  g310
  (
    n263,
    n73
  );


  buf
  g311
  (
    n165,
    n82
  );


  not
  g312
  (
    n200,
    n56
  );


  buf
  g313
  (
    n309,
    n49
  );


  not
  g314
  (
    n420,
    n106
  );


  buf
  g315
  (
    n326,
    n100
  );


  buf
  g316
  (
    n413,
    n52
  );


  buf
  g317
  (
    n395,
    n76
  );


  not
  g318
  (
    n340,
    n71
  );


  buf
  g319
  (
    n423,
    n69
  );


  buf
  g320
  (
    KeyWire_0_29,
    n90
  );


  buf
  g321
  (
    n399,
    n34
  );


  not
  g322
  (
    n354,
    n50
  );


  not
  g323
  (
    n294,
    n78
  );


  buf
  g324
  (
    n248,
    n69
  );


  buf
  g325
  (
    KeyWire_0_21,
    n40
  );


  not
  g326
  (
    n412,
    n84
  );


  not
  g327
  (
    n421,
    n34
  );


  buf
  g328
  (
    n203,
    n45
  );


  buf
  g329
  (
    n383,
    n99
  );


  buf
  g330
  (
    n293,
    n107
  );


  buf
  g331
  (
    n456,
    n52
  );


  buf
  g332
  (
    n425,
    n87
  );


  buf
  g333
  (
    n443,
    n104
  );


  not
  g334
  (
    n396,
    n89
  );


  not
  g335
  (
    n434,
    n76
  );


  not
  g336
  (
    n242,
    n92
  );


  not
  g337
  (
    n297,
    n84
  );


  not
  g338
  (
    n247,
    n70
  );


  buf
  g339
  (
    n246,
    n66
  );


  not
  g340
  (
    n368,
    n37
  );


  not
  g341
  (
    n217,
    n96
  );


  not
  g342
  (
    n166,
    n55
  );


  not
  g343
  (
    KeyWire_0_55,
    n94
  );


  buf
  g344
  (
    n433,
    n62
  );


  not
  g345
  (
    n439,
    n44
  );


  not
  g346
  (
    n449,
    n33
  );


  not
  g347
  (
    KeyWire_0_42,
    n85
  );


  buf
  g348
  (
    n348,
    n83
  );


  not
  g349
  (
    KeyWire_0_32,
    n63
  );


  not
  g350
  (
    n442,
    n88
  );


  not
  g351
  (
    n264,
    n95
  );


  buf
  g352
  (
    n234,
    n92
  );


  buf
  g353
  (
    n384,
    n86
  );


  buf
  g354
  (
    n180,
    n36
  );


  buf
  g355
  (
    n455,
    n95
  );


  not
  g356
  (
    n265,
    n69
  );


  buf
  g357
  (
    n367,
    n73
  );


  not
  g358
  (
    n336,
    n95
  );


  buf
  g359
  (
    n291,
    n85
  );


  not
  g360
  (
    n355,
    n77
  );


  not
  g361
  (
    n252,
    n104
  );


  buf
  g362
  (
    n350,
    n97
  );


  buf
  g363
  (
    n321,
    n110
  );


  buf
  g364
  (
    n438,
    n43
  );


  not
  g365
  (
    n258,
    n67
  );


  buf
  g366
  (
    n287,
    n91
  );


  buf
  g367
  (
    n391,
    n98
  );


  not
  g368
  (
    n214,
    n39
  );


  buf
  g369
  (
    n204,
    n53
  );


  not
  g370
  (
    n219,
    n75
  );


  buf
  g371
  (
    n292,
    n89
  );


  not
  g372
  (
    KeyWire_0_45,
    n35
  );


  buf
  g373
  (
    n268,
    n82
  );


  buf
  g374
  (
    n450,
    n42
  );


  buf
  g375
  (
    n311,
    n81
  );


  not
  g376
  (
    n299,
    n56
  );


  not
  g377
  (
    n303,
    n60
  );


  not
  g378
  (
    n322,
    n93
  );


  not
  g379
  (
    n345,
    n67
  );


  buf
  g380
  (
    n374,
    n61
  );


  not
  g381
  (
    n357,
    n71
  );


  not
  g382
  (
    n236,
    n101
  );


  not
  g383
  (
    n416,
    n72
  );


  not
  g384
  (
    KeyWire_0_3,
    n86
  );


  not
  g385
  (
    n386,
    n68
  );


  not
  g386
  (
    n254,
    n108
  );


  not
  g387
  (
    n290,
    n62
  );


  buf
  g388
  (
    n231,
    n63
  );


  buf
  g389
  (
    n460,
    n66
  );


  buf
  g390
  (
    n315,
    n51
  );


  not
  g391
  (
    n238,
    n36
  );


  not
  g392
  (
    n431,
    n90
  );


  buf
  g393
  (
    n337,
    n68
  );


  buf
  g394
  (
    n370,
    n54
  );


  buf
  g395
  (
    n267,
    n47
  );


  not
  g396
  (
    n296,
    n77
  );


  not
  g397
  (
    n253,
    n59
  );


  not
  g398
  (
    n183,
    n52
  );


  buf
  g399
  (
    n211,
    n107
  );


  buf
  g400
  (
    n459,
    n75
  );


  buf
  g401
  (
    n295,
    n59
  );


  not
  g402
  (
    n378,
    n109
  );


  not
  g403
  (
    n398,
    n70
  );


  buf
  g404
  (
    n469,
    n88
  );


  not
  g405
  (
    n397,
    n77
  );


  buf
  g406
  (
    n353,
    n91
  );


  not
  g407
  (
    n344,
    n52
  );


  not
  g408
  (
    n444,
    n59
  );


  buf
  g409
  (
    n281,
    n101
  );


  buf
  g410
  (
    n387,
    n95
  );


  not
  g411
  (
    n411,
    n85
  );


  not
  g412
  (
    n375,
    n50
  );


  buf
  g413
  (
    n451,
    n81
  );


  buf
  g414
  (
    n352,
    n70
  );


  buf
  g415
  (
    KeyWire_0_31,
    n56
  );


  buf
  g416
  (
    n364,
    n97
  );


  not
  g417
  (
    n187,
    n75
  );


  not
  g418
  (
    n280,
    n80
  );


  not
  g419
  (
    n172,
    n41
  );


  buf
  g420
  (
    n191,
    n64
  );


  buf
  g421
  (
    n347,
    n65
  );


  not
  g422
  (
    n277,
    n53
  );


  buf
  g423
  (
    n323,
    n57
  );


  buf
  g424
  (
    n363,
    n59
  );


  buf
  g425
  (
    n218,
    n105
  );


  buf
  g426
  (
    n359,
    n38
  );


  not
  g427
  (
    n454,
    n97
  );


  buf
  g428
  (
    n261,
    n33
  );


  buf
  g429
  (
    n331,
    n49
  );


  not
  g430
  (
    KeyWire_0_28,
    n47
  );


  not
  g431
  (
    n422,
    n74
  );


  buf
  g432
  (
    n307,
    n82
  );


  buf
  g433
  (
    n381,
    n64
  );


  not
  g434
  (
    n286,
    n46
  );


  buf
  g435
  (
    n301,
    n111
  );


  not
  g436
  (
    n212,
    n42
  );


  buf
  g437
  (
    n464,
    n79
  );


  not
  g438
  (
    n325,
    n48
  );


  not
  g439
  (
    n215,
    n39
  );


  not
  g440
  (
    n408,
    n62
  );


  buf
  g441
  (
    n484,
    n188
  );


  not
  g442
  (
    n486,
    n183
  );


  buf
  g443
  (
    n498,
    n177
  );


  buf
  g444
  (
    n476,
    n185
  );


  not
  g445
  (
    n489,
    n182
  );


  buf
  g446
  (
    n488,
    n173
  );


  buf
  g447
  (
    KeyWire_0_63,
    n174
  );


  buf
  g448
  (
    n480,
    n161
  );


  not
  g449
  (
    n487,
    n170
  );


  buf
  g450
  (
    n485,
    n167
  );


  not
  g451
  (
    n483,
    n178
  );


  not
  g452
  (
    n495,
    n168
  );


  not
  g453
  (
    n482,
    n184
  );


  not
  g454
  (
    n496,
    n186
  );


  not
  g455
  (
    n494,
    n189
  );


  not
  g456
  (
    n497,
    n165
  );


  buf
  g457
  (
    n479,
    n164
  );


  buf
  g458
  (
    n474,
    n176
  );


  buf
  g459
  (
    n481,
    n166
  );


  not
  g460
  (
    n475,
    n162
  );


  not
  g461
  (
    n477,
    n179
  );


  buf
  g462
  (
    n490,
    n171
  );


  not
  g463
  (
    n493,
    n175
  );


  buf
  g464
  (
    KeyWire_0_12,
    n190
  );


  buf
  g465
  (
    n499,
    n181
  );


  not
  g466
  (
    n500,
    n187
  );


  xnor
  g467
  (
    n501,
    n172,
    n169
  );


  or
  g468
  (
    n478,
    n180,
    n163
  );


  buf
  g469
  (
    n531,
    n117
  );


  buf
  g470
  (
    n511,
    n131
  );


  buf
  g471
  (
    n516,
    n115
  );


  buf
  g472
  (
    n558,
    n144
  );


  buf
  g473
  (
    n527,
    n127
  );


  buf
  g474
  (
    n507,
    n501
  );


  not
  g475
  (
    n519,
    n482
  );


  not
  g476
  (
    n553,
    n138
  );


  nor
  g477
  (
    n513,
    n475,
    n123,
    n113,
    n496
  );


  and
  g478
  (
    n508,
    n495,
    n118,
    n192,
    n132
  );


  nand
  g479
  (
    n533,
    n501,
    n126,
    n138,
    n139
  );


  nor
  g480
  (
    n517,
    n117,
    n139,
    n499,
    n201
  );


  and
  g481
  (
    n520,
    n144,
    n142,
    n121,
    n497
  );


  nor
  g482
  (
    n518,
    n119,
    n493,
    n487,
    n121
  );


  nand
  g483
  (
    n525,
    n121,
    n129,
    n122
  );


  xor
  g484
  (
    n556,
    n477,
    n140,
    n136,
    n474
  );


  xnor
  g485
  (
    n523,
    n143,
    n491,
    n114,
    n123
  );


  nand
  g486
  (
    n522,
    n500,
    n129,
    n124,
    n134
  );


  and
  g487
  (
    n503,
    n134,
    n493,
    n143,
    n481
  );


  or
  g488
  (
    n512,
    n494,
    n498,
    n120,
    n485
  );


  and
  g489
  (
    n552,
    n492,
    n128,
    n113,
    n120
  );


  xnor
  g490
  (
    n543,
    n112,
    n499,
    n135,
    n495
  );


  xnor
  g491
  (
    n559,
    n134,
    n496,
    n116,
    n140
  );


  nand
  g492
  (
    n551,
    n143,
    n120,
    n131,
    n144
  );


  nand
  g493
  (
    n555,
    n126,
    n125,
    n492,
    n122
  );


  or
  g494
  (
    n509,
    n138,
    n130,
    n133,
    n195
  );


  xor
  g495
  (
    n524,
    n116,
    n136,
    n122,
    n128
  );


  nor
  g496
  (
    n536,
    n116,
    n492,
    n498,
    n112
  );


  nand
  g497
  (
    n539,
    n498,
    n497,
    n478,
    n489
  );


  and
  g498
  (
    n545,
    n498,
    n124,
    n136,
    n141
  );


  and
  g499
  (
    n538,
    n493,
    n115,
    n117,
    n202
  );


  nand
  g500
  (
    n542,
    n493,
    n143,
    n198,
    n116
  );


  nor
  g501
  (
    n532,
    n145,
    n133,
    n142
  );


  or
  g502
  (
    KeyWire_0_2,
    n111,
    n114,
    n124,
    n486
  );


  nand
  g503
  (
    KeyWire_0_35,
    n199,
    n127,
    n130,
    n118
  );


  xor
  g504
  (
    n506,
    n113,
    n119,
    n112
  );


  or
  g505
  (
    n526,
    n128,
    n194,
    n132,
    n200
  );


  and
  g506
  (
    n537,
    n115,
    n114,
    n495,
    n120
  );


  xnor
  g507
  (
    n502,
    n500,
    n141,
    n135,
    n483
  );


  nand
  g508
  (
    n547,
    n118,
    n121,
    n494,
    n196
  );


  xor
  g509
  (
    n544,
    n494,
    n111,
    n128,
    n134
  );


  and
  g510
  (
    n540,
    n142,
    n480,
    n139,
    n127
  );


  nor
  g511
  (
    KeyWire_0_4,
    n123,
    n137,
    n132,
    n145
  );


  and
  g512
  (
    n557,
    n484,
    n133,
    n136,
    n500
  );


  nor
  g513
  (
    n549,
    n494,
    n488,
    n112,
    n140
  );


  xnor
  g514
  (
    n528,
    n132,
    n124,
    n137,
    n497
  );


  and
  g515
  (
    n554,
    n496,
    n479,
    n141,
    n144
  );


  or
  g516
  (
    n529,
    n119,
    n135,
    n130,
    n133
  );


  nor
  g517
  (
    n535,
    n495,
    n122,
    n139,
    n126
  );


  xor
  g518
  (
    n548,
    n499,
    n123,
    n135,
    n131
  );


  nand
  g519
  (
    n514,
    n492,
    n130,
    n127,
    n118
  );


  and
  g520
  (
    n541,
    n137,
    n113,
    n131,
    n499
  );


  xor
  g521
  (
    n504,
    n126,
    n193,
    n501,
    n137
  );


  or
  g522
  (
    n546,
    n197,
    n125,
    n501,
    n140
  );


  xor
  g523
  (
    n521,
    n497,
    n500,
    n125,
    n145
  );


  or
  g524
  (
    n534,
    n490,
    n115,
    n191,
    n125
  );


  and
  g525
  (
    n510,
    n114,
    n138,
    n141,
    n476
  );


  nand
  g526
  (
    n550,
    n496,
    n111,
    n117,
    n129
  );


  buf
  g527
  (
    n785,
    n147
  );


  buf
  g528
  (
    n686,
    n503
  );


  buf
  g529
  (
    n692,
    n531
  );


  buf
  g530
  (
    n595,
    n516
  );


  not
  g531
  (
    n772,
    n550
  );


  buf
  g532
  (
    n777,
    n156
  );


  buf
  g533
  (
    n721,
    n537
  );


  not
  g534
  (
    n663,
    n517
  );


  buf
  g535
  (
    KeyWire_0_14,
    n524
  );


  not
  g536
  (
    n791,
    n512
  );


  buf
  g537
  (
    n766,
    n550
  );


  buf
  g538
  (
    n742,
    n558
  );


  not
  g539
  (
    n617,
    n513
  );


  not
  g540
  (
    n580,
    n214
  );


  buf
  g541
  (
    n734,
    n555
  );


  not
  g542
  (
    n591,
    n559
  );


  not
  g543
  (
    n572,
    n507
  );


  buf
  g544
  (
    n653,
    n547
  );


  buf
  g545
  (
    KeyWire_0_13,
    n535
  );


  buf
  g546
  (
    n612,
    n146
  );


  buf
  g547
  (
    n751,
    n556
  );


  buf
  g548
  (
    n672,
    n149
  );


  not
  g549
  (
    n724,
    n148
  );


  not
  g550
  (
    n630,
    n555
  );


  not
  g551
  (
    n626,
    n528
  );


  buf
  g552
  (
    n589,
    n216
  );


  buf
  g553
  (
    n763,
    n250
  );


  buf
  g554
  (
    n631,
    n554
  );


  buf
  g555
  (
    n670,
    n545
  );


  buf
  g556
  (
    n671,
    n535
  );


  buf
  g557
  (
    n750,
    n515
  );


  buf
  g558
  (
    n654,
    n552
  );


  not
  g559
  (
    n741,
    n151
  );


  not
  g560
  (
    n752,
    n502
  );


  buf
  g561
  (
    n584,
    n152
  );


  not
  g562
  (
    KeyWire_0_23,
    n242
  );


  buf
  g563
  (
    n786,
    n543
  );


  buf
  g564
  (
    n638,
    n158
  );


  not
  g565
  (
    n702,
    n156
  );


  buf
  g566
  (
    KeyWire_0_43,
    n548
  );


  not
  g567
  (
    n790,
    n551
  );


  not
  g568
  (
    n652,
    n542
  );


  buf
  g569
  (
    n755,
    n530
  );


  buf
  g570
  (
    n603,
    n552
  );


  not
  g571
  (
    n743,
    n527
  );


  not
  g572
  (
    n758,
    n249
  );


  buf
  g573
  (
    n634,
    n526
  );


  not
  g574
  (
    n677,
    n245
  );


  buf
  g575
  (
    n737,
    n504
  );


  buf
  g576
  (
    n636,
    n228
  );


  buf
  g577
  (
    n602,
    n531
  );


  not
  g578
  (
    n695,
    n506
  );


  not
  g579
  (
    n687,
    n502
  );


  not
  g580
  (
    n649,
    n516
  );


  not
  g581
  (
    n756,
    n515
  );


  not
  g582
  (
    n712,
    n146
  );


  buf
  g583
  (
    n637,
    n505
  );


  buf
  g584
  (
    n749,
    n514
  );


  not
  g585
  (
    n604,
    n238
  );


  buf
  g586
  (
    n633,
    n522
  );


  not
  g587
  (
    n757,
    n536
  );


  not
  g588
  (
    n764,
    n153
  );


  not
  g589
  (
    n629,
    n510
  );


  buf
  g590
  (
    n662,
    n517
  );


  buf
  g591
  (
    n658,
    n155
  );


  buf
  g592
  (
    n568,
    n224
  );


  buf
  g593
  (
    n641,
    n528
  );


  not
  g594
  (
    n588,
    n240
  );


  buf
  g595
  (
    n646,
    n241
  );


  not
  g596
  (
    n779,
    n154
  );


  buf
  g597
  (
    n709,
    n527
  );


  buf
  g598
  (
    n661,
    n541
  );


  buf
  g599
  (
    n645,
    n540
  );


  buf
  g600
  (
    n600,
    n531
  );


  not
  g601
  (
    KeyWire_0_53,
    n212
  );


  buf
  g602
  (
    n625,
    n523
  );


  not
  g603
  (
    n780,
    n235
  );


  not
  g604
  (
    n620,
    n544
  );


  buf
  g605
  (
    n583,
    n545
  );


  buf
  g606
  (
    n747,
    n156
  );


  not
  g607
  (
    n782,
    n514
  );


  buf
  g608
  (
    n674,
    n548
  );


  buf
  g609
  (
    n697,
    n523
  );


  buf
  g610
  (
    n570,
    n237
  );


  not
  g611
  (
    n759,
    n219
  );


  buf
  g612
  (
    n754,
    n530
  );


  buf
  g613
  (
    n628,
    n203
  );


  not
  g614
  (
    n680,
    n155
  );


  not
  g615
  (
    n726,
    n159
  );


  not
  g616
  (
    n691,
    n513
  );


  not
  g617
  (
    n593,
    n511
  );


  buf
  g618
  (
    n668,
    n157
  );


  not
  g619
  (
    n562,
    n518
  );


  buf
  g620
  (
    n567,
    n541
  );


  not
  g621
  (
    n725,
    n152
  );


  not
  g622
  (
    n784,
    n150
  );


  buf
  g623
  (
    n770,
    n511
  );


  buf
  g624
  (
    n748,
    n555
  );


  buf
  g625
  (
    n738,
    n510
  );


  not
  g626
  (
    n616,
    n553
  );


  buf
  g627
  (
    KeyWire_0_41,
    n559
  );


  not
  g628
  (
    n566,
    n536
  );


  buf
  g629
  (
    n615,
    n524
  );


  not
  g630
  (
    n673,
    n521
  );


  not
  g631
  (
    n710,
    n513
  );


  buf
  g632
  (
    n699,
    n540
  );


  not
  g633
  (
    n746,
    n525
  );


  buf
  g634
  (
    n598,
    n538
  );


  buf
  g635
  (
    n611,
    n502
  );


  buf
  g636
  (
    n703,
    n523
  );


  not
  g637
  (
    n582,
    n222
  );


  buf
  g638
  (
    n643,
    n149
  );


  not
  g639
  (
    n719,
    n538
  );


  buf
  g640
  (
    n675,
    n557
  );


  buf
  g641
  (
    n592,
    n543
  );


  not
  g642
  (
    n660,
    n531
  );


  buf
  g643
  (
    n635,
    n514
  );


  not
  g644
  (
    n561,
    n248
  );


  buf
  g645
  (
    n594,
    n529
  );


  buf
  g646
  (
    n723,
    n508
  );


  not
  g647
  (
    n607,
    n160
  );


  buf
  g648
  (
    n745,
    n160
  );


  buf
  g649
  (
    n619,
    n538
  );


  buf
  g650
  (
    n676,
    n150
  );


  buf
  g651
  (
    n585,
    n157
  );


  buf
  g652
  (
    n605,
    n555
  );


  not
  g653
  (
    n655,
    n146
  );


  not
  g654
  (
    n560,
    n149
  );


  buf
  g655
  (
    n573,
    n151
  );


  buf
  g656
  (
    n776,
    n251
  );


  not
  g657
  (
    n621,
    n509
  );


  not
  g658
  (
    n656,
    n556
  );


  buf
  g659
  (
    n774,
    n520
  );


  not
  g660
  (
    n760,
    n537
  );


  buf
  g661
  (
    n733,
    n543
  );


  buf
  g662
  (
    n720,
    n551
  );


  buf
  g663
  (
    n578,
    n530
  );


  buf
  g664
  (
    n575,
    n558
  );


  not
  g665
  (
    n684,
    n232
  );


  buf
  g666
  (
    n762,
    n148
  );


  not
  g667
  (
    n704,
    n146
  );


  buf
  g668
  (
    KeyWire_0_47,
    n511
  );


  not
  g669
  (
    n648,
    n521
  );


  not
  g670
  (
    n627,
    n148
  );


  buf
  g671
  (
    n681,
    n151
  );


  buf
  g672
  (
    n576,
    n151
  );


  not
  g673
  (
    n647,
    n506
  );


  buf
  g674
  (
    n775,
    n532
  );


  buf
  g675
  (
    n640,
    n158
  );


  buf
  g676
  (
    n773,
    n522
  );


  not
  g677
  (
    n783,
    n549
  );


  buf
  g678
  (
    n728,
    n544
  );


  not
  g679
  (
    n688,
    n147
  );


  not
  g680
  (
    n744,
    n547
  );


  not
  g681
  (
    n606,
    n210
  );


  buf
  g682
  (
    n644,
    n523
  );


  not
  g683
  (
    n609,
    n230
  );


  buf
  g684
  (
    n669,
    n550
  );


  not
  g685
  (
    n608,
    n507
  );


  not
  g686
  (
    n642,
    n145
  );


  not
  g687
  (
    n665,
    n160
  );


  buf
  g688
  (
    KeyWire_0_61,
    n533
  );


  not
  g689
  (
    n711,
    n508
  );


  buf
  g690
  (
    n659,
    n533
  );


  buf
  g691
  (
    n761,
    n233
  );


  not
  g692
  (
    n736,
    n551
  );


  buf
  g693
  (
    n618,
    n534
  );


  not
  g694
  (
    n706,
    n532
  );


  not
  g695
  (
    n622,
    n517
  );


  buf
  g696
  (
    KeyWire_0_37,
    n505
  );


  buf
  g697
  (
    n767,
    n205
  );


  not
  g698
  (
    n693,
    n217
  );


  not
  g699
  (
    n678,
    n521
  );


  not
  g700
  (
    n624,
    n503
  );


  buf
  g701
  (
    n732,
    n544
  );


  buf
  g702
  (
    n666,
    n553
  );


  buf
  g703
  (
    n700,
    n518
  );


  not
  g704
  (
    n613,
    n553
  );


  not
  g705
  (
    n667,
    n528
  );


  not
  g706
  (
    n694,
    n503
  );


  buf
  g707
  (
    n718,
    n559
  );


  not
  g708
  (
    n739,
    n211
  );


  not
  g709
  (
    KeyWire_0_27,
    n534
  );


  buf
  g710
  (
    n587,
    n512
  );


  buf
  g711
  (
    n597,
    n504
  );


  buf
  g712
  (
    n564,
    n208
  );


  not
  g713
  (
    n586,
    n554
  );


  not
  g714
  (
    n565,
    n544
  );


  not
  g715
  (
    n651,
    n541
  );


  buf
  g716
  (
    n731,
    n158
  );


  buf
  g717
  (
    n596,
    n150
  );


  not
  g718
  (
    n610,
    n559
  );


  not
  g719
  (
    n753,
    n524
  );


  not
  g720
  (
    n788,
    n505
  );


  not
  g721
  (
    n715,
    n527
  );


  xor
  g722
  (
    n735,
    n502,
    n510,
    n507,
    n529
  );


  or
  g723
  (
    n571,
    n534,
    n517,
    n231,
    n156
  );


  xnor
  g724
  (
    n730,
    n155,
    n519,
    n512
  );


  nand
  g725
  (
    n789,
    n550,
    n546,
    n558,
    n518
  );


  nor
  g726
  (
    n664,
    n551,
    n158,
    n243,
    n503
  );


  xnor
  g727
  (
    n690,
    n508,
    n549,
    n227,
    n160
  );


  or
  g728
  (
    n614,
    n547,
    n540,
    n539,
    n252
  );


  xnor
  g729
  (
    n696,
    n525,
    n539,
    n218,
    n507
  );


  or
  g730
  (
    n771,
    n556,
    n244,
    n518,
    n509
  );


  xnor
  g731
  (
    KeyWire_0_1,
    n526,
    n533,
    n553,
    n530
  );


  xnor
  g732
  (
    n590,
    n504,
    n508,
    n221,
    n209
  );


  nor
  g733
  (
    n705,
    n215,
    n539,
    n510,
    n148
  );


  nand
  g734
  (
    KeyWire_0_44,
    n557,
    n529,
    n556,
    n225
  );


  xnor
  g735
  (
    n701,
    n520,
    n548,
    n528,
    n153
  );


  nand
  g736
  (
    n729,
    n532,
    n504,
    n152,
    n534
  );


  xnor
  g737
  (
    n740,
    n526,
    n557,
    n525,
    n154
  );


  and
  g738
  (
    n716,
    n226,
    n509,
    n229,
    n505
  );


  xnor
  g739
  (
    n601,
    n239,
    n552,
    n223,
    n546
  );


  nand
  g740
  (
    n682,
    n543,
    n147,
    n515,
    n540
  );


  and
  g741
  (
    n581,
    n236,
    n539,
    n524,
    n537
  );


  or
  g742
  (
    KeyWire_0_36,
    n234,
    n516,
    n204,
    n506
  );


  and
  g743
  (
    n683,
    n536,
    n552,
    n513,
    n549
  );


  xor
  g744
  (
    n577,
    n157,
    n525,
    n511,
    n554
  );


  xnor
  g745
  (
    n778,
    n220,
    n522,
    n154,
    n159
  );


  and
  g746
  (
    n650,
    n159,
    n542,
    n536,
    n546
  );


  xnor
  g747
  (
    n698,
    n527,
    n554,
    n520,
    n247
  );


  or
  g748
  (
    n787,
    n520,
    n542,
    n155,
    n533
  );


  xor
  g749
  (
    n707,
    n516,
    n537,
    n522,
    n150
  );


  nor
  g750
  (
    n722,
    n557,
    n519,
    n207,
    n149
  );


  xor
  g751
  (
    n769,
    n548,
    n515,
    n514,
    n542
  );


  xor
  g752
  (
    n765,
    n519,
    n546,
    n213,
    n549
  );


  or
  g753
  (
    n685,
    n558,
    n509,
    n529,
    n147
  );


  or
  g754
  (
    n569,
    n153,
    n535,
    n154,
    n246
  );


  and
  g755
  (
    n679,
    n545,
    n206,
    n535,
    n159
  );


  nor
  g756
  (
    n717,
    n545,
    n506,
    n547,
    n521
  );


  or
  g757
  (
    n599,
    n519,
    n538,
    n526,
    n532
  );


  and
  g758
  (
    n727,
    n152,
    n157,
    n153,
    n541
  );


  xnor
  g759
  (
    n800,
    n264,
    n267,
    n260,
    n561
  );


  or
  g760
  (
    n798,
    n259,
    n253,
    n261,
    n257
  );


  and
  g761
  (
    n801,
    n562,
    n256,
    n258,
    n281
  );


  xnor
  g762
  (
    n792,
    n255,
    n560,
    n566,
    n282
  );


  xor
  g763
  (
    n794,
    n254,
    n270,
    n567,
    n277
  );


  nor
  g764
  (
    n799,
    n279,
    n568,
    n274,
    n280
  );


  xnor
  g765
  (
    n796,
    n263,
    n276,
    n268,
    n278
  );


  xor
  g766
  (
    n793,
    n563,
    n273,
    n269,
    n266
  );


  nor
  g767
  (
    n797,
    n271,
    n262,
    n265,
    n564
  );


  xnor
  g768
  (
    n795,
    n565,
    n275,
    n272,
    n569
  );


  xnor
  g769
  (
    n802,
    n304,
    n795,
    n793
  );


  nor
  g770
  (
    n807,
    n294,
    n296,
    n285,
    n297
  );


  or
  g771
  (
    n805,
    n797,
    n305,
    n798,
    n299
  );


  xnor
  g772
  (
    n809,
    n283,
    n292,
    n796,
    n290
  );


  nand
  g773
  (
    n808,
    n298,
    n291,
    n792,
    n293
  );


  xnor
  g774
  (
    n804,
    n302,
    n289,
    n288,
    n287
  );


  xor
  g775
  (
    n803,
    n286,
    n295,
    n794,
    n301
  );


  nand
  g776
  (
    n806,
    n284,
    n300,
    n799,
    n303
  );


  and
  g777
  (
    n811,
    n306,
    n804,
    n585
  );


  or
  g778
  (
    n825,
    n584,
    n308,
    n318,
    n588
  );


  or
  g779
  (
    n827,
    n322,
    n598,
    n571,
    n586
  );


  and
  g780
  (
    KeyWire_0_17,
    n806,
    n591,
    n578,
    n594
  );


  nand
  g781
  (
    n823,
    n581,
    n579,
    n328,
    n320
  );


  nand
  g782
  (
    n812,
    n334,
    n333,
    n808,
    n329
  );


  and
  g783
  (
    n828,
    n590,
    n582,
    n600,
    n807
  );


  nand
  g784
  (
    n810,
    n574,
    n592,
    n593,
    n331
  );


  or
  g785
  (
    n821,
    n803,
    n332,
    n583,
    n317
  );


  nor
  g786
  (
    n817,
    n599,
    n325,
    n327,
    n806
  );


  xor
  g787
  (
    n826,
    n806,
    n807,
    n570,
    n804
  );


  nand
  g788
  (
    n819,
    n321,
    n307,
    n573,
    n805
  );


  xor
  g789
  (
    n814,
    n572,
    n802,
    n316,
    n804
  );


  nand
  g790
  (
    n824,
    n326,
    n319,
    n595,
    n597
  );


  nor
  g791
  (
    n820,
    n596,
    n310,
    n309,
    n587
  );


  xor
  g792
  (
    n815,
    n324,
    n311,
    n807,
    n330
  );


  xnor
  g793
  (
    n829,
    n805,
    n575,
    n576,
    n589
  );


  nand
  g794
  (
    KeyWire_0_9,
    n807,
    n315,
    n580,
    n314
  );


  and
  g795
  (
    n813,
    n806,
    n312,
    n577,
    n805
  );


  xnor
  g796
  (
    n822,
    n805,
    n323,
    n808,
    n313
  );


  buf
  g797
  (
    n835,
    n815
  );


  xnor
  g798
  (
    n832,
    n606,
    n601,
    n816
  );


  or
  g799
  (
    n834,
    n617,
    n613,
    n811,
    n615
  );


  xnor
  g800
  (
    n833,
    n814,
    n614,
    n612,
    n602
  );


  or
  g801
  (
    n830,
    n813,
    n609,
    n604,
    n603
  );


  nand
  g802
  (
    n836,
    n611,
    n605,
    n812,
    n610
  );


  nor
  g803
  (
    n831,
    n607,
    n810,
    n616,
    n608
  );


  or
  g804
  (
    n839,
    n359,
    n360,
    n414,
    n832
  );


  xnor
  g805
  (
    n863,
    n378,
    n830,
    n356,
    n382
  );


  xnor
  g806
  (
    n849,
    n396,
    n366,
    n835,
    n349
  );


  and
  g807
  (
    n842,
    n833,
    n836,
    n363,
    n348
  );


  nand
  g808
  (
    n855,
    n834,
    n834,
    n833,
    n402
  );


  or
  g809
  (
    n840,
    n338,
    n370,
    n388,
    n834
  );


  nand
  g810
  (
    n860,
    n832,
    n397,
    n835,
    n409
  );


  nor
  g811
  (
    n841,
    n369,
    n413,
    n350,
    n410
  );


  nor
  g812
  (
    n862,
    n831,
    n368,
    n383,
    n830
  );


  xor
  g813
  (
    n853,
    n358,
    n800,
    n831,
    n833
  );


  or
  g814
  (
    n846,
    n400,
    n381,
    n354,
    n362
  );


  nand
  g815
  (
    n854,
    n830,
    n618,
    n833,
    n365
  );


  and
  g816
  (
    n838,
    n831,
    n391,
    n364,
    n340
  );


  and
  g817
  (
    n858,
    n836,
    n386,
    n385,
    n404
  );


  xnor
  g818
  (
    n850,
    n373,
    n387,
    n412,
    n336
  );


  nor
  g819
  (
    n861,
    n380,
    n415,
    n394,
    n344
  );


  and
  g820
  (
    n847,
    n367,
    n384,
    n343,
    n353
  );


  or
  g821
  (
    n859,
    n361,
    n830,
    n832,
    n372
  );


  and
  g822
  (
    n843,
    n379,
    n836,
    n403
  );


  and
  g823
  (
    n844,
    n347,
    n835,
    n374,
    n834
  );


  nand
  g824
  (
    n852,
    n339,
    n352,
    n351,
    n389
  );


  nor
  g825
  (
    n845,
    n393,
    n371,
    n406,
    n831
  );


  nand
  g826
  (
    n857,
    n345,
    n832,
    n405,
    n355
  );


  xnor
  g827
  (
    n837,
    n408,
    n407,
    n375,
    n411
  );


  nand
  g828
  (
    n864,
    n337,
    n357,
    n335,
    n342
  );


  and
  g829
  (
    n856,
    n395,
    n399,
    n346,
    n377
  );


  nand
  g830
  (
    n851,
    n341,
    n392,
    n398,
    n390
  );


  xnor
  g831
  (
    n848,
    n801,
    n835,
    n376,
    n401
  );


  buf
  g832
  (
    n888,
    n668
  );


  nor
  g833
  (
    n918,
    n852,
    n631,
    n862
  );


  nand
  g834
  (
    n874,
    n718,
    n720,
    n749,
    n748
  );


  xor
  g835
  (
    n928,
    n630,
    n844,
    n750,
    n768
  );


  xnor
  g836
  (
    n909,
    n681,
    n773,
    n623,
    n420
  );


  nand
  g837
  (
    n919,
    n688,
    n767,
    n847,
    n427
  );


  nor
  g838
  (
    n956,
    n771,
    n762,
    n663,
    n637
  );


  or
  g839
  (
    n923,
    n864,
    n652,
    n849,
    n698
  );


  nor
  g840
  (
    n887,
    n762,
    n849,
    n640,
    n847
  );


  nand
  g841
  (
    n945,
    n856,
    n706,
    n862,
    n778
  );


  xor
  g842
  (
    n878,
    n662,
    n430,
    n771,
    n763
  );


  xnor
  g843
  (
    n957,
    n753,
    n840,
    n767,
    n778
  );


  nand
  g844
  (
    n898,
    n638,
    n808,
    n757
  );


  and
  g845
  (
    n910,
    n765,
    n762,
    n861,
    n703
  );


  xnor
  g846
  (
    n911,
    n633,
    n809,
    n770,
    n844
  );


  nor
  g847
  (
    n867,
    n723,
    n848,
    n760,
    n851
  );


  and
  g848
  (
    n931,
    n766,
    n656,
    n719,
    n624
  );


  or
  g849
  (
    n950,
    n851,
    n678,
    n657,
    n727
  );


  xnor
  g850
  (
    n866,
    n855,
    n845,
    n758,
    n632
  );


  nor
  g851
  (
    n944,
    n849,
    n748,
    n765,
    n661
  );


  xnor
  g852
  (
    n873,
    n760,
    n772,
    n858
  );


  or
  g853
  (
    n881,
    n680,
    n839,
    n682,
    n725
  );


  or
  g854
  (
    n930,
    n691,
    n772,
    n841,
    n416
  );


  xnor
  g855
  (
    n953,
    n643,
    n686,
    n672,
    n635
  );


  or
  g856
  (
    n902,
    n837,
    n844,
    n847,
    n753
  );


  and
  g857
  (
    n871,
    n759,
    n709,
    n626,
    n847
  );


  xor
  g858
  (
    n872,
    n694,
    n679,
    n646,
    n757
  );


  or
  g859
  (
    n883,
    n736,
    n738,
    n621,
    n619
  );


  or
  g860
  (
    n924,
    n728,
    n751,
    n642,
    n809
  );


  nor
  g861
  (
    n954,
    n735,
    n622,
    n777,
    n852
  );


  nand
  g862
  (
    n940,
    n775,
    n761,
    n770,
    n717
  );


  xnor
  g863
  (
    n896,
    n756,
    n769,
    n763,
    n740
  );


  xnor
  g864
  (
    KeyWire_0_51,
    n850,
    n864,
    n849,
    n726
  );


  xor
  g865
  (
    n899,
    n685,
    n776,
    n750,
    n739
  );


  and
  g866
  (
    n958,
    n846,
    n846,
    n701,
    n714
  );


  nand
  g867
  (
    n886,
    n757,
    n855,
    n628,
    n863
  );


  xor
  g868
  (
    n939,
    n705,
    n673,
    n751,
    n766
  );


  xnor
  g869
  (
    n891,
    n721,
    n687,
    n754,
    n434
  );


  nand
  g870
  (
    n885,
    n843,
    n425,
    n754,
    n692
  );


  xor
  g871
  (
    n935,
    n857,
    n764,
    n854,
    n752
  );


  nand
  g872
  (
    n892,
    n711,
    n629,
    n771,
    n755
  );


  nor
  g873
  (
    n920,
    n861,
    n649,
    n751,
    n423
  );


  and
  g874
  (
    n869,
    n763,
    n857,
    n733,
    n848
  );


  nor
  g875
  (
    KeyWire_0_34,
    n860,
    n859,
    n732,
    n704
  );


  or
  g876
  (
    KeyWire_0_7,
    n737,
    n758,
    n775,
    n769
  );


  or
  g877
  (
    n941,
    n845,
    n752,
    n769,
    n665
  );


  nor
  g878
  (
    n903,
    n856,
    n734,
    n660,
    n677
  );


  xnor
  g879
  (
    n922,
    n693,
    n777,
    n776,
    n764
  );


  nand
  g880
  (
    KeyWire_0_59,
    n641,
    n761,
    n684,
    n730
  );


  or
  g881
  (
    n908,
    n855,
    n758,
    n772,
    n417
  );


  nor
  g882
  (
    n895,
    n432,
    n768,
    n857,
    n696
  );


  xnor
  g883
  (
    n936,
    n777,
    n647,
    n750,
    n770
  );


  and
  g884
  (
    n925,
    n759,
    n761,
    n861,
    n757
  );


  or
  g885
  (
    n929,
    n770,
    n765,
    n846,
    n858
  );


  nand
  g886
  (
    n915,
    n768,
    n683,
    n748,
    n852
  );


  and
  g887
  (
    n875,
    n418,
    n864,
    n855,
    n653
  );


  nor
  g888
  (
    n949,
    n860,
    n856,
    n748,
    n774
  );


  nand
  g889
  (
    n877,
    n851,
    n743,
    n861,
    n722
  );


  xor
  g890
  (
    n890,
    n775,
    n741,
    n854,
    n769
  );


  and
  g891
  (
    n947,
    n809,
    n716,
    n843,
    n671
  );


  nor
  g892
  (
    n894,
    n654,
    n670,
    n854,
    n777
  );


  nor
  g893
  (
    n943,
    n845,
    n710,
    n772,
    n773
  );


  nor
  g894
  (
    n897,
    n700,
    n754,
    n699,
    n859
  );


  nor
  g895
  (
    n948,
    n659,
    n724,
    n667,
    n856
  );


  xor
  g896
  (
    n893,
    n763,
    n766,
    n863,
    n697
  );


  or
  g897
  (
    n951,
    n774,
    n774,
    n745,
    n854
  );


  nand
  g898
  (
    n932,
    n753,
    n676,
    n848,
    n634
  );


  or
  g899
  (
    n955,
    n429,
    n755,
    n845,
    n858
  );


  xnor
  g900
  (
    n905,
    n674,
    n636,
    n752,
    n755
  );


  nor
  g901
  (
    KeyWire_0_8,
    n760,
    n753,
    n853,
    n729
  );


  nor
  g902
  (
    KeyWire_0_60,
    n862,
    n707,
    n666,
    n744
  );


  xnor
  g903
  (
    n879,
    n695,
    n768,
    n850,
    n746
  );


  or
  g904
  (
    KeyWire_0_33,
    n860,
    n435,
    n863,
    n433
  );


  or
  g905
  (
    n942,
    n859,
    n760,
    n644,
    n648
  );


  and
  g906
  (
    n901,
    n842,
    n689,
    n690,
    n852
  );


  xor
  g907
  (
    n946,
    n431,
    n759,
    n771,
    n419
  );


  nor
  g908
  (
    n907,
    n421,
    n766,
    n853,
    n843
  );


  nor
  g909
  (
    n917,
    n863,
    n850,
    n761,
    n715
  );


  xor
  g910
  (
    n876,
    n620,
    n625,
    n860,
    n655
  );


  xor
  g911
  (
    n906,
    n756,
    n756,
    n750,
    n762
  );


  nor
  g912
  (
    n952,
    n742,
    n639,
    n749,
    n775
  );


  nand
  g913
  (
    n933,
    n731,
    n747,
    n658,
    n764
  );


  nor
  g914
  (
    KeyWire_0_18,
    n756,
    n759,
    n651,
    n708
  );


  xnor
  g915
  (
    n882,
    n749,
    n754,
    n645,
    n426
  );


  nand
  g916
  (
    n865,
    n853,
    n857,
    n755,
    n422
  );


  nand
  g917
  (
    n884,
    n774,
    n838,
    n424,
    n851
  );


  and
  g918
  (
    n934,
    n848,
    n853,
    n767,
    n864
  );


  nand
  g919
  (
    n926,
    n767,
    n773,
    n752,
    n844
  );


  nor
  g920
  (
    n921,
    n749,
    n712,
    n751,
    n669
  );


  xnor
  g921
  (
    n904,
    n664,
    n627,
    n843,
    n773
  );


  xor
  g922
  (
    n927,
    n778,
    n859,
    n765,
    n713
  );


  xnor
  g923
  (
    n870,
    n702,
    n428,
    n776,
    n764
  );


  nand
  g924
  (
    n938,
    n758,
    n776,
    n675,
    n809
  );


  xnor
  g925
  (
    n889,
    n846,
    n650,
    n862,
    n850
  );


  xnor
  g926
  (
    n962,
    n888,
    n823,
    n779,
    n819
  );


  and
  g927
  (
    n971,
    n886,
    n865,
    n873,
    n827
  );


  and
  g928
  (
    n985,
    n781,
    n820,
    n889,
    n875
  );


  xor
  g929
  (
    n981,
    n828,
    n785,
    n781,
    n823
  );


  xor
  g930
  (
    n966,
    n867,
    n871,
    n877,
    n827
  );


  xor
  g931
  (
    n976,
    n821,
    n779,
    n892,
    n818
  );


  and
  g932
  (
    n961,
    n783,
    n820,
    n822,
    n829
  );


  or
  g933
  (
    n984,
    n782,
    n780,
    n826,
    n883
  );


  nand
  g934
  (
    KeyWire_0_15,
    n825,
    n822,
    n878,
    n828
  );


  and
  g935
  (
    n964,
    n780,
    n782,
    n868,
    n872
  );


  xor
  g936
  (
    n975,
    n782,
    n784,
    n780
  );


  xnor
  g937
  (
    n982,
    n881,
    n825,
    n887,
    n828
  );


  xor
  g938
  (
    n973,
    n826,
    n869,
    n866,
    n885
  );


  and
  g939
  (
    n963,
    n825,
    n829,
    n779,
    n824
  );


  xor
  g940
  (
    KeyWire_0_48,
    n819,
    n820,
    n825,
    n778
  );


  and
  g941
  (
    n972,
    n821,
    n827,
    n786,
    n785
  );


  xor
  g942
  (
    n980,
    n876,
    n819,
    n781,
    n829
  );


  or
  g943
  (
    n978,
    n826,
    n824,
    n870,
    n786
  );


  or
  g944
  (
    n965,
    n817,
    n822,
    n820,
    n874
  );


  xnor
  g945
  (
    n960,
    n882,
    n824,
    n784,
    n786
  );


  or
  g946
  (
    n959,
    n824,
    n879,
    n819,
    n785
  );


  or
  g947
  (
    n983,
    n782,
    n783,
    n880,
    n784
  );


  nor
  g948
  (
    n967,
    n821,
    n884,
    n829,
    n828
  );


  xor
  g949
  (
    n969,
    n780,
    n783,
    n821,
    n890
  );


  nor
  g950
  (
    n977,
    n827,
    n779,
    n823,
    n781
  );


  or
  g951
  (
    n979,
    n826,
    n785,
    n891,
    n818
  );


  xnor
  g952
  (
    n968,
    n783,
    n823,
    n817,
    n822
  );


  nor
  g953
  (
    n991,
    n983,
    n789,
    n790,
    n791
  );


  and
  g954
  (
    n988,
    n790,
    n979,
    n787,
    n786
  );


  nand
  g955
  (
    KeyWire_0_11,
    n985,
    n984,
    n788,
    n787
  );


  and
  g956
  (
    n990,
    n790,
    n789,
    n788
  );


  xnor
  g957
  (
    n992,
    n787,
    n982,
    n790,
    n789
  );


  nor
  g958
  (
    n986,
    n787,
    n791,
    n981
  );


  or
  g959
  (
    n987,
    n789,
    n980,
    n791,
    n788
  );


  nor
  g960
  (
    n1010,
    n934,
    n473,
    n443,
    n988
  );


  and
  g961
  (
    n1001,
    n918,
    n902,
    n932,
    n990
  );


  xor
  g962
  (
    n1016,
    n469,
    n906,
    n927,
    n466
  );


  xnor
  g963
  (
    KeyWire_0_16,
    n447,
    n921,
    n450,
    n436
  );


  xnor
  g964
  (
    n1020,
    n438,
    n897,
    n986,
    n903
  );


  xor
  g965
  (
    n998,
    n938,
    n445,
    n454,
    n456
  );


  nand
  g966
  (
    n1008,
    n444,
    n989,
    n933,
    n987
  );


  or
  g967
  (
    n1014,
    n931,
    n986,
    n928,
    n452
  );


  or
  g968
  (
    n1013,
    n458,
    n987,
    n909,
    n913
  );


  xor
  g969
  (
    KeyWire_0_10,
    n992,
    n929,
    n900,
    n989
  );


  xor
  g970
  (
    n996,
    n992,
    n907,
    n926,
    n914
  );


  or
  g971
  (
    n1004,
    n895,
    n908,
    n453,
    n990
  );


  xnor
  g972
  (
    n1012,
    n986,
    n460,
    n440,
    n449
  );


  xor
  g973
  (
    n1009,
    n471,
    n991,
    n463,
    n457
  );


  or
  g974
  (
    n1000,
    n904,
    n922,
    n461,
    n992
  );


  nand
  g975
  (
    n994,
    n924,
    n989,
    n893,
    n990
  );


  nand
  g976
  (
    n1006,
    n991,
    n935,
    n451,
    n894
  );


  and
  g977
  (
    n1005,
    n986,
    n910,
    n465,
    n464
  );


  or
  g978
  (
    n997,
    n448,
    n916,
    n988,
    n919
  );


  xor
  g979
  (
    n995,
    n930,
    n467,
    n472,
    n988
  );


  nor
  g980
  (
    n1015,
    n987,
    n920,
    n437,
    n901
  );


  nand
  g981
  (
    n1007,
    n991,
    n468,
    n992,
    n459
  );


  nor
  g982
  (
    n1002,
    n989,
    n462,
    n470,
    n899
  );


  or
  g983
  (
    n1011,
    n915,
    n898,
    n991,
    n987
  );


  nor
  g984
  (
    n1003,
    n911,
    n442,
    n936,
    n990
  );


  xor
  g985
  (
    n1018,
    n912,
    n937,
    n439,
    n455
  );


  xor
  g986
  (
    n1017,
    n441,
    n925,
    n988,
    n446
  );


  nor
  g987
  (
    KeyWire_0_52,
    n923,
    n917,
    n896,
    n905
  );


  xor
  g988
  (
    KeyWire_0_49,
    n1002,
    n1012,
    n939,
    n949
  );


  or
  g989
  (
    n1023,
    n1020,
    n999,
    n1015,
    n1009
  );


  xor
  g990
  (
    n1024,
    n1018,
    n1011,
    n997,
    n947
  );


  nand
  g991
  (
    n1026,
    n993,
    n995,
    n943,
    n1019
  );


  nand
  g992
  (
    n1029,
    n953,
    n1014,
    n1004,
    n955
  );


  and
  g993
  (
    n1028,
    n1003,
    n1007,
    n944,
    n956
  );


  xnor
  g994
  (
    n1030,
    n1010,
    n940,
    n946,
    n941
  );


  xor
  g995
  (
    n1025,
    n996,
    n1006,
    n1008,
    n950
  );


  xnor
  g996
  (
    n1031,
    n1001,
    n945,
    n958,
    n948
  );


  xor
  g997
  (
    n1021,
    n998,
    n954,
    n994,
    n1017
  );


  nand
  g998
  (
    n1027,
    n1013,
    n1005,
    n1016,
    n951
  );


  nand
  g999
  (
    n1032,
    n1000,
    n957,
    n952,
    n942
  );


  xor
  KeyGate_0_0
  (
    n125,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n714,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n530,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n240,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n515,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n77,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n205,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n900,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n913,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n818,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n999,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n989,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n491,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n781,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n563,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n970,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n1019,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n816,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n880,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n272,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n465,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n466,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n71,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n632,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n44,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n43,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    n196,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n713,
    keyIn_0_27,
    KeyWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n401,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n274,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n49,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n249,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    n436,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n868,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n914,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n505,
    KeyNOTWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n579,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n768,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n118,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n334,
    KeyNOTWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n92,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n574,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    n371,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    n657,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n639,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n312,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n429,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n623,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n974,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n1022,
    KeyNOTWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    n366,
    keyIn_0_50,
    KeyWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n912,
    KeyNOTWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n993,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n708,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n232,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n330,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n278,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n458,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n275,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n916,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    n937,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n689,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n250,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n492,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

