

module Stat_1000_106
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1025,
  n1015,
  n1017,
  n1011,
  n1001,
  n1003,
  n1016,
  n1012,
  n1028,
  n1014,
  n1029,
  n1018,
  n1021,
  n1008,
  n1010,
  n1030,
  n1002,
  n1019,
  n1031,
  n1023,
  n1005,
  n1022,
  n1027,
  n1020,
  n1024,
  n1007,
  n1004,
  n1009,
  n1013,
  n1006,
  n1026,
  n1032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1025;output n1015;output n1017;output n1011;output n1001;output n1003;output n1016;output n1012;output n1028;output n1014;output n1029;output n1018;output n1021;output n1008;output n1010;output n1030;output n1002;output n1019;output n1031;output n1023;output n1005;output n1022;output n1027;output n1020;output n1024;output n1007;output n1004;output n1009;output n1013;output n1006;output n1026;output n1032;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyNOTWire_0_19;wire KeyWire_0_20;wire KeyNOTWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyNOTWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyNOTWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyNOTWire_0_27;wire KeyWire_0_28;wire KeyNOTWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyNOTWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  not
  g0
  (
    n83,
    n2
  );


  buf
  g1
  (
    n131,
    n27
  );


  not
  g2
  (
    n91,
    n5
  );


  not
  g3
  (
    n58,
    n14
  );


  not
  g4
  (
    n43,
    n25
  );


  buf
  g5
  (
    n112,
    n17
  );


  not
  g6
  (
    KeyWire_0_9,
    n24
  );


  buf
  g7
  (
    n74,
    n11
  );


  buf
  g8
  (
    n96,
    n16
  );


  not
  g9
  (
    n108,
    n5
  );


  not
  g10
  (
    n113,
    n4
  );


  buf
  g11
  (
    KeyWire_0_3,
    n18
  );


  not
  g12
  (
    n73,
    n10
  );


  buf
  g13
  (
    n82,
    n10
  );


  buf
  g14
  (
    n56,
    n9
  );


  buf
  g15
  (
    n98,
    n17
  );


  not
  g16
  (
    n38,
    n24
  );


  not
  g17
  (
    n125,
    n24
  );


  not
  g18
  (
    n88,
    n27
  );


  buf
  g19
  (
    n89,
    n3
  );


  buf
  g20
  (
    n84,
    n7
  );


  buf
  g21
  (
    n57,
    n21
  );


  buf
  g22
  (
    n50,
    n7
  );


  buf
  g23
  (
    n41,
    n18
  );


  not
  g24
  (
    n128,
    n23
  );


  not
  g25
  (
    n51,
    n4
  );


  not
  g26
  (
    n69,
    n1
  );


  not
  g27
  (
    n134,
    n25
  );


  buf
  g28
  (
    n42,
    n8
  );


  not
  g29
  (
    n92,
    n13
  );


  buf
  g30
  (
    n48,
    n9
  );


  buf
  g31
  (
    n85,
    n18
  );


  buf
  g32
  (
    n103,
    n25
  );


  buf
  g33
  (
    n52,
    n24
  );


  not
  g34
  (
    n126,
    n10
  );


  not
  g35
  (
    n70,
    n17
  );


  buf
  g36
  (
    n121,
    n5
  );


  buf
  g37
  (
    n100,
    n16
  );


  not
  g38
  (
    n127,
    n12
  );


  not
  g39
  (
    n101,
    n14
  );


  not
  g40
  (
    n35,
    n2
  );


  buf
  g41
  (
    n132,
    n9
  );


  not
  g42
  (
    n117,
    n6
  );


  not
  g43
  (
    n60,
    n18
  );


  buf
  g44
  (
    n63,
    n13
  );


  buf
  g45
  (
    n118,
    n7
  );


  not
  g46
  (
    n40,
    n22
  );


  not
  g47
  (
    n75,
    n19
  );


  buf
  g48
  (
    n95,
    n11
  );


  not
  g49
  (
    n93,
    n20
  );


  buf
  g50
  (
    n80,
    n26
  );


  buf
  g51
  (
    n122,
    n15
  );


  buf
  g52
  (
    n94,
    n10
  );


  not
  g53
  (
    n46,
    n26
  );


  not
  g54
  (
    KeyWire_0_8,
    n20
  );


  buf
  g55
  (
    n49,
    n5
  );


  buf
  g56
  (
    KeyWire_0_10,
    n6
  );


  buf
  g57
  (
    n55,
    n23
  );


  not
  g58
  (
    n107,
    n8
  );


  buf
  g59
  (
    n130,
    n2
  );


  buf
  g60
  (
    n54,
    n26
  );


  not
  g61
  (
    n36,
    n11
  );


  buf
  g62
  (
    n136,
    n1
  );


  not
  g63
  (
    n45,
    n14
  );


  not
  g64
  (
    n33,
    n14
  );


  buf
  g65
  (
    n62,
    n13
  );


  not
  g66
  (
    n138,
    n3
  );


  not
  g67
  (
    n116,
    n17
  );


  buf
  g68
  (
    n64,
    n1
  );


  buf
  g69
  (
    n99,
    n6
  );


  buf
  g70
  (
    n72,
    n21
  );


  not
  g71
  (
    n78,
    n9
  );


  buf
  g72
  (
    n71,
    n15
  );


  not
  g73
  (
    n97,
    n22
  );


  buf
  g74
  (
    n123,
    n20
  );


  buf
  g75
  (
    n104,
    n7
  );


  not
  g76
  (
    n53,
    n6
  );


  not
  g77
  (
    n44,
    n3
  );


  not
  g78
  (
    n90,
    n22
  );


  not
  g79
  (
    n87,
    n8
  );


  buf
  g80
  (
    n137,
    n1
  );


  not
  g81
  (
    n115,
    n12
  );


  not
  g82
  (
    n34,
    n22
  );


  buf
  g83
  (
    KeyWire_0_17,
    n16
  );


  not
  g84
  (
    n119,
    n3
  );


  not
  g85
  (
    n59,
    n16
  );


  not
  g86
  (
    n133,
    n19
  );


  not
  g87
  (
    n105,
    n8
  );


  not
  g88
  (
    n77,
    n11
  );


  not
  g89
  (
    n66,
    n12
  );


  not
  g90
  (
    n114,
    n26
  );


  buf
  g91
  (
    n135,
    n21
  );


  buf
  g92
  (
    n47,
    n4
  );


  buf
  g93
  (
    n124,
    n13
  );


  buf
  g94
  (
    n102,
    n19
  );


  buf
  g95
  (
    n37,
    n27
  );


  not
  g96
  (
    n129,
    n15
  );


  buf
  g97
  (
    n86,
    n12
  );


  buf
  g98
  (
    n81,
    n19
  );


  buf
  g99
  (
    n109,
    n2
  );


  not
  g100
  (
    n111,
    n4
  );


  buf
  g101
  (
    n79,
    n20
  );


  not
  g102
  (
    n76,
    n25
  );


  not
  g103
  (
    n39,
    n15
  );


  buf
  g104
  (
    n139,
    n23
  );


  buf
  g105
  (
    n120,
    n23
  );


  not
  g106
  (
    n110,
    n21
  );


  not
  g107
  (
    n243,
    n59
  );


  buf
  g108
  (
    n256,
    n67
  );


  not
  g109
  (
    n250,
    n39
  );


  not
  g110
  (
    n192,
    n43
  );


  buf
  g111
  (
    n206,
    n49
  );


  buf
  g112
  (
    n236,
    n48
  );


  buf
  g113
  (
    n194,
    n44
  );


  buf
  g114
  (
    n176,
    n66
  );


  buf
  g115
  (
    n159,
    n39
  );


  not
  g116
  (
    n254,
    n59
  );


  buf
  g117
  (
    n149,
    n62
  );


  not
  g118
  (
    n252,
    n34
  );


  buf
  g119
  (
    n189,
    n47
  );


  not
  g120
  (
    n269,
    n42
  );


  buf
  g121
  (
    n185,
    n61
  );


  not
  g122
  (
    n188,
    n51
  );


  not
  g123
  (
    n164,
    n48
  );


  not
  g124
  (
    n181,
    n50
  );


  not
  g125
  (
    n230,
    n56
  );


  buf
  g126
  (
    n210,
    n45
  );


  not
  g127
  (
    n268,
    n54
  );


  not
  g128
  (
    n169,
    n51
  );


  not
  g129
  (
    n179,
    n34
  );


  not
  g130
  (
    n193,
    n60
  );


  buf
  g131
  (
    n251,
    n63
  );


  not
  g132
  (
    n270,
    n55
  );


  buf
  g133
  (
    n148,
    n38
  );


  not
  g134
  (
    n143,
    n60
  );


  buf
  g135
  (
    n224,
    n50
  );


  buf
  g136
  (
    n258,
    n51
  );


  not
  g137
  (
    n240,
    n47
  );


  buf
  g138
  (
    n198,
    n59
  );


  not
  g139
  (
    n233,
    n41
  );


  not
  g140
  (
    n196,
    n62
  );


  not
  g141
  (
    n219,
    n61
  );


  buf
  g142
  (
    n199,
    n42
  );


  not
  g143
  (
    n271,
    n37
  );


  buf
  g144
  (
    n190,
    n66
  );


  not
  g145
  (
    n223,
    n33
  );


  buf
  g146
  (
    n217,
    n63
  );


  not
  g147
  (
    n226,
    n45
  );


  not
  g148
  (
    n182,
    n43
  );


  not
  g149
  (
    n204,
    n33
  );


  buf
  g150
  (
    n225,
    n38
  );


  not
  g151
  (
    n142,
    n43
  );


  not
  g152
  (
    n170,
    n44
  );


  not
  g153
  (
    n153,
    n35
  );


  buf
  g154
  (
    n146,
    n57
  );


  buf
  g155
  (
    n231,
    n49
  );


  buf
  g156
  (
    n178,
    n63
  );


  buf
  g157
  (
    n241,
    n35
  );


  buf
  g158
  (
    n168,
    n57
  );


  buf
  g159
  (
    n274,
    n53
  );


  buf
  g160
  (
    n202,
    n34
  );


  buf
  g161
  (
    n266,
    n58
  );


  buf
  g162
  (
    n247,
    n52
  );


  not
  g163
  (
    n200,
    n59
  );


  buf
  g164
  (
    n261,
    n62
  );


  not
  g165
  (
    KeyWire_0_27,
    n55
  );


  buf
  g166
  (
    n175,
    n36
  );


  buf
  g167
  (
    n228,
    n36
  );


  buf
  g168
  (
    n141,
    n49
  );


  not
  g169
  (
    n272,
    n53
  );


  buf
  g170
  (
    n155,
    n64
  );


  buf
  g171
  (
    n215,
    n52
  );


  not
  g172
  (
    n246,
    n45
  );


  buf
  g173
  (
    n201,
    n61
  );


  buf
  g174
  (
    n203,
    n39
  );


  buf
  g175
  (
    n197,
    n46
  );


  buf
  g176
  (
    n151,
    n62
  );


  buf
  g177
  (
    n145,
    n40
  );


  buf
  g178
  (
    n187,
    n58
  );


  buf
  g179
  (
    n273,
    n38
  );


  not
  g180
  (
    n162,
    n61
  );


  buf
  g181
  (
    n275,
    n33
  );


  not
  g182
  (
    n173,
    n36
  );


  not
  g183
  (
    n158,
    n42
  );


  buf
  g184
  (
    n166,
    n56
  );


  not
  g185
  (
    n213,
    n51
  );


  buf
  g186
  (
    n232,
    n35
  );


  not
  g187
  (
    n220,
    n55
  );


  buf
  g188
  (
    KeyWire_0_12,
    n53
  );


  buf
  g189
  (
    n238,
    n39
  );


  not
  g190
  (
    n237,
    n56
  );


  not
  g191
  (
    n174,
    n37
  );


  not
  g192
  (
    n244,
    n53
  );


  buf
  g193
  (
    n234,
    n54
  );


  buf
  g194
  (
    n257,
    n54
  );


  buf
  g195
  (
    n160,
    n34
  );


  buf
  g196
  (
    n183,
    n64
  );


  buf
  g197
  (
    n191,
    n35
  );


  not
  g198
  (
    n267,
    n33
  );


  not
  g199
  (
    n264,
    n65
  );


  buf
  g200
  (
    n150,
    n64
  );


  buf
  g201
  (
    n209,
    n67
  );


  not
  g202
  (
    n156,
    n50
  );


  not
  g203
  (
    n195,
    n55
  );


  buf
  g204
  (
    n205,
    n46
  );


  not
  g205
  (
    n140,
    n52
  );


  not
  g206
  (
    n180,
    n41
  );


  not
  g207
  (
    n255,
    n64
  );


  not
  g208
  (
    n227,
    n42
  );


  buf
  g209
  (
    n157,
    n66
  );


  buf
  g210
  (
    n167,
    n44
  );


  buf
  g211
  (
    n242,
    n46
  );


  buf
  g212
  (
    n212,
    n36
  );


  not
  g213
  (
    n260,
    n57
  );


  buf
  g214
  (
    n249,
    n38
  );


  buf
  g215
  (
    n265,
    n58
  );


  not
  g216
  (
    n184,
    n52
  );


  buf
  g217
  (
    n154,
    n40
  );


  not
  g218
  (
    n207,
    n60
  );


  buf
  g219
  (
    n177,
    n47
  );


  buf
  g220
  (
    n239,
    n47
  );


  not
  g221
  (
    n259,
    n63
  );


  buf
  g222
  (
    n263,
    n65
  );


  buf
  g223
  (
    n253,
    n56
  );


  not
  g224
  (
    n171,
    n57
  );


  buf
  g225
  (
    n161,
    n65
  );


  buf
  g226
  (
    n163,
    n45
  );


  not
  g227
  (
    n211,
    n46
  );


  buf
  g228
  (
    n218,
    n48
  );


  buf
  g229
  (
    n147,
    n41
  );


  buf
  g230
  (
    n222,
    n43
  );


  buf
  g231
  (
    n245,
    n40
  );


  buf
  g232
  (
    n186,
    n44
  );


  not
  g233
  (
    n208,
    n41
  );


  buf
  g234
  (
    n248,
    n37
  );


  buf
  g235
  (
    n172,
    n66
  );


  buf
  g236
  (
    n235,
    n40
  );


  buf
  g237
  (
    n216,
    n54
  );


  buf
  g238
  (
    n221,
    n48
  );


  not
  g239
  (
    n276,
    n37
  );


  not
  g240
  (
    n144,
    n50
  );


  buf
  g241
  (
    n214,
    n49
  );


  buf
  g242
  (
    n277,
    n67
  );


  buf
  g243
  (
    n229,
    n67
  );


  nand
  g244
  (
    n165,
    n60,
    n65,
    n58
  );


  not
  g245
  (
    n346,
    n190
  );


  buf
  g246
  (
    n293,
    n140
  );


  not
  g247
  (
    n378,
    n197
  );


  buf
  g248
  (
    n440,
    n155
  );


  buf
  g249
  (
    n425,
    n199
  );


  buf
  g250
  (
    n287,
    n201
  );


  buf
  g251
  (
    n393,
    n195
  );


  buf
  g252
  (
    n380,
    n175
  );


  buf
  g253
  (
    n381,
    n143
  );


  buf
  g254
  (
    n323,
    n167
  );


  not
  g255
  (
    n412,
    n171
  );


  not
  g256
  (
    n288,
    n184
  );


  buf
  g257
  (
    n413,
    n222
  );


  not
  g258
  (
    n354,
    n223
  );


  buf
  g259
  (
    n309,
    n213
  );


  not
  g260
  (
    n329,
    n201
  );


  not
  g261
  (
    n363,
    n164
  );


  buf
  g262
  (
    n297,
    n213
  );


  not
  g263
  (
    n321,
    n207
  );


  not
  g264
  (
    n331,
    n207
  );


  not
  g265
  (
    n342,
    n177
  );


  buf
  g266
  (
    n372,
    n198
  );


  not
  g267
  (
    n326,
    n162
  );


  buf
  g268
  (
    n348,
    n182
  );


  buf
  g269
  (
    n357,
    n202
  );


  not
  g270
  (
    n295,
    n210
  );


  not
  g271
  (
    n285,
    n170
  );


  buf
  g272
  (
    n324,
    n207
  );


  buf
  g273
  (
    n399,
    n143
  );


  buf
  g274
  (
    n286,
    n166
  );


  not
  g275
  (
    n426,
    n218
  );


  not
  g276
  (
    n401,
    n163
  );


  buf
  g277
  (
    n396,
    n144
  );


  not
  g278
  (
    n388,
    n195
  );


  not
  g279
  (
    n435,
    n166
  );


  buf
  g280
  (
    KeyWire_0_14,
    n214
  );


  not
  g281
  (
    n402,
    n205
  );


  buf
  g282
  (
    n283,
    n208
  );


  buf
  g283
  (
    n409,
    n174
  );


  not
  g284
  (
    n289,
    n161
  );


  buf
  g285
  (
    n300,
    n177
  );


  not
  g286
  (
    n368,
    n219
  );


  not
  g287
  (
    n345,
    n208
  );


  buf
  g288
  (
    n392,
    n169
  );


  buf
  g289
  (
    n318,
    n206
  );


  buf
  g290
  (
    n296,
    n195
  );


  buf
  g291
  (
    n405,
    n178
  );


  buf
  g292
  (
    n379,
    n202
  );


  not
  g293
  (
    n366,
    n147
  );


  not
  g294
  (
    n386,
    n151
  );


  buf
  g295
  (
    n374,
    n218
  );


  buf
  g296
  (
    n410,
    n143
  );


  buf
  g297
  (
    n391,
    n175
  );


  buf
  g298
  (
    n437,
    n168
  );


  buf
  g299
  (
    n302,
    n211
  );


  not
  g300
  (
    n427,
    n206
  );


  buf
  g301
  (
    n330,
    n178
  );


  not
  g302
  (
    n433,
    n183
  );


  buf
  g303
  (
    n281,
    n141
  );


  buf
  g304
  (
    n347,
    n170
  );


  not
  g305
  (
    n404,
    n171
  );


  buf
  g306
  (
    n403,
    n172
  );


  not
  g307
  (
    n284,
    n164
  );


  not
  g308
  (
    n350,
    n205
  );


  not
  g309
  (
    n279,
    n159
  );


  buf
  g310
  (
    n290,
    n169
  );


  buf
  g311
  (
    n292,
    n186
  );


  buf
  g312
  (
    n304,
    n209
  );


  not
  g313
  (
    n351,
    n191
  );


  buf
  g314
  (
    n317,
    n198
  );


  not
  g315
  (
    n428,
    n146
  );


  not
  g316
  (
    n398,
    n215
  );


  not
  g317
  (
    n438,
    n215
  );


  buf
  g318
  (
    n308,
    n200
  );


  buf
  g319
  (
    n387,
    n224
  );


  not
  g320
  (
    n430,
    n151
  );


  buf
  g321
  (
    n316,
    n210
  );


  not
  g322
  (
    KeyWire_0_4,
    n153
  );


  not
  g323
  (
    n376,
    n149
  );


  buf
  g324
  (
    n422,
    n204
  );


  not
  g325
  (
    n360,
    n176
  );


  buf
  g326
  (
    n307,
    n207
  );


  not
  g327
  (
    n335,
    n167
  );


  buf
  g328
  (
    n334,
    n199
  );


  not
  g329
  (
    KeyWire_0_0,
    n155
  );


  not
  g330
  (
    n406,
    n192
  );


  not
  g331
  (
    n312,
    n141
  );


  not
  g332
  (
    n358,
    n153
  );


  buf
  g333
  (
    n371,
    n190
  );


  buf
  g334
  (
    n408,
    n143
  );


  buf
  g335
  (
    n315,
    n158
  );


  buf
  g336
  (
    n415,
    n184
  );


  buf
  g337
  (
    n336,
    n189
  );


  not
  g338
  (
    n414,
    n185
  );


  not
  g339
  (
    n299,
    n159
  );


  buf
  g340
  (
    KeyWire_0_19,
    n174
  );


  buf
  g341
  (
    n337,
    n176
  );


  buf
  g342
  (
    n306,
    n140
  );


  buf
  g343
  (
    n352,
    n216
  );


  not
  g344
  (
    n361,
    n153
  );


  not
  g345
  (
    n322,
    n170
  );


  not
  g346
  (
    n369,
    n191
  );


  not
  g347
  (
    n384,
    n219
  );


  not
  g348
  (
    n441,
    n169
  );


  buf
  g349
  (
    n349,
    n210
  );


  and
  g350
  (
    n390,
    n214,
    n172,
    n142,
    n160
  );


  nor
  g351
  (
    n340,
    n161,
    n223,
    n173,
    n189
  );


  xor
  g352
  (
    n421,
    n145,
    n175,
    n217,
    n167
  );


  nor
  g353
  (
    n434,
    n156,
    n141,
    n168,
    n167
  );


  nor
  g354
  (
    n431,
    n215,
    n163,
    n180,
    n192
  );


  or
  g355
  (
    n355,
    n216,
    n185,
    n158,
    n194
  );


  or
  g356
  (
    KeyWire_0_16,
    n148,
    n174,
    n180
  );


  xor
  g357
  (
    n278,
    n162,
    n166,
    n142,
    n221
  );


  xnor
  g358
  (
    n389,
    n209,
    n205,
    n169,
    n204
  );


  nand
  g359
  (
    KeyWire_0_22,
    n218,
    n178,
    n212,
    n163
  );


  xnor
  g360
  (
    n432,
    n190,
    n162,
    n177,
    n205
  );


  xnor
  g361
  (
    n400,
    n221,
    n217,
    n197,
    n220
  );


  xnor
  g362
  (
    n377,
    n199,
    n213,
    n186,
    n194
  );


  xor
  g363
  (
    n375,
    n212,
    n140,
    n171,
    n190
  );


  and
  g364
  (
    n301,
    n200,
    n146,
    n151,
    n224
  );


  nand
  g365
  (
    KeyWire_0_2,
    n164,
    n224,
    n218,
    n148
  );


  nor
  g366
  (
    n310,
    n188,
    n196,
    n183
  );


  or
  g367
  (
    n436,
    n144,
    n188,
    n154,
    n165
  );


  nand
  g368
  (
    n294,
    n224,
    n188,
    n163,
    n221
  );


  xor
  g369
  (
    n311,
    n200,
    n181,
    n206,
    n144
  );


  or
  g370
  (
    n344,
    n211,
    n185,
    n177
  );


  and
  g371
  (
    n423,
    n145,
    n179,
    n152,
    n172
  );


  nand
  g372
  (
    n338,
    n141,
    n161,
    n225,
    n220
  );


  xor
  g373
  (
    n327,
    n198,
    n217,
    n159,
    n154
  );


  xnor
  g374
  (
    n418,
    n223,
    n145,
    n157,
    n156
  );


  and
  g375
  (
    n407,
    n196,
    n151,
    n192,
    n154
  );


  xor
  g376
  (
    n411,
    n159,
    n173,
    n211,
    n181
  );


  and
  g377
  (
    n319,
    n222,
    n176,
    n158,
    n208
  );


  xor
  g378
  (
    n439,
    n150,
    n179,
    n201,
    n152
  );


  nor
  g379
  (
    n314,
    n217,
    n183,
    n155,
    n158
  );


  nor
  g380
  (
    n373,
    n216,
    n204,
    n154,
    n165
  );


  or
  g381
  (
    n429,
    n219,
    n161,
    n146,
    n170
  );


  nor
  g382
  (
    n320,
    n212,
    n187,
    n209,
    n175
  );


  and
  g383
  (
    n365,
    n146,
    n214,
    n165,
    n193
  );


  xor
  g384
  (
    n332,
    n142,
    n199,
    n182,
    n193
  );


  xnor
  g385
  (
    n328,
    n165,
    n219,
    n220,
    n203
  );


  or
  g386
  (
    n280,
    n179,
    n197,
    n149,
    n187
  );


  nor
  g387
  (
    n353,
    n194,
    n194,
    n142,
    n157
  );


  nor
  g388
  (
    n416,
    n208,
    n168,
    n150
  );


  and
  g389
  (
    n367,
    n225,
    n179,
    n168,
    n203
  );


  and
  g390
  (
    n305,
    n181,
    n153,
    n222,
    n186
  );


  nand
  g391
  (
    n370,
    n209,
    n164,
    n192,
    n204
  );


  nor
  g392
  (
    n364,
    n213,
    n223,
    n176,
    n160
  );


  xor
  g393
  (
    n385,
    n187,
    n182,
    n166,
    n160
  );


  and
  g394
  (
    n382,
    n184,
    n195,
    n173,
    n156
  );


  and
  g395
  (
    n313,
    n203,
    n172,
    n201,
    n145
  );


  nor
  g396
  (
    n397,
    n152,
    n221,
    n156,
    n174
  );


  or
  g397
  (
    n303,
    n171,
    n203,
    n197,
    n150
  );


  nor
  g398
  (
    n417,
    n140,
    n188,
    n196,
    n215
  );


  xnor
  g399
  (
    n362,
    n152,
    n149,
    n202,
    n220
  );


  xor
  g400
  (
    n424,
    n157,
    n144,
    n147,
    n206
  );


  xnor
  g401
  (
    n282,
    n222,
    n182,
    n155,
    n225
  );


  nand
  g402
  (
    n359,
    n212,
    n200,
    n193,
    n191
  );


  nor
  g403
  (
    n341,
    n148,
    n226,
    n181,
    n157
  );


  xnor
  g404
  (
    KeyWire_0_28,
    n210,
    n160,
    n211,
    n180
  );


  or
  g405
  (
    n325,
    n198,
    n216,
    n147,
    n202
  );


  nand
  g406
  (
    n420,
    n178,
    n193,
    n225,
    n189
  );


  xnor
  g407
  (
    n339,
    n183,
    n187,
    n147,
    n186
  );


  nand
  g408
  (
    n383,
    n149,
    n162,
    n173,
    n148
  );


  xnor
  g409
  (
    n298,
    n191,
    n189,
    n184,
    n214
  );


  buf
  g410
  (
    n449,
    n279
  );


  buf
  g411
  (
    n447,
    n280
  );


  buf
  g412
  (
    n452,
    n283
  );


  buf
  g413
  (
    n451,
    n281
  );


  buf
  g414
  (
    n444,
    n279
  );


  not
  g415
  (
    n450,
    n281
  );


  nand
  g416
  (
    n445,
    n278,
    n283
  );


  xnor
  g417
  (
    n454,
    n281,
    n280,
    n282,
    n284
  );


  xnor
  g418
  (
    n446,
    n279,
    n283,
    n278,
    n284
  );


  nand
  g419
  (
    n448,
    n279,
    n284,
    n281,
    n278
  );


  xnor
  g420
  (
    n453,
    n282,
    n278,
    n280
  );


  xor
  g421
  (
    n443,
    n282,
    n282,
    n284,
    n283
  );


  not
  g422
  (
    n500,
    n447
  );


  not
  g423
  (
    n483,
    n449
  );


  buf
  g424
  (
    n480,
    n451
  );


  not
  g425
  (
    n460,
    n445
  );


  buf
  g426
  (
    n495,
    n444
  );


  buf
  g427
  (
    n501,
    n448
  );


  not
  g428
  (
    n468,
    n444
  );


  buf
  g429
  (
    n466,
    n450
  );


  not
  g430
  (
    KeyWire_0_26,
    n446
  );


  not
  g431
  (
    n467,
    n451
  );


  buf
  g432
  (
    n462,
    n454
  );


  not
  g433
  (
    n490,
    n448
  );


  not
  g434
  (
    KeyWire_0_21,
    n454
  );


  not
  g435
  (
    n482,
    n444
  );


  not
  g436
  (
    n472,
    n445
  );


  not
  g437
  (
    n463,
    n447
  );


  not
  g438
  (
    n461,
    n454
  );


  buf
  g439
  (
    n479,
    n450
  );


  buf
  g440
  (
    n469,
    n450
  );


  buf
  g441
  (
    n494,
    n452
  );


  buf
  g442
  (
    n478,
    n453
  );


  buf
  g443
  (
    n470,
    n446
  );


  not
  g444
  (
    n458,
    n445
  );


  not
  g445
  (
    n456,
    n443
  );


  not
  g446
  (
    n485,
    n447
  );


  buf
  g447
  (
    n457,
    n452
  );


  buf
  g448
  (
    n496,
    n446
  );


  not
  g449
  (
    n491,
    n448
  );


  not
  g450
  (
    n459,
    n449
  );


  not
  g451
  (
    n473,
    n449
  );


  not
  g452
  (
    n489,
    n443
  );


  not
  g453
  (
    n499,
    n451
  );


  buf
  g454
  (
    n486,
    n453
  );


  buf
  g455
  (
    n465,
    n447
  );


  not
  g456
  (
    n475,
    n448
  );


  buf
  g457
  (
    n464,
    n453
  );


  not
  g458
  (
    n484,
    n445
  );


  not
  g459
  (
    KeyWire_0_1,
    n443
  );


  buf
  g460
  (
    n498,
    n446
  );


  not
  g461
  (
    n493,
    n451
  );


  buf
  g462
  (
    n502,
    n452
  );


  buf
  g463
  (
    n476,
    n444
  );


  not
  g464
  (
    n488,
    n450
  );


  buf
  g465
  (
    n474,
    n453
  );


  not
  g466
  (
    n487,
    n454
  );


  not
  g467
  (
    n455,
    n452
  );


  not
  g468
  (
    n481,
    n449
  );


  not
  g469
  (
    n492,
    n443
  );


  or
  g470
  (
    n511,
    n297,
    n456,
    n381,
    n473
  );


  and
  g471
  (
    n677,
    n461,
    n358,
    n382,
    n399
  );


  or
  g472
  (
    n669,
    n349,
    n327,
    n468,
    n489
  );


  and
  g473
  (
    n565,
    n378,
    n465,
    n489,
    n391
  );


  nand
  g474
  (
    n660,
    n324,
    n378,
    n379,
    n356
  );


  nand
  g475
  (
    n693,
    n387,
    n368,
    n498,
    n420
  );


  xor
  g476
  (
    n662,
    n328,
    n482,
    n300,
    n404
  );


  or
  g477
  (
    n563,
    n298,
    n410,
    n288,
    n348
  );


  and
  g478
  (
    n685,
    n425,
    n488,
    n292,
    n377
  );


  nor
  g479
  (
    n658,
    n416,
    n370,
    n393,
    n337
  );


  xor
  g480
  (
    n626,
    n335,
    n390,
    n397,
    n465
  );


  xor
  g481
  (
    n672,
    n408,
    n312,
    n369,
    n372
  );


  nand
  g482
  (
    n525,
    n467,
    n322,
    n482,
    n410
  );


  xnor
  g483
  (
    n536,
    n387,
    n318,
    n334,
    n412
  );


  xor
  g484
  (
    n668,
    n387,
    n287,
    n497,
    n399
  );


  xor
  g485
  (
    n692,
    n354,
    n411,
    n457,
    n405
  );


  xor
  g486
  (
    n583,
    n460,
    n422,
    n417,
    n311
  );


  xor
  g487
  (
    n684,
    n327,
    n325,
    n350,
    n304
  );


  nor
  g488
  (
    n593,
    n482,
    n455,
    n419,
    n489
  );


  and
  g489
  (
    n682,
    n373,
    n352,
    n381,
    n426
  );


  xnor
  g490
  (
    n575,
    n500,
    n416,
    n423,
    n358
  );


  and
  g491
  (
    n554,
    n392,
    n478,
    n373,
    n405
  );


  or
  g492
  (
    n582,
    n309,
    n325,
    n318,
    n413
  );


  and
  g493
  (
    n592,
    n293,
    n480,
    n493,
    n364
  );


  nand
  g494
  (
    n504,
    n331,
    n481,
    n415,
    n459
  );


  xnor
  g495
  (
    n671,
    n410,
    n334,
    n302,
    n348
  );


  and
  g496
  (
    n581,
    n371,
    n359,
    n410,
    n415
  );


  nand
  g497
  (
    KeyWire_0_18,
    n485,
    n459,
    n334,
    n303
  );


  and
  g498
  (
    n580,
    n379,
    n478,
    n475
  );


  and
  g499
  (
    n683,
    n343,
    n400,
    n377,
    n305
  );


  nand
  g500
  (
    n674,
    n378,
    n390,
    n350,
    n363
  );


  xor
  g501
  (
    n609,
    n287,
    n396,
    n369,
    n388
  );


  xor
  g502
  (
    n527,
    n414,
    n404,
    n418,
    n317
  );


  xor
  g503
  (
    n624,
    n414,
    n402,
    n383,
    n487
  );


  nand
  g504
  (
    n586,
    n466,
    n460,
    n413,
    n294
  );


  or
  g505
  (
    n577,
    n380,
    n317,
    n340,
    n498
  );


  xnor
  g506
  (
    n571,
    n357,
    n316,
    n427,
    n313
  );


  or
  g507
  (
    KeyWire_0_20,
    n292,
    n386,
    n391,
    n392
  );


  or
  g508
  (
    n566,
    n289,
    n420,
    n455,
    n490
  );


  and
  g509
  (
    n572,
    n300,
    n331,
    n330,
    n359
  );


  xor
  g510
  (
    n646,
    n331,
    n411,
    n409,
    n367
  );


  nand
  g511
  (
    n588,
    n477,
    n491,
    n333,
    n362
  );


  xor
  g512
  (
    n618,
    n477,
    n295,
    n297,
    n476
  );


  nor
  g513
  (
    n568,
    n455,
    n390,
    n298,
    n480
  );


  nand
  g514
  (
    KeyWire_0_30,
    n491,
    n394,
    n360,
    n401
  );


  xnor
  g515
  (
    n616,
    n472,
    n344,
    n301,
    n363
  );


  and
  g516
  (
    n515,
    n365,
    n345,
    n481,
    n323
  );


  nor
  g517
  (
    n613,
    n468,
    n398,
    n353,
    n470
  );


  xor
  g518
  (
    n644,
    n307,
    n461,
    n285,
    n496
  );


  or
  g519
  (
    n679,
    n474,
    n343,
    n425,
    n389
  );


  or
  g520
  (
    n555,
    n375,
    n317,
    n495,
    n365
  );


  and
  g521
  (
    n610,
    n403,
    n377,
    n292,
    n476
  );


  xnor
  g522
  (
    n622,
    n358,
    n472,
    n400,
    n323
  );


  nor
  g523
  (
    n558,
    n294,
    n322,
    n290,
    n339
  );


  nand
  g524
  (
    n638,
    n291,
    n346,
    n333,
    n377
  );


  nor
  g525
  (
    n600,
    n499,
    n456,
    n459,
    n358
  );


  nand
  g526
  (
    n508,
    n412,
    n427,
    n476,
    n479
  );


  xor
  g527
  (
    n512,
    n299,
    n380,
    n296,
    n499
  );


  or
  g528
  (
    n579,
    n402,
    n404,
    n341,
    n348
  );


  nor
  g529
  (
    n510,
    n492,
    n419,
    n479,
    n413
  );


  xor
  g530
  (
    n604,
    n318,
    n341,
    n325,
    n285
  );


  and
  g531
  (
    n630,
    n311,
    n466,
    n490,
    n363
  );


  nor
  g532
  (
    n559,
    n399,
    n473,
    n497
  );


  nand
  g533
  (
    n547,
    n493,
    n355,
    n471,
    n408
  );


  nand
  g534
  (
    n553,
    n361,
    n294,
    n380,
    n463
  );


  or
  g535
  (
    n657,
    n473,
    n320,
    n313,
    n456
  );


  or
  g536
  (
    n631,
    n301,
    n288,
    n374,
    n332
  );


  and
  g537
  (
    n540,
    n361,
    n291,
    n344,
    n401
  );


  nand
  g538
  (
    n544,
    n501,
    n475,
    n320,
    n288
  );


  xnor
  g539
  (
    n615,
    n481,
    n495,
    n389,
    n295
  );


  and
  g540
  (
    n552,
    n298,
    n326,
    n486,
    n398
  );


  nand
  g541
  (
    n584,
    n455,
    n401,
    n311,
    n352
  );


  nand
  g542
  (
    n641,
    n462,
    n375,
    n285,
    n314
  );


  xnor
  g543
  (
    n594,
    n467,
    n360,
    n352,
    n424
  );


  nand
  g544
  (
    n590,
    n367,
    n496,
    n493,
    n321
  );


  xor
  g545
  (
    n611,
    n390,
    n492,
    n471,
    n402
  );


  nand
  g546
  (
    n526,
    n353,
    n461,
    n296,
    n308
  );


  nand
  g547
  (
    n620,
    n344,
    n406,
    n322,
    n494
  );


  nor
  g548
  (
    n561,
    n332,
    n314,
    n350,
    n329
  );


  and
  g549
  (
    n680,
    n495,
    n458,
    n344,
    n469
  );


  nand
  g550
  (
    n601,
    n327,
    n287,
    n341,
    n357
  );


  xor
  g551
  (
    n654,
    n498,
    n313,
    n286,
    n428
  );


  or
  g552
  (
    n509,
    n391,
    n366,
    n502,
    n465
  );


  xnor
  g553
  (
    n567,
    n500,
    n303,
    n308,
    n357
  );


  xor
  g554
  (
    n614,
    n312,
    n367,
    n345,
    n328
  );


  or
  g555
  (
    n517,
    n362,
    n423,
    n336,
    n408
  );


  nand
  g556
  (
    n545,
    n343,
    n306,
    n468,
    n302
  );


  xor
  g557
  (
    n607,
    n476,
    n488,
    n414,
    n368
  );


  nand
  g558
  (
    n661,
    n343,
    n412,
    n428,
    n491
  );


  or
  g559
  (
    n689,
    n371,
    n466,
    n424,
    n384
  );


  xor
  g560
  (
    n681,
    n287,
    n335,
    n502,
    n480
  );


  nand
  g561
  (
    n656,
    n320,
    n400,
    n473,
    n341
  );


  and
  g562
  (
    n647,
    n411,
    n424,
    n347,
    n381
  );


  nor
  g563
  (
    n522,
    n332,
    n499,
    n346,
    n406
  );


  xnor
  g564
  (
    n538,
    n425,
    n316,
    n417,
    n383
  );


  or
  g565
  (
    n650,
    n329,
    n315,
    n309,
    n349
  );


  xnor
  g566
  (
    n691,
    n370,
    n398,
    n286,
    n484
  );


  nand
  g567
  (
    n539,
    n394,
    n318,
    n310,
    n316
  );


  xor
  g568
  (
    n560,
    n383,
    n464,
    n426,
    n313
  );


  xnor
  g569
  (
    n587,
    n376,
    n486,
    n342,
    n400
  );


  nand
  g570
  (
    KeyWire_0_7,
    n463,
    n457,
    n346,
    n416
  );


  or
  g571
  (
    n535,
    n486,
    n485,
    n286,
    n409
  );


  nor
  g572
  (
    n597,
    n383,
    n371,
    n349,
    n470
  );


  and
  g573
  (
    n534,
    n396,
    n290,
    n350,
    n324
  );


  and
  g574
  (
    n557,
    n363,
    n354,
    n496,
    n339
  );


  or
  g575
  (
    n546,
    n376,
    n464,
    n501,
    n365
  );


  nor
  g576
  (
    n632,
    n426,
    n373,
    n397,
    n409
  );


  or
  g577
  (
    n688,
    n291,
    n303,
    n502,
    n368
  );


  xnor
  g578
  (
    n542,
    n356,
    n310,
    n467,
    n418
  );


  xnor
  g579
  (
    n506,
    n405,
    n310,
    n361,
    n418
  );


  xnor
  g580
  (
    n676,
    n388,
    n492,
    n326,
    n366
  );


  nand
  g581
  (
    n663,
    n309,
    n338,
    n315,
    n502
  );


  xor
  g582
  (
    n603,
    n305,
    n392,
    n290,
    n375
  );


  nand
  g583
  (
    n556,
    n484,
    n319,
    n465,
    n474
  );


  or
  g584
  (
    n591,
    n333,
    n384,
    n407,
    n427
  );


  xor
  g585
  (
    n629,
    n342,
    n319,
    n315,
    n393
  );


  nor
  g586
  (
    n628,
    n291,
    n304,
    n345,
    n379
  );


  nand
  g587
  (
    n530,
    n361,
    n332,
    n293,
    n330
  );


  xnor
  g588
  (
    n617,
    n325,
    n305,
    n386,
    n336
  );


  xnor
  g589
  (
    n642,
    n406,
    n388,
    n491,
    n371
  );


  xnor
  g590
  (
    n667,
    n301,
    n362,
    n498
  );


  or
  g591
  (
    n549,
    n327,
    n373,
    n286,
    n319
  );


  xor
  g592
  (
    n537,
    n423,
    n405,
    n347,
    n501
  );


  nor
  g593
  (
    n653,
    n289,
    n360,
    n475,
    n379
  );


  or
  g594
  (
    n520,
    n389,
    n484,
    n469,
    n409
  );


  xor
  g595
  (
    n621,
    n345,
    n299,
    n305,
    n300
  );


  xor
  g596
  (
    n673,
    n355,
    n323,
    n356,
    n324
  );


  nand
  g597
  (
    n652,
    n369,
    n385,
    n488,
    n289
  );


  nor
  g598
  (
    n569,
    n427,
    n408,
    n492,
    n484
  );


  nor
  g599
  (
    n598,
    n297,
    n482,
    n333,
    n407
  );


  nor
  g600
  (
    n570,
    n494,
    n300,
    n337,
    n353
  );


  and
  g601
  (
    n605,
    n304,
    n328,
    n422,
    n428
  );


  or
  g602
  (
    n665,
    n469,
    n415,
    n312,
    n338
  );


  xnor
  g603
  (
    n659,
    n348,
    n285,
    n464,
    n299
  );


  xor
  g604
  (
    n532,
    n412,
    n296,
    n297,
    n370
  );


  or
  g605
  (
    n516,
    n330,
    n421,
    n354,
    n407
  );


  nand
  g606
  (
    n655,
    n419,
    n351,
    n381,
    n466
  );


  xnor
  g607
  (
    n528,
    n331,
    n337,
    n328,
    n398
  );


  nand
  g608
  (
    n531,
    n459,
    n423,
    n372,
    n401
  );


  or
  g609
  (
    n649,
    n485,
    n386,
    n397,
    n395
  );


  or
  g610
  (
    n548,
    n387,
    n354,
    n296,
    n366
  );


  and
  g611
  (
    n670,
    n374,
    n372,
    n396,
    n339
  );


  and
  g612
  (
    n627,
    n470,
    n468,
    n403,
    n396
  );


  xnor
  g613
  (
    n533,
    n372,
    n340,
    n462,
    n395
  );


  and
  g614
  (
    n690,
    n386,
    n310,
    n288,
    n425
  );


  xnor
  g615
  (
    n606,
    n330,
    n299,
    n306,
    n394
  );


  xnor
  g616
  (
    n576,
    n422,
    n303,
    n320,
    n487
  );


  or
  g617
  (
    n541,
    n397,
    n351,
    n471,
    n475
  );


  or
  g618
  (
    n514,
    n494,
    n329,
    n340,
    n321
  );


  xor
  g619
  (
    n578,
    n421,
    n483,
    n467,
    n460
  );


  nor
  g620
  (
    n599,
    n488,
    n486,
    n335,
    n393
  );


  and
  g621
  (
    n643,
    n374,
    n416,
    n295,
    n376
  );


  xnor
  g622
  (
    n524,
    n463,
    n464,
    n478,
    n315
  );


  or
  g623
  (
    n585,
    n338,
    n340,
    n334,
    n359
  );


  and
  g624
  (
    n651,
    n357,
    n500,
    n369,
    n385
  );


  xor
  g625
  (
    n639,
    n295,
    n302,
    n347,
    n388
  );


  xnor
  g626
  (
    n518,
    n421,
    n403,
    n314,
    n339
  );


  nor
  g627
  (
    n551,
    n326,
    n326,
    n366,
    n469
  );


  xnor
  g628
  (
    n612,
    n292,
    n316,
    n337,
    n490
  );


  nor
  g629
  (
    n619,
    n298,
    n319,
    n306,
    n364
  );


  nor
  g630
  (
    n562,
    n457,
    n393,
    n462,
    n422
  );


  or
  g631
  (
    n625,
    n347,
    n294,
    n500,
    n499
  );


  and
  g632
  (
    n636,
    n353,
    n417,
    n497
  );


  xor
  g633
  (
    n589,
    n428,
    n489,
    n477,
    n474
  );


  or
  g634
  (
    n687,
    n355,
    n342,
    n308,
    n314
  );


  xnor
  g635
  (
    n596,
    n317,
    n420,
    n321,
    n367
  );


  xnor
  g636
  (
    n513,
    n395,
    n324,
    n480,
    n458
  );


  and
  g637
  (
    n573,
    n463,
    n404,
    n352,
    n481
  );


  xnor
  g638
  (
    n648,
    n392,
    n374,
    n308,
    n380
  );


  or
  g639
  (
    n521,
    n462,
    n483,
    n351
  );


  xnor
  g640
  (
    n529,
    n360,
    n490,
    n359,
    n307
  );


  xnor
  g641
  (
    n694,
    n471,
    n302,
    n395,
    n384
  );


  nand
  g642
  (
    n633,
    n307,
    n458,
    n322,
    n336
  );


  xor
  g643
  (
    n666,
    n494,
    n335,
    n419,
    n457
  );


  xor
  g644
  (
    n637,
    n290,
    n474,
    n311,
    n306
  );


  xnor
  g645
  (
    n564,
    n385,
    n456,
    n389,
    n382
  );


  xnor
  g646
  (
    n503,
    n329,
    n472,
    n293,
    n402
  );


  nor
  g647
  (
    n523,
    n356,
    n414,
    n321,
    n312
  );


  xor
  g648
  (
    n634,
    n375,
    n364,
    n487,
    n378
  );


  xnor
  g649
  (
    n640,
    n426,
    n338,
    n460,
    n406
  );


  xor
  g650
  (
    n602,
    n382,
    n342,
    n289,
    n376
  );


  nor
  g651
  (
    n507,
    n304,
    n323,
    n424,
    n470
  );


  xnor
  g652
  (
    n675,
    n384,
    n370,
    n501,
    n479
  );


  xor
  g653
  (
    n678,
    n309,
    n461,
    n472,
    n293
  );


  nor
  g654
  (
    n645,
    n394,
    n411,
    n385,
    n487
  );


  nor
  g655
  (
    n686,
    n382,
    n364,
    n479,
    n349
  );


  nand
  g656
  (
    n505,
    n418,
    n413,
    n307,
    n483
  );


  and
  g657
  (
    n623,
    n336,
    n458,
    n407,
    n346
  );


  nand
  g658
  (
    n550,
    n415,
    n365,
    n495,
    n403
  );


  nor
  g659
  (
    n635,
    n399,
    n301,
    n420,
    n368
  );


  or
  g660
  (
    n574,
    n477,
    n355,
    n391,
    n493
  );


  nand
  g661
  (
    n608,
    n421,
    n496,
    n351,
    n485
  );


  nand
  g662
  (
    n728,
    n512,
    n614,
    n657,
    n638
  );


  nor
  g663
  (
    n705,
    n610,
    n691,
    n612,
    n676
  );


  nand
  g664
  (
    KeyWire_0_31,
    n662,
    n627,
    n674,
    n636
  );


  or
  g665
  (
    n715,
    n558,
    n618,
    n642,
    n694
  );


  xor
  g666
  (
    n778,
    n663,
    n660,
    n555,
    n653
  );


  and
  g667
  (
    n725,
    n551,
    n623,
    n606,
    n602
  );


  or
  g668
  (
    n701,
    n571,
    n579,
    n572,
    n621
  );


  or
  g669
  (
    n739,
    n31,
    n623,
    n606,
    n634
  );


  nor
  g670
  (
    n802,
    n664,
    n643,
    n613,
    n593
  );


  and
  g671
  (
    n797,
    n611,
    n635,
    n631
  );


  nand
  g672
  (
    n714,
    n632,
    n608,
    n675,
    n536
  );


  or
  g673
  (
    n817,
    n688,
    n521,
    n596,
    n633
  );


  xnor
  g674
  (
    n818,
    n682,
    n595,
    n693,
    n577
  );


  and
  g675
  (
    n805,
    n553,
    n679,
    n580,
    n609
  );


  xor
  g676
  (
    n792,
    n618,
    n694,
    n556,
    n560
  );


  nand
  g677
  (
    n811,
    n682,
    n667,
    n623,
    n652
  );


  xnor
  g678
  (
    n770,
    n602,
    n615,
    n638,
    n620
  );


  xor
  g679
  (
    n730,
    n626,
    n653,
    n617,
    n557
  );


  nand
  g680
  (
    n777,
    n672,
    n685,
    n617,
    n607
  );


  or
  g681
  (
    n809,
    n656,
    n654,
    n663,
    n506
  );


  nand
  g682
  (
    n812,
    n672,
    n565,
    n575,
    n621
  );


  nand
  g683
  (
    n779,
    n569,
    n659,
    n636,
    n676
  );


  nand
  g684
  (
    n726,
    n640,
    n591,
    n564,
    n664
  );


  nand
  g685
  (
    n700,
    n635,
    n643,
    n515,
    n655
  );


  xor
  g686
  (
    n787,
    n674,
    n691,
    n661,
    n689
  );


  xor
  g687
  (
    n708,
    n686,
    n678,
    n665,
    n504
  );


  nand
  g688
  (
    n710,
    n683,
    n692,
    n668,
    n639
  );


  xnor
  g689
  (
    n761,
    n690,
    n672,
    n590,
    n600
  );


  xnor
  g690
  (
    n791,
    n652,
    n32,
    n639,
    n610
  );


  and
  g691
  (
    n719,
    n637,
    n597,
    n647,
    n687
  );


  and
  g692
  (
    n731,
    n691,
    n559,
    n617,
    n634
  );


  and
  g693
  (
    n727,
    n605,
    n666,
    n30,
    n608
  );


  nand
  g694
  (
    KeyWire_0_25,
    n657,
    n671,
    n648,
    n543
  );


  and
  g695
  (
    n768,
    n692,
    n29,
    n639,
    n647
  );


  xnor
  g696
  (
    n707,
    n651,
    n604,
    n635,
    n637
  );


  nor
  g697
  (
    n807,
    n673,
    n669,
    n662,
    n628
  );


  xor
  g698
  (
    n713,
    n520,
    n647,
    n642,
    n533
  );


  nand
  g699
  (
    n773,
    n681,
    n573,
    n667,
    n658
  );


  xor
  g700
  (
    n815,
    n614,
    n505,
    n644,
    n634
  );


  or
  g701
  (
    n711,
    n603,
    n532,
    n683,
    n609
  );


  xor
  g702
  (
    n737,
    n680,
    n678,
    n648,
    n503
  );


  xnor
  g703
  (
    n733,
    n644,
    n574,
    n661,
    n629
  );


  nor
  g704
  (
    n729,
    n693,
    n626,
    n609,
    n688
  );


  and
  g705
  (
    n767,
    n29,
    n664,
    n607,
    n592
  );


  or
  g706
  (
    n801,
    n644,
    n511,
    n578,
    n616
  );


  or
  g707
  (
    n800,
    n668,
    n28,
    n642,
    n689
  );


  and
  g708
  (
    n755,
    n656,
    n660,
    n688,
    n561
  );


  and
  g709
  (
    n764,
    n646,
    n629,
    n605,
    n688
  );


  xor
  g710
  (
    n716,
    n28,
    n634,
    n624,
    n632
  );


  and
  g711
  (
    n756,
    n685,
    n534,
    n633,
    n613
  );


  nor
  g712
  (
    n794,
    n687,
    n616,
    n610,
    n627
  );


  xor
  g713
  (
    n793,
    n677,
    n668,
    n641,
    n690
  );


  and
  g714
  (
    n738,
    n530,
    n568,
    n664,
    n594
  );


  or
  g715
  (
    n762,
    n608,
    n606,
    n675,
    n619
  );


  nand
  g716
  (
    n740,
    n613,
    n677,
    n612,
    n650
  );


  xor
  g717
  (
    n781,
    n645,
    n603,
    n563,
    n650
  );


  or
  g718
  (
    n724,
    n687,
    n673,
    n649,
    n508
  );


  nand
  g719
  (
    n741,
    n601,
    n619,
    n671,
    n638
  );


  xor
  g720
  (
    n720,
    n648,
    n620,
    n655,
    n676
  );


  nor
  g721
  (
    n732,
    n624,
    n660,
    n669,
    n685
  );


  and
  g722
  (
    n772,
    n645,
    n648,
    n669,
    n28
  );


  nor
  g723
  (
    n744,
    n611,
    n673,
    n661,
    n621
  );


  xor
  g724
  (
    n747,
    n637,
    n615,
    n674,
    n666
  );


  or
  g725
  (
    n814,
    n624,
    n631,
    n649,
    n671
  );


  or
  g726
  (
    n717,
    n614,
    n602,
    n656,
    n684
  );


  and
  g727
  (
    n782,
    n680,
    n612,
    n646,
    n542
  );


  nor
  g728
  (
    n748,
    n682,
    n636,
    n604,
    n680
  );


  xor
  g729
  (
    n749,
    n601,
    n625,
    n581,
    n665
  );


  and
  g730
  (
    n786,
    n537,
    n630,
    n624,
    n519
  );


  or
  g731
  (
    n796,
    n518,
    n586,
    n622,
    n651
  );


  and
  g732
  (
    n799,
    n585,
    n32,
    n611,
    n652
  );


  nor
  g733
  (
    KeyWire_0_15,
    n552,
    n670,
    n641
  );


  or
  g734
  (
    n784,
    n675,
    n625,
    n690,
    n598
  );


  xor
  g735
  (
    n766,
    n686,
    n628,
    n627,
    n625
  );


  and
  g736
  (
    n709,
    n655,
    n694,
    n522,
    n603
  );


  xnor
  g737
  (
    n723,
    n608,
    n570,
    n630,
    n29
  );


  or
  g738
  (
    n760,
    n673,
    n681,
    n545,
    n636
  );


  nor
  g739
  (
    n699,
    n677,
    n675,
    n562,
    n613
  );


  or
  g740
  (
    n798,
    n672,
    n629,
    n589,
    n540
  );


  nand
  g741
  (
    n816,
    n646,
    n630,
    n523,
    n550
  );


  xnor
  g742
  (
    KeyWire_0_13,
    n627,
    n686,
    n601,
    n626
  );


  and
  g743
  (
    n774,
    n670,
    n604,
    n601,
    n610
  );


  xor
  g744
  (
    n785,
    n692,
    n646,
    n602,
    n544
  );


  nand
  g745
  (
    n759,
    n607,
    n693,
    n609,
    n679
  );


  xor
  g746
  (
    n718,
    n31,
    n662,
    n684,
    n658
  );


  xor
  g747
  (
    n788,
    n618,
    n32,
    n649,
    n667
  );


  nor
  g748
  (
    n742,
    n654,
    n510,
    n631,
    n682
  );


  and
  g749
  (
    n771,
    n605,
    n628,
    n660,
    n641
  );


  nor
  g750
  (
    n697,
    n587,
    n685,
    n639,
    n662
  );


  xor
  g751
  (
    n753,
    n679,
    n583,
    n683,
    n661
  );


  xor
  g752
  (
    n752,
    n677,
    n620,
    n640
  );


  and
  g753
  (
    n763,
    n621,
    n567,
    n643,
    n584
  );


  or
  g754
  (
    n746,
    n606,
    n546,
    n666,
    n626
  );


  xor
  g755
  (
    n735,
    n616,
    n548,
    n547,
    n30
  );


  xnor
  g756
  (
    n790,
    n666,
    n31,
    n651,
    n690
  );


  or
  g757
  (
    n751,
    n676,
    n681,
    n684,
    n659
  );


  xor
  g758
  (
    n776,
    n655,
    n645,
    n668,
    n650
  );


  xnor
  g759
  (
    n808,
    n527,
    n663,
    n652,
    n607
  );


  nor
  g760
  (
    n712,
    n641,
    n680,
    n30,
    n611
  );


  nor
  g761
  (
    n696,
    n28,
    n615,
    n539,
    n622
  );


  xor
  g762
  (
    n757,
    n509,
    n657,
    n689,
    n653
  );


  or
  g763
  (
    n804,
    n679,
    n647,
    n517,
    n526
  );


  xor
  g764
  (
    n704,
    n681,
    n538,
    n665,
    n630
  );


  xnor
  g765
  (
    n803,
    n693,
    n642,
    n513,
    n654
  );


  nor
  g766
  (
    n810,
    n32,
    n616,
    n549,
    n566
  );


  nor
  g767
  (
    n795,
    n529,
    n659,
    n656,
    n669
  );


  xnor
  g768
  (
    n780,
    n582,
    n599,
    n514,
    n633
  );


  or
  g769
  (
    n695,
    n653,
    n657,
    n665,
    n678
  );


  nand
  g770
  (
    n806,
    n640,
    n633,
    n629,
    n654
  );


  or
  g771
  (
    n754,
    n524,
    n614,
    n588,
    n638
  );


  xnor
  g772
  (
    n769,
    n667,
    n605,
    n670,
    n689
  );


  xor
  g773
  (
    n698,
    n671,
    n617,
    n643,
    n619
  );


  and
  g774
  (
    n789,
    n692,
    n29,
    n658,
    n507
  );


  and
  g775
  (
    n703,
    n632,
    n623,
    n659,
    n612
  );


  nor
  g776
  (
    n758,
    n625,
    n429,
    n525,
    n603
  );


  and
  g777
  (
    n745,
    n658,
    n650,
    n619,
    n644
  );


  nand
  g778
  (
    n765,
    n640,
    n535,
    n674,
    n576
  );


  and
  g779
  (
    n721,
    n528,
    n615,
    n678,
    n686
  );


  and
  g780
  (
    n722,
    n628,
    n649,
    n531,
    n635
  );


  nor
  g781
  (
    n702,
    n30,
    n691,
    n618,
    n622
  );


  nand
  g782
  (
    n750,
    n683,
    n516,
    n27,
    n687
  );


  nand
  g783
  (
    n734,
    n541,
    n622,
    n651,
    n554
  );


  nor
  g784
  (
    n783,
    n604,
    n645,
    n663,
    n694
  );


  nand
  g785
  (
    n775,
    n637,
    n31,
    n632,
    n684
  );


  xor
  g786
  (
    n902,
    n777,
    n81,
    n716,
    n69
  );


  xnor
  g787
  (
    n828,
    n750,
    n105,
    n80,
    n109
  );


  nand
  g788
  (
    n883,
    n784,
    n804,
    n731,
    n115
  );


  nand
  g789
  (
    n829,
    n725,
    n113,
    n806,
    n705
  );


  nor
  g790
  (
    n872,
    n126,
    n81,
    n89,
    n697
  );


  xnor
  g791
  (
    n911,
    n92,
    n114,
    n94,
    n765
  );


  or
  g792
  (
    n869,
    n740,
    n79,
    n69,
    n767
  );


  xor
  g793
  (
    n918,
    n135,
    n108,
    n717,
    n115
  );


  or
  g794
  (
    n843,
    n758,
    n100,
    n748,
    n759
  );


  xor
  g795
  (
    n859,
    n779,
    n109,
    n102,
    n68
  );


  nand
  g796
  (
    n916,
    n105,
    n103,
    n80,
    n85
  );


  nand
  g797
  (
    n897,
    n723,
    n128,
    n124,
    n79
  );


  xor
  g798
  (
    n870,
    n714,
    n132,
    n121,
    n71
  );


  nor
  g799
  (
    n823,
    n743,
    n83,
    n118,
    n700
  );


  xnor
  g800
  (
    n827,
    n106,
    n116,
    n118,
    n99
  );


  xnor
  g801
  (
    n865,
    n123,
    n770,
    n73,
    n703
  );


  xnor
  g802
  (
    n906,
    n741,
    n102,
    n131,
    n808
  );


  and
  g803
  (
    n839,
    n702,
    n789,
    n128,
    n82
  );


  nor
  g804
  (
    n904,
    n122,
    n122,
    n734,
    n788
  );


  and
  g805
  (
    n896,
    n68,
    n801,
    n135,
    n774
  );


  or
  g806
  (
    n882,
    n813,
    n131,
    n756,
    n124
  );


  nand
  g807
  (
    n867,
    n139,
    n133,
    n707,
    n109
  );


  xor
  g808
  (
    n912,
    n95,
    n78,
    n107,
    n104
  );


  xnor
  g809
  (
    n881,
    n722,
    n772,
    n97,
    n735
  );


  or
  g810
  (
    n830,
    n783,
    n72,
    n786,
    n101
  );


  nand
  g811
  (
    n855,
    n120,
    n89,
    n128,
    n112
  );


  nor
  g812
  (
    KeyWire_0_11,
    n768,
    n781,
    n129,
    n101
  );


  or
  g813
  (
    n876,
    n136,
    n84,
    n79,
    n119
  );


  nor
  g814
  (
    n871,
    n70,
    n807,
    n72,
    n105
  );


  nor
  g815
  (
    n880,
    n724,
    n102,
    n110,
    n696
  );


  nor
  g816
  (
    n893,
    n125,
    n96,
    n129,
    n117
  );


  or
  g817
  (
    n884,
    n792,
    n137,
    n747,
    n811
  );


  nand
  g818
  (
    n837,
    n136,
    n111,
    n721,
    n712
  );


  nand
  g819
  (
    n845,
    n86,
    n809,
    n125,
    n69
  );


  nand
  g820
  (
    n894,
    n125,
    n69,
    n120,
    n803
  );


  xor
  g821
  (
    n889,
    n85,
    n114,
    n89,
    n119
  );


  xor
  g822
  (
    n866,
    n128,
    n130,
    n124,
    n790
  );


  nand
  g823
  (
    n888,
    n709,
    n800,
    n132,
    n104
  );


  or
  g824
  (
    n910,
    n812,
    n732,
    n86
  );


  nor
  g825
  (
    n908,
    n88,
    n116,
    n76,
    n75
  );


  nor
  g826
  (
    n868,
    n726,
    n98,
    n95,
    n138
  );


  nor
  g827
  (
    n831,
    n751,
    n715,
    n117,
    n74
  );


  and
  g828
  (
    n840,
    n126,
    n138,
    n120,
    n785
  );


  nor
  g829
  (
    n848,
    n97,
    n127,
    n113,
    n742
  );


  xor
  g830
  (
    n820,
    n134,
    n761,
    n112,
    n91
  );


  nand
  g831
  (
    n885,
    n730,
    n134,
    n91,
    n90
  );


  nand
  g832
  (
    n909,
    n76,
    n103,
    n794,
    n136
  );


  nor
  g833
  (
    n878,
    n75,
    n766,
    n95,
    n97
  );


  and
  g834
  (
    n853,
    n814,
    n708,
    n798,
    n136
  );


  or
  g835
  (
    n917,
    n96,
    n106,
    n746,
    n110
  );


  nand
  g836
  (
    n900,
    n87,
    n87,
    n94,
    n771
  );


  nor
  g837
  (
    n834,
    n93,
    n103,
    n754,
    n76
  );


  xor
  g838
  (
    n851,
    n94,
    n87,
    n139,
    n755
  );


  or
  g839
  (
    n861,
    n737,
    n84,
    n701,
    n93
  );


  xnor
  g840
  (
    n847,
    n129,
    n695,
    n85,
    n83
  );


  nand
  g841
  (
    n886,
    n817,
    n101,
    n105,
    n102
  );


  xnor
  g842
  (
    n905,
    n79,
    n97,
    n84
  );


  and
  g843
  (
    n913,
    n99,
    n77,
    n71,
    n115
  );


  and
  g844
  (
    KeyWire_0_5,
    n77,
    n71,
    n118,
    n88
  );


  nand
  g845
  (
    n826,
    n773,
    n74,
    n88,
    n96
  );


  or
  g846
  (
    n860,
    n73,
    n124,
    n80,
    n89
  );


  and
  g847
  (
    n857,
    n719,
    n791,
    n70,
    n137
  );


  xor
  g848
  (
    n850,
    n711,
    n91,
    n133,
    n123
  );


  nand
  g849
  (
    n852,
    n121,
    n122,
    n780,
    n816
  );


  nor
  g850
  (
    n844,
    n129,
    n126,
    n132,
    n108
  );


  or
  g851
  (
    n841,
    n769,
    n775,
    n116,
    n117
  );


  nand
  g852
  (
    n903,
    n99,
    n753,
    n104,
    n778
  );


  or
  g853
  (
    n898,
    n752,
    n793,
    n744,
    n83
  );


  xnor
  g854
  (
    n879,
    n119,
    n83,
    n762,
    n135
  );


  nor
  g855
  (
    n892,
    n117,
    n132,
    n68,
    n115
  );


  nor
  g856
  (
    n919,
    n127,
    n81,
    n114,
    n78
  );


  or
  g857
  (
    KeyWire_0_6,
    n82,
    n100,
    n121,
    n81
  );


  nor
  g858
  (
    n875,
    n127,
    n134,
    n98,
    n130
  );


  nand
  g859
  (
    n846,
    n787,
    n109,
    n764,
    n72
  );


  xor
  g860
  (
    n891,
    n77,
    n137,
    n82,
    n706
  );


  xnor
  g861
  (
    n832,
    n130,
    n93,
    n776,
    n106
  );


  or
  g862
  (
    n849,
    n73,
    n727,
    n113,
    n125
  );


  xor
  g863
  (
    n907,
    n123,
    n805,
    n110,
    n108
  );


  xor
  g864
  (
    n914,
    n107,
    n127,
    n122,
    n718
  );


  and
  g865
  (
    n825,
    n733,
    n101,
    n116,
    n138
  );


  xor
  g866
  (
    n821,
    n796,
    n82,
    n728,
    n118
  );


  or
  g867
  (
    n874,
    n92,
    n134,
    n818,
    n713
  );


  xnor
  g868
  (
    n890,
    n99,
    n107,
    n78,
    n749
  );


  nor
  g869
  (
    n864,
    n815,
    n98,
    n92,
    n131
  );


  nor
  g870
  (
    n833,
    n710,
    n108,
    n760,
    n111
  );


  nor
  g871
  (
    n887,
    n704,
    n123,
    n74,
    n729
  );


  xor
  g872
  (
    n819,
    n795,
    n106,
    n71,
    n90
  );


  and
  g873
  (
    n901,
    n699,
    n133,
    n736,
    n757
  );


  and
  g874
  (
    n920,
    n745,
    n72,
    n68,
    n75
  );


  nand
  g875
  (
    n838,
    n112,
    n113,
    n74,
    n138
  );


  or
  g876
  (
    n863,
    n139,
    n111,
    n739,
    n76
  );


  xor
  g877
  (
    n877,
    n100,
    n133,
    n98,
    n110
  );


  xor
  g878
  (
    n895,
    n810,
    n93,
    n120,
    n698
  );


  and
  g879
  (
    n921,
    n90,
    n91,
    n799,
    n70
  );


  nor
  g880
  (
    n899,
    n90,
    n130,
    n763,
    n135
  );


  or
  g881
  (
    n842,
    n107,
    n85,
    n137,
    n797
  );


  nor
  g882
  (
    n822,
    n126,
    n87,
    n738,
    n114
  );


  xnor
  g883
  (
    n856,
    n75,
    n78,
    n86,
    n104
  );


  xnor
  g884
  (
    n858,
    n139,
    n100,
    n88,
    n95
  );


  nand
  g885
  (
    n862,
    n96,
    n782,
    n94,
    n111
  );


  xor
  g886
  (
    n824,
    n720,
    n80,
    n112,
    n70
  );


  nand
  g887
  (
    n836,
    n92,
    n802,
    n77,
    n131
  );


  or
  g888
  (
    n873,
    n121,
    n103,
    n119,
    n73
  );


  nand
  g889
  (
    n998,
    n822,
    n259,
    n235
  );


  nand
  g890
  (
    n979,
    n254,
    n276,
    n260,
    n228
  );


  or
  g891
  (
    n960,
    n920,
    n843,
    n261,
    n253
  );


  nand
  g892
  (
    n983,
    n896,
    n864,
    n244,
    n867
  );


  or
  g893
  (
    n966,
    n259,
    n269,
    n911,
    n267
  );


  xor
  g894
  (
    n930,
    n892,
    n839,
    n915,
    n255
  );


  xor
  g895
  (
    n992,
    n912,
    n236,
    n275,
    n903
  );


  and
  g896
  (
    n963,
    n264,
    n820,
    n269,
    n429
  );


  or
  g897
  (
    n956,
    n253,
    n238,
    n233,
    n272
  );


  and
  g898
  (
    n944,
    n876,
    n232,
    n273,
    n249
  );


  or
  g899
  (
    n928,
    n857,
    n852,
    n226,
    n244
  );


  or
  g900
  (
    n999,
    n230,
    n828,
    n250,
    n236
  );


  xor
  g901
  (
    n939,
    n239,
    n256,
    n893,
    n910
  );


  or
  g902
  (
    n994,
    n242,
    n257,
    n243,
    n238
  );


  xor
  g903
  (
    n923,
    n231,
    n228,
    n919,
    n901
  );


  nor
  g904
  (
    n962,
    n274,
    n831,
    n846,
    n271
  );


  and
  g905
  (
    n926,
    n266,
    n838,
    n227,
    n909
  );


  nand
  g906
  (
    KeyWire_0_24,
    n841,
    n250,
    n837,
    n851
  );


  xor
  g907
  (
    n985,
    n235,
    n885,
    n269,
    n905
  );


  or
  g908
  (
    n959,
    n250,
    n253,
    n241,
    n261
  );


  xor
  g909
  (
    n925,
    n890,
    n237,
    n826,
    n888
  );


  or
  g910
  (
    n969,
    n886,
    n277,
    n228,
    n819
  );


  or
  g911
  (
    n929,
    n274,
    n255,
    n883,
    n258
  );


  nor
  g912
  (
    n977,
    n258,
    n887,
    n921,
    n874
  );


  xor
  g913
  (
    n947,
    n258,
    n821,
    n272,
    n917
  );


  nand
  g914
  (
    n927,
    n832,
    n245,
    n275,
    n246
  );


  nand
  g915
  (
    n965,
    n273,
    n261,
    n235,
    n861
  );


  or
  g916
  (
    n955,
    n241,
    n239,
    n242,
    n273
  );


  xor
  g917
  (
    n984,
    n244,
    n850,
    n262,
    n245
  );


  xor
  g918
  (
    n972,
    n904,
    n900,
    n877,
    n239
  );


  xnor
  g919
  (
    n996,
    n246,
    n227,
    n829,
    n252
  );


  xor
  g920
  (
    KeyWire_0_29,
    n231,
    n842,
    n863,
    n226
  );


  xor
  g921
  (
    n986,
    n248,
    n233,
    n251,
    n847
  );


  xnor
  g922
  (
    n934,
    n227,
    n246,
    n263,
    n260
  );


  xnor
  g923
  (
    n993,
    n229,
    n231,
    n273,
    n267
  );


  xnor
  g924
  (
    n938,
    n261,
    n274,
    n880,
    n236
  );


  nor
  g925
  (
    n951,
    n881,
    n872,
    n253,
    n247
  );


  xor
  g926
  (
    n981,
    n247,
    n241,
    n268,
    n259
  );


  nand
  g927
  (
    n932,
    n266,
    n875,
    n259,
    n267
  );


  and
  g928
  (
    n961,
    n256,
    n836,
    n265,
    n245
  );


  and
  g929
  (
    n967,
    n244,
    n265,
    n270,
    n240
  );


  nor
  g930
  (
    n982,
    n825,
    n835,
    n234,
    n250
  );


  or
  g931
  (
    n940,
    n871,
    n263,
    n234,
    n232
  );


  and
  g932
  (
    n946,
    n429,
    n243,
    n849,
    n233
  );


  xor
  g933
  (
    n936,
    n271,
    n242,
    n237,
    n246
  );


  and
  g934
  (
    n975,
    n845,
    n902,
    n248,
    n265
  );


  nand
  g935
  (
    n987,
    n254,
    n899,
    n233,
    n827
  );


  or
  g936
  (
    n941,
    n248,
    n891,
    n275,
    n226
  );


  xor
  g937
  (
    n953,
    n270,
    n248,
    n858,
    n275
  );


  nor
  g938
  (
    n997,
    n430,
    n855,
    n247,
    n249
  );


  or
  g939
  (
    n931,
    n264,
    n271,
    n895,
    n234
  );


  nand
  g940
  (
    n933,
    n274,
    n237,
    n257,
    n914
  );


  and
  g941
  (
    n990,
    n824,
    n251,
    n277
  );


  or
  g942
  (
    n935,
    n906,
    n860,
    n898,
    n865
  );


  xnor
  g943
  (
    n978,
    n245,
    n249,
    n232,
    n236
  );


  xor
  g944
  (
    n970,
    n243,
    n884,
    n897,
    n241
  );


  and
  g945
  (
    n924,
    n830,
    n269,
    n229,
    n227
  );


  xor
  g946
  (
    n971,
    n266,
    n276,
    n854,
    n240
  );


  and
  g947
  (
    n988,
    n866,
    n270,
    n862,
    n238
  );


  xnor
  g948
  (
    n991,
    n263,
    n268,
    n251,
    n243
  );


  and
  g949
  (
    n968,
    n429,
    n276,
    n430,
    n264
  );


  and
  g950
  (
    n954,
    n254,
    n265,
    n262,
    n232
  );


  or
  g951
  (
    n958,
    n252,
    n268,
    n238
  );


  and
  g952
  (
    n980,
    n240,
    n272,
    n260,
    n266
  );


  nor
  g953
  (
    n937,
    n247,
    n262,
    n255,
    n856
  );


  nand
  g954
  (
    n973,
    n894,
    n844,
    n853,
    n913
  );


  xnor
  g955
  (
    n945,
    n263,
    n258,
    n229,
    n276
  );


  or
  g956
  (
    n942,
    n270,
    n916,
    n254,
    n257
  );


  nand
  g957
  (
    n1000,
    n272,
    n859,
    n230,
    n239
  );


  nor
  g958
  (
    n952,
    n234,
    n242,
    n834,
    n228
  );


  xor
  g959
  (
    n949,
    n252,
    n264,
    n879,
    n907
  );


  and
  g960
  (
    n976,
    n868,
    n256,
    n833,
    n873
  );


  and
  g961
  (
    n989,
    n229,
    n840,
    n823,
    n231
  );


  nor
  g962
  (
    n995,
    n257,
    n255,
    n878,
    n869
  );


  or
  g963
  (
    n948,
    n848,
    n889,
    n237,
    n256
  );


  nand
  g964
  (
    n950,
    n230,
    n271,
    n260,
    n918
  );


  and
  g965
  (
    n974,
    n430,
    n277,
    n882
  );


  and
  g966
  (
    n964,
    n262,
    n908,
    n240,
    n267
  );


  xor
  g967
  (
    KeyWire_0_23,
    n870,
    n252,
    n249,
    n230
  );


  and
  g968
  (
    n1007,
    n437,
    n945,
    n962,
    n998
  );


  and
  g969
  (
    n1004,
    n924,
    n987,
    n981,
    n963
  );


  and
  g970
  (
    n1029,
    n977,
    n922,
    n997,
    n432
  );


  nand
  g971
  (
    n1020,
    n995,
    n437,
    n970,
    n950
  );


  xor
  g972
  (
    n1013,
    n432,
    n439,
    n433,
    n961
  );


  and
  g973
  (
    n1021,
    n440,
    n937,
    n433,
    n960
  );


  xnor
  g974
  (
    n1015,
    n931,
    n438,
    n434,
    n440
  );


  nand
  g975
  (
    n1023,
    n431,
    n927,
    n442,
    n438
  );


  and
  g976
  (
    n1024,
    n967,
    n442,
    n434,
    n431
  );


  xnor
  g977
  (
    n1002,
    n442,
    n435,
    n975,
    n988
  );


  nand
  g978
  (
    n1011,
    n955,
    n438,
    n935,
    n938
  );


  nor
  g979
  (
    n1019,
    n991,
    n437,
    n956,
    n936
  );


  xnor
  g980
  (
    n1003,
    n972,
    n954,
    n437,
    n434
  );


  nand
  g981
  (
    n1028,
    n957,
    n979,
    n951,
    n982
  );


  nor
  g982
  (
    n1025,
    n992,
    n973,
    n984,
    n959
  );


  and
  g983
  (
    n1030,
    n433,
    n933,
    n983,
    n940
  );


  or
  g984
  (
    n1001,
    n989,
    n441,
    n928,
    n929
  );


  or
  g985
  (
    n1026,
    n435,
    n440,
    n930,
    n925
  );


  or
  g986
  (
    n1017,
    n932,
    n436,
    n434,
    n440
  );


  or
  g987
  (
    n1016,
    n432,
    n948,
    n941,
    n442
  );


  and
  g988
  (
    n1012,
    n949,
    n436,
    n432,
    n976
  );


  nand
  g989
  (
    n1022,
    n964,
    n943,
    n435,
    n436
  );


  nor
  g990
  (
    n1032,
    n999,
    n953,
    n439,
    n947
  );


  nand
  g991
  (
    n1005,
    n980,
    n433,
    n435,
    n996
  );


  nand
  g992
  (
    n1010,
    n993,
    n994,
    n438,
    n978
  );


  nand
  g993
  (
    n1014,
    n939,
    n971,
    n969,
    n431
  );


  xnor
  g994
  (
    n1006,
    n944,
    n942,
    n966,
    n974
  );


  nand
  g995
  (
    n1018,
    n439,
    n441,
    n990,
    n430
  );


  or
  g996
  (
    n1008,
    n923,
    n965,
    n985,
    n1000
  );


  xor
  g997
  (
    n1031,
    n946,
    n441,
    n958,
    n431
  );


  xor
  g998
  (
    n1027,
    n968,
    n952,
    n986,
    n439
  );


  xor
  g999
  (
    n1009,
    n926,
    n436,
    n934,
    n441
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n395,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n471,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n356,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n61,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n291,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n854,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n915,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n543,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n68,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n65,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n106,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n835,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n262,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n813,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n394,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n743,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n419,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n67,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n519,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n333,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n664,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n477,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n442,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n957,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n943,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n706,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n497,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n152,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n343,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n922,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n595,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n736,
    KeyNOTWire_0_31
  );


endmodule

