

module Stat_736_2431
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n718,
  n721,
  n699,
  n697,
  n694,
  n695,
  n715,
  n717,
  n705,
  n719,
  n727,
  n711,
  n706,
  n712,
  n716,
  n713,
  n726,
  n707,
  n698,
  n696,
  n730,
  n753,
  n754,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n718;
  output n721;
  output n699;
  output n697;
  output n694;
  output n695;
  output n715;
  output n717;
  output n705;
  output n719;
  output n727;
  output n711;
  output n706;
  output n712;
  output n716;
  output n713;
  output n726;
  output n707;
  output n698;
  output n696;
  output n730;
  output n753;
  output n754;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n708;
  wire n709;
  wire n710;
  wire n714;
  wire n720;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n728;
  wire n729;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;

  not
  g0
  (
    n20,
    n2
  );


  buf
  g1
  (
    n26,
    n1
  );


  buf
  g2
  (
    n22,
    n2
  );


  buf
  g3
  (
    n21,
    n1
  );


  buf
  g4
  (
    n25,
    n3
  );


  not
  g5
  (
    n27,
    n1
  );


  not
  g6
  (
    n24,
    n2
  );


  not
  g7
  (
    n19,
    n2
  );


  buf
  g8
  (
    n23,
    n1
  );


  not
  g9
  (
    n46,
    n20
  );


  buf
  g10
  (
    n51,
    n27
  );


  not
  g11
  (
    n53,
    n25
  );


  not
  g12
  (
    n39,
    n27
  );


  buf
  g13
  (
    n42,
    n23
  );


  buf
  g14
  (
    n61,
    n24
  );


  buf
  g15
  (
    n31,
    n25
  );


  not
  g16
  (
    n59,
    n25
  );


  not
  g17
  (
    n36,
    n19
  );


  not
  g18
  (
    n30,
    n19
  );


  buf
  g19
  (
    n56,
    n23
  );


  buf
  g20
  (
    n55,
    n19
  );


  not
  g21
  (
    n52,
    n22
  );


  not
  g22
  (
    n49,
    n20
  );


  not
  g23
  (
    n41,
    n19
  );


  not
  g24
  (
    n47,
    n24
  );


  not
  g25
  (
    n62,
    n21
  );


  buf
  g26
  (
    n38,
    n23
  );


  buf
  g27
  (
    n32,
    n26
  );


  buf
  g28
  (
    n60,
    n27
  );


  not
  g29
  (
    n37,
    n26
  );


  not
  g30
  (
    n43,
    n22
  );


  not
  g31
  (
    n40,
    n27
  );


  not
  g32
  (
    n28,
    n20
  );


  not
  g33
  (
    n35,
    n26
  );


  buf
  g34
  (
    n33,
    n24
  );


  not
  g35
  (
    n50,
    n22
  );


  buf
  g36
  (
    n29,
    n24
  );


  not
  g37
  (
    n48,
    n26
  );


  not
  g38
  (
    n44,
    n21
  );


  not
  g39
  (
    n58,
    n20
  );


  not
  g40
  (
    n54,
    n21
  );


  not
  g41
  (
    n63,
    n25
  );


  buf
  g42
  (
    n45,
    n22
  );


  not
  g43
  (
    n34,
    n23
  );


  buf
  g44
  (
    n57,
    n21
  );


  buf
  g45
  (
    n170,
    n52
  );


  not
  g46
  (
    n80,
    n61
  );


  buf
  g47
  (
    n100,
    n15
  );


  buf
  g48
  (
    n109,
    n18
  );


  buf
  g49
  (
    n162,
    n54
  );


  not
  g50
  (
    n197,
    n7
  );


  not
  g51
  (
    n91,
    n46
  );


  buf
  g52
  (
    n112,
    n5
  );


  buf
  g53
  (
    n117,
    n37
  );


  buf
  g54
  (
    n186,
    n5
  );


  buf
  g55
  (
    n166,
    n35
  );


  not
  g56
  (
    n147,
    n58
  );


  not
  g57
  (
    n159,
    n31
  );


  buf
  g58
  (
    n187,
    n33
  );


  not
  g59
  (
    n87,
    n9
  );


  buf
  g60
  (
    n198,
    n41
  );


  buf
  g61
  (
    n121,
    n45
  );


  not
  g62
  (
    n131,
    n17
  );


  not
  g63
  (
    n125,
    n60
  );


  not
  g64
  (
    n71,
    n38
  );


  not
  g65
  (
    n70,
    n35
  );


  not
  g66
  (
    n74,
    n10
  );


  buf
  g67
  (
    n156,
    n39
  );


  buf
  g68
  (
    n86,
    n35
  );


  not
  g69
  (
    n191,
    n45
  );


  buf
  g70
  (
    n184,
    n43
  );


  not
  g71
  (
    n92,
    n55
  );


  buf
  g72
  (
    n76,
    n30
  );


  buf
  g73
  (
    n154,
    n38
  );


  buf
  g74
  (
    n102,
    n3
  );


  buf
  g75
  (
    n153,
    n29
  );


  not
  g76
  (
    n78,
    n56
  );


  not
  g77
  (
    n124,
    n10
  );


  buf
  g78
  (
    n106,
    n61
  );


  buf
  g79
  (
    n133,
    n60
  );


  buf
  g80
  (
    n122,
    n37
  );


  buf
  g81
  (
    n146,
    n37
  );


  not
  g82
  (
    n150,
    n28
  );


  not
  g83
  (
    n96,
    n60
  );


  buf
  g84
  (
    n176,
    n42
  );


  buf
  g85
  (
    n110,
    n46
  );


  not
  g86
  (
    n199,
    n35
  );


  not
  g87
  (
    n88,
    n31
  );


  buf
  g88
  (
    n160,
    n50
  );


  not
  g89
  (
    n175,
    n34
  );


  not
  g90
  (
    n168,
    n15
  );


  not
  g91
  (
    n101,
    n56
  );


  buf
  g92
  (
    n161,
    n9
  );


  buf
  g93
  (
    n193,
    n54
  );


  not
  g94
  (
    n132,
    n4
  );


  buf
  g95
  (
    n142,
    n55
  );


  buf
  g96
  (
    n192,
    n12
  );


  buf
  g97
  (
    n67,
    n52
  );


  buf
  g98
  (
    n126,
    n11
  );


  not
  g99
  (
    n195,
    n52
  );


  not
  g100
  (
    n152,
    n32
  );


  buf
  g101
  (
    n183,
    n16
  );


  not
  g102
  (
    KeyWire_0_7,
    n59
  );


  not
  g103
  (
    n113,
    n9
  );


  buf
  g104
  (
    n158,
    n34
  );


  not
  g105
  (
    n83,
    n37
  );


  not
  g106
  (
    n115,
    n16
  );


  buf
  g107
  (
    n185,
    n40
  );


  not
  g108
  (
    n68,
    n14
  );


  buf
  g109
  (
    n155,
    n48
  );


  not
  g110
  (
    n81,
    n61
  );


  not
  g111
  (
    n65,
    n62
  );


  not
  g112
  (
    n196,
    n49
  );


  not
  g113
  (
    n194,
    n57
  );


  buf
  g114
  (
    n104,
    n31
  );


  not
  g115
  (
    n202,
    n47
  );


  buf
  g116
  (
    n179,
    n33
  );


  not
  g117
  (
    n128,
    n51
  );


  not
  g118
  (
    n94,
    n13
  );


  not
  g119
  (
    n75,
    n32
  );


  not
  g120
  (
    n182,
    n8
  );


  not
  g121
  (
    n157,
    n50
  );


  buf
  g122
  (
    n139,
    n7
  );


  buf
  g123
  (
    n173,
    n52
  );


  buf
  g124
  (
    n144,
    n49
  );


  buf
  g125
  (
    n123,
    n6
  );


  buf
  g126
  (
    n120,
    n48
  );


  not
  g127
  (
    n167,
    n56
  );


  not
  g128
  (
    n95,
    n28
  );


  not
  g129
  (
    n69,
    n11
  );


  not
  g130
  (
    n93,
    n14
  );


  not
  g131
  (
    n140,
    n58
  );


  buf
  g132
  (
    n138,
    n12
  );


  not
  g133
  (
    n73,
    n5
  );


  buf
  g134
  (
    n99,
    n28
  );


  not
  g135
  (
    n79,
    n17
  );


  buf
  g136
  (
    n178,
    n49
  );


  not
  g137
  (
    n163,
    n12
  );


  not
  g138
  (
    n97,
    n50
  );


  not
  g139
  (
    n107,
    n51
  );


  buf
  g140
  (
    n84,
    n41
  );


  not
  g141
  (
    n137,
    n44
  );


  not
  g142
  (
    n72,
    n38
  );


  buf
  g143
  (
    n148,
    n36
  );


  buf
  g144
  (
    n108,
    n36
  );


  buf
  g145
  (
    n64,
    n60
  );


  buf
  g146
  (
    n119,
    n18
  );


  not
  g147
  (
    n177,
    n46
  );


  buf
  g148
  (
    KeyWire_0_1,
    n53
  );


  buf
  g149
  (
    n85,
    n12
  );


  not
  g150
  (
    n136,
    n31
  );


  not
  g151
  (
    n66,
    n32
  );


  not
  g152
  (
    n89,
    n54
  );


  buf
  g153
  (
    n171,
    n14
  );


  buf
  g154
  (
    n103,
    n55
  );


  not
  g155
  (
    n151,
    n62
  );


  not
  g156
  (
    n143,
    n36
  );


  not
  g157
  (
    n201,
    n50
  );


  buf
  g158
  (
    n130,
    n51
  );


  buf
  g159
  (
    n127,
    n18
  );


  not
  g160
  (
    n134,
    n47
  );


  buf
  g161
  (
    n188,
    n54
  );


  xnor
  g162
  (
    n169,
    n7,
    n63,
    n58
  );


  or
  g163
  (
    n174,
    n46,
    n47,
    n48,
    n3
  );


  and
  g164
  (
    n172,
    n56,
    n6,
    n57,
    n40
  );


  xnor
  g165
  (
    n90,
    n30,
    n34,
    n42,
    n15
  );


  nor
  g166
  (
    n129,
    n10,
    n42,
    n6,
    n39
  );


  nand
  g167
  (
    n111,
    n11,
    n43,
    n14,
    n9
  );


  nor
  g168
  (
    n181,
    n57,
    n45,
    n7,
    n11
  );


  xor
  g169
  (
    n190,
    n40,
    n62,
    n4,
    n39
  );


  xor
  g170
  (
    n149,
    n49,
    n28,
    n57,
    n8
  );


  nor
  g171
  (
    n135,
    n4,
    n48,
    n29,
    n47
  );


  or
  g172
  (
    n118,
    n59,
    n33,
    n8,
    n44
  );


  nand
  g173
  (
    n180,
    n29,
    n59,
    n5,
    n30
  );


  xnor
  g174
  (
    n189,
    n18,
    n41,
    n4,
    n15
  );


  nand
  g175
  (
    n114,
    n43,
    n58,
    n45,
    n40
  );


  or
  g176
  (
    n82,
    n33,
    n13,
    n29,
    n39
  );


  xnor
  g177
  (
    n116,
    n62,
    n42,
    n53,
    n43
  );


  nand
  g178
  (
    n141,
    n30,
    n53,
    n13,
    n55
  );


  nor
  g179
  (
    n77,
    n53,
    n32,
    n44,
    n16
  );


  nor
  g180
  (
    n98,
    n34,
    n3,
    n13,
    n10
  );


  nor
  g181
  (
    KeyWire_0_8,
    n17,
    n41,
    n59,
    n16
  );


  or
  g182
  (
    n164,
    n51,
    n44,
    n17,
    n38
  );


  xor
  g183
  (
    n105,
    n61,
    n36,
    n8,
    n6
  );


  not
  g184
  (
    n204,
    n64
  );


  not
  g185
  (
    n203,
    n65
  );


  not
  g186
  (
    n211,
    n204
  );


  not
  g187
  (
    n210,
    n204
  );


  buf
  g188
  (
    n212,
    n63
  );


  not
  g189
  (
    n207,
    n204
  );


  not
  g190
  (
    n209,
    n203
  );


  buf
  g191
  (
    n205,
    n203
  );


  not
  g192
  (
    n208,
    n203
  );


  or
  g193
  (
    n206,
    n203,
    n63,
    n204
  );


  and
  g194
  (
    n215,
    n210,
    n94,
    n212,
    n114
  );


  xor
  g195
  (
    n220,
    n101,
    n74,
    n73,
    n80
  );


  nand
  g196
  (
    n224,
    n104,
    n112,
    n101,
    n103
  );


  and
  g197
  (
    n233,
    n207,
    n104,
    n102,
    n86
  );


  or
  g198
  (
    KeyWire_0_2,
    n106,
    n207,
    n114,
    n99
  );


  nor
  g199
  (
    n228,
    n107,
    n212,
    n102,
    n84
  );


  xnor
  g200
  (
    n244,
    n97,
    n101,
    n212,
    n110
  );


  nor
  g201
  (
    n243,
    n111,
    n110,
    n106,
    n208
  );


  or
  g202
  (
    n240,
    n87,
    n93,
    n113,
    n81
  );


  nand
  g203
  (
    n236,
    n72,
    n211,
    n91,
    n114
  );


  xnor
  g204
  (
    n238,
    n209,
    n209,
    n112,
    n115
  );


  nand
  g205
  (
    n234,
    n205,
    n88,
    n104,
    n115
  );


  xor
  g206
  (
    n237,
    n210,
    n102,
    n100,
    n90
  );


  xnor
  g207
  (
    n226,
    n106,
    n208,
    n205,
    n75
  );


  xnor
  g208
  (
    n219,
    n205,
    n100,
    n109,
    n111
  );


  nor
  g209
  (
    n222,
    n114,
    n98,
    n79,
    n211
  );


  nor
  g210
  (
    n217,
    n100,
    n206,
    n110,
    n85
  );


  or
  g211
  (
    n242,
    n70,
    n110,
    n103,
    n111
  );


  and
  g212
  (
    n214,
    n105,
    n105,
    n207,
    n100
  );


  and
  g213
  (
    n239,
    n95,
    n109,
    n108,
    n83
  );


  xor
  g214
  (
    n235,
    n205,
    n106,
    n210,
    n108
  );


  xnor
  g215
  (
    n225,
    n82,
    n96,
    n211,
    n67
  );


  and
  g216
  (
    n229,
    n108,
    n109,
    n103,
    n113
  );


  xnor
  g217
  (
    n221,
    n68,
    n207,
    n107
  );


  xnor
  g218
  (
    n216,
    n109,
    n103,
    n92,
    n111
  );


  xor
  g219
  (
    n227,
    n206,
    n206,
    n209,
    n112
  );


  nor
  g220
  (
    n230,
    n206,
    n108,
    n113,
    n89
  );


  nand
  g221
  (
    n223,
    n105,
    n101,
    n102,
    n77
  );


  xor
  g222
  (
    n232,
    n113,
    n107,
    n69,
    n208
  );


  xor
  g223
  (
    n213,
    n212,
    n209,
    n71,
    n208
  );


  xor
  g224
  (
    n218,
    n66,
    n210,
    n76,
    n78
  );


  xnor
  g225
  (
    n241,
    n104,
    n105,
    n211,
    n112
  );


  not
  g226
  (
    n249,
    n216
  );


  buf
  g227
  (
    n247,
    n214
  );


  buf
  g228
  (
    n250,
    n219
  );


  not
  g229
  (
    n246,
    n115
  );


  buf
  g230
  (
    n251,
    n116
  );


  nand
  g231
  (
    n248,
    n218,
    n215,
    n213,
    n116
  );


  xor
  g232
  (
    n245,
    n217,
    n116,
    n115
  );


  not
  g233
  (
    n260,
    n119
  );


  buf
  g234
  (
    n274,
    n251
  );


  buf
  g235
  (
    n265,
    n122
  );


  buf
  g236
  (
    KeyWire_0_10,
    n249
  );


  not
  g237
  (
    n273,
    n122
  );


  buf
  g238
  (
    n267,
    n248
  );


  buf
  g239
  (
    n269,
    n117
  );


  buf
  g240
  (
    n255,
    n250
  );


  buf
  g241
  (
    n276,
    n123
  );


  not
  g242
  (
    n259,
    n121
  );


  buf
  g243
  (
    n252,
    n117
  );


  xnor
  g244
  (
    n272,
    n120,
    n247,
    n123
  );


  or
  g245
  (
    n268,
    n248,
    n120,
    n121
  );


  xnor
  g246
  (
    n277,
    n118,
    n117,
    n119
  );


  nand
  g247
  (
    n261,
    n246,
    n120,
    n122
  );


  xnor
  g248
  (
    n253,
    n246,
    n119,
    n247
  );


  and
  g249
  (
    n266,
    n249,
    n250,
    n247
  );


  or
  g250
  (
    n258,
    n251,
    n248,
    n246
  );


  nand
  g251
  (
    n263,
    n118,
    n245,
    n122
  );


  xnor
  g252
  (
    n256,
    n123,
    n118,
    n245
  );


  or
  g253
  (
    n270,
    n251,
    n117,
    n120
  );


  nand
  g254
  (
    n262,
    n124,
    n249,
    n123
  );


  nor
  g255
  (
    n254,
    n250,
    n121
  );


  or
  g256
  (
    n264,
    n249,
    n124,
    n251
  );


  nand
  g257
  (
    n275,
    n118,
    n246,
    n119
  );


  and
  g258
  (
    n257,
    n247,
    n250,
    n248
  );


  not
  g259
  (
    n333,
    n143
  );


  buf
  g260
  (
    n331,
    n141
  );


  buf
  g261
  (
    n346,
    n130
  );


  buf
  g262
  (
    n324,
    n130
  );


  not
  g263
  (
    n348,
    n252
  );


  not
  g264
  (
    n310,
    n266
  );


  buf
  g265
  (
    n292,
    n145
  );


  not
  g266
  (
    n349,
    n266
  );


  not
  g267
  (
    n369,
    n259
  );


  not
  g268
  (
    n364,
    n273
  );


  not
  g269
  (
    n361,
    n264
  );


  buf
  g270
  (
    n284,
    n135
  );


  not
  g271
  (
    n315,
    n270
  );


  not
  g272
  (
    n343,
    n124
  );


  buf
  g273
  (
    n353,
    n142
  );


  buf
  g274
  (
    n347,
    n267
  );


  buf
  g275
  (
    n357,
    n238
  );


  buf
  g276
  (
    n325,
    n267
  );


  buf
  g277
  (
    n293,
    n137
  );


  buf
  g278
  (
    n359,
    n139
  );


  buf
  g279
  (
    n354,
    n254
  );


  buf
  g280
  (
    n278,
    n234
  );


  buf
  g281
  (
    n320,
    n226
  );


  not
  g282
  (
    n290,
    n144
  );


  not
  g283
  (
    n296,
    n236
  );


  not
  g284
  (
    n306,
    n239
  );


  not
  g285
  (
    n304,
    n127
  );


  not
  g286
  (
    n335,
    n131
  );


  buf
  g287
  (
    n336,
    n128
  );


  buf
  g288
  (
    n326,
    n222
  );


  not
  g289
  (
    n367,
    n228
  );


  not
  g290
  (
    n339,
    n269
  );


  nor
  g291
  (
    n332,
    n258,
    n131,
    n137
  );


  xnor
  g292
  (
    n297,
    n241,
    n259,
    n260
  );


  xor
  g293
  (
    n281,
    n131,
    n256,
    n127
  );


  or
  g294
  (
    n329,
    n142,
    n271,
    n272
  );


  and
  g295
  (
    KeyWire_0_6,
    n134,
    n257,
    n267
  );


  or
  g296
  (
    n371,
    n244,
    n253,
    n268
  );


  nor
  g297
  (
    KeyWire_0_12,
    n275,
    n252,
    n225
  );


  or
  g298
  (
    n365,
    n273,
    n140,
    n242
  );


  xor
  g299
  (
    n305,
    n136,
    n237,
    n270
  );


  or
  g300
  (
    n298,
    n236,
    n271,
    n227
  );


  nand
  g301
  (
    n286,
    n270,
    n261,
    n254
  );


  nor
  g302
  (
    n317,
    n130,
    n133,
    n220
  );


  nor
  g303
  (
    n344,
    n274,
    n125,
    n275
  );


  xor
  g304
  (
    n285,
    n262,
    n258,
    n238
  );


  nand
  g305
  (
    n288,
    n244,
    n255,
    n258
  );


  nor
  g306
  (
    n372,
    n260,
    n261,
    n266
  );


  and
  g307
  (
    n341,
    n240,
    n142,
    n275
  );


  nor
  g308
  (
    n308,
    n235,
    n256,
    n139
  );


  xor
  g309
  (
    n360,
    n242,
    n138,
    n255
  );


  xnor
  g310
  (
    n300,
    n263,
    n128,
    n231
  );


  xor
  g311
  (
    n283,
    n242,
    n127,
    n272
  );


  xor
  g312
  (
    n295,
    n143,
    n259,
    n274
  );


  nand
  g313
  (
    n309,
    n129,
    n271,
    n270
  );


  xnor
  g314
  (
    n318,
    n263,
    n136,
    n274
  );


  nor
  g315
  (
    n338,
    n265,
    n125,
    n271
  );


  nand
  g316
  (
    n313,
    n145,
    n144,
    n269
  );


  nor
  g317
  (
    n280,
    n257,
    n259,
    n232
  );


  nor
  g318
  (
    n350,
    n138,
    n260,
    n257
  );


  xnor
  g319
  (
    n302,
    n265,
    n260,
    n241
  );


  or
  g320
  (
    n323,
    n233,
    n243,
    n140
  );


  nand
  g321
  (
    n303,
    n244,
    n136,
    n241
  );


  or
  g322
  (
    n307,
    n143,
    n135,
    n126
  );


  nor
  g323
  (
    n299,
    n132,
    n268,
    n255
  );


  xnor
  g324
  (
    n351,
    n141,
    n243,
    n240
  );


  xor
  g325
  (
    n312,
    n137,
    n141,
    n134
  );


  nand
  g326
  (
    n366,
    n264,
    n263,
    n261
  );


  and
  g327
  (
    n321,
    n266,
    n143,
    n134
  );


  xnor
  g328
  (
    n356,
    n134,
    n267,
    n274
  );


  and
  g329
  (
    n319,
    n273,
    n224,
    n124
  );


  xnor
  g330
  (
    n328,
    n130,
    n258,
    n133
  );


  and
  g331
  (
    n287,
    n133,
    n256,
    n229
  );


  nor
  g332
  (
    n294,
    n129,
    n141,
    n126
  );


  and
  g333
  (
    n291,
    n253,
    n223,
    n252
  );


  and
  g334
  (
    n282,
    n129,
    n262,
    n257
  );


  and
  g335
  (
    n342,
    n262,
    n230,
    n132
  );


  nand
  g336
  (
    n368,
    n139,
    n221,
    n135
  );


  or
  g337
  (
    n301,
    n127,
    n261,
    n269
  );


  or
  g338
  (
    n358,
    n142,
    n273,
    n132
  );


  or
  g339
  (
    n327,
    n135,
    n237,
    n145
  );


  nor
  g340
  (
    n362,
    n243,
    n125,
    n138
  );


  xor
  g341
  (
    n316,
    n144,
    n265,
    n256
  );


  nor
  g342
  (
    n330,
    n275,
    n262,
    n131
  );


  xor
  g343
  (
    n370,
    n239,
    n268,
    n144
  );


  nor
  g344
  (
    n373,
    n272,
    n145,
    n265
  );


  or
  g345
  (
    n352,
    n268,
    n126,
    n263
  );


  xnor
  g346
  (
    n289,
    n264,
    n244,
    n254
  );


  nand
  g347
  (
    n311,
    n242,
    n129,
    n137
  );


  xnor
  g348
  (
    n355,
    n125,
    n132,
    n243
  );


  xor
  g349
  (
    n314,
    n139,
    n253,
    n136
  );


  xor
  g350
  (
    n363,
    n254,
    n138,
    n128
  );


  and
  g351
  (
    n279,
    n133,
    n252,
    n269
  );


  nor
  g352
  (
    n334,
    n253,
    n140,
    n272
  );


  nand
  g353
  (
    n345,
    n241,
    n126,
    n128
  );


  and
  g354
  (
    n322,
    n264,
    n255,
    n140
  );


  xor
  g355
  (
    n411,
    n284,
    n331,
    n359,
    n332
  );


  xnor
  g356
  (
    n403,
    n332,
    n321,
    n339,
    n335
  );


  xor
  g357
  (
    n409,
    n351,
    n312,
    n283,
    n358
  );


  or
  g358
  (
    n376,
    n341,
    n301,
    n342,
    n332
  );


  and
  g359
  (
    n406,
    n290,
    n345,
    n299,
    n335
  );


  nor
  g360
  (
    n444,
    n324,
    n349,
    n313,
    n348
  );


  and
  g361
  (
    n401,
    n345,
    n338,
    n342,
    n303
  );


  xnor
  g362
  (
    n435,
    n355,
    n287,
    n304,
    n318
  );


  nand
  g363
  (
    n384,
    n306,
    n323,
    n315,
    n330
  );


  xor
  g364
  (
    n386,
    n344,
    n315,
    n337,
    n347
  );


  nor
  g365
  (
    n441,
    n328,
    n341,
    n316,
    n282
  );


  nor
  g366
  (
    n414,
    n316,
    n346,
    n313,
    n320
  );


  xnor
  g367
  (
    n394,
    n293,
    n302,
    n281,
    n326
  );


  or
  g368
  (
    n379,
    n329,
    n327,
    n334,
    n350
  );


  nand
  g369
  (
    n419,
    n287,
    n296,
    n302,
    n306
  );


  and
  g370
  (
    n415,
    n285,
    n312,
    n348,
    n334
  );


  xor
  g371
  (
    n385,
    n282,
    n339,
    n321,
    n324
  );


  nor
  g372
  (
    n442,
    n310,
    n290,
    n295,
    n317
  );


  and
  g373
  (
    n383,
    n354,
    n326,
    n279,
    n353
  );


  xor
  g374
  (
    n454,
    n311,
    n292,
    n333,
    n334
  );


  xnor
  g375
  (
    n421,
    n354,
    n288,
    n355,
    n312
  );


  and
  g376
  (
    n408,
    n308,
    n287,
    n283,
    n291
  );


  or
  g377
  (
    n377,
    n346,
    n297,
    n315,
    n289
  );


  nor
  g378
  (
    n378,
    n299,
    n357,
    n316,
    n305
  );


  nand
  g379
  (
    n429,
    n287,
    n333,
    n307,
    n299
  );


  nand
  g380
  (
    n433,
    n294,
    n293,
    n308,
    n325
  );


  and
  g381
  (
    n405,
    n322,
    n285,
    n323,
    n304
  );


  nor
  g382
  (
    n423,
    n336,
    n278,
    n330,
    n360
  );


  nor
  g383
  (
    n450,
    n289,
    n279,
    n288,
    n338
  );


  xnor
  g384
  (
    n380,
    n322,
    n324,
    n303,
    n326
  );


  xnor
  g385
  (
    n390,
    n341,
    n291,
    n290,
    n298
  );


  nand
  g386
  (
    n393,
    n296,
    n310,
    n300,
    n281
  );


  or
  g387
  (
    n396,
    n319,
    n344,
    n298,
    n353
  );


  nor
  g388
  (
    n381,
    n338,
    n360,
    n340,
    n346
  );


  or
  g389
  (
    n446,
    n301,
    n339,
    n359,
    n357
  );


  and
  g390
  (
    n447,
    n314,
    n334,
    n320,
    n295
  );


  nor
  g391
  (
    n426,
    n356,
    n279,
    n350,
    n285
  );


  nand
  g392
  (
    n434,
    n355,
    n354,
    n328,
    n313
  );


  nand
  g393
  (
    n374,
    n302,
    n355,
    n326,
    n323
  );


  xor
  g394
  (
    KeyWire_0_0,
    n301,
    n342,
    n283,
    n288
  );


  xor
  g395
  (
    n456,
    n328,
    n343,
    n280,
    n311
  );


  xor
  g396
  (
    n445,
    n359,
    n341,
    n339,
    n342
  );


  or
  g397
  (
    n438,
    n305,
    n320,
    n315,
    n344
  );


  nand
  g398
  (
    n440,
    n350,
    n286,
    n329,
    n357
  );


  xor
  g399
  (
    n425,
    n313,
    n286,
    n332,
    n349
  );


  and
  g400
  (
    n413,
    n357,
    n349,
    n280,
    n358
  );


  or
  g401
  (
    n375,
    n318,
    n300,
    n325,
    n351
  );


  or
  g402
  (
    n439,
    n353,
    n288,
    n327,
    n304
  );


  xnor
  g403
  (
    n422,
    n314,
    n284,
    n331,
    n297
  );


  xor
  g404
  (
    n418,
    n359,
    n282,
    n343,
    n356
  );


  and
  g405
  (
    n416,
    n281,
    n310,
    n327,
    n280
  );


  nand
  g406
  (
    n398,
    n340,
    n297,
    n292,
    n338
  );


  and
  g407
  (
    n388,
    n309,
    n319,
    n337,
    n360
  );


  or
  g408
  (
    n404,
    n328,
    n279,
    n304,
    n289
  );


  and
  g409
  (
    n412,
    n300,
    n345,
    n352
  );


  xnor
  g410
  (
    n407,
    n356,
    n337,
    n286,
    n347
  );


  and
  g411
  (
    n397,
    n308,
    n333,
    n291,
    n335
  );


  xor
  g412
  (
    n420,
    n336,
    n350,
    n302,
    n280
  );


  nor
  g413
  (
    n410,
    n283,
    n330,
    n317,
    n289
  );


  xor
  g414
  (
    n402,
    n310,
    n295,
    n278,
    n285
  );


  nand
  g415
  (
    n389,
    n344,
    n294,
    n297,
    n305
  );


  xnor
  g416
  (
    n455,
    n343,
    n336,
    n281,
    n348
  );


  xor
  g417
  (
    n417,
    n335,
    n329,
    n293,
    n343
  );


  nand
  g418
  (
    KeyWire_0_3,
    n309,
    n323,
    n358,
    n352
  );


  or
  g419
  (
    n428,
    n330,
    n345,
    n331,
    n306
  );


  and
  g420
  (
    n391,
    n337,
    n346,
    n294,
    n308
  );


  or
  g421
  (
    n449,
    n290,
    n296,
    n298,
    n348
  );


  nand
  g422
  (
    n387,
    n322,
    n351,
    n327,
    n349
  );


  nor
  g423
  (
    n395,
    n293,
    n305,
    n347,
    n278
  );


  nand
  g424
  (
    n437,
    n336,
    n286,
    n319,
    n353
  );


  and
  g425
  (
    n436,
    n278,
    n295,
    n312,
    n294
  );


  or
  g426
  (
    n400,
    n352,
    n309,
    n354,
    n298
  );


  nand
  g427
  (
    n443,
    n316,
    n325,
    n296,
    n340
  );


  nor
  g428
  (
    n382,
    n292,
    n358,
    n319,
    n321
  );


  nor
  g429
  (
    n399,
    n321,
    n300,
    n291,
    n303
  );


  and
  g430
  (
    n448,
    n318,
    n314,
    n329,
    n306
  );


  xor
  g431
  (
    n431,
    n309,
    n340,
    n318,
    n356
  );


  or
  g432
  (
    n392,
    n292,
    n324,
    n331,
    n303
  );


  nor
  g433
  (
    n430,
    n307,
    n322,
    n311,
    n360
  );


  xor
  g434
  (
    n427,
    n320,
    n299,
    n351,
    n314
  );


  xor
  g435
  (
    n453,
    n284,
    n284,
    n307,
    n333
  );


  nor
  g436
  (
    n451,
    n311,
    n347,
    n307,
    n301
  );


  xnor
  g437
  (
    n424,
    n325,
    n282,
    n317
  );


  not
  g438
  (
    n464,
    n390
  );


  buf
  g439
  (
    n471,
    n382
  );


  buf
  g440
  (
    n459,
    n377
  );


  not
  g441
  (
    n477,
    n381
  );


  not
  g442
  (
    n472,
    n379
  );


  buf
  g443
  (
    n467,
    n395
  );


  not
  g444
  (
    n461,
    n380
  );


  buf
  g445
  (
    n476,
    n392
  );


  buf
  g446
  (
    n460,
    n386
  );


  not
  g447
  (
    n468,
    n374
  );


  buf
  g448
  (
    n466,
    n384
  );


  buf
  g449
  (
    n470,
    n385
  );


  not
  g450
  (
    n474,
    n376
  );


  buf
  g451
  (
    n469,
    n375
  );


  buf
  g452
  (
    n473,
    n387
  );


  buf
  g453
  (
    n462,
    n394
  );


  not
  g454
  (
    n458,
    n391
  );


  not
  g455
  (
    n478,
    n383
  );


  buf
  g456
  (
    n465,
    n378
  );


  buf
  g457
  (
    n475,
    n393
  );


  not
  g458
  (
    n457,
    n389
  );


  buf
  g459
  (
    n463,
    n388
  );


  nor
  g460
  (
    n481,
    n361,
    n369,
    n371,
    n460
  );


  xor
  g461
  (
    n479,
    n362,
    n459,
    n368,
    n457
  );


  nor
  g462
  (
    n483,
    n457,
    n363
  );


  xnor
  g463
  (
    n480,
    n461,
    n459,
    n365,
    n369
  );


  xnor
  g464
  (
    n482,
    n364,
    n365,
    n460,
    n368
  );


  nor
  g465
  (
    n494,
    n457,
    n372,
    n367,
    n364
  );


  xnor
  g466
  (
    n486,
    n458,
    n371,
    n459
  );


  or
  g467
  (
    n495,
    n366,
    n373,
    n370
  );


  nor
  g468
  (
    n490,
    n367,
    n372,
    n365,
    n371
  );


  or
  g469
  (
    n492,
    n458,
    n457,
    n459,
    n370
  );


  xor
  g470
  (
    n485,
    n368,
    n368,
    n370,
    n372
  );


  nand
  g471
  (
    n487,
    n458,
    n361,
    n366
  );


  and
  g472
  (
    n488,
    n369,
    n364,
    n361,
    n365
  );


  xnor
  g473
  (
    n484,
    n364,
    n363,
    n458,
    n362
  );


  and
  g474
  (
    n489,
    n366,
    n362,
    n369
  );


  or
  g475
  (
    n491,
    n373,
    n460,
    n367,
    n370
  );


  and
  g476
  (
    n493,
    n367,
    n361,
    n372,
    n460
  );


  not
  g477
  (
    n510,
    n494
  );


  buf
  g478
  (
    n511,
    n481
  );


  not
  g479
  (
    n507,
    n480
  );


  not
  g480
  (
    n503,
    n483
  );


  not
  g481
  (
    n504,
    n482
  );


  not
  g482
  (
    n506,
    n485
  );


  buf
  g483
  (
    n497,
    n484
  );


  buf
  g484
  (
    n496,
    n486
  );


  buf
  g485
  (
    n505,
    n493
  );


  buf
  g486
  (
    n502,
    n490
  );


  not
  g487
  (
    n508,
    n479
  );


  buf
  g488
  (
    n500,
    n487
  );


  buf
  g489
  (
    n499,
    n489
  );


  not
  g490
  (
    n501,
    n488
  );


  buf
  g491
  (
    n498,
    n491
  );


  buf
  g492
  (
    n509,
    n492
  );


  nor
  g493
  (
    n513,
    n473,
    n463,
    n399,
    n423
  );


  nor
  g494
  (
    n540,
    n472,
    n499,
    n464,
    n400
  );


  xnor
  g495
  (
    n538,
    n469,
    n476,
    n427,
    n500
  );


  or
  g496
  (
    n547,
    n474,
    n503,
    n404
  );


  nor
  g497
  (
    n536,
    n442,
    n475,
    n424,
    n499
  );


  xnor
  g498
  (
    n550,
    n406,
    n471,
    n412,
    n497
  );


  xnor
  g499
  (
    n548,
    n422,
    n468,
    n436,
    n475
  );


  xnor
  g500
  (
    n521,
    n431,
    n428,
    n498,
    n506
  );


  nor
  g501
  (
    n522,
    n461,
    n438,
    n473,
    n470
  );


  or
  g502
  (
    n552,
    n496,
    n472,
    n441,
    n466
  );


  xor
  g503
  (
    KeyWire_0_5,
    n502,
    n467,
    n430,
    n417
  );


  and
  g504
  (
    n524,
    n476,
    n476,
    n464,
    n477
  );


  xor
  g505
  (
    n516,
    n439,
    n466,
    n501
  );


  and
  g506
  (
    n545,
    n465,
    n469,
    n435,
    n146
  );


  nand
  g507
  (
    n528,
    n462,
    n463,
    n461,
    n474
  );


  or
  g508
  (
    n526,
    n500,
    n469,
    n402,
    n398
  );


  xor
  g509
  (
    n543,
    n476,
    n401,
    n465,
    n475
  );


  nor
  g510
  (
    n518,
    n501,
    n478,
    n500,
    n433
  );


  nand
  g511
  (
    n541,
    n405,
    n470,
    n429,
    n502
  );


  xor
  g512
  (
    n542,
    n503,
    n415,
    n474,
    n408
  );


  xor
  g513
  (
    n554,
    n465,
    n462,
    n496,
    n475
  );


  or
  g514
  (
    KeyWire_0_11,
    n478,
    n472,
    n464,
    n447
  );


  nand
  g515
  (
    n544,
    n468,
    n413,
    n471,
    n497
  );


  nor
  g516
  (
    n535,
    n414,
    n506,
    n501,
    n146
  );


  xnor
  g517
  (
    n515,
    n470,
    n498,
    n499,
    n373
  );


  and
  g518
  (
    n517,
    n473,
    n478,
    n461,
    n467
  );


  and
  g519
  (
    n531,
    n496,
    n463,
    n409,
    n446
  );


  nor
  g520
  (
    n546,
    n416,
    n462,
    n504
  );


  xnor
  g521
  (
    n527,
    n465,
    n462,
    n505,
    n146
  );


  xor
  g522
  (
    n512,
    n418,
    n467,
    n505,
    n498
  );


  xor
  g523
  (
    n537,
    n443,
    n471,
    n407
  );


  nor
  g524
  (
    n523,
    n499,
    n397,
    n468,
    n496
  );


  xnor
  g525
  (
    n534,
    n477,
    n421,
    n146,
    n432
  );


  nand
  g526
  (
    n530,
    n506,
    n466,
    n467,
    n464
  );


  nand
  g527
  (
    n533,
    n504,
    n498,
    n478,
    n437
  );


  nand
  g528
  (
    n520,
    n500,
    n420,
    n473,
    n468
  );


  or
  g529
  (
    n514,
    n426,
    n410,
    n469,
    n445
  );


  xor
  g530
  (
    n549,
    n403,
    n505,
    n497,
    n440
  );


  nor
  g531
  (
    n529,
    n505,
    n472,
    n504,
    n470
  );


  and
  g532
  (
    n551,
    n411,
    n502,
    n503,
    n425
  );


  nand
  g533
  (
    n553,
    n466,
    n497,
    n396,
    n448
  );


  xor
  g534
  (
    n525,
    n434,
    n502,
    n444,
    n419
  );


  nand
  g535
  (
    n539,
    n477,
    n477,
    n474,
    n463
  );


  nand
  g536
  (
    n556,
    n183,
    n526,
    n149,
    n170
  );


  nand
  g537
  (
    n597,
    n152,
    n151,
    n526,
    n169
  );


  or
  g538
  (
    n592,
    n149,
    n177,
    n520,
    n170
  );


  nand
  g539
  (
    n583,
    n166,
    n190,
    n514,
    n184
  );


  xnor
  g540
  (
    n566,
    n518,
    n158,
    n167,
    n168
  );


  nand
  g541
  (
    n579,
    n179,
    n173,
    n155,
    n160
  );


  nor
  g542
  (
    n555,
    n512,
    n155,
    n522,
    n154
  );


  and
  g543
  (
    n557,
    n191,
    n188,
    n154,
    n163
  );


  and
  g544
  (
    n582,
    n181,
    n186,
    n167,
    n174
  );


  nor
  g545
  (
    n601,
    n162,
    n162,
    n188,
    n512
  );


  nor
  g546
  (
    n599,
    n525,
    n523,
    n150,
    n147
  );


  nand
  g547
  (
    n571,
    n175,
    n165,
    n154,
    n520
  );


  or
  g548
  (
    n567,
    n147,
    n526,
    n156,
    n184
  );


  xor
  g549
  (
    n585,
    n180,
    n524,
    n152
  );


  xnor
  g550
  (
    n568,
    n521,
    n169,
    n185,
    n184
  );


  nand
  g551
  (
    n598,
    n178,
    n514,
    n516,
    n515
  );


  xor
  g552
  (
    n581,
    n166,
    n156,
    n171
  );


  or
  g553
  (
    n564,
    n157,
    n517,
    n187,
    n495
  );


  and
  g554
  (
    n558,
    n169,
    n171,
    n161,
    n160
  );


  nand
  g555
  (
    n580,
    n525,
    n166,
    n172,
    n520
  );


  nand
  g556
  (
    n609,
    n170,
    n167,
    n153,
    n174
  );


  nor
  g557
  (
    n586,
    n162,
    n190,
    n158,
    n515
  );


  xor
  g558
  (
    n562,
    n157,
    n190,
    n150,
    n191
  );


  xor
  g559
  (
    n591,
    n519,
    n526,
    n517
  );


  and
  g560
  (
    n600,
    n519,
    n159,
    n163,
    n157
  );


  or
  g561
  (
    n603,
    n186,
    n159,
    n521,
    n185
  );


  xor
  g562
  (
    n615,
    n177,
    n149,
    n165,
    n519
  );


  nand
  g563
  (
    n606,
    n183,
    n523,
    n190,
    n169
  );


  xnor
  g564
  (
    n578,
    n166,
    n184,
    n178,
    n180
  );


  and
  g565
  (
    n574,
    n156,
    n148,
    n161,
    n160
  );


  nor
  g566
  (
    n614,
    n177,
    n523,
    n516,
    n515
  );


  xor
  g567
  (
    n576,
    n518,
    n149,
    n185,
    n172
  );


  xor
  g568
  (
    n604,
    n191,
    n179,
    n176,
    n164
  );


  nor
  g569
  (
    n589,
    n150,
    n513,
    n182,
    n192
  );


  nand
  g570
  (
    n611,
    n514,
    n182,
    n191,
    n517
  );


  and
  g571
  (
    n590,
    n516,
    n168,
    n152,
    n175
  );


  nand
  g572
  (
    n572,
    n192,
    n174,
    n173,
    n524
  );


  or
  g573
  (
    n570,
    n178,
    n171,
    n177,
    n186
  );


  and
  g574
  (
    n596,
    n182,
    n164,
    n513,
    n151
  );


  and
  g575
  (
    n608,
    n181,
    n519,
    n155,
    n158
  );


  xnor
  g576
  (
    n569,
    n524,
    n522,
    n188,
    n163
  );


  or
  g577
  (
    n560,
    n153,
    n161,
    n525,
    n176
  );


  or
  g578
  (
    n612,
    n165,
    n189,
    n148,
    n512
  );


  or
  g579
  (
    n613,
    n179,
    n527,
    n172,
    n170
  );


  xor
  g580
  (
    n565,
    n160,
    n522,
    n185,
    n162
  );


  and
  g581
  (
    n573,
    n174,
    n159,
    n173,
    n525
  );


  or
  g582
  (
    n602,
    n522,
    n172,
    n521,
    n153
  );


  nand
  g583
  (
    n607,
    n178,
    n188,
    n521,
    n150
  );


  xor
  g584
  (
    n575,
    n514,
    n175,
    n154,
    n512
  );


  or
  g585
  (
    KeyWire_0_15,
    n158,
    n183,
    n167,
    n164
  );


  nand
  g586
  (
    n593,
    n523,
    n520,
    n189,
    n516
  );


  nand
  g587
  (
    n587,
    n186,
    n518,
    n187,
    n147
  );


  or
  g588
  (
    n584,
    n164,
    n151,
    n518,
    n180
  );


  nor
  g589
  (
    n561,
    n153,
    n165,
    n147,
    n176
  );


  nor
  g590
  (
    n563,
    n183,
    n513,
    n181
  );


  nor
  g591
  (
    n595,
    n187,
    n163,
    n515,
    n173
  );


  xor
  g592
  (
    n588,
    n159,
    n189,
    n155,
    n152
  );


  and
  g593
  (
    n605,
    n176,
    n187,
    n180,
    n156
  );


  nor
  g594
  (
    n559,
    n157,
    n182,
    n168,
    n148
  );


  nor
  g595
  (
    n594,
    n151,
    n148,
    n168,
    n189
  );


  xnor
  g596
  (
    n577,
    n161,
    n179,
    n175,
    n513
  );


  or
  g597
  (
    n669,
    n594,
    n570,
    n557,
    n593
  );


  nor
  g598
  (
    n684,
    n575,
    n558,
    n599,
    n571
  );


  or
  g599
  (
    n674,
    n615,
    n450,
    n562,
    n567
  );


  or
  g600
  (
    n651,
    n588,
    n602,
    n573
  );


  or
  g601
  (
    n676,
    n605,
    n603,
    n199,
    n198
  );


  and
  g602
  (
    n632,
    n593,
    n573,
    n193,
    n612
  );


  xor
  g603
  (
    n667,
    n506,
    n590,
    n193,
    n561
  );


  nand
  g604
  (
    n685,
    n510,
    n198,
    n563,
    n574
  );


  or
  g605
  (
    n627,
    n585,
    n601,
    n590,
    n599
  );


  nor
  g606
  (
    n658,
    n589,
    n198,
    n197,
    n194
  );


  xnor
  g607
  (
    n660,
    n589,
    n615,
    n194,
    n201
  );


  xnor
  g608
  (
    n645,
    n455,
    n584,
    n596,
    n566
  );


  nor
  g609
  (
    n647,
    n579,
    n578,
    n613,
    n608
  );


  and
  g610
  (
    n654,
    n586,
    n558,
    n510,
    n559
  );


  nor
  g611
  (
    n673,
    n586,
    n606,
    n582,
    n508
  );


  nor
  g612
  (
    n665,
    n611,
    n507,
    n574,
    n195
  );


  nor
  g613
  (
    n671,
    n583,
    n200,
    n507,
    n563
  );


  xnor
  g614
  (
    n664,
    n195,
    n570,
    n192,
    n562
  );


  or
  g615
  (
    n686,
    n602,
    n597,
    n615,
    n599
  );


  nand
  g616
  (
    n631,
    n591,
    n194,
    n577,
    n600
  );


  and
  g617
  (
    n634,
    n197,
    n510,
    n611,
    n606
  );


  nor
  g618
  (
    n657,
    n585,
    n200,
    n608,
    n594
  );


  xor
  g619
  (
    n656,
    n569,
    n566,
    n603,
    n588
  );


  nor
  g620
  (
    n663,
    n580,
    n600,
    n592,
    n583
  );


  xnor
  g621
  (
    n668,
    n563,
    n451,
    n576,
    n564
  );


  xnor
  g622
  (
    n633,
    n575,
    n605,
    n612,
    n609
  );


  xor
  g623
  (
    n643,
    n599,
    n575,
    n511,
    n564
  );


  nor
  g624
  (
    n661,
    n558,
    n508,
    n588,
    n576
  );


  nor
  g625
  (
    n689,
    n573,
    n576,
    n567
  );


  nand
  g626
  (
    n680,
    n614,
    n596,
    n564,
    n507
  );


  or
  g627
  (
    n644,
    n580,
    n508,
    n571,
    n558
  );


  xnor
  g628
  (
    n630,
    n587,
    n202,
    n564,
    n509
  );


  and
  g629
  (
    n629,
    n611,
    n596,
    n562,
    n600
  );


  nor
  g630
  (
    n659,
    n614,
    n595,
    n591,
    n578
  );


  and
  g631
  (
    n662,
    n598,
    n604,
    n585,
    n581
  );


  or
  g632
  (
    n638,
    n582,
    n584,
    n601,
    n511
  );


  or
  g633
  (
    n677,
    n566,
    n605,
    n615,
    n593
  );


  and
  g634
  (
    n681,
    n562,
    n201,
    n567,
    n608
  );


  or
  g635
  (
    n652,
    n597,
    n613,
    n596,
    n576
  );


  nand
  g636
  (
    n655,
    n585,
    n509,
    n595,
    n201
  );


  nor
  g637
  (
    n628,
    n578,
    n586,
    n588,
    n570
  );


  xnor
  g638
  (
    KeyWire_0_9,
    n557,
    n597,
    n572,
    n574
  );


  nand
  g639
  (
    n623,
    n598,
    n607,
    n565,
    n571
  );


  or
  g640
  (
    n636,
    n559,
    n590,
    n579,
    n581
  );


  or
  g641
  (
    n653,
    n196,
    n589,
    n199,
    n193
  );


  or
  g642
  (
    n640,
    n509,
    n196,
    n197,
    n508
  );


  xnor
  g643
  (
    n691,
    n559,
    n507,
    n566,
    n583
  );


  nor
  g644
  (
    n635,
    n587,
    n579,
    n200,
    n201
  );


  nor
  g645
  (
    n646,
    n613,
    n577,
    n607,
    n561
  );


  and
  g646
  (
    n624,
    n572,
    n595,
    n560,
    n556
  );


  and
  g647
  (
    n625,
    n195,
    n591,
    n608,
    n561
  );


  or
  g648
  (
    n648,
    n563,
    n589,
    n569
  );


  xnor
  g649
  (
    n639,
    n449,
    n610,
    n194,
    n592
  );


  nor
  g650
  (
    n690,
    n577,
    n610,
    n584,
    n580
  );


  nor
  g651
  (
    n649,
    n565,
    n560,
    n609,
    n510
  );


  nor
  g652
  (
    n641,
    n452,
    n453,
    n560,
    n602
  );


  and
  g653
  (
    n688,
    n197,
    n594,
    n565,
    n196
  );


  or
  g654
  (
    n682,
    n587,
    n195,
    n511,
    n603
  );


  xnor
  g655
  (
    n626,
    n606,
    n582,
    n200,
    n614
  );


  xnor
  g656
  (
    n616,
    n601,
    n590,
    n573,
    n582
  );


  xnor
  g657
  (
    n622,
    n601,
    n609,
    n598,
    n568
  );


  xor
  g658
  (
    n672,
    n559,
    n196,
    n612,
    n610
  );


  or
  g659
  (
    n678,
    n198,
    n509,
    n569,
    n606
  );


  xor
  g660
  (
    n621,
    n577,
    n612,
    n610,
    n586
  );


  nand
  g661
  (
    n679,
    n604,
    n592,
    n192,
    n583
  );


  xnor
  g662
  (
    n617,
    n575,
    n611,
    n603,
    n454
  );


  or
  g663
  (
    n618,
    n572,
    n555,
    n609,
    n580
  );


  nor
  g664
  (
    n675,
    n511,
    n604,
    n613,
    n592
  );


  xnor
  g665
  (
    n620,
    n607,
    n605,
    n199,
    n568
  );


  and
  g666
  (
    n619,
    n199,
    n595,
    n572,
    n584
  );


  and
  g667
  (
    n637,
    n581,
    n598,
    n593,
    n561
  );


  nor
  g668
  (
    n683,
    n571,
    n565,
    n581,
    n614
  );


  xnor
  g669
  (
    n670,
    n607,
    n560,
    n587,
    n456
  );


  nor
  g670
  (
    n642,
    n600,
    n193,
    n594,
    n568
  );


  nor
  g671
  (
    n650,
    n597,
    n570,
    n574,
    n578
  );


  and
  g672
  (
    n666,
    n579,
    n604,
    n591,
    n568
  );


  xor
  g673
  (
    n713,
    n553,
    n532,
    n528,
    n622
  );


  and
  g674
  (
    n702,
    n530,
    n648,
    n546,
    n642
  );


  nor
  g675
  (
    n726,
    n535,
    n625,
    n546,
    n542
  );


  or
  g676
  (
    n693,
    n544,
    n651,
    n532,
    n542
  );


  xnor
  g677
  (
    n715,
    n551,
    n616,
    n532,
    n623
  );


  nor
  g678
  (
    n694,
    n542,
    n537,
    n548,
    n531
  );


  or
  g679
  (
    n706,
    n554,
    n636,
    n530,
    n529
  );


  and
  g680
  (
    n723,
    n542,
    n632,
    n629,
    n553
  );


  xor
  g681
  (
    n728,
    n534,
    n541,
    n545,
    n549
  );


  or
  g682
  (
    n709,
    n527,
    n540,
    n547,
    n534
  );


  nor
  g683
  (
    n707,
    n529,
    n533,
    n537,
    n552
  );


  or
  g684
  (
    n712,
    n531,
    n535,
    n534,
    n638
  );


  and
  g685
  (
    n697,
    n553,
    n548,
    n545,
    n551
  );


  or
  g686
  (
    n701,
    n635,
    n543,
    n545,
    n539
  );


  and
  g687
  (
    n722,
    n538,
    n631,
    n551,
    n537
  );


  nor
  g688
  (
    n692,
    n538,
    n543,
    n548,
    n533
  );


  xnor
  g689
  (
    KeyWire_0_4,
    n628,
    n536,
    n550,
    n549
  );


  and
  g690
  (
    n721,
    n546,
    n545,
    n533,
    n536
  );


  or
  g691
  (
    n696,
    n554,
    n550,
    n553,
    n640
  );


  and
  g692
  (
    n708,
    n548,
    n528,
    n645
  );


  xnor
  g693
  (
    n698,
    n634,
    n540,
    n527,
    n554
  );


  xor
  g694
  (
    n703,
    n539,
    n549,
    n619,
    n532
  );


  xnor
  g695
  (
    n695,
    n547,
    n530,
    n626,
    n550
  );


  and
  g696
  (
    n700,
    n652,
    n650,
    n530,
    n546
  );


  nor
  g697
  (
    n727,
    n543,
    n641,
    n649,
    n643
  );


  nand
  g698
  (
    n724,
    n536,
    n541,
    n535,
    n550
  );


  xnor
  g699
  (
    n714,
    n549,
    n528,
    n544,
    n539
  );


  xor
  g700
  (
    n719,
    n527,
    n543,
    n639,
    n547
  );


  xnor
  g701
  (
    n718,
    n534,
    n617,
    n552,
    n633
  );


  nand
  g702
  (
    n716,
    n538,
    n541,
    n624,
    n620
  );


  xnor
  g703
  (
    n717,
    n627,
    n630,
    n644,
    n621
  );


  xnor
  g704
  (
    n725,
    n552,
    n540,
    n618
  );


  or
  g705
  (
    n711,
    n539,
    n537,
    n531,
    n544
  );


  nand
  g706
  (
    n705,
    n551,
    n646,
    n647,
    n541
  );


  nand
  g707
  (
    n704,
    n538,
    n533,
    n536,
    n637
  );


  nand
  g708
  (
    n710,
    n531,
    n547,
    n529,
    n535
  );


  or
  g709
  (
    n720,
    n552,
    n554,
    n544,
    n529
  );


  buf
  g710
  (
    n729,
    n713
  );


  not
  g711
  (
    KeyWire_0_13,
    n712
  );


  nor
  g712
  (
    n731,
    n655,
    n653,
    n730,
    n654
  );


  or
  g713
  (
    n733,
    n717,
    n731,
    n724,
    n715
  );


  nand
  g714
  (
    n734,
    n716,
    n731,
    n722,
    n723
  );


  nand
  g715
  (
    n735,
    n721,
    n718,
    n720,
    n725
  );


  nand
  g716
  (
    n732,
    n719,
    n731,
    n714
  );


  xor
  g717
  (
    n739,
    n656,
    n661,
    n672,
    n735
  );


  nand
  g718
  (
    n738,
    n671,
    n660,
    n735,
    n679
  );


  xnor
  g719
  (
    n742,
    n678,
    n664,
    n734,
    n662
  );


  xor
  g720
  (
    n740,
    n673,
    n733,
    n735
  );


  or
  g721
  (
    n736,
    n657,
    n663,
    n676,
    n675
  );


  xnor
  g722
  (
    n743,
    n734,
    n668,
    n670,
    n677
  );


  and
  g723
  (
    n741,
    n667,
    n658,
    n732,
    n674
  );


  nand
  g724
  (
    n737,
    n659,
    n665,
    n669,
    n666
  );


  nand
  g725
  (
    n745,
    n688,
    n738,
    n685,
    n681
  );


  or
  g726
  (
    n744,
    n739,
    n691,
    n682,
    n683
  );


  nor
  g727
  (
    n747,
    n689,
    n687,
    n680,
    n737
  );


  nor
  g728
  (
    n746,
    n686,
    n690,
    n684,
    n736
  );


  xnor
  g729
  (
    n751,
    n276,
    n727,
    n746,
    n747
  );


  and
  g730
  (
    n748,
    n276,
    n277,
    n728,
    n740
  );


  nand
  g731
  (
    n749,
    n277,
    n276,
    n202
  );


  nor
  g732
  (
    KeyWire_0_14,
    n744,
    n202,
    n277,
    n747
  );


  and
  g733
  (
    n750,
    n726,
    n745,
    n277,
    n202
  );


  nand
  g734
  (
    n753,
    n752,
    n750,
    n742,
    n751
  );


  nor
  g735
  (
    n754,
    n743,
    n741,
    n749,
    n748
  );


  xor
  KeyGate_0_0
  (
    n452,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n145,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n231,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n432,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n699,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n532,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n337,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n200,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n165,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n687,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n271,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n519,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n340,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n730,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n752,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n610,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule

