

module Stat_2916_29_2
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n2802,
  n2805,
  n2799,
  n2816,
  n2800,
  n2810,
  n2796,
  n2811,
  n2814,
  n2794,
  n2815,
  n2797,
  n2817,
  n2801,
  n2798,
  n2793,
  n2806,
  n2808,
  n2818,
  n2809,
  n2804,
  n2803,
  n2807,
  n2812,
  n2820,
  n2822,
  n2821,
  n2826,
  n2825,
  n2849,
  n2850,
  n2851,
  n2852,
  n2854,
  n2848,
  n2853,
  n2914,
  n2943,
  n2939,
  n2944,
  n2945,
  n2942,
  n2941,
  n2936,
  n2946,
  n2938,
  n2937,
  n2940,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;
  output n2802;output n2805;output n2799;output n2816;output n2800;output n2810;output n2796;output n2811;output n2814;output n2794;output n2815;output n2797;output n2817;output n2801;output n2798;output n2793;output n2806;output n2808;output n2818;output n2809;output n2804;output n2803;output n2807;output n2812;output n2820;output n2822;output n2821;output n2826;output n2825;output n2849;output n2850;output n2851;output n2852;output n2854;output n2848;output n2853;output n2914;output n2943;output n2939;output n2944;output n2945;output n2942;output n2941;output n2936;output n2946;output n2938;output n2937;output n2940;
  wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2795;wire n2813;wire n2819;wire n2823;wire n2824;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n31,
    n5
  );


  buf
  g1
  (
    n76,
    n12
  );


  buf
  g2
  (
    n68,
    n16
  );


  buf
  g3
  (
    n33,
    n19
  );


  buf
  g4
  (
    n105,
    n20
  );


  buf
  g5
  (
    n113,
    n9
  );


  buf
  g6
  (
    n67,
    n15
  );


  not
  g7
  (
    n89,
    n7
  );


  buf
  g8
  (
    n83,
    n1
  );


  buf
  g9
  (
    n102,
    n5
  );


  buf
  g10
  (
    n36,
    n12
  );


  not
  g11
  (
    n84,
    n4
  );


  buf
  g12
  (
    n35,
    n12
  );


  buf
  g13
  (
    n79,
    n18
  );


  not
  g14
  (
    n52,
    n25
  );


  buf
  g15
  (
    n112,
    n9
  );


  not
  g16
  (
    n122,
    n11
  );


  buf
  g17
  (
    n42,
    n1
  );


  not
  g18
  (
    n37,
    n18
  );


  not
  g19
  (
    n63,
    n13
  );


  buf
  g20
  (
    n51,
    n3
  );


  not
  g21
  (
    n41,
    n21
  );


  not
  g22
  (
    n45,
    n15
  );


  not
  g23
  (
    n88,
    n7
  );


  buf
  g24
  (
    n98,
    n12
  );


  buf
  g25
  (
    n53,
    n23
  );


  buf
  g26
  (
    n49,
    n9
  );


  buf
  g27
  (
    n32,
    n13
  );


  buf
  g28
  (
    n97,
    n14
  );


  buf
  g29
  (
    n104,
    n14
  );


  buf
  g30
  (
    n66,
    n21
  );


  buf
  g31
  (
    n71,
    n6
  );


  not
  g32
  (
    n62,
    n4
  );


  not
  g33
  (
    n50,
    n24
  );


  buf
  g34
  (
    n77,
    n13
  );


  not
  g35
  (
    n110,
    n19
  );


  buf
  g36
  (
    n100,
    n7
  );


  not
  g37
  (
    n108,
    n24
  );


  not
  g38
  (
    n61,
    n23
  );


  buf
  g39
  (
    n120,
    n10
  );


  not
  g40
  (
    n46,
    n22
  );


  not
  g41
  (
    n44,
    n14
  );


  not
  g42
  (
    n109,
    n1
  );


  buf
  g43
  (
    n54,
    n17
  );


  not
  g44
  (
    n57,
    n15
  );


  not
  g45
  (
    n118,
    n10
  );


  buf
  g46
  (
    n91,
    n25
  );


  buf
  g47
  (
    n124,
    n4
  );


  not
  g48
  (
    n72,
    n3
  );


  not
  g49
  (
    n60,
    n17
  );


  buf
  g50
  (
    n48,
    n17
  );


  buf
  g51
  (
    n75,
    n16
  );


  buf
  g52
  (
    n127,
    n22
  );


  not
  g53
  (
    n55,
    n19
  );


  not
  g54
  (
    n43,
    n24
  );


  not
  g55
  (
    n81,
    n9
  );


  buf
  g56
  (
    n34,
    n24
  );


  not
  g57
  (
    n74,
    n20
  );


  buf
  g58
  (
    n80,
    n20
  );


  buf
  g59
  (
    n90,
    n11
  );


  not
  g60
  (
    n82,
    n1
  );


  not
  g61
  (
    n65,
    n21
  );


  not
  g62
  (
    n121,
    n5
  );


  buf
  g63
  (
    n115,
    n15
  );


  buf
  g64
  (
    n101,
    n16
  );


  not
  g65
  (
    n128,
    n2
  );


  not
  g66
  (
    n116,
    n2
  );


  buf
  g67
  (
    n40,
    n23
  );


  buf
  g68
  (
    n93,
    n20
  );


  buf
  g69
  (
    n117,
    n11
  );


  buf
  g70
  (
    n38,
    n21
  );


  not
  g71
  (
    n125,
    n5
  );


  buf
  g72
  (
    n70,
    n2
  );


  buf
  g73
  (
    n114,
    n22
  );


  buf
  g74
  (
    n99,
    n17
  );


  not
  g75
  (
    n96,
    n13
  );


  buf
  g76
  (
    n69,
    n6
  );


  not
  g77
  (
    n56,
    n4
  );


  not
  g78
  (
    n73,
    n3
  );


  buf
  g79
  (
    n106,
    n7
  );


  buf
  g80
  (
    n103,
    n18
  );


  buf
  g81
  (
    n126,
    n10
  );


  buf
  g82
  (
    n94,
    n2
  );


  buf
  g83
  (
    n78,
    n6
  );


  buf
  g84
  (
    n95,
    n10
  );


  not
  g85
  (
    n92,
    n8
  );


  buf
  g86
  (
    n111,
    n3
  );


  buf
  g87
  (
    n85,
    n11
  );


  not
  g88
  (
    n107,
    n19
  );


  buf
  g89
  (
    n86,
    n14
  );


  buf
  g90
  (
    n64,
    n8
  );


  not
  g91
  (
    n58,
    n8
  );


  not
  g92
  (
    n47,
    n6
  );


  not
  g93
  (
    n87,
    n8
  );


  buf
  g94
  (
    n59,
    n18
  );


  buf
  g95
  (
    n39,
    n22
  );


  buf
  g96
  (
    n123,
    n16
  );


  buf
  g97
  (
    n119,
    n23
  );


  buf
  g98
  (
    n304,
    n41
  );


  not
  g99
  (
    n414,
    n86
  );


  not
  g100
  (
    n212,
    n34
  );


  buf
  g101
  (
    n276,
    n96
  );


  buf
  g102
  (
    n146,
    n80
  );


  not
  g103
  (
    n292,
    n83
  );


  not
  g104
  (
    n373,
    n110
  );


  buf
  g105
  (
    n162,
    n49
  );


  buf
  g106
  (
    n176,
    n107
  );


  not
  g107
  (
    n231,
    n41
  );


  buf
  g108
  (
    n403,
    n59
  );


  buf
  g109
  (
    n199,
    n65
  );


  buf
  g110
  (
    n299,
    n102
  );


  buf
  g111
  (
    n213,
    n53
  );


  not
  g112
  (
    n468,
    n107
  );


  not
  g113
  (
    n413,
    n36
  );


  not
  g114
  (
    n281,
    n32
  );


  not
  g115
  (
    n138,
    n78
  );


  buf
  g116
  (
    n238,
    n71
  );


  buf
  g117
  (
    n228,
    n81
  );


  not
  g118
  (
    n283,
    n37
  );


  buf
  g119
  (
    n423,
    n46
  );


  buf
  g120
  (
    n322,
    n89
  );


  buf
  g121
  (
    n369,
    n85
  );


  not
  g122
  (
    n394,
    n69
  );


  buf
  g123
  (
    n151,
    n83
  );


  buf
  g124
  (
    n298,
    n82
  );


  buf
  g125
  (
    n421,
    n80
  );


  not
  g126
  (
    n415,
    n99
  );


  not
  g127
  (
    n189,
    n32
  );


  not
  g128
  (
    n132,
    n97
  );


  buf
  g129
  (
    n380,
    n62
  );


  buf
  g130
  (
    n224,
    n36
  );


  buf
  g131
  (
    n181,
    n63
  );


  buf
  g132
  (
    n220,
    n104
  );


  not
  g133
  (
    n156,
    n54
  );


  buf
  g134
  (
    n437,
    n81
  );


  not
  g135
  (
    n412,
    n51
  );


  not
  g136
  (
    n195,
    n57
  );


  buf
  g137
  (
    n260,
    n58
  );


  buf
  g138
  (
    n161,
    n79
  );


  buf
  g139
  (
    n432,
    n89
  );


  not
  g140
  (
    n426,
    n104
  );


  buf
  g141
  (
    n411,
    n94
  );


  not
  g142
  (
    n257,
    n72
  );


  buf
  g143
  (
    n433,
    n35
  );


  not
  g144
  (
    n417,
    n66
  );


  not
  g145
  (
    n191,
    n111
  );


  buf
  g146
  (
    n297,
    n49
  );


  buf
  g147
  (
    n172,
    n77
  );


  not
  g148
  (
    n274,
    n40
  );


  not
  g149
  (
    n234,
    n72
  );


  buf
  g150
  (
    n321,
    n115
  );


  buf
  g151
  (
    n319,
    n86
  );


  buf
  g152
  (
    n177,
    n62
  );


  buf
  g153
  (
    n392,
    n44
  );


  not
  g154
  (
    n353,
    n110
  );


  buf
  g155
  (
    n150,
    n56
  );


  not
  g156
  (
    n210,
    n42
  );


  buf
  g157
  (
    n402,
    n108
  );


  not
  g158
  (
    n337,
    n106
  );


  buf
  g159
  (
    n160,
    n87
  );


  not
  g160
  (
    n266,
    n107
  );


  buf
  g161
  (
    n280,
    n52
  );


  buf
  g162
  (
    n350,
    n55
  );


  buf
  g163
  (
    n331,
    n37
  );


  buf
  g164
  (
    n452,
    n104
  );


  buf
  g165
  (
    n342,
    n88
  );


  not
  g166
  (
    n371,
    n58
  );


  buf
  g167
  (
    n334,
    n97
  );


  not
  g168
  (
    n448,
    n34
  );


  buf
  g169
  (
    n435,
    n95
  );


  not
  g170
  (
    n378,
    n71
  );


  buf
  g171
  (
    n209,
    n72
  );


  not
  g172
  (
    n307,
    n106
  );


  buf
  g173
  (
    n262,
    n114
  );


  buf
  g174
  (
    n460,
    n102
  );


  buf
  g175
  (
    n236,
    n45
  );


  not
  g176
  (
    n301,
    n43
  );


  not
  g177
  (
    n186,
    n74
  );


  buf
  g178
  (
    n436,
    n78
  );


  not
  g179
  (
    n393,
    n74
  );


  buf
  g180
  (
    n259,
    n47
  );


  not
  g181
  (
    n287,
    n50
  );


  buf
  g182
  (
    n453,
    n108
  );


  not
  g183
  (
    n290,
    n55
  );


  buf
  g184
  (
    n286,
    n38
  );


  not
  g185
  (
    n279,
    n79
  );


  not
  g186
  (
    n187,
    n33
  );


  not
  g187
  (
    n370,
    n104
  );


  buf
  g188
  (
    n400,
    n51
  );


  not
  g189
  (
    n357,
    n53
  );


  buf
  g190
  (
    n250,
    n66
  );


  buf
  g191
  (
    n193,
    n63
  );


  not
  g192
  (
    n142,
    n51
  );


  not
  g193
  (
    n316,
    n35
  );


  not
  g194
  (
    n246,
    n57
  );


  not
  g195
  (
    n243,
    n44
  );


  not
  g196
  (
    n149,
    n109
  );


  not
  g197
  (
    n340,
    n36
  );


  buf
  g198
  (
    n382,
    n112
  );


  not
  g199
  (
    n227,
    n39
  );


  buf
  g200
  (
    n196,
    n39
  );


  buf
  g201
  (
    n406,
    n83
  );


  not
  g202
  (
    n404,
    n76
  );


  not
  g203
  (
    n291,
    n102
  );


  buf
  g204
  (
    n133,
    n48
  );


  buf
  g205
  (
    n444,
    n101
  );


  not
  g206
  (
    n140,
    n37
  );


  buf
  g207
  (
    n129,
    n71
  );


  buf
  g208
  (
    n467,
    n113
  );


  buf
  g209
  (
    n205,
    n86
  );


  not
  g210
  (
    n339,
    n57
  );


  not
  g211
  (
    n441,
    n114
  );


  not
  g212
  (
    n325,
    n98
  );


  not
  g213
  (
    n416,
    n75
  );


  not
  g214
  (
    n200,
    n101
  );


  buf
  g215
  (
    n459,
    n56
  );


  buf
  g216
  (
    n364,
    n46
  );


  buf
  g217
  (
    n390,
    n60
  );


  buf
  g218
  (
    n247,
    n82
  );


  buf
  g219
  (
    n285,
    n48
  );


  not
  g220
  (
    n447,
    n69
  );


  not
  g221
  (
    n363,
    n77
  );


  not
  g222
  (
    n130,
    n86
  );


  not
  g223
  (
    n208,
    n35
  );


  buf
  g224
  (
    n389,
    n45
  );


  buf
  g225
  (
    n253,
    n103
  );


  not
  g226
  (
    n248,
    n48
  );


  buf
  g227
  (
    n320,
    n105
  );


  not
  g228
  (
    n451,
    n38
  );


  not
  g229
  (
    n282,
    n109
  );


  buf
  g230
  (
    n273,
    n63
  );


  not
  g231
  (
    n343,
    n60
  );


  buf
  g232
  (
    n445,
    n67
  );


  buf
  g233
  (
    n410,
    n91
  );


  not
  g234
  (
    n134,
    n115
  );


  buf
  g235
  (
    n314,
    n93
  );


  not
  g236
  (
    n173,
    n67
  );


  buf
  g237
  (
    n249,
    n77
  );


  not
  g238
  (
    n336,
    n95
  );


  buf
  g239
  (
    n230,
    n111
  );


  not
  g240
  (
    n137,
    n58
  );


  buf
  g241
  (
    n143,
    n76
  );


  buf
  g242
  (
    n296,
    n92
  );


  not
  g243
  (
    n333,
    n64
  );


  buf
  g244
  (
    n135,
    n101
  );


  not
  g245
  (
    n399,
    n44
  );


  buf
  g246
  (
    n308,
    n50
  );


  buf
  g247
  (
    n409,
    n37
  );


  buf
  g248
  (
    n275,
    n42
  );


  not
  g249
  (
    n207,
    n31
  );


  buf
  g250
  (
    n241,
    n59
  );


  buf
  g251
  (
    n198,
    n69
  );


  buf
  g252
  (
    n192,
    n68
  );


  buf
  g253
  (
    n365,
    n89
  );


  buf
  g254
  (
    n157,
    n110
  );


  not
  g255
  (
    n217,
    n65
  );


  not
  g256
  (
    n235,
    n93
  );


  buf
  g257
  (
    n376,
    n40
  );


  not
  g258
  (
    n313,
    n55
  );


  not
  g259
  (
    n255,
    n84
  );


  not
  g260
  (
    n405,
    n31
  );


  buf
  g261
  (
    n152,
    n40
  );


  not
  g262
  (
    n461,
    n50
  );


  not
  g263
  (
    n202,
    n61
  );


  not
  g264
  (
    n449,
    n56
  );


  buf
  g265
  (
    n377,
    n33
  );


  not
  g266
  (
    n396,
    n61
  );


  buf
  g267
  (
    n182,
    n92
  );


  not
  g268
  (
    n375,
    n114
  );


  buf
  g269
  (
    n465,
    n64
  );


  not
  g270
  (
    n215,
    n103
  );


  not
  g271
  (
    n163,
    n85
  );


  not
  g272
  (
    n167,
    n95
  );


  not
  g273
  (
    n427,
    n88
  );


  buf
  g274
  (
    n263,
    n47
  );


  buf
  g275
  (
    n456,
    n101
  );


  buf
  g276
  (
    n216,
    n65
  );


  buf
  g277
  (
    n359,
    n73
  );


  not
  g278
  (
    n261,
    n42
  );


  not
  g279
  (
    n211,
    n57
  );


  buf
  g280
  (
    n315,
    n67
  );


  not
  g281
  (
    n131,
    n39
  );


  not
  g282
  (
    n317,
    n106
  );


  not
  g283
  (
    n289,
    n61
  );


  not
  g284
  (
    n366,
    n66
  );


  not
  g285
  (
    n148,
    n108
  );


  buf
  g286
  (
    n218,
    n113
  );


  buf
  g287
  (
    n225,
    n64
  );


  not
  g288
  (
    n425,
    n43
  );


  not
  g289
  (
    n344,
    n64
  );


  not
  g290
  (
    n221,
    n91
  );


  buf
  g291
  (
    n244,
    n39
  );


  buf
  g292
  (
    n312,
    n67
  );


  not
  g293
  (
    n306,
    n92
  );


  not
  g294
  (
    n190,
    n88
  );


  not
  g295
  (
    n240,
    n58
  );


  not
  g296
  (
    n352,
    n93
  );


  not
  g297
  (
    n345,
    n66
  );


  not
  g298
  (
    n430,
    n115
  );


  not
  g299
  (
    n226,
    n90
  );


  not
  g300
  (
    n391,
    n45
  );


  buf
  g301
  (
    n395,
    n55
  );


  not
  g302
  (
    n332,
    n100
  );


  not
  g303
  (
    n251,
    n94
  );


  not
  g304
  (
    n164,
    n54
  );


  buf
  g305
  (
    n464,
    n92
  );


  not
  g306
  (
    n168,
    n38
  );


  not
  g307
  (
    n328,
    n79
  );


  buf
  g308
  (
    n442,
    n111
  );


  not
  g309
  (
    n374,
    n91
  );


  not
  g310
  (
    n158,
    n105
  );


  buf
  g311
  (
    n431,
    n61
  );


  not
  g312
  (
    n326,
    n68
  );


  buf
  g313
  (
    n397,
    n47
  );


  buf
  g314
  (
    n136,
    n103
  );


  buf
  g315
  (
    n258,
    n106
  );


  not
  g316
  (
    n381,
    n105
  );


  buf
  g317
  (
    n311,
    n100
  );


  buf
  g318
  (
    n141,
    n112
  );


  not
  g319
  (
    n457,
    n42
  );


  not
  g320
  (
    n154,
    n81
  );


  not
  g321
  (
    n302,
    n98
  );


  buf
  g322
  (
    n153,
    n33
  );


  buf
  g323
  (
    n348,
    n36
  );


  not
  g324
  (
    n300,
    n33
  );


  not
  g325
  (
    n324,
    n84
  );


  buf
  g326
  (
    n358,
    n59
  );


  not
  g327
  (
    n145,
    n43
  );


  buf
  g328
  (
    n418,
    n90
  );


  buf
  g329
  (
    n194,
    n40
  );


  buf
  g330
  (
    n310,
    n73
  );


  not
  g331
  (
    n166,
    n34
  );


  not
  g332
  (
    n455,
    n113
  );


  buf
  g333
  (
    n183,
    n84
  );


  buf
  g334
  (
    n450,
    n112
  );


  buf
  g335
  (
    n165,
    n56
  );


  buf
  g336
  (
    n434,
    n49
  );


  not
  g337
  (
    n269,
    n91
  );


  not
  g338
  (
    n303,
    n53
  );


  buf
  g339
  (
    n171,
    n109
  );


  not
  g340
  (
    n367,
    n110
  );


  not
  g341
  (
    n178,
    n87
  );


  buf
  g342
  (
    n385,
    n114
  );


  not
  g343
  (
    n139,
    n78
  );


  buf
  g344
  (
    n159,
    n103
  );


  buf
  g345
  (
    n346,
    n79
  );


  buf
  g346
  (
    n422,
    n34
  );


  not
  g347
  (
    n245,
    n54
  );


  buf
  g348
  (
    n169,
    n68
  );


  not
  g349
  (
    n454,
    n84
  );


  not
  g350
  (
    n271,
    n98
  );


  buf
  g351
  (
    n268,
    n35
  );


  not
  g352
  (
    n278,
    n77
  );


  buf
  g353
  (
    n419,
    n93
  );


  not
  g354
  (
    n323,
    n99
  );


  not
  g355
  (
    n458,
    n75
  );


  not
  g356
  (
    n188,
    n85
  );


  not
  g357
  (
    n284,
    n89
  );


  buf
  g358
  (
    n293,
    n95
  );


  buf
  g359
  (
    n204,
    n102
  );


  buf
  g360
  (
    n439,
    n69
  );


  not
  g361
  (
    n233,
    n70
  );


  buf
  g362
  (
    n408,
    n98
  );


  not
  g363
  (
    n318,
    n32
  );


  buf
  g364
  (
    n254,
    n52
  );


  not
  g365
  (
    n175,
    n74
  );


  not
  g366
  (
    n428,
    n87
  );


  buf
  g367
  (
    n256,
    n70
  );


  buf
  g368
  (
    n179,
    n80
  );


  not
  g369
  (
    n351,
    n78
  );


  buf
  g370
  (
    n362,
    n50
  );


  not
  g371
  (
    n294,
    n38
  );


  buf
  g372
  (
    n252,
    n73
  );


  buf
  g373
  (
    n264,
    n44
  );


  not
  g374
  (
    n368,
    n76
  );


  buf
  g375
  (
    n354,
    n52
  );


  not
  g376
  (
    n401,
    n115
  );


  buf
  g377
  (
    n360,
    n82
  );


  not
  g378
  (
    n466,
    n90
  );


  buf
  g379
  (
    n420,
    n97
  );


  buf
  g380
  (
    n407,
    n88
  );


  buf
  g381
  (
    n277,
    n63
  );


  buf
  g382
  (
    n438,
    n112
  );


  not
  g383
  (
    n327,
    n43
  );


  not
  g384
  (
    n185,
    n80
  );


  not
  g385
  (
    n361,
    n65
  );


  buf
  g386
  (
    n201,
    n113
  );


  not
  g387
  (
    n372,
    n52
  );


  buf
  g388
  (
    n388,
    n59
  );


  not
  g389
  (
    n265,
    n75
  );


  buf
  g390
  (
    n356,
    n82
  );


  not
  g391
  (
    n272,
    n90
  );


  not
  g392
  (
    n446,
    n96
  );


  not
  g393
  (
    n329,
    n96
  );


  buf
  g394
  (
    n347,
    n85
  );


  not
  g395
  (
    n229,
    n51
  );


  buf
  g396
  (
    n232,
    n94
  );


  buf
  g397
  (
    n239,
    n62
  );


  not
  g398
  (
    n270,
    n71
  );


  buf
  g399
  (
    n144,
    n94
  );


  buf
  g400
  (
    n309,
    n111
  );


  not
  g401
  (
    n398,
    n81
  );


  not
  g402
  (
    n267,
    n46
  );


  buf
  g403
  (
    n440,
    n99
  );


  not
  g404
  (
    n288,
    n47
  );


  buf
  g405
  (
    n443,
    n74
  );


  buf
  g406
  (
    n330,
    n83
  );


  not
  g407
  (
    n147,
    n41
  );


  buf
  g408
  (
    n384,
    n60
  );


  buf
  g409
  (
    n184,
    n72
  );


  not
  g410
  (
    n237,
    n109
  );


  not
  g411
  (
    n429,
    n31
  );


  not
  g412
  (
    n462,
    n107
  );


  buf
  g413
  (
    n222,
    n60
  );


  buf
  g414
  (
    n305,
    n32
  );


  buf
  g415
  (
    n386,
    n105
  );


  buf
  g416
  (
    n335,
    n62
  );


  not
  g417
  (
    n155,
    n46
  );


  not
  g418
  (
    n383,
    n73
  );


  not
  g419
  (
    n424,
    n31
  );


  buf
  g420
  (
    n341,
    n99
  );


  not
  g421
  (
    n197,
    n70
  );


  buf
  g422
  (
    n174,
    n97
  );


  buf
  g423
  (
    n463,
    n100
  );


  buf
  g424
  (
    n387,
    n45
  );


  buf
  g425
  (
    n219,
    n53
  );


  buf
  g426
  (
    n338,
    n68
  );


  not
  g427
  (
    n214,
    n96
  );


  not
  g428
  (
    n206,
    n75
  );


  buf
  g429
  (
    n223,
    n108
  );


  buf
  g430
  (
    n170,
    n70
  );


  buf
  g431
  (
    n379,
    n100
  );


  not
  g432
  (
    n242,
    n48
  );


  buf
  g433
  (
    n295,
    n76
  );


  buf
  g434
  (
    n180,
    n87
  );


  buf
  g435
  (
    n349,
    n49
  );


  buf
  g436
  (
    n355,
    n54
  );


  not
  g437
  (
    n203,
    n41
  );


  buf
  g438
  (
    n963,
    n454
  );


  buf
  g439
  (
    n1149,
    n275
  );


  not
  g440
  (
    n592,
    n210
  );


  buf
  g441
  (
    n791,
    n277
  );


  not
  g442
  (
    n1548,
    n138
  );


  not
  g443
  (
    n1670,
    n443
  );


  buf
  g444
  (
    n821,
    n415
  );


  not
  g445
  (
    n997,
    n407
  );


  not
  g446
  (
    n1355,
    n162
  );


  buf
  g447
  (
    n1439,
    n355
  );


  not
  g448
  (
    n1265,
    n207
  );


  not
  g449
  (
    n1567,
    n305
  );


  buf
  g450
  (
    n902,
    n345
  );


  buf
  g451
  (
    n1672,
    n150
  );


  not
  g452
  (
    n1135,
    n372
  );


  not
  g453
  (
    n813,
    n185
  );


  not
  g454
  (
    n629,
    n330
  );


  not
  g455
  (
    n1660,
    n255
  );


  buf
  g456
  (
    n1302,
    n414
  );


  buf
  g457
  (
    n1239,
    n442
  );


  not
  g458
  (
    n1631,
    n453
  );


  buf
  g459
  (
    n1738,
    n427
  );


  not
  g460
  (
    n612,
    n309
  );


  not
  g461
  (
    n870,
    n330
  );


  not
  g462
  (
    n556,
    n391
  );


  not
  g463
  (
    n599,
    n231
  );


  buf
  g464
  (
    n1572,
    n457
  );


  buf
  g465
  (
    n1075,
    n391
  );


  buf
  g466
  (
    n1577,
    n233
  );


  buf
  g467
  (
    n721,
    n283
  );


  buf
  g468
  (
    n898,
    n215
  );


  not
  g469
  (
    n936,
    n288
  );


  not
  g470
  (
    n640,
    n308
  );


  buf
  g471
  (
    n1196,
    n273
  );


  buf
  g472
  (
    n1167,
    n397
  );


  not
  g473
  (
    n1399,
    n397
  );


  not
  g474
  (
    n1383,
    n173
  );


  buf
  g475
  (
    n535,
    n394
  );


  buf
  g476
  (
    n1369,
    n181
  );


  buf
  g477
  (
    n486,
    n149
  );


  not
  g478
  (
    n1676,
    n172
  );


  not
  g479
  (
    n1626,
    n134
  );


  not
  g480
  (
    n733,
    n418
  );


  buf
  g481
  (
    n1415,
    n259
  );


  buf
  g482
  (
    n1730,
    n368
  );


  buf
  g483
  (
    n1744,
    n357
  );


  not
  g484
  (
    n708,
    n280
  );


  not
  g485
  (
    n1463,
    n447
  );


  buf
  g486
  (
    n940,
    n293
  );


  buf
  g487
  (
    n690,
    n392
  );


  buf
  g488
  (
    n1291,
    n129
  );


  buf
  g489
  (
    n675,
    n381
  );


  not
  g490
  (
    n653,
    n377
  );


  not
  g491
  (
    n1034,
    n407
  );


  not
  g492
  (
    n1137,
    n403
  );


  buf
  g493
  (
    n469,
    n242
  );


  not
  g494
  (
    n1320,
    n146
  );


  not
  g495
  (
    n1185,
    n223
  );


  not
  g496
  (
    n603,
    n168
  );


  buf
  g497
  (
    n927,
    n422
  );


  not
  g498
  (
    n687,
    n379
  );


  not
  g499
  (
    n879,
    n414
  );


  not
  g500
  (
    n1124,
    n370
  );


  buf
  g501
  (
    n738,
    n180
  );


  buf
  g502
  (
    n1554,
    n392
  );


  buf
  g503
  (
    n1059,
    n209
  );


  not
  g504
  (
    n515,
    n328
  );


  buf
  g505
  (
    n673,
    n401
  );


  not
  g506
  (
    n1243,
    n278
  );


  not
  g507
  (
    n667,
    n159
  );


  buf
  g508
  (
    n845,
    n430
  );


  buf
  g509
  (
    n1125,
    n133
  );


  not
  g510
  (
    n1552,
    n316
  );


  not
  g511
  (
    n1371,
    n254
  );


  buf
  g512
  (
    n606,
    n226
  );


  not
  g513
  (
    n1594,
    n283
  );


  buf
  g514
  (
    n814,
    n445
  );


  buf
  g515
  (
    n1664,
    n224
  );


  buf
  g516
  (
    n1236,
    n138
  );


  buf
  g517
  (
    n490,
    n274
  );


  buf
  g518
  (
    n881,
    n436
  );


  not
  g519
  (
    n684,
    n257
  );


  not
  g520
  (
    n1639,
    n244
  );


  buf
  g521
  (
    n555,
    n148
  );


  not
  g522
  (
    n974,
    n221
  );


  not
  g523
  (
    n1413,
    n197
  );


  not
  g524
  (
    n771,
    n423
  );


  not
  g525
  (
    n529,
    n358
  );


  not
  g526
  (
    n1301,
    n181
  );


  buf
  g527
  (
    n1556,
    n440
  );


  not
  g528
  (
    n1347,
    n267
  );


  buf
  g529
  (
    n532,
    n180
  );


  buf
  g530
  (
    n1665,
    n199
  );


  not
  g531
  (
    n1433,
    n269
  );


  not
  g532
  (
    n1614,
    n325
  );


  not
  g533
  (
    n750,
    n446
  );


  buf
  g534
  (
    n985,
    n271
  );


  buf
  g535
  (
    n596,
    n431
  );


  buf
  g536
  (
    n1218,
    n323
  );


  not
  g537
  (
    n875,
    n269
  );


  buf
  g538
  (
    n1314,
    n285
  );


  buf
  g539
  (
    n948,
    n424
  );


  not
  g540
  (
    n1398,
    n387
  );


  buf
  g541
  (
    n1742,
    n261
  );


  not
  g542
  (
    n1328,
    n450
  );


  not
  g543
  (
    n649,
    n333
  );


  not
  g544
  (
    n1654,
    n266
  );


  not
  g545
  (
    n1526,
    n404
  );


  not
  g546
  (
    n1411,
    n160
  );


  not
  g547
  (
    n1465,
    n282
  );


  not
  g548
  (
    n1254,
    n327
  );


  not
  g549
  (
    n1106,
    n307
  );


  buf
  g550
  (
    n1166,
    n393
  );


  not
  g551
  (
    n626,
    n292
  );


  not
  g552
  (
    n892,
    n377
  );


  not
  g553
  (
    n1242,
    n245
  );


  not
  g554
  (
    n672,
    n150
  );


  buf
  g555
  (
    n1268,
    n136
  );


  buf
  g556
  (
    n1017,
    n310
  );


  buf
  g557
  (
    n832,
    n171
  );


  buf
  g558
  (
    n1388,
    n230
  );


  not
  g559
  (
    n582,
    n340
  );


  not
  g560
  (
    n1560,
    n326
  );


  buf
  g561
  (
    n1653,
    n155
  );


  buf
  g562
  (
    n836,
    n405
  );


  buf
  g563
  (
    n1157,
    n401
  );


  not
  g564
  (
    n1686,
    n378
  );


  not
  g565
  (
    n1066,
    n175
  );


  not
  g566
  (
    n1495,
    n313
  );


  buf
  g567
  (
    n1512,
    n215
  );


  not
  g568
  (
    n843,
    n269
  );


  not
  g569
  (
    n876,
    n291
  );


  not
  g570
  (
    n573,
    n188
  );


  buf
  g571
  (
    n1354,
    n221
  );


  buf
  g572
  (
    n664,
    n443
  );


  not
  g573
  (
    n803,
    n217
  );


  buf
  g574
  (
    n546,
    n452
  );


  buf
  g575
  (
    n1055,
    n277
  );


  not
  g576
  (
    n1698,
    n417
  );


  buf
  g577
  (
    n1531,
    n402
  );


  not
  g578
  (
    n1104,
    n242
  );


  buf
  g579
  (
    n1726,
    n158
  );


  not
  g580
  (
    n481,
    n388
  );


  not
  g581
  (
    n557,
    n456
  );


  not
  g582
  (
    n671,
    n327
  );


  buf
  g583
  (
    n1128,
    n359
  );


  not
  g584
  (
    n1276,
    n179
  );


  not
  g585
  (
    n1256,
    n400
  );


  not
  g586
  (
    n1522,
    n240
  );


  buf
  g587
  (
    n888,
    n239
  );


  not
  g588
  (
    n1561,
    n172
  );


  buf
  g589
  (
    n1624,
    n406
  );


  buf
  g590
  (
    n987,
    n403
  );


  buf
  g591
  (
    n1083,
    n253
  );


  not
  g592
  (
    n1656,
    n227
  );


  buf
  g593
  (
    n1538,
    n188
  );


  buf
  g594
  (
    n809,
    n363
  );


  buf
  g595
  (
    n1629,
    n281
  );


  buf
  g596
  (
    n1138,
    n266
  );


  buf
  g597
  (
    n1337,
    n192
  );


  not
  g598
  (
    n907,
    n142
  );


  buf
  g599
  (
    n1400,
    n148
  );


  not
  g600
  (
    n967,
    n147
  );


  not
  g601
  (
    n1005,
    n278
  );


  buf
  g602
  (
    n470,
    n367
  );


  buf
  g603
  (
    n1012,
    n419
  );


  not
  g604
  (
    n552,
    n430
  );


  not
  g605
  (
    n1559,
    n455
  );


  not
  g606
  (
    n758,
    n388
  );


  not
  g607
  (
    n1309,
    n385
  );


  buf
  g608
  (
    n729,
    n327
  );


  not
  g609
  (
    n1693,
    n429
  );


  not
  g610
  (
    n790,
    n217
  );


  not
  g611
  (
    n1036,
    n168
  );


  not
  g612
  (
    n1273,
    n240
  );


  not
  g613
  (
    n577,
    n413
  );


  not
  g614
  (
    n1246,
    n417
  );


  buf
  g615
  (
    n1035,
    n184
  );


  buf
  g616
  (
    n954,
    n386
  );


  not
  g617
  (
    n1436,
    n203
  );


  not
  g618
  (
    n884,
    n233
  );


  not
  g619
  (
    n1651,
    n202
  );


  not
  g620
  (
    n585,
    n254
  );


  buf
  g621
  (
    n1638,
    n391
  );


  not
  g622
  (
    n937,
    n298
  );


  not
  g623
  (
    n1148,
    n338
  );


  not
  g624
  (
    n1504,
    n307
  );


  buf
  g625
  (
    n1487,
    n326
  );


  buf
  g626
  (
    n1683,
    n289
  );


  buf
  g627
  (
    n1192,
    n325
  );


  buf
  g628
  (
    n1620,
    n185
  );


  buf
  g629
  (
    n1011,
    n438
  );


  buf
  g630
  (
    n1304,
    n295
  );


  not
  g631
  (
    n982,
    n334
  );


  buf
  g632
  (
    n678,
    n244
  );


  not
  g633
  (
    n613,
    n195
  );


  not
  g634
  (
    n639,
    n364
  );


  buf
  g635
  (
    n831,
    n434
  );


  buf
  g636
  (
    n1645,
    n231
  );


  not
  g637
  (
    n784,
    n286
  );


  buf
  g638
  (
    n1222,
    n429
  );


  buf
  g639
  (
    n568,
    n425
  );


  buf
  g640
  (
    n1249,
    n145
  );


  not
  g641
  (
    n1384,
    n448
  );


  buf
  g642
  (
    n1370,
    n392
  );


  buf
  g643
  (
    n901,
    n408
  );


  not
  g644
  (
    n1311,
    n189
  );


  not
  g645
  (
    n1679,
    n306
  );


  not
  g646
  (
    n736,
    n327
  );


  buf
  g647
  (
    n1003,
    n442
  );


  not
  g648
  (
    n1119,
    n273
  );


  not
  g649
  (
    n610,
    n351
  );


  not
  g650
  (
    n1220,
    n362
  );


  buf
  g651
  (
    n1736,
    n290
  );


  not
  g652
  (
    n1392,
    n261
  );


  buf
  g653
  (
    n842,
    n174
  );


  not
  g654
  (
    n540,
    n351
  );


  not
  g655
  (
    n1533,
    n317
  );


  not
  g656
  (
    n949,
    n313
  );


  buf
  g657
  (
    n1326,
    n211
  );


  not
  g658
  (
    n754,
    n251
  );


  buf
  g659
  (
    n1032,
    n212
  );


  buf
  g660
  (
    n880,
    n422
  );


  not
  g661
  (
    n579,
    n174
  );


  buf
  g662
  (
    n972,
    n435
  );


  buf
  g663
  (
    n638,
    n191
  );


  not
  g664
  (
    n1093,
    n230
  );


  buf
  g665
  (
    n1122,
    n317
  );


  not
  g666
  (
    n1351,
    n441
  );


  buf
  g667
  (
    n893,
    n412
  );


  buf
  g668
  (
    n1727,
    n202
  );


  buf
  g669
  (
    n652,
    n325
  );


  buf
  g670
  (
    n1356,
    n268
  );


  not
  g671
  (
    n1159,
    n251
  );


  not
  g672
  (
    n1091,
    n344
  );


  not
  g673
  (
    n1745,
    n339
  );


  buf
  g674
  (
    n1600,
    n387
  );


  buf
  g675
  (
    n1402,
    n212
  );


  buf
  g676
  (
    n666,
    n239
  );


  buf
  g677
  (
    n781,
    n210
  );


  not
  g678
  (
    n1688,
    n274
  );


  not
  g679
  (
    n1366,
    n234
  );


  buf
  g680
  (
    n1330,
    n154
  );


  not
  g681
  (
    n1061,
    n209
  );


  not
  g682
  (
    n1168,
    n395
  );


  not
  g683
  (
    n1016,
    n379
  );


  not
  g684
  (
    n1608,
    n238
  );


  not
  g685
  (
    n1345,
    n332
  );


  buf
  g686
  (
    n1110,
    n314
  );


  buf
  g687
  (
    n1004,
    n372
  );


  buf
  g688
  (
    n897,
    n407
  );


  buf
  g689
  (
    n669,
    n433
  );


  buf
  g690
  (
    n586,
    n244
  );


  buf
  g691
  (
    n1596,
    n302
  );


  not
  g692
  (
    n913,
    n268
  );


  buf
  g693
  (
    n659,
    n251
  );


  not
  g694
  (
    n524,
    n428
  );


  buf
  g695
  (
    n1000,
    n198
  );


  not
  g696
  (
    n1696,
    n256
  );


  buf
  g697
  (
    n740,
    n335
  );


  not
  g698
  (
    n1597,
    n288
  );


  not
  g699
  (
    n1292,
    n448
  );


  not
  g700
  (
    n1283,
    n293
  );


  not
  g701
  (
    n977,
    n320
  );


  not
  g702
  (
    n1549,
    n437
  );


  buf
  g703
  (
    n1027,
    n347
  );


  buf
  g704
  (
    n602,
    n361
  );


  not
  g705
  (
    n1432,
    n133
  );


  not
  g706
  (
    n1606,
    n336
  );


  buf
  g707
  (
    n822,
    n357
  );


  buf
  g708
  (
    n1146,
    n444
  );


  not
  g709
  (
    n642,
    n260
  );


  not
  g710
  (
    n844,
    n350
  );


  not
  g711
  (
    n1532,
    n303
  );


  not
  g712
  (
    n550,
    n195
  );


  not
  g713
  (
    n1096,
    n193
  );


  not
  g714
  (
    n973,
    n410
  );


  not
  g715
  (
    n1340,
    n414
  );


  buf
  g716
  (
    n1281,
    n234
  );


  not
  g717
  (
    n1113,
    n432
  );


  buf
  g718
  (
    n724,
    n141
  );


  not
  g719
  (
    n979,
    n403
  );


  buf
  g720
  (
    n1617,
    n403
  );


  not
  g721
  (
    n595,
    n310
  );


  not
  g722
  (
    n489,
    n165
  );


  buf
  g723
  (
    n1461,
    n321
  );


  not
  g724
  (
    n800,
    n356
  );


  buf
  g725
  (
    n1257,
    n344
  );


  not
  g726
  (
    n1587,
    n167
  );


  buf
  g727
  (
    n565,
    n157
  );


  buf
  g728
  (
    n1018,
    n334
  );


  buf
  g729
  (
    n852,
    n150
  );


  not
  g730
  (
    n864,
    n401
  );


  buf
  g731
  (
    n1107,
    n181
  );


  buf
  g732
  (
    n525,
    n205
  );


  not
  g733
  (
    n1460,
    n186
  );


  not
  g734
  (
    n655,
    n427
  );


  not
  g735
  (
    n1476,
    n352
  );


  buf
  g736
  (
    n1408,
    n317
  );


  not
  g737
  (
    n995,
    n455
  );


  buf
  g738
  (
    n1490,
    n431
  );


  buf
  g739
  (
    n1178,
    n345
  );


  not
  g740
  (
    n663,
    n407
  );


  buf
  g741
  (
    n543,
    n355
  );


  buf
  g742
  (
    n1485,
    n221
  );


  not
  g743
  (
    n1618,
    n216
  );


  not
  g744
  (
    n1247,
    n288
  );


  not
  g745
  (
    n946,
    n333
  );


  buf
  g746
  (
    n1735,
    n250
  );


  not
  g747
  (
    n1214,
    n224
  );


  not
  g748
  (
    n1267,
    n426
  );


  buf
  g749
  (
    n922,
    n433
  );


  buf
  g750
  (
    n1278,
    n149
  );


  buf
  g751
  (
    n956,
    n276
  );


  buf
  g752
  (
    n633,
    n413
  );


  buf
  g753
  (
    n1636,
    n421
  );


  not
  g754
  (
    n915,
    n341
  );


  buf
  g755
  (
    n707,
    n450
  );


  not
  g756
  (
    n763,
    n195
  );


  buf
  g757
  (
    n1725,
    n268
  );


  not
  g758
  (
    n700,
    n240
  );


  buf
  g759
  (
    n1667,
    n426
  );


  buf
  g760
  (
    n1643,
    n146
  );


  not
  g761
  (
    n628,
    n319
  );


  not
  g762
  (
    n1628,
    n416
  );


  not
  g763
  (
    n850,
    n267
  );


  not
  g764
  (
    n1103,
    n160
  );


  not
  g765
  (
    n1502,
    n171
  );


  buf
  g766
  (
    n1129,
    n265
  );


  not
  g767
  (
    n651,
    n376
  );


  not
  g768
  (
    n780,
    n137
  );


  not
  g769
  (
    n709,
    n137
  );


  not
  g770
  (
    n676,
    n311
  );


  not
  g771
  (
    n1286,
    n329
  );


  not
  g772
  (
    n1358,
    n300
  );


  not
  g773
  (
    n1090,
    n200
  );


  buf
  g774
  (
    n1139,
    n250
  );


  buf
  g775
  (
    n1458,
    n129
  );


  not
  g776
  (
    n1553,
    n138
  );


  not
  g777
  (
    n984,
    n142
  );


  not
  g778
  (
    n1648,
    n130
  );


  buf
  g779
  (
    n1322,
    n349
  );


  not
  g780
  (
    n1321,
    n243
  );


  not
  g781
  (
    n919,
    n303
  );


  buf
  g782
  (
    n912,
    n236
  );


  not
  g783
  (
    n597,
    n373
  );


  not
  g784
  (
    n559,
    n282
  );


  buf
  g785
  (
    n742,
    n412
  );


  not
  g786
  (
    n894,
    n275
  );


  not
  g787
  (
    n1662,
    n428
  );


  buf
  g788
  (
    n816,
    n399
  );


  not
  g789
  (
    n522,
    n248
  );


  not
  g790
  (
    n1423,
    n215
  );


  buf
  g791
  (
    n959,
    n359
  );


  buf
  g792
  (
    n1422,
    n204
  );


  not
  g793
  (
    n1380,
    n197
  );


  buf
  g794
  (
    n1069,
    n164
  );


  buf
  g795
  (
    n620,
    n314
  );


  buf
  g796
  (
    n1344,
    n212
  );


  not
  g797
  (
    n615,
    n220
  );


  not
  g798
  (
    n1068,
    n421
  );


  not
  g799
  (
    n1456,
    n256
  );


  buf
  g800
  (
    n1447,
    n382
  );


  not
  g801
  (
    n662,
    n386
  );


  not
  g802
  (
    n1682,
    n226
  );


  not
  g803
  (
    n957,
    n262
  );


  buf
  g804
  (
    n699,
    n339
  );


  buf
  g805
  (
    n1428,
    n411
  );


  not
  g806
  (
    n1047,
    n435
  );


  buf
  g807
  (
    n1573,
    n343
  );


  not
  g808
  (
    n862,
    n296
  );


  not
  g809
  (
    n874,
    n191
  );


  not
  g810
  (
    n768,
    n366
  );


  buf
  g811
  (
    n773,
    n354
  );


  not
  g812
  (
    n1255,
    n178
  );


  buf
  g813
  (
    n1227,
    n360
  );


  not
  g814
  (
    n1101,
    n156
  );


  not
  g815
  (
    n1316,
    n367
  );


  buf
  g816
  (
    n1580,
    n350
  );


  buf
  g817
  (
    n1374,
    n277
  );


  buf
  g818
  (
    n1472,
    n223
  );


  not
  g819
  (
    n1073,
    n170
  );


  not
  g820
  (
    n1510,
    n419
  );


  not
  g821
  (
    n1611,
    n217
  );


  buf
  g822
  (
    n1026,
    n342
  );


  not
  g823
  (
    n1607,
    n254
  );


  buf
  g824
  (
    n1590,
    n163
  );


  not
  g825
  (
    n1082,
    n382
  );


  not
  g826
  (
    n1063,
    n161
  );


  not
  g827
  (
    n507,
    n249
  );


  not
  g828
  (
    n1202,
    n345
  );


  not
  g829
  (
    n1058,
    n390
  );


  buf
  g830
  (
    n1045,
    n247
  );


  not
  g831
  (
    n1712,
    n422
  );


  buf
  g832
  (
    n970,
    n325
  );


  buf
  g833
  (
    n1571,
    n417
  );


  not
  g834
  (
    n1443,
    n356
  );


  buf
  g835
  (
    n1747,
    n226
  );


  not
  g836
  (
    n1695,
    n164
  );


  buf
  g837
  (
    n1713,
    n131
  );


  buf
  g838
  (
    n718,
    n176
  );


  not
  g839
  (
    n583,
    n139
  );


  not
  g840
  (
    n1563,
    n316
  );


  buf
  g841
  (
    n794,
    n175
  );


  buf
  g842
  (
    n934,
    n261
  );


  buf
  g843
  (
    n1241,
    n378
  );


  buf
  g844
  (
    n1332,
    n170
  );


  not
  g845
  (
    n1352,
    n280
  );


  not
  g846
  (
    n1453,
    n277
  );


  buf
  g847
  (
    n472,
    n301
  );


  buf
  g848
  (
    n925,
    n144
  );


  buf
  g849
  (
    n1537,
    n134
  );


  not
  g850
  (
    n1235,
    n132
  );


  buf
  g851
  (
    n731,
    n398
  );


  not
  g852
  (
    n1405,
    n208
  );


  not
  g853
  (
    n795,
    n439
  );


  not
  g854
  (
    n1444,
    n428
  );


  not
  g855
  (
    n1038,
    n418
  );


  buf
  g856
  (
    n1467,
    n147
  );


  not
  g857
  (
    n1494,
    n314
  );


  buf
  g858
  (
    n968,
    n309
  );


  not
  g859
  (
    n576,
    n431
  );


  not
  g860
  (
    n1030,
    n225
  );


  buf
  g861
  (
    n1165,
    n197
  );


  buf
  g862
  (
    n834,
    n432
  );


  not
  g863
  (
    n1550,
    n350
  );


  not
  g864
  (
    n752,
    n252
  );


  buf
  g865
  (
    n826,
    n419
  );


  buf
  g866
  (
    n562,
    n416
  );


  not
  g867
  (
    n1566,
    n371
  );


  not
  g868
  (
    n1293,
    n375
  );


  not
  g869
  (
    n1655,
    n382
  );


  not
  g870
  (
    n1529,
    n164
  );


  buf
  g871
  (
    n1395,
    n320
  );


  not
  g872
  (
    n593,
    n316
  );


  buf
  g873
  (
    n1622,
    n371
  );


  not
  g874
  (
    n1592,
    n179
  );


  not
  g875
  (
    n847,
    n436
  );


  buf
  g876
  (
    n1394,
    n449
  );


  buf
  g877
  (
    n846,
    n152
  );


  buf
  g878
  (
    n644,
    n208
  );


  buf
  g879
  (
    n1290,
    n241
  );


  not
  g880
  (
    n1440,
    n190
  );


  buf
  g881
  (
    n473,
    n437
  );


  not
  g882
  (
    n1640,
    n283
  );


  not
  g883
  (
    n820,
    n426
  );


  not
  g884
  (
    n726,
    n281
  );


  not
  g885
  (
    n1717,
    n355
  );


  not
  g886
  (
    n1603,
    n324
  );


  buf
  g887
  (
    n520,
    n451
  );


  buf
  g888
  (
    n1240,
    n432
  );


  not
  g889
  (
    n1248,
    n213
  );


  not
  g890
  (
    n591,
    n425
  );


  not
  g891
  (
    n1387,
    n278
  );


  buf
  g892
  (
    n1479,
    n137
  );


  buf
  g893
  (
    n1085,
    n234
  );


  not
  g894
  (
    n1363,
    n284
  );


  not
  g895
  (
    n746,
    n279
  );


  not
  g896
  (
    n1642,
    n324
  );


  not
  g897
  (
    n939,
    n402
  );


  buf
  g898
  (
    n830,
    n245
  );


  buf
  g899
  (
    n1739,
    n224
  );


  buf
  g900
  (
    n770,
    n131
  );


  buf
  g901
  (
    n1051,
    n291
  );


  buf
  g902
  (
    n1019,
    n306
  );


  buf
  g903
  (
    n1279,
    n448
  );


  buf
  g904
  (
    n1033,
    n224
  );


  buf
  g905
  (
    n483,
    n129
  );


  buf
  g906
  (
    n825,
    n177
  );


  buf
  g907
  (
    n1427,
    n334
  );


  not
  g908
  (
    n1591,
    n409
  );


  not
  g909
  (
    n1732,
    n316
  );


  buf
  g910
  (
    n1703,
    n191
  );


  buf
  g911
  (
    n514,
    n158
  );


  not
  g912
  (
    n1177,
    n172
  );


  not
  g913
  (
    n561,
    n243
  );


  buf
  g914
  (
    n1435,
    n260
  );


  buf
  g915
  (
    n1212,
    n315
  );


  not
  g916
  (
    n737,
    n250
  );


  not
  g917
  (
    n1724,
    n404
  );


  buf
  g918
  (
    n744,
    n190
  );


  not
  g919
  (
    n503,
    n447
  );


  not
  g920
  (
    n1517,
    n307
  );


  not
  g921
  (
    n786,
    n364
  );


  not
  g922
  (
    n1039,
    n133
  );


  not
  g923
  (
    n1111,
    n248
  );


  not
  g924
  (
    n779,
    n205
  );


  buf
  g925
  (
    n1353,
    n435
  );


  not
  g926
  (
    n1403,
    n235
  );


  buf
  g927
  (
    n1277,
    n256
  );


  not
  g928
  (
    n1300,
    n227
  );


  not
  g929
  (
    n767,
    n430
  );


  buf
  g930
  (
    n716,
    n258
  );


  not
  g931
  (
    n1540,
    n292
  );


  not
  g932
  (
    n857,
    n298
  );


  not
  g933
  (
    n1275,
    n286
  );


  not
  g934
  (
    n1515,
    n343
  );


  not
  g935
  (
    n528,
    n348
  );


  buf
  g936
  (
    n928,
    n372
  );


  not
  g937
  (
    n1306,
    n228
  );


  not
  g938
  (
    n908,
    n252
  );


  buf
  g939
  (
    n1327,
    n380
  );


  buf
  g940
  (
    n777,
    n337
  );


  not
  g941
  (
    n1610,
    n247
  );


  not
  g942
  (
    n1489,
    n204
  );


  not
  g943
  (
    n537,
    n286
  );


  buf
  g944
  (
    n637,
    n143
  );


  not
  g945
  (
    n978,
    n141
  );


  buf
  g946
  (
    n965,
    n404
  );


  buf
  g947
  (
    n1547,
    n135
  );


  not
  g948
  (
    n1224,
    n214
  );


  buf
  g949
  (
    n1378,
    n287
  );


  buf
  g950
  (
    n534,
    n343
  );


  buf
  g951
  (
    n1579,
    n436
  );


  not
  g952
  (
    n553,
    n441
  );


  buf
  g953
  (
    n588,
    n378
  );


  not
  g954
  (
    n1117,
    n335
  );


  not
  g955
  (
    n506,
    n450
  );


  not
  g956
  (
    n933,
    n335
  );


  not
  g957
  (
    n635,
    n406
  );


  not
  g958
  (
    n1635,
    n219
  );


  buf
  g959
  (
    n1743,
    n182
  );


  not
  g960
  (
    n578,
    n383
  );


  not
  g961
  (
    n1261,
    n159
  );


  not
  g962
  (
    n622,
    n203
  );


  buf
  g963
  (
    n802,
    n166
  );


  buf
  g964
  (
    n885,
    n165
  );


  buf
  g965
  (
    n871,
    n456
  );


  buf
  g966
  (
    n1086,
    n353
  );


  not
  g967
  (
    n1022,
    n186
  );


  buf
  g968
  (
    n835,
    n152
  );


  not
  g969
  (
    n854,
    n429
  );


  not
  g970
  (
    n1109,
    n445
  );


  not
  g971
  (
    n1060,
    n368
  );


  not
  g972
  (
    n1718,
    n306
  );


  buf
  g973
  (
    n491,
    n360
  );


  buf
  g974
  (
    n1583,
    n293
  );


  not
  g975
  (
    n1194,
    n229
  );


  buf
  g976
  (
    n1084,
    n178
  );


  not
  g977
  (
    n1315,
    n359
  );


  not
  g978
  (
    n1652,
    n384
  );


  not
  g979
  (
    n683,
    n142
  );


  not
  g980
  (
    n1514,
    n180
  );


  not
  g981
  (
    n1262,
    n300
  );


  not
  g982
  (
    n1015,
    n222
  );


  not
  g983
  (
    n1731,
    n217
  );


  buf
  g984
  (
    n1710,
    n233
  );


  buf
  g985
  (
    n1496,
    n238
  );


  buf
  g986
  (
    n866,
    n269
  );


  buf
  g987
  (
    n1681,
    n358
  );


  buf
  g988
  (
    n1187,
    n445
  );


  not
  g989
  (
    n1163,
    n332
  );


  buf
  g990
  (
    n658,
    n242
  );


  buf
  g991
  (
    n960,
    n404
  );


  buf
  g992
  (
    n551,
    n361
  );


  not
  g993
  (
    n1287,
    n323
  );


  buf
  g994
  (
    n1649,
    n324
  );


  buf
  g995
  (
    n488,
    n295
  );


  not
  g996
  (
    n523,
    n207
  );


  buf
  g997
  (
    n1335,
    n357
  );


  buf
  g998
  (
    n1729,
    n353
  );


  not
  g999
  (
    n1438,
    n188
  );


  not
  g1000
  (
    n1336,
    n364
  );


  buf
  g1001
  (
    n1269,
    n411
  );


  buf
  g1002
  (
    n1329,
    n370
  );


  buf
  g1003
  (
    n1143,
    n204
  );


  buf
  g1004
  (
    n600,
    n249
  );


  not
  g1005
  (
    n882,
    n374
  );


  not
  g1006
  (
    n1357,
    n154
  );


  not
  g1007
  (
    n1014,
    n362
  );


  not
  g1008
  (
    n1521,
    n144
  );


  not
  g1009
  (
    n604,
    n337
  );


  buf
  g1010
  (
    n1633,
    n387
  );


  buf
  g1011
  (
    n650,
    n238
  );


  buf
  g1012
  (
    n964,
    n236
  );


  not
  g1013
  (
    n1154,
    n423
  );


  not
  g1014
  (
    n765,
    n208
  );


  buf
  g1015
  (
    n656,
    n265
  );


  not
  g1016
  (
    n1367,
    n396
  );


  buf
  g1017
  (
    n1132,
    n275
  );


  buf
  g1018
  (
    n828,
    n409
  );


  buf
  g1019
  (
    n1072,
    n389
  );


  not
  g1020
  (
    n545,
    n405
  );


  not
  g1021
  (
    n1716,
    n218
  );


  buf
  g1022
  (
    n1260,
    n229
  );


  not
  g1023
  (
    n1190,
    n220
  );


  buf
  g1024
  (
    n1152,
    n360
  );


  buf
  g1025
  (
    n1312,
    n216
  );


  not
  g1026
  (
    n1570,
    n227
  );


  buf
  g1027
  (
    n677,
    n435
  );


  not
  g1028
  (
    n1062,
    n389
  );


  not
  g1029
  (
    n858,
    n142
  );


  buf
  g1030
  (
    n778,
    n207
  );


  not
  g1031
  (
    n722,
    n317
  );


  buf
  g1032
  (
    n587,
    n423
  );


  buf
  g1033
  (
    n1155,
    n167
  );


  not
  g1034
  (
    n646,
    n287
  );


  not
  g1035
  (
    n1215,
    n220
  );


  not
  g1036
  (
    n1721,
    n167
  );


  buf
  g1037
  (
    n911,
    n252
  );


  buf
  g1038
  (
    n1244,
    n342
  );


  not
  g1039
  (
    n1595,
    n132
  );


  not
  g1040
  (
    n1418,
    n456
  );


  buf
  g1041
  (
    n1581,
    n153
  );


  buf
  g1042
  (
    n1604,
    n156
  );


  not
  g1043
  (
    n533,
    n393
  );


  not
  g1044
  (
    n833,
    n408
  );


  not
  g1045
  (
    n1709,
    n376
  );


  buf
  g1046
  (
    n921,
    n441
  );


  buf
  g1047
  (
    n906,
    n159
  );


  buf
  g1048
  (
    n1404,
    n157
  );


  not
  g1049
  (
    n688,
    n231
  );


  buf
  g1050
  (
    n547,
    n294
  );


  not
  g1051
  (
    n1021,
    n297
  );


  buf
  g1052
  (
    n1714,
    n204
  );


  buf
  g1053
  (
    n558,
    n457
  );


  not
  g1054
  (
    n1705,
    n162
  );


  not
  g1055
  (
    n717,
    n299
  );


  not
  g1056
  (
    n1054,
    n200
  );


  not
  g1057
  (
    n829,
    n453
  );


  not
  g1058
  (
    n1223,
    n374
  );


  buf
  g1059
  (
    n668,
    n156
  );


  not
  g1060
  (
    n1341,
    n330
  );


  buf
  g1061
  (
    n903,
    n447
  );


  not
  g1062
  (
    n789,
    n263
  );


  buf
  g1063
  (
    n886,
    n437
  );


  not
  g1064
  (
    n945,
    n199
  );


  buf
  g1065
  (
    n1174,
    n140
  );


  buf
  g1066
  (
    n1585,
    n299
  );


  buf
  g1067
  (
    n1195,
    n421
  );


  buf
  g1068
  (
    n1448,
    n393
  );


  not
  g1069
  (
    n1131,
    n356
  );


  not
  g1070
  (
    n872,
    n350
  );


  buf
  g1071
  (
    n914,
    n146
  );


  not
  g1072
  (
    n1518,
    n430
  );


  not
  g1073
  (
    n544,
    n155
  );


  buf
  g1074
  (
    n1067,
    n348
  );


  buf
  g1075
  (
    n1612,
    n300
  );


  buf
  g1076
  (
    n1719,
    n225
  );


  buf
  g1077
  (
    n989,
    n420
  );


  buf
  g1078
  (
    n743,
    n135
  );


  buf
  g1079
  (
    n1179,
    n424
  );


  buf
  g1080
  (
    n999,
    n451
  );


  buf
  g1081
  (
    n804,
    n433
  );


  not
  g1082
  (
    n538,
    n176
  );


  buf
  g1083
  (
    n1233,
    n363
  );


  buf
  g1084
  (
    n787,
    n397
  );


  buf
  g1085
  (
    n680,
    n361
  );


  not
  g1086
  (
    n807,
    n337
  );


  buf
  g1087
  (
    n1040,
    n340
  );


  not
  g1088
  (
    n1150,
    n191
  );


  not
  g1089
  (
    n679,
    n209
  );


  not
  g1090
  (
    n1305,
    n190
  );


  not
  g1091
  (
    n1468,
    n311
  );


  buf
  g1092
  (
    n670,
    n239
  );


  buf
  g1093
  (
    n1115,
    n390
  );


  not
  g1094
  (
    n776,
    n178
  );


  not
  g1095
  (
    n1412,
    n197
  );


  buf
  g1096
  (
    n519,
    n374
  );


  not
  g1097
  (
    n1114,
    n288
  );


  buf
  g1098
  (
    n1420,
    n363
  );


  buf
  g1099
  (
    n900,
    n410
  );


  not
  g1100
  (
    n1704,
    n230
  );


  not
  g1101
  (
    n1361,
    n214
  );


  not
  g1102
  (
    n792,
    n358
  );


  buf
  g1103
  (
    n703,
    n230
  );


  not
  g1104
  (
    n909,
    n290
  );


  not
  g1105
  (
    n1543,
    n201
  );


  buf
  g1106
  (
    n1258,
    n171
  );


  not
  g1107
  (
    n480,
    n272
  );


  buf
  g1108
  (
    n760,
    n222
  );


  not
  g1109
  (
    n856,
    n309
  );


  buf
  g1110
  (
    n788,
    n454
  );


  not
  g1111
  (
    n1689,
    n381
  );


  buf
  g1112
  (
    n1230,
    n366
  );


  not
  g1113
  (
    n1508,
    n352
  );


  not
  g1114
  (
    n1541,
    n253
  );


  buf
  g1115
  (
    n1271,
    n398
  );


  not
  g1116
  (
    n1284,
    n149
  );


  buf
  g1117
  (
    n574,
    n399
  );


  buf
  g1118
  (
    n1441,
    n384
  );


  not
  g1119
  (
    n855,
    n347
  );


  not
  g1120
  (
    n1459,
    n427
  );


  buf
  g1121
  (
    n810,
    n396
  );


  buf
  g1122
  (
    n861,
    n377
  );


  buf
  g1123
  (
    n1081,
    n331
  );


  not
  g1124
  (
    n1574,
    n272
  );


  buf
  g1125
  (
    n951,
    n201
  );


  buf
  g1126
  (
    n1625,
    n373
  );


  not
  g1127
  (
    n1050,
    n381
  );


  buf
  g1128
  (
    n713,
    n280
  );


  buf
  g1129
  (
    n1098,
    n418
  );


  not
  g1130
  (
    n1406,
    n349
  );


  buf
  g1131
  (
    n1551,
    n215
  );


  buf
  g1132
  (
    n1048,
    n155
  );


  buf
  g1133
  (
    n1160,
    n341
  );


  not
  g1134
  (
    n747,
    n285
  );


  buf
  g1135
  (
    n818,
    n318
  );


  not
  g1136
  (
    n1052,
    n158
  );


  buf
  g1137
  (
    n1094,
    n183
  );


  not
  g1138
  (
    n571,
    n301
  );


  not
  g1139
  (
    n1501,
    n184
  );


  buf
  g1140
  (
    n504,
    n205
  );


  buf
  g1141
  (
    n971,
    n388
  );


  buf
  g1142
  (
    n1484,
    n443
  );


  not
  g1143
  (
    n931,
    n378
  );


  not
  g1144
  (
    n1706,
    n394
  );


  buf
  g1145
  (
    n1319,
    n408
  );


  not
  g1146
  (
    n1497,
    n202
  );


  buf
  g1147
  (
    n1201,
    n356
  );


  buf
  g1148
  (
    n1070,
    n302
  );


  buf
  g1149
  (
    n723,
    n418
  );


  buf
  g1150
  (
    n1020,
    n246
  );


  not
  g1151
  (
    n1498,
    n263
  );


  not
  g1152
  (
    n705,
    n342
  );


  not
  g1153
  (
    n609,
    n322
  );


  buf
  g1154
  (
    n1360,
    n346
  );


  buf
  g1155
  (
    n1041,
    n263
  );


  buf
  g1156
  (
    n567,
    n216
  );


  not
  g1157
  (
    n623,
    n369
  );


  buf
  g1158
  (
    n1707,
    n360
  );


  not
  g1159
  (
    n1417,
    n194
  );


  not
  g1160
  (
    n1671,
    n233
  );


  buf
  g1161
  (
    n1006,
    n380
  );


  buf
  g1162
  (
    n1362,
    n226
  );


  not
  g1163
  (
    n950,
    n346
  );


  not
  g1164
  (
    n1282,
    n311
  );


  buf
  g1165
  (
    n887,
    n135
  );


  not
  g1166
  (
    n1375,
    n318
  );


  buf
  g1167
  (
    n1697,
    n371
  );


  not
  g1168
  (
    n1049,
    n139
  );


  not
  g1169
  (
    n1564,
    n397
  );


  not
  g1170
  (
    n1527,
    n422
  );


  buf
  g1171
  (
    n479,
    n443
  );


  buf
  g1172
  (
    n494,
    n145
  );


  buf
  g1173
  (
    n527,
    n136
  );


  buf
  g1174
  (
    n1430,
    n182
  );


  not
  g1175
  (
    n1650,
    n164
  );


  buf
  g1176
  (
    n1621,
    n177
  );


  not
  g1177
  (
    n1516,
    n312
  );


  buf
  g1178
  (
    n797,
    n361
  );


  not
  g1179
  (
    n1274,
    n300
  );


  buf
  g1180
  (
    n1557,
    n218
  );


  not
  g1181
  (
    n1184,
    n349
  );


  buf
  g1182
  (
    n863,
    n315
  );


  buf
  g1183
  (
    n1701,
    n284
  );


  not
  g1184
  (
    n1659,
    n134
  );


  buf
  g1185
  (
    n840,
    n256
  );


  not
  g1186
  (
    n1080,
    n219
  );


  buf
  g1187
  (
    n630,
    n452
  );


  buf
  g1188
  (
    n1044,
    n434
  );


  buf
  g1189
  (
    n1372,
    n292
  );


  buf
  g1190
  (
    n1525,
    n302
  );


  not
  g1191
  (
    n753,
    n185
  );


  not
  g1192
  (
    n1627,
    n424
  );


  buf
  g1193
  (
    n1333,
    n447
  );


  buf
  g1194
  (
    n1619,
    n249
  );


  not
  g1195
  (
    n890,
    n319
  );


  buf
  g1196
  (
    n654,
    n250
  );


  buf
  g1197
  (
    n1191,
    n183
  );


  not
  g1198
  (
    n1507,
    n222
  );


  not
  g1199
  (
    n1295,
    n149
  );


  not
  g1200
  (
    n873,
    n267
  );


  buf
  g1201
  (
    n634,
    n131
  );


  buf
  g1202
  (
    n1429,
    n211
  );


  not
  g1203
  (
    n499,
    n237
  );


  buf
  g1204
  (
    n918,
    n189
  );


  buf
  g1205
  (
    n1368,
    n200
  );


  buf
  g1206
  (
    n766,
    n190
  );


  buf
  g1207
  (
    n1386,
    n270
  );


  buf
  g1208
  (
    n1634,
    n332
  );


  buf
  g1209
  (
    n1171,
    n284
  );


  not
  g1210
  (
    n966,
    n238
  );


  buf
  g1211
  (
    n1409,
    n258
  );


  not
  g1212
  (
    n1449,
    n246
  );


  buf
  g1213
  (
    n1087,
    n307
  );


  buf
  g1214
  (
    n1466,
    n401
  );


  buf
  g1215
  (
    n1410,
    n272
  );


  not
  g1216
  (
    n1569,
    n342
  );


  buf
  g1217
  (
    n572,
    n203
  );


  buf
  g1218
  (
    n696,
    n184
  );


  not
  g1219
  (
    n1700,
    n196
  );


  buf
  g1220
  (
    n1488,
    n453
  );


  buf
  g1221
  (
    n1173,
    n229
  );


  buf
  g1222
  (
    n869,
    n266
  );


  buf
  g1223
  (
    n1147,
    n346
  );


  not
  g1224
  (
    n619,
    n296
  );


  buf
  g1225
  (
    n1234,
    n452
  );


  buf
  g1226
  (
    n1646,
    n257
  );


  not
  g1227
  (
    n1013,
    n264
  );


  buf
  g1228
  (
    n899,
    n236
  );


  buf
  g1229
  (
    n1506,
    n334
  );


  not
  g1230
  (
    n487,
    n332
  );


  buf
  g1231
  (
    n848,
    n240
  );


  buf
  g1232
  (
    n607,
    n206
  );


  buf
  g1233
  (
    n1545,
    n157
  );


  not
  g1234
  (
    n720,
    n170
  );


  buf
  g1235
  (
    n513,
    n151
  );


  buf
  g1236
  (
    n799,
    n370
  );


  buf
  g1237
  (
    n1346,
    n366
  );


  buf
  g1238
  (
    n1535,
    n137
  );


  buf
  g1239
  (
    n660,
    n144
  );


  buf
  g1240
  (
    n1140,
    n365
  );


  buf
  g1241
  (
    n590,
    n223
  );


  not
  g1242
  (
    n476,
    n262
  );


  buf
  g1243
  (
    n841,
    n322
  );


  not
  g1244
  (
    n1180,
    n167
  );


  buf
  g1245
  (
    n1396,
    n209
  );


  buf
  g1246
  (
    n958,
    n154
  );


  not
  g1247
  (
    n1511,
    n365
  );


  buf
  g1248
  (
    n618,
    n283
  );


  buf
  g1249
  (
    n549,
    n297
  );


  buf
  g1250
  (
    n811,
    n259
  );


  buf
  g1251
  (
    n1684,
    n331
  );


  buf
  g1252
  (
    n1377,
    n402
  );


  not
  g1253
  (
    n859,
    n305
  );


  buf
  g1254
  (
    n824,
    n187
  );


  not
  g1255
  (
    n701,
    n134
  );


  buf
  g1256
  (
    n1715,
    n176
  );


  buf
  g1257
  (
    n1199,
    n210
  );


  buf
  g1258
  (
    n748,
    n439
  );


  buf
  g1259
  (
    n878,
    n273
  );


  buf
  g1260
  (
    n1740,
    n232
  );


  not
  g1261
  (
    n983,
    n414
  );


  buf
  g1262
  (
    n1324,
    n415
  );


  not
  g1263
  (
    n1568,
    n276
  );


  not
  g1264
  (
    n1161,
    n349
  );


  buf
  g1265
  (
    n1325,
    n308
  );


  not
  g1266
  (
    n605,
    n391
  );


  buf
  g1267
  (
    n1723,
    n399
  );


  not
  g1268
  (
    n570,
    n244
  );


  not
  g1269
  (
    n1089,
    n321
  );


  not
  g1270
  (
    n1385,
    n389
  );


  not
  g1271
  (
    n926,
    n390
  );


  buf
  g1272
  (
    n478,
    n415
  );


  buf
  g1273
  (
    n1741,
    n259
  );


  buf
  g1274
  (
    n1042,
    n173
  );


  buf
  g1275
  (
    n976,
    n417
  );


  not
  g1276
  (
    n1289,
    n427
  );


  buf
  g1277
  (
    n785,
    n442
  );


  buf
  g1278
  (
    n657,
    n214
  );


  not
  g1279
  (
    n1452,
    n260
  );


  not
  g1280
  (
    n1605,
    n241
  );


  not
  g1281
  (
    n647,
    n166
  );


  not
  g1282
  (
    n493,
    n365
  );


  buf
  g1283
  (
    n575,
    n438
  );


  buf
  g1284
  (
    n942,
    n441
  );


  buf
  g1285
  (
    n661,
    n379
  );


  buf
  g1286
  (
    n1037,
    n336
  );


  not
  g1287
  (
    n1520,
    n304
  );


  buf
  g1288
  (
    n1342,
    n372
  );


  not
  g1289
  (
    n932,
    n130
  );


  buf
  g1290
  (
    n739,
    n211
  );


  not
  g1291
  (
    n484,
    n437
  );


  not
  g1292
  (
    n756,
    n328
  );


  buf
  g1293
  (
    n806,
    n232
  );


  buf
  g1294
  (
    n1365,
    n235
  );


  not
  g1295
  (
    n1505,
    n146
  );


  buf
  g1296
  (
    n497,
    n295
  );


  not
  g1297
  (
    n775,
    n318
  );


  not
  g1298
  (
    n1349,
    n409
  );


  buf
  g1299
  (
    n1211,
    n141
  );


  buf
  g1300
  (
    n1317,
    n150
  );


  buf
  g1301
  (
    n904,
    n425
  );


  buf
  g1302
  (
    n796,
    n312
  );


  not
  g1303
  (
    n627,
    n148
  );


  not
  g1304
  (
    n1088,
    n319
  );


  buf
  g1305
  (
    n1156,
    n210
  );


  buf
  g1306
  (
    n1539,
    n299
  );


  not
  g1307
  (
    n1593,
    n145
  );


  not
  g1308
  (
    n517,
    n206
  );


  not
  g1309
  (
    n1623,
    n242
  );


  not
  g1310
  (
    n1102,
    n140
  );


  not
  g1311
  (
    n827,
    n248
  );


  buf
  g1312
  (
    n501,
    n129
  );


  not
  g1313
  (
    n1555,
    n337
  );


  buf
  g1314
  (
    n1127,
    n314
  );


  buf
  g1315
  (
    n682,
    n151
  );


  buf
  g1316
  (
    n1121,
    n439
  );


  buf
  g1317
  (
    n631,
    n279
  );


  buf
  g1318
  (
    n521,
    n294
  );


  not
  g1319
  (
    n560,
    n153
  );


  buf
  g1320
  (
    n943,
    n410
  );


  not
  g1321
  (
    n1024,
    n312
  );


  not
  g1322
  (
    n1499,
    n400
  );


  not
  g1323
  (
    n793,
    n411
  );


  not
  g1324
  (
    n981,
    n371
  );


  not
  g1325
  (
    n530,
    n305
  );


  not
  g1326
  (
    n495,
    n442
  );


  not
  g1327
  (
    n1205,
    n444
  );


  buf
  g1328
  (
    n757,
    n291
  );


  buf
  g1329
  (
    n812,
    n153
  );


  not
  g1330
  (
    n891,
    n237
  );


  not
  g1331
  (
    n1112,
    n373
  );


  not
  g1332
  (
    n865,
    n286
  );


  not
  g1333
  (
    n636,
    n280
  );


  not
  g1334
  (
    n772,
    n412
  );


  buf
  g1335
  (
    n1523,
    n385
  );


  buf
  g1336
  (
    n1264,
    n295
  );


  not
  g1337
  (
    n617,
    n169
  );


  buf
  g1338
  (
    n526,
    n136
  );


  buf
  g1339
  (
    n1226,
    n237
  );


  not
  g1340
  (
    n1181,
    n264
  );


  not
  g1341
  (
    n1582,
    n231
  );


  buf
  g1342
  (
    n1450,
    n303
  );


  not
  g1343
  (
    n1172,
    n232
  );


  buf
  g1344
  (
    n1419,
    n154
  );


  not
  g1345
  (
    n1451,
    n161
  );


  buf
  g1346
  (
    n714,
    n161
  );


  not
  g1347
  (
    n1270,
    n143
  );


  buf
  g1348
  (
    n1661,
    n362
  );


  buf
  g1349
  (
    n764,
    n415
  );


  not
  g1350
  (
    n1382,
    n276
  );


  not
  g1351
  (
    n474,
    n382
  );


  not
  g1352
  (
    n1252,
    n383
  );


  not
  g1353
  (
    n1296,
    n213
  );


  not
  g1354
  (
    n761,
    n194
  );


  not
  g1355
  (
    n1421,
    n194
  );


  buf
  g1356
  (
    n1100,
    n308
  );


  buf
  g1357
  (
    n641,
    n258
  );


  not
  g1358
  (
    n910,
    n398
  );


  buf
  g1359
  (
    n719,
    n348
  );


  buf
  g1360
  (
    n920,
    n179
  );


  not
  g1361
  (
    n1307,
    n304
  );


  buf
  g1362
  (
    n1397,
    n302
  );


  buf
  g1363
  (
    n1480,
    n396
  );


  not
  g1364
  (
    n1133,
    n305
  );


  buf
  g1365
  (
    n986,
    n183
  );


  buf
  g1366
  (
    n563,
    n299
  );


  not
  g1367
  (
    n1188,
    n174
  );


  buf
  g1368
  (
    n1464,
    n309
  );


  buf
  g1369
  (
    n769,
    n411
  );


  buf
  g1370
  (
    n632,
    n368
  );


  not
  g1371
  (
    n692,
    n396
  );


  not
  g1372
  (
    n711,
    n261
  );


  not
  g1373
  (
    n580,
    n416
  );


  buf
  g1374
  (
    n1092,
    n384
  );


  buf
  g1375
  (
    n935,
    n180
  );


  not
  g1376
  (
    n704,
    n289
  );


  buf
  g1377
  (
    n1746,
    n338
  );


  buf
  g1378
  (
    n755,
    n381
  );


  buf
  g1379
  (
    n1546,
    n406
  );


  buf
  g1380
  (
    n1071,
    n446
  );


  not
  g1381
  (
    n975,
    n168
  );


  not
  g1382
  (
    n1250,
    n303
  );


  buf
  g1383
  (
    n1134,
    n220
  );


  buf
  g1384
  (
    n710,
    n424
  );


  buf
  g1385
  (
    n1391,
    n395
  );


  buf
  g1386
  (
    n1737,
    n394
  );


  buf
  g1387
  (
    n1426,
    n448
  );


  buf
  g1388
  (
    n1217,
    n390
  );


  buf
  g1389
  (
    n1434,
    n270
  );


  not
  g1390
  (
    n1208,
    n421
  );


  buf
  g1391
  (
    n1158,
    n282
  );


  not
  g1392
  (
    n895,
    n173
  );


  buf
  g1393
  (
    n1477,
    n405
  );


  buf
  g1394
  (
    n930,
    n330
  );


  buf
  g1395
  (
    n838,
    n301
  );


  not
  g1396
  (
    n1562,
    n400
  );


  not
  g1397
  (
    n1145,
    n301
  );


  not
  g1398
  (
    n1457,
    n431
  );


  not
  g1399
  (
    n998,
    n130
  );


  not
  g1400
  (
    n1198,
    n357
  );


  not
  g1401
  (
    n1280,
    n387
  );


  buf
  g1402
  (
    n1674,
    n192
  );


  not
  g1403
  (
    n730,
    n218
  );


  not
  g1404
  (
    n749,
    n153
  );


  buf
  g1405
  (
    n759,
    n152
  );


  buf
  g1406
  (
    n1641,
    n251
  );


  buf
  g1407
  (
    n851,
    n194
  );


  buf
  g1408
  (
    n1303,
    n354
  );


  not
  g1409
  (
    n608,
    n198
  );


  not
  g1410
  (
    n1373,
    n255
  );


  not
  g1411
  (
    n1077,
    n166
  );


  buf
  g1412
  (
    n1065,
    n304
  );


  buf
  g1413
  (
    n1474,
    n341
  );


  not
  g1414
  (
    n1666,
    n320
  );


  not
  g1415
  (
    n1001,
    n274
  );


  not
  g1416
  (
    n1609,
    n257
  );


  not
  g1417
  (
    n508,
    n132
  );


  not
  g1418
  (
    n990,
    n284
  );


  not
  g1419
  (
    n674,
    n227
  );


  not
  g1420
  (
    n1079,
    n436
  );


  buf
  g1421
  (
    n1031,
    n239
  );


  not
  g1422
  (
    n1692,
    n151
  );


  not
  g1423
  (
    n685,
    n169
  );


  buf
  g1424
  (
    n1513,
    n420
  );


  buf
  g1425
  (
    n896,
    n323
  );


  buf
  g1426
  (
    n702,
    n399
  );


  not
  g1427
  (
    n1007,
    n368
  );


  buf
  g1428
  (
    n518,
    n440
  );


  not
  g1429
  (
    n598,
    n450
  );


  not
  g1430
  (
    n996,
    n287
  );


  not
  g1431
  (
    n1722,
    n322
  );


  buf
  g1432
  (
    n712,
    n170
  );


  buf
  g1433
  (
    n1470,
    n336
  );


  buf
  g1434
  (
    n961,
    n144
  );


  buf
  g1435
  (
    n1598,
    n290
  );


  not
  g1436
  (
    n815,
    n241
  );


  not
  g1437
  (
    n994,
    n205
  );


  buf
  g1438
  (
    n992,
    n189
  );


  buf
  g1439
  (
    n471,
    n175
  );


  buf
  g1440
  (
    n1095,
    n193
  );


  not
  g1441
  (
    n1334,
    n338
  );


  not
  g1442
  (
    n1204,
    n219
  );


  buf
  g1443
  (
    n1206,
    n355
  );


  buf
  g1444
  (
    n1126,
    n165
  );


  not
  g1445
  (
    n485,
    n255
  );


  buf
  g1446
  (
    n1685,
    n446
  );


  buf
  g1447
  (
    n924,
    n193
  );


  buf
  g1448
  (
    n1266,
    n248
  );


  not
  g1449
  (
    n1616,
    n402
  );


  not
  g1450
  (
    n1478,
    n457
  );


  buf
  g1451
  (
    n849,
    n163
  );


  not
  g1452
  (
    n993,
    n264
  );


  buf
  g1453
  (
    n1483,
    n329
  );


  not
  g1454
  (
    n1182,
    n321
  );


  buf
  g1455
  (
    n1219,
    n165
  );


  not
  g1456
  (
    n1099,
    n344
  );


  not
  g1457
  (
    n698,
    n216
  );


  buf
  g1458
  (
    n686,
    n380
  );


  buf
  g1459
  (
    n531,
    n369
  );


  not
  g1460
  (
    n1169,
    n428
  );


  buf
  g1461
  (
    n1379,
    n147
  );


  buf
  g1462
  (
    n1711,
    n308
  );


  not
  g1463
  (
    n1690,
    n429
  );


  buf
  g1464
  (
    n1338,
    n409
  );


  not
  g1465
  (
    n1339,
    n444
  );


  buf
  g1466
  (
    n1144,
    n212
  );


  buf
  g1467
  (
    n1097,
    n221
  );


  not
  g1468
  (
    n1694,
    n393
  );


  buf
  g1469
  (
    n1200,
    n183
  );


  not
  g1470
  (
    n1294,
    n340
  );


  not
  g1471
  (
    n732,
    n206
  );


  buf
  g1472
  (
    n1108,
    n162
  );


  buf
  g1473
  (
    n512,
    n339
  );


  buf
  g1474
  (
    n1437,
    n201
  );


  not
  g1475
  (
    n1228,
    n331
  );


  buf
  g1476
  (
    n1285,
    n432
  );


  not
  g1477
  (
    n917,
    n187
  );


  not
  g1478
  (
    n782,
    n265
  );


  not
  g1479
  (
    n1599,
    n320
  );


  not
  g1480
  (
    n1588,
    n410
  );


  not
  g1481
  (
    n944,
    n298
  );


  not
  g1482
  (
    n1118,
    n354
  );


  not
  g1483
  (
    n1602,
    n446
  );


  not
  g1484
  (
    n625,
    n369
  );


  not
  g1485
  (
    n1424,
    n200
  );


  buf
  g1486
  (
    n883,
    n294
  );


  not
  g1487
  (
    n539,
    n152
  );


  buf
  g1488
  (
    n839,
    n262
  );


  not
  g1489
  (
    n665,
    n161
  );


  not
  g1490
  (
    n1238,
    n207
  );


  not
  g1491
  (
    n548,
    n265
  );


  not
  g1492
  (
    n751,
    n139
  );


  buf
  g1493
  (
    n1584,
    n365
  );


  buf
  g1494
  (
    n1542,
    n351
  );


  buf
  g1495
  (
    n1078,
    n285
  );


  not
  g1496
  (
    n541,
    n434
  );


  not
  g1497
  (
    n889,
    n196
  );


  not
  g1498
  (
    n1677,
    n324
  );


  buf
  g1499
  (
    n1313,
    n246
  );


  buf
  g1500
  (
    n1162,
    n136
  );


  not
  g1501
  (
    n783,
    n438
  );


  buf
  g1502
  (
    n1210,
    n343
  );


  not
  g1503
  (
    n1544,
    n352
  );


  buf
  g1504
  (
    n808,
    n247
  );


  buf
  g1505
  (
    n1272,
    n285
  );


  not
  g1506
  (
    n805,
    n329
  );


  buf
  g1507
  (
    n1183,
    n243
  );


  buf
  g1508
  (
    n1232,
    n333
  );


  not
  g1509
  (
    n1130,
    n143
  );


  buf
  g1510
  (
    n1010,
    n198
  );


  buf
  g1511
  (
    n916,
    n370
  );


  not
  g1512
  (
    n819,
    n271
  );


  buf
  g1513
  (
    n798,
    n353
  );


  buf
  g1514
  (
    n1348,
    n438
  );


  buf
  g1515
  (
    n905,
    n193
  );


  not
  g1516
  (
    n566,
    n198
  );


  buf
  g1517
  (
    n1657,
    n385
  );


  buf
  g1518
  (
    n1630,
    n232
  );


  not
  g1519
  (
    n1136,
    n419
  );


  not
  g1520
  (
    n734,
    n340
  );


  not
  g1521
  (
    n1350,
    n253
  );


  not
  g1522
  (
    n1046,
    n175
  );


  buf
  g1523
  (
    n745,
    n158
  );


  buf
  g1524
  (
    n1455,
    n281
  );


  buf
  g1525
  (
    n1389,
    n263
  );


  not
  g1526
  (
    n801,
    n336
  );


  not
  g1527
  (
    n1297,
    n169
  );


  buf
  g1528
  (
    n1028,
    n328
  );


  buf
  g1529
  (
    n505,
    n169
  );


  buf
  g1530
  (
    n694,
    n182
  );


  not
  g1531
  (
    n477,
    n367
  );


  buf
  g1532
  (
    n554,
    n449
  );


  buf
  g1533
  (
    n1720,
    n386
  );


  not
  g1534
  (
    n1359,
    n259
  );


  buf
  g1535
  (
    n511,
    n266
  );


  buf
  g1536
  (
    n643,
    n177
  );


  not
  g1537
  (
    n594,
    n440
  );


  buf
  g1538
  (
    n1503,
    n420
  );


  buf
  g1539
  (
    n1637,
    n345
  );


  not
  g1540
  (
    n1376,
    n275
  );


  not
  g1541
  (
    n853,
    n313
  );


  not
  g1542
  (
    n1493,
    n452
  );


  not
  g1543
  (
    n1414,
    n258
  );


  not
  g1544
  (
    n1364,
    n426
  );


  not
  g1545
  (
    n727,
    n278
  );


  not
  g1546
  (
    n1601,
    n172
  );


  not
  g1547
  (
    n955,
    n133
  );


  buf
  g1548
  (
    n1442,
    n412
  );


  buf
  g1549
  (
    n1647,
    n174
  );


  buf
  g1550
  (
    n1644,
    n384
  );


  buf
  g1551
  (
    n1023,
    n306
  );


  buf
  g1552
  (
    n953,
    n139
  );


  not
  g1553
  (
    n1469,
    n454
  );


  buf
  g1554
  (
    n1216,
    n143
  );


  buf
  g1555
  (
    n1475,
    n388
  );


  not
  g1556
  (
    n1142,
    n246
  );


  buf
  g1557
  (
    n1586,
    n176
  );


  buf
  g1558
  (
    n1105,
    n185
  );


  buf
  g1559
  (
    n929,
    n339
  );


  not
  g1560
  (
    n475,
    n416
  );


  not
  g1561
  (
    n648,
    n179
  );


  not
  g1562
  (
    n1310,
    n444
  );


  not
  g1563
  (
    n1056,
    n297
  );


  not
  g1564
  (
    n616,
    n228
  );


  buf
  g1565
  (
    n510,
    n228
  );


  buf
  g1566
  (
    n1209,
    n189
  );


  buf
  g1567
  (
    n1390,
    n440
  );


  not
  g1568
  (
    n1323,
    n385
  );


  buf
  g1569
  (
    n1534,
    n377
  );


  buf
  g1570
  (
    n969,
    n223
  );


  buf
  g1571
  (
    n877,
    n383
  );


  not
  g1572
  (
    n988,
    n214
  );


  not
  g1573
  (
    n1471,
    n234
  );


  buf
  g1574
  (
    n1675,
    n413
  );


  buf
  g1575
  (
    n697,
    n182
  );


  not
  g1576
  (
    n589,
    n160
  );


  not
  g1577
  (
    n1253,
    n255
  );


  buf
  g1578
  (
    n1189,
    n203
  );


  not
  g1579
  (
    n1733,
    n455
  );


  not
  g1580
  (
    n1008,
    n400
  );


  not
  g1581
  (
    n509,
    n321
  );


  buf
  g1582
  (
    n735,
    n359
  );


  not
  g1583
  (
    n1632,
    n351
  );


  not
  g1584
  (
    n645,
    n235
  );


  not
  g1585
  (
    n1245,
    n130
  );


  not
  g1586
  (
    n1029,
    n171
  );


  not
  g1587
  (
    n1691,
    n293
  );


  not
  g1588
  (
    n1530,
    n184
  );


  buf
  g1589
  (
    n1678,
    n222
  );


  buf
  g1590
  (
    n502,
    n206
  );


  not
  g1591
  (
    n1053,
    n148
  );


  not
  g1592
  (
    n492,
    n241
  );


  buf
  g1593
  (
    n1416,
    n318
  );


  not
  g1594
  (
    n1445,
    n264
  );


  not
  g1595
  (
    n947,
    n151
  );


  not
  g1596
  (
    n1576,
    n310
  );


  buf
  g1597
  (
    n1237,
    n439
  );


  buf
  g1598
  (
    n741,
    n298
  );


  not
  g1599
  (
    n1708,
    n173
  );


  buf
  g1600
  (
    n1197,
    n376
  );


  buf
  g1601
  (
    n1728,
    n453
  );


  not
  g1602
  (
    n1203,
    n290
  );


  buf
  g1603
  (
    n860,
    n257
  );


  buf
  g1604
  (
    n1299,
    n353
  );


  buf
  g1605
  (
    n1318,
    n289
  );


  not
  g1606
  (
    n1578,
    n236
  );


  not
  g1607
  (
    n1193,
    n333
  );


  buf
  g1608
  (
    n1431,
    n274
  );


  not
  g1609
  (
    n695,
    n347
  );


  buf
  g1610
  (
    n1064,
    n352
  );


  not
  g1611
  (
    n762,
    n272
  );


  buf
  g1612
  (
    n725,
    n252
  );


  buf
  g1613
  (
    n1151,
    n281
  );


  not
  g1614
  (
    n1473,
    n260
  );


  not
  g1615
  (
    n1509,
    n408
  );


  buf
  g1616
  (
    n1298,
    n451
  );


  not
  g1617
  (
    n1425,
    n211
  );


  not
  g1618
  (
    n482,
    n392
  );


  buf
  g1619
  (
    n1702,
    n156
  );


  not
  g1620
  (
    n693,
    n271
  );


  not
  g1621
  (
    n1668,
    n449
  );


  not
  g1622
  (
    n1565,
    n196
  );


  not
  g1623
  (
    n1221,
    n287
  );


  not
  g1624
  (
    n938,
    n196
  );


  not
  g1625
  (
    n952,
    n282
  );


  buf
  g1626
  (
    n1025,
    n326
  );


  not
  g1627
  (
    n991,
    n451
  );


  not
  g1628
  (
    n516,
    n254
  );


  not
  g1629
  (
    n1401,
    n208
  );


  not
  g1630
  (
    n498,
    n406
  );


  buf
  g1631
  (
    n728,
    n145
  );


  not
  g1632
  (
    n1393,
    n228
  );


  not
  g1633
  (
    n1481,
    n131
  );


  not
  g1634
  (
    n1486,
    n315
  );


  not
  g1635
  (
    n1658,
    n379
  );


  not
  g1636
  (
    n1558,
    n389
  );


  buf
  g1637
  (
    n1500,
    n383
  );


  not
  g1638
  (
    n1454,
    n237
  );


  not
  g1639
  (
    n1673,
    n373
  );


  not
  g1640
  (
    n1669,
    n270
  );


  not
  g1641
  (
    n1492,
    n358
  );


  not
  g1642
  (
    n1288,
    n186
  );


  buf
  g1643
  (
    n1524,
    n374
  );


  buf
  g1644
  (
    n1589,
    n341
  );


  not
  g1645
  (
    n1536,
    n375
  );


  not
  g1646
  (
    n1680,
    n163
  );


  buf
  g1647
  (
    n1009,
    n394
  );


  not
  g1648
  (
    n1057,
    n425
  );


  buf
  g1649
  (
    n1002,
    n376
  );


  not
  g1650
  (
    n1613,
    n296
  );


  not
  g1651
  (
    n624,
    n243
  );


  not
  g1652
  (
    n689,
    n147
  );


  buf
  g1653
  (
    n1381,
    n445
  );


  not
  g1654
  (
    n1491,
    n201
  );


  buf
  g1655
  (
    n1170,
    n367
  );


  not
  g1656
  (
    n691,
    n186
  );


  not
  g1657
  (
    n1153,
    n335
  );


  not
  g1658
  (
    n1259,
    n328
  );


  buf
  g1659
  (
    n1263,
    n319
  );


  buf
  g1660
  (
    n1251,
    n187
  );


  not
  g1661
  (
    n496,
    n289
  );


  buf
  g1662
  (
    n817,
    n225
  );


  not
  g1663
  (
    n1407,
    n188
  );


  buf
  g1664
  (
    n941,
    n178
  );


  buf
  g1665
  (
    n980,
    n346
  );


  buf
  g1666
  (
    n1229,
    n218
  );


  not
  g1667
  (
    n611,
    n245
  );


  not
  g1668
  (
    n1343,
    n273
  );


  not
  g1669
  (
    n500,
    n229
  );


  buf
  g1670
  (
    n1225,
    n262
  );


  buf
  g1671
  (
    n1231,
    n140
  );


  not
  g1672
  (
    n1462,
    n268
  );


  not
  g1673
  (
    n1687,
    n354
  );


  not
  g1674
  (
    n1175,
    n270
  );


  buf
  g1675
  (
    n962,
    n163
  );


  buf
  g1676
  (
    n1164,
    n331
  );


  not
  g1677
  (
    n542,
    n157
  );


  buf
  g1678
  (
    n614,
    n279
  );


  buf
  g1679
  (
    n1176,
    n132
  );


  buf
  g1680
  (
    n823,
    n433
  );


  buf
  g1681
  (
    n1528,
    n344
  );


  buf
  g1682
  (
    n1446,
    n311
  );


  buf
  g1683
  (
    n1663,
    n292
  );


  buf
  g1684
  (
    n1615,
    n195
  );


  buf
  g1685
  (
    n1331,
    n449
  );


  not
  g1686
  (
    n1734,
    n294
  );


  not
  g1687
  (
    n1575,
    n168
  );


  buf
  g1688
  (
    n1308,
    n225
  );


  buf
  g1689
  (
    n1519,
    n366
  );


  not
  g1690
  (
    n536,
    n159
  );


  not
  g1691
  (
    n774,
    n456
  );


  not
  g1692
  (
    n715,
    n375
  );


  not
  g1693
  (
    n584,
    n279
  );


  buf
  g1694
  (
    n1186,
    n375
  );


  buf
  g1695
  (
    n1120,
    n454
  );


  not
  g1696
  (
    n569,
    n326
  );


  not
  g1697
  (
    n681,
    n315
  );


  buf
  g1698
  (
    n1043,
    n267
  );


  not
  g1699
  (
    n1699,
    n363
  );


  buf
  g1700
  (
    n837,
    n192
  );


  not
  g1701
  (
    n1076,
    n138
  );


  not
  g1702
  (
    n867,
    n271
  );


  not
  g1703
  (
    n1123,
    n304
  );


  buf
  g1704
  (
    n706,
    n386
  );


  nand
  g1705
  (
    n581,
    n162,
    n155,
    n245,
    n253
  );


  xnor
  g1706
  (
    n1116,
    n199,
    n291,
    n313,
    n420
  );


  or
  g1707
  (
    n868,
    n166,
    n322,
    n310,
    n249
  );


  and
  g1708
  (
    n564,
    n312,
    n160,
    n219,
    n398
  );


  xnor
  g1709
  (
    n1213,
    n247,
    n181,
    n202,
    n395
  );


  or
  g1710
  (
    n1207,
    n413,
    n364,
    n141,
    n192
  );


  nor
  g1711
  (
    n1482,
    n362,
    n338,
    n140,
    n395
  );


  xnor
  g1712
  (
    n923,
    n213,
    n347,
    n329,
    n187
  );


  xor
  g1713
  (
    n1074,
    n348,
    n380,
    n135,
    n213
  );


  or
  g1714
  (
    n601,
    n199,
    n235,
    n405,
    n434
  );


  and
  g1715
  (
    n621,
    n323,
    n423,
    n177,
    n276
  );


  nand
  g1716
  (
    n1141,
    n455,
    n297,
    n369,
    n296
  );


  or
  g1717
  (
    n2238,
    n1472,
    n1585,
    n1001,
    n845
  );


  nand
  g1718
  (
    n2256,
    n836,
    n482,
    n679,
    n882
  );


  or
  g1719
  (
    n1791,
    n1623,
    n1611,
    n1710,
    n1618
  );


  nor
  g1720
  (
    n2188,
    n1072,
    n1706,
    n861,
    n1456
  );


  xor
  g1721
  (
    n2348,
    n1140,
    n862,
    n1135,
    n1438
  );


  or
  g1722
  (
    n2416,
    n642,
    n522,
    n1579,
    n1244
  );


  nand
  g1723
  (
    n1768,
    n1445,
    n1241,
    n1108,
    n1179
  );


  xnor
  g1724
  (
    n2296,
    n1733,
    n1647,
    n1175,
    n1007
  );


  xnor
  g1725
  (
    n1985,
    n608,
    n1736,
    n1532,
    n1030
  );


  nand
  g1726
  (
    n2065,
    n533,
    n1009,
    n1365,
    n473
  );


  or
  g1727
  (
    n2066,
    n799,
    n1108,
    n1519,
    n568
  );


  nand
  g1728
  (
    n2428,
    n1694,
    n1595,
    n1419,
    n1593
  );


  xor
  g1729
  (
    n1848,
    n1597,
    n1511,
    n1447,
    n1719
  );


  nand
  g1730
  (
    n1999,
    n507,
    n1546,
    n1495,
    n1483
  );


  or
  g1731
  (
    n1808,
    n1458,
    n1367,
    n1579,
    n1592
  );


  nor
  g1732
  (
    n1824,
    n1632,
    n1431,
    n1002,
    n1437
  );


  and
  g1733
  (
    n2353,
    n828,
    n1122,
    n1455,
    n667
  );


  xor
  g1734
  (
    n1752,
    n118,
    n1024,
    n1354,
    n1154
  );


  nor
  g1735
  (
    n1872,
    n1405,
    n1436,
    n1418,
    n1068
  );


  and
  g1736
  (
    n1947,
    n1454,
    n880,
    n939,
    n1200
  );


  and
  g1737
  (
    n2490,
    n1320,
    n1164,
    n1070,
    n1635
  );


  xnor
  g1738
  (
    n2317,
    n1296,
    n1627,
    n846,
    n1696
  );


  xor
  g1739
  (
    n2278,
    n1508,
    n1371,
    n666,
    n755
  );


  xor
  g1740
  (
    n2447,
    n1203,
    n1554,
    n1578,
    n1351
  );


  or
  g1741
  (
    n2090,
    n1628,
    n985,
    n652,
    n1367
  );


  xor
  g1742
  (
    n2425,
    n1059,
    n1000,
    n772,
    n600
  );


  nor
  g1743
  (
    n2133,
    n1331,
    n1569,
    n1403,
    n1346
  );


  and
  g1744
  (
    n2089,
    n1494,
    n1123,
    n991,
    n1599
  );


  and
  g1745
  (
    n2212,
    n1067,
    n1265,
    n1111,
    n1256
  );


  nand
  g1746
  (
    n1760,
    n499,
    n1683,
    n1326,
    n526
  );


  nor
  g1747
  (
    n2041,
    n1079,
    n487,
    n1575,
    n1482
  );


  or
  g1748
  (
    n2149,
    n1674,
    n1534,
    n1488,
    n1088
  );


  and
  g1749
  (
    n2372,
    n1419,
    n1681,
    n668,
    n697
  );


  xor
  g1750
  (
    n2075,
    n1185,
    n1511,
    n1207,
    n1625
  );


  nand
  g1751
  (
    n1935,
    n905,
    n1405,
    n573,
    n921
  );


  or
  g1752
  (
    n2327,
    n515,
    n1656,
    n1345,
    n1230
  );


  nor
  g1753
  (
    n2032,
    n1180,
    n1605,
    n1091,
    n589
  );


  xor
  g1754
  (
    n1827,
    n1653,
    n1025,
    n674,
    n1644
  );


  nand
  g1755
  (
    n2034,
    n1333,
    n694,
    n713,
    n1178
  );


  xor
  g1756
  (
    n2030,
    n860,
    n1512,
    n1230,
    n1558
  );


  and
  g1757
  (
    n2422,
    n611,
    n1280,
    n1695,
    n1070
  );


  xor
  g1758
  (
    n1829,
    n1332,
    n1300,
    n1271,
    n1623
  );


  or
  g1759
  (
    n2499,
    n122,
    n1360,
    n1377,
    n834
  );


  and
  g1760
  (
    n2057,
    n1711,
    n1730,
    n1644,
    n689
  );


  nand
  g1761
  (
    n1860,
    n1658,
    n1684,
    n1378,
    n687
  );


  nand
  g1762
  (
    n1930,
    n1286,
    n1308,
    n1577,
    n719
  );


  xor
  g1763
  (
    n2087,
    n1370,
    n1290,
    n1408,
    n764
  );


  nor
  g1764
  (
    n2373,
    n1699,
    n121,
    n1028,
    n943
  );


  xnor
  g1765
  (
    n2001,
    n508,
    n1672,
    n1717,
    n1656
  );


  nor
  g1766
  (
    n1822,
    n766,
    n652,
    n572,
    n686
  );


  nand
  g1767
  (
    n2158,
    n527,
    n621,
    n1436,
    n1724
  );


  or
  g1768
  (
    n2292,
    n521,
    n1237,
    n1146,
    n117
  );


  or
  g1769
  (
    n2224,
    n593,
    n1497,
    n1642,
    n751
  );


  xnor
  g1770
  (
    n2011,
    n511,
    n1141,
    n485,
    n814
  );


  or
  g1771
  (
    n2421,
    n823,
    n1590,
    n1533,
    n1234
  );


  xnor
  g1772
  (
    n2022,
    n769,
    n1600,
    n1343,
    n1643
  );


  xnor
  g1773
  (
    n2406,
    n1215,
    n1708,
    n831,
    n1560
  );


  nor
  g1774
  (
    n1799,
    n1308,
    n1055,
    n1736,
    n1107
  );


  and
  g1775
  (
    n1987,
    n807,
    n1565,
    n1549,
    n1687
  );


  and
  g1776
  (
    n1815,
    n1543,
    n1435,
    n1235,
    n1507
  );


  nand
  g1777
  (
    n2398,
    n701,
    n497,
    n1310,
    n646
  );


  or
  g1778
  (
    n2483,
    n1182,
    n1223,
    n911,
    n1685
  );


  nand
  g1779
  (
    n2216,
    n558,
    n510,
    n1373,
    n1333
  );


  or
  g1780
  (
    n2247,
    n1574,
    n862,
    n1077,
    n1122
  );


  xor
  g1781
  (
    n2467,
    n1501,
    n727,
    n1663,
    n1173
  );


  xnor
  g1782
  (
    n2080,
    n934,
    n1349,
    n1402,
    n1464
  );


  xor
  g1783
  (
    n2272,
    n783,
    n495,
    n1017,
    n610
  );


  or
  g1784
  (
    n1883,
    n636,
    n1504,
    n866,
    n851
  );


  xnor
  g1785
  (
    n2309,
    n1010,
    n738,
    n1679,
    n949
  );


  xor
  g1786
  (
    n2246,
    n1712,
    n570,
    n124,
    n1137
  );


  and
  g1787
  (
    n2162,
    n615,
    n1532,
    n1411,
    n1516
  );


  xnor
  g1788
  (
    n2378,
    n1284,
    n544,
    n748,
    n1147
  );


  or
  g1789
  (
    n2319,
    n672,
    n1572,
    n741,
    n1571
  );


  or
  g1790
  (
    n2337,
    n826,
    n1255,
    n1666,
    n629
  );


  and
  g1791
  (
    n2314,
    n1256,
    n1671,
    n123,
    n654
  );


  and
  g1792
  (
    n1769,
    n1302,
    n1415,
    n1434,
    n1073
  );


  nor
  g1793
  (
    n2167,
    n1464,
    n1079,
    n562,
    n1530
  );


  and
  g1794
  (
    n1767,
    n1584,
    n117,
    n587,
    n1501
  );


  or
  g1795
  (
    n1776,
    n1589,
    n785,
    n120,
    n1632
  );


  nor
  g1796
  (
    n1846,
    n955,
    n1015,
    n871,
    n1378
  );


  and
  g1797
  (
    n2244,
    n1503,
    n1468,
    n545,
    n1094
  );


  nand
  g1798
  (
    n1979,
    n710,
    n1395,
    n1018,
    n823
  );


  nand
  g1799
  (
    n1803,
    n694,
    n1625,
    n1046,
    n1042
  );


  and
  g1800
  (
    n2449,
    n1655,
    n695,
    n1566,
    n1044
  );


  xor
  g1801
  (
    n2475,
    n502,
    n669,
    n1098,
    n1640
  );


  xor
  g1802
  (
    n2138,
    n1318,
    n522,
    n763,
    n516
  );


  and
  g1803
  (
    n2276,
    n682,
    n799,
    n118,
    n1461
  );


  xor
  g1804
  (
    n2484,
    n1527,
    n683,
    n495,
    n503
  );


  and
  g1805
  (
    n2488,
    n750,
    n1272,
    n541,
    n1282
  );


  or
  g1806
  (
    n1871,
    n916,
    n1658,
    n1369,
    n1313
  );


  nor
  g1807
  (
    n2496,
    n125,
    n548,
    n472,
    n1090
  );


  xnor
  g1808
  (
    n2443,
    n1497,
    n1295,
    n1731,
    n740
  );


  xor
  g1809
  (
    n1782,
    n1054,
    n1551,
    n1640,
    n1522
  );


  nand
  g1810
  (
    n2038,
    n529,
    n1679,
    n1506,
    n1257
  );


  xor
  g1811
  (
    n1789,
    n1110,
    n1306,
    n1395,
    n479
  );


  xnor
  g1812
  (
    n2286,
    n1319,
    n1651,
    n1610,
    n511
  );


  xnor
  g1813
  (
    n1939,
    n1526,
    n668,
    n1518,
    n1673
  );


  xnor
  g1814
  (
    n2017,
    n1637,
    n1324,
    n1075,
    n1532
  );


  xor
  g1815
  (
    n2052,
    n948,
    n975,
    n1083,
    n671
  );


  and
  g1816
  (
    n2086,
    n587,
    n1658,
    n1500,
    n1485
  );


  nand
  g1817
  (
    n2144,
    n1562,
    n1229,
    n491,
    n570
  );


  nor
  g1818
  (
    n2186,
    n512,
    n1310,
    n1707,
    n560
  );


  nand
  g1819
  (
    n1798,
    n1218,
    n1469,
    n123,
    n1715
  );


  xor
  g1820
  (
    n2179,
    n897,
    n947,
    n1688,
    n853
  );


  xor
  g1821
  (
    n1832,
    n1303,
    n801,
    n1565,
    n671
  );


  and
  g1822
  (
    n2503,
    n1556,
    n1287,
    n1709,
    n609
  );


  xnor
  g1823
  (
    n2344,
    n1691,
    n1112,
    n1423,
    n1630
  );


  nor
  g1824
  (
    n2438,
    n1174,
    n1594,
    n1184,
    n588
  );


  xor
  g1825
  (
    n1790,
    n1294,
    n673,
    n705,
    n1605
  );


  nand
  g1826
  (
    n2178,
    n1175,
    n1561,
    n526,
    n1483
  );


  nand
  g1827
  (
    n2334,
    n1339,
    n1213,
    n1553,
    n617
  );


  xnor
  g1828
  (
    n2318,
    n653,
    n630,
    n814,
    n1566
  );


  and
  g1829
  (
    n2287,
    n860,
    n1320,
    n528,
    n1704
  );


  and
  g1830
  (
    n1771,
    n1681,
    n1587,
    n507,
    n1693
  );


  xor
  g1831
  (
    n1854,
    n634,
    n1418,
    n542,
    n1685
  );


  nor
  g1832
  (
    n1925,
    n1295,
    n1277,
    n1570,
    n857
  );


  nand
  g1833
  (
    n1857,
    n662,
    n120,
    n1612,
    n1542
  );


  xnor
  g1834
  (
    n2120,
    n1431,
    n1441,
    n553,
    n1351
  );


  xnor
  g1835
  (
    n2199,
    n876,
    n632,
    n1380,
    n1446
  );


  nand
  g1836
  (
    n2050,
    n1294,
    n680,
    n1158,
    n942
  );


  xor
  g1837
  (
    n2265,
    n891,
    n1647,
    n1514,
    n1301
  );


  or
  g1838
  (
    n1775,
    n1202,
    n1386,
    n1332,
    n1606
  );


  xor
  g1839
  (
    n2331,
    n836,
    n1719,
    n653,
    n830
  );


  nand
  g1840
  (
    n2027,
    n1655,
    n1352,
    n533,
    n1735
  );


  xor
  g1841
  (
    n2401,
    n928,
    n584,
    n1299,
    n1181
  );


  and
  g1842
  (
    n2237,
    n471,
    n1553,
    n1649,
    n1484
  );


  or
  g1843
  (
    n1755,
    n1145,
    n1164,
    n1721,
    n1648
  );


  xor
  g1844
  (
    n2270,
    n916,
    n1491,
    n1707,
    n705
  );


  nand
  g1845
  (
    n1835,
    n1011,
    n503,
    n659,
    n1245
  );


  nand
  g1846
  (
    n1934,
    n490,
    n1540,
    n1355,
    n1132
  );


  xnor
  g1847
  (
    n2129,
    n1265,
    n1210,
    n628,
    n866
  );


  or
  g1848
  (
    n2448,
    n1349,
    n1522,
    n760,
    n1626
  );


  or
  g1849
  (
    n2194,
    n1169,
    n1104,
    n1358,
    n1505
  );


  nand
  g1850
  (
    n1788,
    n1243,
    n1031,
    n1654,
    n523
  );


  xnor
  g1851
  (
    n2501,
    n1336,
    n612,
    n625,
    n564
  );


  and
  g1852
  (
    n2409,
    n650,
    n1442,
    n614,
    n874
  );


  or
  g1853
  (
    n2157,
    n1692,
    n1094,
    n1733,
    n1689
  );


  xnor
  g1854
  (
    n2350,
    n1723,
    n1588,
    n970,
    n551
  );


  xnor
  g1855
  (
    n2143,
    n1450,
    n1596,
    n1688,
    n1400
  );


  nand
  g1856
  (
    n2431,
    n539,
    n1193,
    n1085,
    n709
  );


  xor
  g1857
  (
    n2035,
    n1466,
    n1668,
    n730,
    n687
  );


  xnor
  g1858
  (
    n2430,
    n877,
    n548,
    n599,
    n778
  );


  or
  g1859
  (
    n2232,
    n1168,
    n1605,
    n890,
    n1347
  );


  xor
  g1860
  (
    n1764,
    n987,
    n1571,
    n1249,
    n1408
  );


  nor
  g1861
  (
    n1965,
    n1700,
    n755,
    n1661,
    n675
  );


  xnor
  g1862
  (
    n2197,
    n1385,
    n1580,
    n1439,
    n517
  );


  or
  g1863
  (
    n2259,
    n1309,
    n1205,
    n767,
    n1376
  );


  nand
  g1864
  (
    n2081,
    n1334,
    n1686,
    n1065,
    n1630
  );


  nor
  g1865
  (
    n1904,
    n1629,
    n1248,
    n1642,
    n800
  );


  and
  g1866
  (
    n1864,
    n1534,
    n995,
    n1634,
    n1291
  );


  and
  g1867
  (
    n2083,
    n1445,
    n1214,
    n941,
    n1082
  );


  xor
  g1868
  (
    n1914,
    n1255,
    n1103,
    n837,
    n1462
  );


  xor
  g1869
  (
    n2055,
    n1466,
    n1575,
    n1306,
    n861
  );


  nor
  g1870
  (
    n1950,
    n1261,
    n1655,
    n1067,
    n610
  );


  xnor
  g1871
  (
    n2069,
    n1187,
    n1682,
    n603,
    n856
  );


  nor
  g1872
  (
    n1865,
    n1462,
    n1410,
    n994,
    n1369
  );


  xor
  g1873
  (
    n1858,
    n1499,
    n1358,
    n1257,
    n566
  );


  nand
  g1874
  (
    n2137,
    n1016,
    n644,
    n1385,
    n1622
  );


  and
  g1875
  (
    n2374,
    n752,
    n923,
    n1350,
    n1581
  );


  xnor
  g1876
  (
    n2504,
    n1512,
    n711,
    n1399,
    n927
  );


  xor
  g1877
  (
    n2367,
    n761,
    n1644,
    n983,
    n1202
  );


  and
  g1878
  (
    n2397,
    n1142,
    n488,
    n1377,
    n1567
  );


  nand
  g1879
  (
    n1876,
    n954,
    n1384,
    n1026,
    n901
  );


  nand
  g1880
  (
    n2347,
    n1420,
    n1515,
    n1176,
    n1403
  );


  xnor
  g1881
  (
    n2400,
    n1387,
    n573,
    n1504,
    n1649
  );


  xor
  g1882
  (
    n2067,
    n1454,
    n1475,
    n1602,
    n1559
  );


  nand
  g1883
  (
    n1792,
    n693,
    n1100,
    n1339,
    n602
  );


  and
  g1884
  (
    n2062,
    n1544,
    n1432,
    n1704,
    n751
  );


  nand
  g1885
  (
    n2285,
    n1628,
    n1360,
    n1492,
    n1000
  );


  nand
  g1886
  (
    n2248,
    n724,
    n1698,
    n884,
    n987
  );


  and
  g1887
  (
    n2181,
    n1435,
    n1390,
    n549,
    n1624
  );


  nor
  g1888
  (
    n2392,
    n576,
    n1362,
    n840,
    n802
  );


  xnor
  g1889
  (
    n1875,
    n1668,
    n1287,
    n1415,
    n713
  );


  xor
  g1890
  (
    n2171,
    n1307,
    n1497,
    n117,
    n1047
  );


  nand
  g1891
  (
    n1919,
    n1023,
    n722,
    n1087,
    n1625
  );


  xnor
  g1892
  (
    n2176,
    n1168,
    n1238,
    n1159,
    n1711
  );


  nand
  g1893
  (
    n2415,
    n1240,
    n1667,
    n787,
    n1152
  );


  and
  g1894
  (
    n2433,
    n1433,
    n737,
    n1700,
    n1061
  );


  nor
  g1895
  (
    n2105,
    n496,
    n1113,
    n1650,
    n519
  );


  xnor
  g1896
  (
    n1915,
    n1105,
    n1038,
    n606,
    n1279
  );


  and
  g1897
  (
    n2380,
    n1388,
    n1051,
    n971,
    n1432
  );


  and
  g1898
  (
    n1809,
    n1467,
    n670,
    n1269,
    n1309
  );


  nor
  g1899
  (
    n1825,
    n1728,
    n480,
    n605,
    n1463
  );


  and
  g1900
  (
    n2304,
    n1192,
    n1084,
    n1509,
    n1447
  );


  xnor
  g1901
  (
    n2210,
    n918,
    n1552,
    n857,
    n1071
  );


  nand
  g1902
  (
    n2354,
    n740,
    n886,
    n1374,
    n859
  );


  nand
  g1903
  (
    n2349,
    n909,
    n1721,
    n1665,
    n1688
  );


  xor
  g1904
  (
    n1820,
    n715,
    n1363,
    n1710,
    n1336
  );


  xor
  g1905
  (
    n2366,
    n556,
    n725,
    n747,
    n492
  );


  xor
  g1906
  (
    n2469,
    n1172,
    n1429,
    n1463,
    n516
  );


  nor
  g1907
  (
    n1795,
    n784,
    n1614,
    n1429,
    n566
  );


  xor
  g1908
  (
    n2170,
    n986,
    n476,
    n521,
    n746
  );


  or
  g1909
  (
    n1960,
    n1645,
    n1721,
    n885,
    n1473
  );


  nor
  g1910
  (
    n1772,
    n842,
    n1672,
    n647,
    n1557
  );


  xor
  g1911
  (
    n2260,
    n1027,
    n1099,
    n1434,
    n1357
  );


  or
  g1912
  (
    n2436,
    n1297,
    n1061,
    n896,
    n501
  );


  and
  g1913
  (
    n1982,
    n493,
    n1726,
    n1599,
    n1320
  );


  nor
  g1914
  (
    n2111,
    n1338,
    n730,
    n1327,
    n748
  );


  xor
  g1915
  (
    n1951,
    n1125,
    n749,
    n887,
    n732
  );


  nand
  g1916
  (
    n2126,
    n1428,
    n912,
    n945,
    n119
  );


  xor
  g1917
  (
    n2253,
    n942,
    n475,
    n1539,
    n117
  );


  and
  g1918
  (
    n1912,
    n1155,
    n1323,
    n1093,
    n1697
  );


  nor
  g1919
  (
    n1845,
    n1397,
    n878,
    n1132,
    n1578
  );


  nor
  g1920
  (
    n2071,
    n1521,
    n886,
    n695,
    n1391
  );


  and
  g1921
  (
    n2115,
    n1160,
    n1670,
    n810,
    n1404
  );


  nand
  g1922
  (
    n1969,
    n1054,
    n1685,
    n657,
    n821
  );


  xor
  g1923
  (
    n2320,
    n1314,
    n514,
    n905,
    n1553
  );


  nor
  g1924
  (
    n2482,
    n1347,
    n591,
    n1299,
    n514
  );


  xor
  g1925
  (
    n2487,
    n953,
    n763,
    n1595,
    n535
  );


  xor
  g1926
  (
    n2472,
    n509,
    n1558,
    n1523,
    n982
  );


  xor
  g1927
  (
    n2474,
    n578,
    n677,
    n567,
    n1425
  );


  xnor
  g1928
  (
    n1765,
    n1174,
    n731,
    n1615,
    n969
  );


  nand
  g1929
  (
    n2339,
    n699,
    n1348,
    n1472,
    n1562
  );


  and
  g1930
  (
    n2355,
    n800,
    n777,
    n1628,
    n593
  );


  xor
  g1931
  (
    n2411,
    n1353,
    n1001,
    n1178,
    n1201
  );


  xnor
  g1932
  (
    n2413,
    n1305,
    n791,
    n592,
    n122
  );


  nand
  g1933
  (
    n2209,
    n1356,
    n833,
    n1365,
    n769
  );


  xnor
  g1934
  (
    n2236,
    n1547,
    n1357,
    n988,
    n1713
  );


  or
  g1935
  (
    n2310,
    n1563,
    n1069,
    n947,
    n835
  );


  xor
  g1936
  (
    n1866,
    n662,
    n1595,
    n1270,
    n1474
  );


  and
  g1937
  (
    n1888,
    n1592,
    n1292,
    n1236,
    n676
  );


  xnor
  g1938
  (
    n1787,
    n1518,
    n808,
    n762,
    n1247
  );


  nand
  g1939
  (
    n1842,
    n1264,
    n1151,
    n1014,
    n1536
  );


  xor
  g1940
  (
    n1781,
    n794,
    n1449,
    n910,
    n568
  );


  xor
  g1941
  (
    n2121,
    n119,
    n619,
    n1686,
    n591
  );


  nand
  g1942
  (
    n1936,
    n494,
    n858,
    n1198,
    n1566
  );


  nor
  g1943
  (
    n2442,
    n898,
    n896,
    n1130,
    n1527
  );


  xnor
  g1944
  (
    n2031,
    n1500,
    n1697,
    n931,
    n1418
  );


  xnor
  g1945
  (
    n2103,
    n1714,
    n1233,
    n1126,
    n569
  );


  or
  g1946
  (
    n2219,
    n1386,
    n1552,
    n1361,
    n1078
  );


  nand
  g1947
  (
    n2006,
    n579,
    n834,
    n1607,
    n923
  );


  xnor
  g1948
  (
    n2136,
    n1017,
    n899,
    n571,
    n1120
  );


  nor
  g1949
  (
    n2116,
    n996,
    n1382,
    n875,
    n1121
  );


  xnor
  g1950
  (
    n2377,
    n704,
    n1543,
    n1496,
    n482
  );


  or
  g1951
  (
    n1924,
    n624,
    n1428,
    n603,
    n735
  );


  or
  g1952
  (
    n2018,
    n1508,
    n1268,
    n1010,
    n1224
  );


  and
  g1953
  (
    n2315,
    n1417,
    n1416,
    n1376,
    n1120
  );


  nand
  g1954
  (
    n2000,
    n598,
    n1593,
    n1267,
    n1664
  );


  xnor
  g1955
  (
    n2257,
    n1493,
    n919,
    n1488,
    n762
  );


  xnor
  g1956
  (
    n1953,
    n813,
    n914,
    n756,
    n1211
  );


  nand
  g1957
  (
    n2266,
    n1629,
    n790,
    n1457,
    n1656
  );


  nand
  g1958
  (
    n1761,
    n1144,
    n1583,
    n543,
    n984
  );


  nor
  g1959
  (
    n1773,
    n791,
    n1633,
    n972,
    n502
  );


  xnor
  g1960
  (
    n2332,
    n1409,
    n564,
    n636,
    n1027
  );


  xor
  g1961
  (
    n2385,
    n1725,
    n1691,
    n1616,
    n1545
  );


  or
  g1962
  (
    n2074,
    n586,
    n1636,
    n1124,
    n1171
  );


  xor
  g1963
  (
    n1874,
    n1391,
    n1337,
    n882,
    n731
  );


  nand
  g1964
  (
    n1834,
    n1576,
    n582,
    n1706,
    n1183
  );


  nand
  g1965
  (
    n2420,
    n1192,
    n1528,
    n1285,
    n899
  );


  or
  g1966
  (
    n2214,
    n1637,
    n870,
    n1613,
    n669
  );


  xnor
  g1967
  (
    n2383,
    n688,
    n580,
    n760,
    n1332
  );


  nor
  g1968
  (
    n1908,
    n1322,
    n569,
    n1167,
    n1735
  );


  xnor
  g1969
  (
    n2311,
    n818,
    n752,
    n865,
    n1529
  );


  nand
  g1970
  (
    n1911,
    n1049,
    n527,
    n918,
    n1460
  );


  xnor
  g1971
  (
    n2451,
    n1732,
    n1499,
    n1086,
    n933
  );


  xor
  g1972
  (
    n2299,
    n598,
    n966,
    n1643,
    n1468
  );


  nor
  g1973
  (
    n2019,
    n776,
    n1024,
    n1050,
    n1264
  );


  or
  g1974
  (
    n2231,
    n910,
    n1066,
    n1515,
    n508
  );


  xor
  g1975
  (
    n2132,
    n1341,
    n1568,
    n1506,
    n1103
  );


  xor
  g1976
  (
    n2279,
    n1583,
    n1641,
    n1166,
    n1706
  );


  nor
  g1977
  (
    n1971,
    n595,
    n532,
    n820,
    n807
  );


  nand
  g1978
  (
    n2289,
    n1261,
    n1716,
    n660,
    n883
  );


  and
  g1979
  (
    n2282,
    n1482,
    n1232,
    n1351,
    n1314
  );


  xor
  g1980
  (
    n2072,
    n594,
    n1116,
    n504,
    n1219
  );


  or
  g1981
  (
    n1821,
    n1399,
    n1235,
    n989,
    n1215
  );


  xor
  g1982
  (
    n2437,
    n524,
    n1335,
    n1580,
    n1346
  );


  and
  g1983
  (
    n2059,
    n517,
    n1728,
    n765,
    n871
  );


  nor
  g1984
  (
    n1972,
    n1528,
    n1325,
    n584,
    n720
  );


  and
  g1985
  (
    n2432,
    n489,
    n825,
    n1570,
    n1305
  );


  nand
  g1986
  (
    n2131,
    n902,
    n1555,
    n1646,
    n1328
  );


  xor
  g1987
  (
    n2417,
    n1277,
    n1727,
    n781,
    n1053
  );


  xnor
  g1988
  (
    n2439,
    n619,
    n1626,
    n843,
    n1121
  );


  xnor
  g1989
  (
    n1779,
    n1156,
    n690,
    n868,
    n952
  );


  and
  g1990
  (
    n2024,
    n1596,
    n497,
    n602,
    n1162
  );


  nand
  g1991
  (
    n2396,
    n1560,
    n1325,
    n1396,
    n1018
  );


  xor
  g1992
  (
    n1836,
    n691,
    n1483,
    n989,
    n1204
  );


  or
  g1993
  (
    n2140,
    n709,
    n792,
    n1300,
    n902
  );


  xor
  g1994
  (
    n1956,
    n492,
    n1680,
    n1578,
    n475
  );


  nand
  g1995
  (
    n2096,
    n499,
    n1660,
    n661,
    n1398
  );


  nor
  g1996
  (
    n1754,
    n571,
    n775,
    n917,
    n1705
  );


  xnor
  g1997
  (
    n1870,
    n1341,
    n805,
    n1695,
    n1288
  );


  nor
  g1998
  (
    n2164,
    n950,
    n781,
    n782,
    n1638
  );


  xor
  g1999
  (
    n2012,
    n1034,
    n486,
    n1041,
    n733
  );


  xnor
  g2000
  (
    n2056,
    n1674,
    n1324,
    n125,
    n1333
  );


  nor
  g2001
  (
    n2303,
    n1274,
    n1448,
    n1237,
    n1506
  );


  xor
  g2002
  (
    n2395,
    n1669,
    n1304,
    n655,
    n829
  );


  xor
  g2003
  (
    n2127,
    n1356,
    n1099,
    n1315,
    n703
  );


  nand
  g2004
  (
    n1900,
    n1081,
    n1157,
    n1670,
    n959
  );


  and
  g2005
  (
    n1796,
    n1240,
    n1654,
    n1690,
    n1299
  );


  and
  g2006
  (
    n2245,
    n903,
    n934,
    n716,
    n1577
  );


  xor
  g2007
  (
    n2414,
    n1155,
    n1372,
    n540,
    n1130
  );


  xnor
  g2008
  (
    n2091,
    n666,
    n1385,
    n1557,
    n869
  );


  or
  g2009
  (
    n2283,
    n1653,
    n819,
    n1430,
    n734
  );


  and
  g2010
  (
    n2180,
    n562,
    n674,
    n1065,
    n484
  );


  xnor
  g2011
  (
    n2375,
    n1344,
    n952,
    n1379,
    n1085
  );


  nand
  g2012
  (
    n2284,
    n1450,
    n1726,
    n567,
    n1279
  );


  or
  g2013
  (
    n1981,
    n956,
    n1443,
    n1186,
    n1305
  );


  xnor
  g2014
  (
    n2393,
    n1725,
    n1565,
    n1118,
    n491
  );


  xnor
  g2015
  (
    n1996,
    n1602,
    n1285,
    n1530,
    n1220
  );


  and
  g2016
  (
    n1817,
    n1004,
    n1307,
    n1037,
    n931
  );


  nand
  g2017
  (
    n2163,
    n632,
    n1633,
    n935,
    n785
  );


  or
  g2018
  (
    n2218,
    n793,
    n1158,
    n1639,
    n1543
  );


  nand
  g2019
  (
    n1927,
    n1645,
    n718,
    n1547,
    n1668
  );


  and
  g2020
  (
    n2093,
    n1200,
    n1689,
    n855,
    n1567
  );


  nor
  g2021
  (
    n1920,
    n945,
    n1225,
    n1614,
    n1449
  );


  xnor
  g2022
  (
    n1833,
    n936,
    n1469,
    n1702,
    n618
  );


  xnor
  g2023
  (
    n2147,
    n831,
    n924,
    n913,
    n978
  );


  nor
  g2024
  (
    n2429,
    n1275,
    n1369,
    n608,
    n1530
  );


  xnor
  g2025
  (
    n1995,
    n1450,
    n1699,
    n816,
    n1515
  );


  xnor
  g2026
  (
    n1963,
    n756,
    n1584,
    n951,
    n630
  );


  nand
  g2027
  (
    n2346,
    n920,
    n1336,
    n1630,
    n1446
  );


  nor
  g2028
  (
    n1784,
    n1056,
    n1426,
    n1216,
    n1344
  );


  xnor
  g2029
  (
    n2039,
    n1455,
    n596,
    n1063,
    n1493
  );


  nor
  g2030
  (
    n2128,
    n1598,
    n1241,
    n938,
    n1083
  );


  xor
  g2031
  (
    n2407,
    n1338,
    n667,
    n1196,
    n1505
  );


  and
  g2032
  (
    n1991,
    n1129,
    n1477,
    n1550,
    n1609
  );


  nand
  g2033
  (
    n1998,
    n1647,
    n1621,
    n933,
    n1128
  );


  xnor
  g2034
  (
    n1837,
    n665,
    n914,
    n1294,
    n1680
  );


  nor
  g2035
  (
    n2049,
    n1041,
    n645,
    n1291,
    n513
  );


  xnor
  g2036
  (
    n2381,
    n922,
    n528,
    n1150,
    n1189
  );


  xnor
  g2037
  (
    n2312,
    n710,
    n1334,
    n1159,
    n786
  );


  and
  g2038
  (
    n2301,
    n1572,
    n1347,
    n1631,
    n1489
  );


  or
  g2039
  (
    n2227,
    n1293,
    n1594,
    n1393,
    n993
  );


  xor
  g2040
  (
    n1944,
    n749,
    n513,
    n1603,
    n876
  );


  xor
  g2041
  (
    n2264,
    n848,
    n1413,
    n1546,
    n725
  );


  nor
  g2042
  (
    n1763,
    n736,
    n1443,
    n950,
    n605
  );


  xor
  g2043
  (
    n2338,
    n1478,
    n838,
    n868,
    n1639
  );


  and
  g2044
  (
    n2046,
    n775,
    n1429,
    n758,
    n1062
  );


  nor
  g2045
  (
    n2169,
    n885,
    n1195,
    n1290,
    n1406
  );


  xor
  g2046
  (
    n2365,
    n677,
    n811,
    n765,
    n796
  );


  xnor
  g2047
  (
    n2241,
    n1587,
    n743,
    n1480,
    n770
  );


  and
  g2048
  (
    n1994,
    n477,
    n1636,
    n937,
    n1508
  );


  nor
  g2049
  (
    n1898,
    n1525,
    n505,
    n1066,
    n1229
  );


  xor
  g2050
  (
    n1948,
    n726,
    n1153,
    n964,
    n1081
  );


  nor
  g2051
  (
    n2277,
    n1687,
    n849,
    n1715,
    n1610
  );


  xnor
  g2052
  (
    n2003,
    n833,
    n1434,
    n1096,
    n1600
  );


  xnor
  g2053
  (
    n2165,
    n941,
    n1113,
    n770,
    n1245
  );


  xor
  g2054
  (
    n2053,
    n1731,
    n1254,
    n572,
    n474
  );


  nand
  g2055
  (
    n2104,
    n1252,
    n1102,
    n1273,
    n1048
  );


  and
  g2056
  (
    n2119,
    n722,
    n547,
    n1364,
    n1660
  );


  or
  g2057
  (
    n1885,
    n1400,
    n1278,
    n1105,
    n1258
  );


  or
  g2058
  (
    n2193,
    n1636,
    n745,
    n1720,
    n1502
  );


  xnor
  g2059
  (
    n1861,
    n821,
    n1626,
    n1139,
    n639
  );


  or
  g2060
  (
    n2117,
    n1437,
    n927,
    n1542,
    n1672
  );


  and
  g2061
  (
    n2010,
    n1262,
    n1169,
    n979,
    n1381
  );


  and
  g2062
  (
    n2150,
    n881,
    n1696,
    n1280,
    n637
  );


  xor
  g2063
  (
    n2084,
    n1150,
    n692,
    n1641,
    n911
  );


  and
  g2064
  (
    n1831,
    n1502,
    n1538,
    n122,
    n124
  );


  or
  g2065
  (
    n2462,
    n1661,
    n697,
    n1712,
    n1408
  );


  xor
  g2066
  (
    n2368,
    n1708,
    n574,
    n808,
    n841
  );


  and
  g2067
  (
    n2445,
    n1424,
    n1589,
    n1303,
    n537
  );


  xnor
  g2068
  (
    n2328,
    n1492,
    n1292,
    n1002,
    n1317
  );


  xor
  g2069
  (
    n2008,
    n811,
    n1484,
    n555,
    n1163
  );


  nor
  g2070
  (
    n1910,
    n1601,
    n538,
    n878,
    n729
  );


  and
  g2071
  (
    n2228,
    n1249,
    n1734,
    n1703,
    n779
  );


  nor
  g2072
  (
    n1749,
    n1032,
    n1214,
    n604,
    n720
  );


  nand
  g2073
  (
    n2110,
    n1504,
    n827,
    n574,
    n1708
  );


  and
  g2074
  (
    n2047,
    n840,
    n469,
    n1188,
    n1284
  );


  or
  g2075
  (
    n2343,
    n948,
    n1125,
    n1384,
    n1520
  );


  xor
  g2076
  (
    n2048,
    n1667,
    n739,
    n999,
    n1580
  );


  nand
  g2077
  (
    n2118,
    n1574,
    n534,
    n1381,
    n581
  );


  and
  g2078
  (
    n2426,
    n1128,
    n1564,
    n116,
    n745
  );


  xnor
  g2079
  (
    n1880,
    n1665,
    n1541,
    n1597,
    n778
  );


  nor
  g2080
  (
    n1891,
    n536,
    n1119,
    n965,
    n974
  );


  and
  g2081
  (
    n2456,
    n1452,
    n505,
    n1470,
    n1110
  );


  or
  g2082
  (
    n1753,
    n1194,
    n1623,
    n1162,
    n889
  );


  nand
  g2083
  (
    n2242,
    n1126,
    n1013,
    n1288,
    n664
  );


  and
  g2084
  (
    n1955,
    n1714,
    n1362,
    n1498,
    n1263
  );


  nand
  g2085
  (
    n2106,
    n692,
    n1520,
    n1262,
    n1682
  );


  and
  g2086
  (
    n2026,
    n1337,
    n771,
    n663,
    n1693
  );


  or
  g2087
  (
    n2423,
    n515,
    n531,
    n1585,
    n1491
  );


  and
  g2088
  (
    n2098,
    n539,
    n1223,
    n1109,
    n753
  );


  xnor
  g2089
  (
    n2330,
    n1422,
    n1107,
    n1638,
    n971
  );


  or
  g2090
  (
    n1945,
    n1451,
    n641,
    n622,
    n1289
  );


  and
  g2091
  (
    n2495,
    n1031,
    n1260,
    n1469,
    n1561
  );


  nor
  g2092
  (
    n2229,
    n1253,
    n1433,
    n532,
    n890
  );


  xnor
  g2093
  (
    n2094,
    n901,
    n1058,
    n1682,
    n1258
  );


  or
  g2094
  (
    n2280,
    n1377,
    n1331,
    n1452,
    n768
  );


  and
  g2095
  (
    n2427,
    n777,
    n1293,
    n1479,
    n1275
  );


  xor
  g2096
  (
    n1942,
    n1590,
    n1387,
    n1276,
    n1040
  );


  nand
  g2097
  (
    n2435,
    n1650,
    n966,
    n1293,
    n928
  );


  nand
  g2098
  (
    n2300,
    n483,
    n480,
    n1486,
    n921
  );


  xnor
  g2099
  (
    n2016,
    n1300,
    n1567,
    n1454,
    n698
  );


  and
  g2100
  (
    n2183,
    n718,
    n1392,
    n743,
    n1475
  );


  or
  g2101
  (
    n1964,
    n1152,
    n810,
    n1403,
    n559
  );


  xnor
  g2102
  (
    n2113,
    n721,
    n1345,
    n723,
    n1572
  );


  nand
  g2103
  (
    n1800,
    n917,
    n707,
    n1290,
    n1441
  );


  xnor
  g2104
  (
    n2302,
    n1665,
    n1671,
    n535,
    n550
  );


  nand
  g2105
  (
    n2079,
    n926,
    n1422,
    n1640,
    n1517
  );


  or
  g2106
  (
    n2042,
    n1095,
    n1562,
    n1394,
    n759
  );


  nor
  g2107
  (
    n1946,
    n1193,
    n1516,
    n1116,
    n1022
  );


  xnor
  g2108
  (
    n1884,
    n1694,
    n1680,
    n1146,
    n494
  );


  nand
  g2109
  (
    n2271,
    n1563,
    n1349,
    n883,
    n1129
  );


  or
  g2110
  (
    n1777,
    n469,
    n1423,
    n1496,
    n1524
  );


  xor
  g2111
  (
    n1859,
    n1607,
    n1003,
    n651,
    n622
  );


  xnor
  g2112
  (
    n2267,
    n626,
    n1513,
    n1365,
    n754
  );


  nor
  g2113
  (
    n2268,
    n1522,
    n1317,
    n1043,
    n1398
  );


  xnor
  g2114
  (
    n2198,
    n520,
    n870,
    n1576,
    n1327
  );


  xor
  g2115
  (
    n1938,
    n738,
    n1477,
    n1324,
    n498
  );


  and
  g2116
  (
    n2088,
    n1025,
    n804,
    n1371,
    n1573
  );


  nand
  g2117
  (
    n2250,
    n1700,
    n1143,
    n1693,
    n1555
  );


  xor
  g2118
  (
    n2470,
    n977,
    n856,
    n1692,
    n1191
  );


  or
  g2119
  (
    n2481,
    n1526,
    n863,
    n1205,
    n767
  );


  and
  g2120
  (
    n2351,
    n1510,
    n1465,
    n1537,
    n123
  );


  and
  g2121
  (
    n2294,
    n651,
    n1727,
    n1555,
    n1535
  );


  nor
  g2122
  (
    n2340,
    n1318,
    n1716,
    n1076,
    n1250
  );


  nand
  g2123
  (
    n1895,
    n1705,
    n1392,
    n643,
    n1427
  );


  and
  g2124
  (
    n2243,
    n963,
    n1545,
    n592,
    n1052
  );


  nand
  g2125
  (
    n2187,
    n504,
    n1195,
    n1380,
    n1359
  );


  nor
  g2126
  (
    n2155,
    n937,
    n1702,
    n545,
    n536
  );


  nand
  g2127
  (
    n2015,
    n1673,
    n1514,
    n633,
    n1196
  );


  nand
  g2128
  (
    n2073,
    n1427,
    n1319,
    n1494,
    n801
  );


  or
  g2129
  (
    n2389,
    n798,
    n1425,
    n1104,
    n546
  );


  nor
  g2130
  (
    n2200,
    n1165,
    n1609,
    n583,
    n1641
  );


  xnor
  g2131
  (
    n1869,
    n1453,
    n1424,
    n1490,
    n1092
  );


  nand
  g2132
  (
    n2493,
    n1171,
    n1463,
    n712,
    n1343
  );


  xnor
  g2133
  (
    n2263,
    n544,
    n1419,
    n1352,
    n1068
  );


  nand
  g2134
  (
    n2384,
    n1579,
    n120,
    n1045,
    n1516
  );


  or
  g2135
  (
    n2142,
    n579,
    n506,
    n1321,
    n1352
  );


  and
  g2136
  (
    n2325,
    n708,
    n1639,
    n1711,
    n621
  );


  nor
  g2137
  (
    n2100,
    n1021,
    n1101,
    n1209,
    n1662
  );


  xnor
  g2138
  (
    n2473,
    n830,
    n949,
    n698,
    n1381
  );


  nor
  g2139
  (
    n1810,
    n1619,
    n1540,
    n1734,
    n1531
  );


  nand
  g2140
  (
    n2480,
    n1611,
    n696,
    n1425,
    n873
  );


  or
  g2141
  (
    n1983,
    n869,
    n1617,
    n1312,
    n1533
  );


  xnor
  g2142
  (
    n2233,
    n1476,
    n702,
    n685,
    n796
  );


  nand
  g2143
  (
    n1819,
    n1007,
    n1718,
    n553,
    n472
  );


  xor
  g2144
  (
    n2387,
    n716,
    n1153,
    n1412,
    n1390
  );


  nand
  g2145
  (
    n1806,
    n1470,
    n124,
    n1723,
    n1701
  );


  or
  g2146
  (
    n1780,
    n663,
    n1474,
    n585,
    n122
  );


  xor
  g2147
  (
    n2261,
    n1729,
    n1370,
    n547,
    n552
  );


  nand
  g2148
  (
    n2102,
    n1503,
    n1142,
    n907,
    n922
  );


  xor
  g2149
  (
    n2321,
    n819,
    n1677,
    n1398,
    n1048
  );


  nand
  g2150
  (
    n2082,
    n696,
    n1589,
    n1303,
    n1675
  );


  nand
  g2151
  (
    n2173,
    n1709,
    n1486,
    n970,
    n1549
  );


  xor
  g2152
  (
    n2491,
    n1326,
    n1076,
    n1732,
    n795
  );


  xor
  g2153
  (
    n2063,
    n1676,
    n1436,
    n967,
    n631
  );


  nand
  g2154
  (
    n1882,
    n501,
    n1075,
    n1435,
    n1388
  );


  xnor
  g2155
  (
    n1758,
    n559,
    n1393,
    n1499,
    n973
  );


  nand
  g2156
  (
    n2500,
    n1670,
    n1354,
    n1021,
    n1131
  );


  xor
  g2157
  (
    n2444,
    n1495,
    n982,
    n481,
    n1051
  );


  xor
  g2158
  (
    n1847,
    n1667,
    n1047,
    n640,
    n590
  );


  xor
  g2159
  (
    n2450,
    n1380,
    n1611,
    n1593,
    n1063
  );


  nand
  g2160
  (
    n1762,
    n1344,
    n1696,
    n1161,
    n1720
  );


  xnor
  g2161
  (
    n2465,
    n670,
    n824,
    n1426,
    n1559
  );


  nor
  g2162
  (
    n2434,
    n1109,
    n1465,
    n1619,
    n742
  );


  and
  g2163
  (
    n2021,
    n1340,
    n1073,
    n1267,
    n1722
  );


  xnor
  g2164
  (
    n2044,
    n581,
    n1296,
    n483,
    n1413
  );


  nor
  g2165
  (
    n2281,
    n1106,
    n1471,
    n1493,
    n474
  );


  and
  g2166
  (
    n2306,
    n732,
    n1131,
    n1617,
    n1701
  );


  and
  g2167
  (
    n2020,
    n1674,
    n1343,
    n1224,
    n893
  );


  nand
  g2168
  (
    n2002,
    n1401,
    n842,
    n1615,
    n647
  );


  nor
  g2169
  (
    n2004,
    n477,
    n1359,
    n1028,
    n721
  );


  nor
  g2170
  (
    n2478,
    n655,
    n1420,
    n940,
    n894
  );


  xor
  g2171
  (
    n2399,
    n959,
    n589,
    n1198,
    n906
  );


  nor
  g2172
  (
    n1828,
    n1004,
    n805,
    n1561,
    n529
  );


  xor
  g2173
  (
    n2092,
    n1568,
    n1368,
    n963,
    n1100
  );


  and
  g2174
  (
    n2486,
    n485,
    n703,
    n1723,
    n1374
  );


  xor
  g2175
  (
    n2097,
    n1554,
    n1715,
    n616,
    n1481
  );


  xor
  g2176
  (
    n1826,
    n595,
    n711,
    n607,
    n1458
  );


  nand
  g2177
  (
    n1878,
    n1328,
    n1404,
    n665,
    n1587
  );


  nand
  g2178
  (
    n1807,
    n1586,
    n1598,
    n1545,
    n1057
  );


  nor
  g2179
  (
    n1850,
    n1127,
    n124,
    n1559,
    n1646
  );


  or
  g2180
  (
    n2252,
    n798,
    n1087,
    n1728,
    n1414
  );


  xnor
  g2181
  (
    n1756,
    n1372,
    n1537,
    n1394,
    n1102
  );


  nand
  g2182
  (
    n2151,
    n484,
    n1445,
    n116,
    n1362
  );


  or
  g2183
  (
    n1967,
    n1447,
    n1368,
    n1317,
    n1428
  );


  nor
  g2184
  (
    n2419,
    n1439,
    n1417,
    n1112,
    n1480
  );


  or
  g2185
  (
    n2208,
    n978,
    n1474,
    n1157,
    n633
  );


  nor
  g2186
  (
    n2145,
    n1325,
    n1395,
    n980,
    n1213
  );


  and
  g2187
  (
    n2364,
    n1009,
    n1228,
    n999,
    n1691
  );


  nor
  g2188
  (
    n1851,
    n1311,
    n623,
    n1232,
    n1315
  );


  or
  g2189
  (
    n2440,
    n1712,
    n1383,
    n1323,
    n609
  );


  nor
  g2190
  (
    n2077,
    n968,
    n1714,
    n620,
    n1448
  );


  xor
  g2191
  (
    n2184,
    n1629,
    n1226,
    n1577,
    n719
  );


  or
  g2192
  (
    n1954,
    n1620,
    n812,
    n1487,
    n1588
  );


  or
  g2193
  (
    n1868,
    n1727,
    n974,
    n1039,
    n973
  );


  nor
  g2194
  (
    n2477,
    n604,
    n975,
    n1564,
    n759
  );


  nor
  g2195
  (
    n2391,
    n1676,
    n1534,
    n1089,
    n1350
  );


  or
  g2196
  (
    n2037,
    n1618,
    n1302,
    n1481,
    n1149
  );


  xnor
  g2197
  (
    n2479,
    n900,
    n1523,
    n1659,
    n1206
  );


  xor
  g2198
  (
    n2471,
    n997,
    n804,
    n1342,
    n849
  );


  or
  g2199
  (
    n2174,
    n520,
    n802,
    n1456,
    n837
  );


  or
  g2200
  (
    n2109,
    n1111,
    n1459,
    n1458,
    n1539
  );


  xnor
  g2201
  (
    n1959,
    n891,
    n649,
    n1335,
    n844
  );


  nor
  g2202
  (
    n2005,
    n1509,
    n1319,
    n1594,
    n1627
  );


  xnor
  g2203
  (
    n2489,
    n1062,
    n606,
    n854,
    n1308
  );


  xnor
  g2204
  (
    n2189,
    n1190,
    n1657,
    n757,
    n1652
  );


  xor
  g2205
  (
    n2297,
    n1476,
    n614,
    n846,
    n996
  );


  xor
  g2206
  (
    n1881,
    n1342,
    n1117,
    n1368,
    n627
  );


  or
  g2207
  (
    n1748,
    n640,
    n1659,
    n1621,
    n1525
  );


  or
  g2208
  (
    n2191,
    n586,
    n1234,
    n1203,
    n481
  );


  xnor
  g2209
  (
    n2206,
    n1401,
    n618,
    n1217,
    n1355
  );


  or
  g2210
  (
    n2223,
    n1648,
    n1564,
    n1383,
    n1052
  );


  nor
  g2211
  (
    n2101,
    n1238,
    n1244,
    n1459,
    n867
  );


  nand
  g2212
  (
    n1839,
    n1375,
    n969,
    n1340,
    n1233
  );


  and
  g2213
  (
    n1966,
    n1248,
    n1673,
    n1634,
    n939
  );


  xnor
  g2214
  (
    n2459,
    n542,
    n997,
    n844,
    n852
  );


  or
  g2215
  (
    n1793,
    n1250,
    n707,
    n1729,
    n956
  );


  and
  g2216
  (
    n1990,
    n684,
    n1273,
    n693,
    n957
  );


  or
  g2217
  (
    n2226,
    n597,
    n1502,
    n1071,
    n1731
  );


  nor
  g2218
  (
    n1786,
    n1414,
    n1638,
    n806,
    n648
  );


  and
  g2219
  (
    n2195,
    n1520,
    n1652,
    n624,
    n1389
  );


  or
  g2220
  (
    n1941,
    n1199,
    n1379,
    n894,
    n1514
  );


  xor
  g2221
  (
    n2403,
    n1511,
    n903,
    n554,
    n1519
  );


  nor
  g2222
  (
    n2371,
    n1127,
    n1598,
    n1396,
    n601
  );


  xnor
  g2223
  (
    n2333,
    n1189,
    n735,
    n1296,
    n518
  );


  nor
  g2224
  (
    n1977,
    n1460,
    n995,
    n1726,
    n1221
  );


  xnor
  g2225
  (
    n1770,
    n704,
    n1409,
    n1037,
    n541
  );


  or
  g2226
  (
    n2291,
    n682,
    n1289,
    n940,
    n988
  );


  or
  g2227
  (
    n1892,
    n850,
    n1509,
    n1036,
    n1451
  );


  xor
  g2228
  (
    n2201,
    n645,
    n1097,
    n1389,
    n1604
  );


  and
  g2229
  (
    n1867,
    n1393,
    n1371,
    n487,
    n1734
  );


  xor
  g2230
  (
    n2476,
    n524,
    n1003,
    n1735,
    n1346
  );


  xor
  g2231
  (
    n2122,
    n1531,
    n1272,
    n1143,
    n1524
  );


  or
  g2232
  (
    n2159,
    n1357,
    n551,
    n1348,
    n897
  );


  nand
  g2233
  (
    n2172,
    n1397,
    n1526,
    n641,
    n118
  );


  nand
  g2234
  (
    n1813,
    n1662,
    n1407,
    n706,
    n1675
  );


  or
  g2235
  (
    n1906,
    n1335,
    n825,
    n681,
    n1311
  );


  xnor
  g2236
  (
    n1899,
    n1488,
    n1058,
    n1557,
    n1416
  );


  xor
  g2237
  (
    n2014,
    n993,
    n1457,
    n943,
    n599
  );


  nor
  g2238
  (
    n1992,
    n919,
    n1651,
    n887,
    n1383
  );


  xor
  g2239
  (
    n2043,
    n1539,
    n793,
    n1406,
    n1217
  );


  nor
  g2240
  (
    n1759,
    n888,
    n1138,
    n1438,
    n1608
  );


  nor
  g2241
  (
    n2316,
    n1596,
    n628,
    n1148,
    n660
  );


  and
  g2242
  (
    n2390,
    n1304,
    n958,
    n638,
    n1388
  );


  or
  g2243
  (
    n2108,
    n1034,
    n615,
    n1086,
    n1461
  );


  xnor
  g2244
  (
    n2185,
    n1407,
    n1026,
    n1663,
    n1404
  );


  xor
  g2245
  (
    n1855,
    n1251,
    n1620,
    n1039,
    n1457
  );


  nor
  g2246
  (
    n2045,
    n879,
    n1490,
    n1218,
    n590
  );


  xor
  g2247
  (
    n2033,
    n1304,
    n717,
    n1468,
    n1616
  );


  nand
  g2248
  (
    n1863,
    n1134,
    n1246,
    n1176,
    n1529
  );


  or
  g2249
  (
    n1973,
    n1513,
    n1402,
    n1115,
    n790
  );


  xor
  g2250
  (
    n2203,
    n1364,
    n1342,
    n629,
    n1149
  );


  nand
  g2251
  (
    n2405,
    n1420,
    n1642,
    n1519,
    n1732
  );


  and
  g2252
  (
    n2359,
    n688,
    n1179,
    n1269,
    n892
  );


  or
  g2253
  (
    n2123,
    n1610,
    n1338,
    n1632,
    n1634
  );


  xor
  g2254
  (
    n2342,
    n728,
    n794,
    n1367,
    n1057
  );


  nor
  g2255
  (
    n2182,
    n1554,
    n1678,
    n1556,
    n1424
  );


  nand
  g2256
  (
    n2124,
    n992,
    n816,
    n964,
    n795
  );


  and
  g2257
  (
    n2295,
    n977,
    n1430,
    n1612,
    n766
  );


  xnor
  g2258
  (
    n2408,
    n1370,
    n1571,
    n1170,
    n1005
  );


  and
  g2259
  (
    n1794,
    n985,
    n1019,
    n1612,
    n1006
  );


  nand
  g2260
  (
    n1997,
    n924,
    n803,
    n1182,
    n1147
  );


  nor
  g2261
  (
    n2114,
    n1528,
    n1686,
    n1473,
    n518
  );


  xor
  g2262
  (
    n2125,
    n1306,
    n1536,
    n908,
    n853
  );


  nor
  g2263
  (
    n1830,
    n649,
    n490,
    n1703,
    n684
  );


  nand
  g2264
  (
    n2369,
    n685,
    n1156,
    n813,
    n607
  );


  or
  g2265
  (
    n1879,
    n803,
    n558,
    n478,
    n1148
  );


  nor
  g2266
  (
    n2288,
    n839,
    n1208,
    n1013,
    n1276
  );


  nand
  g2267
  (
    n2352,
    n1603,
    n1359,
    n1281,
    n1643
  );


  xor
  g2268
  (
    n2141,
    n560,
    n1533,
    n1432,
    n1423
  );


  nor
  g2269
  (
    n2254,
    n1096,
    n1518,
    n953,
    n1183
  );


  xor
  g2270
  (
    n2345,
    n1414,
    n1581,
    n1510,
    n1716
  );


  xor
  g2271
  (
    n2130,
    n1560,
    n488,
    n1236,
    n838
  );


  nor
  g2272
  (
    n2175,
    n486,
    n1145,
    n1573,
    n683
  );


  xnor
  g2273
  (
    n1873,
    n1092,
    n893,
    n972,
    n1430
  );


  nand
  g2274
  (
    n1889,
    n1050,
    n957,
    n583,
    n1699
  );


  and
  g2275
  (
    n2161,
    n1651,
    n119,
    n1373,
    n646
  );


  or
  g2276
  (
    n2412,
    n575,
    n1460,
    n1088,
    n1212
  );


  nor
  g2277
  (
    n2146,
    n1613,
    n1427,
    n1556,
    n656
  );


  xnor
  g2278
  (
    n2273,
    n1627,
    n1485,
    n1705,
    n979
  );


  nor
  g2279
  (
    n2463,
    n1582,
    n1701,
    n1239,
    n1440
  );


  nand
  g2280
  (
    n2255,
    n983,
    n690,
    n946,
    n1478
  );


  xor
  g2281
  (
    n1823,
    n1660,
    n1453,
    n1620,
    n784
  );


  or
  g2282
  (
    n2029,
    n895,
    n1503,
    n1466,
    n839
  );


  xnor
  g2283
  (
    n2335,
    n575,
    n1144,
    n1710,
    n1353
  );


  and
  g2284
  (
    n1974,
    n625,
    n1456,
    n1591,
    n944
  );


  xor
  g2285
  (
    n2376,
    n728,
    n1321,
    n1470,
    n1177
  );


  and
  g2286
  (
    n2307,
    n1604,
    n1209,
    n471,
    n864
  );


  and
  g2287
  (
    n1962,
    n1093,
    n1576,
    n1600,
    n764
  );


  nand
  g2288
  (
    n2023,
    n1363,
    n788,
    n1392,
    n654
  );


  nor
  g2289
  (
    n2222,
    n1391,
    n1246,
    n1313,
    n1364
  );


  and
  g2290
  (
    n2370,
    n557,
    n881,
    n1402,
    n1206
  );


  or
  g2291
  (
    n2078,
    n1662,
    n737,
    n1375,
    n809
  );


  nand
  g2292
  (
    n1811,
    n1410,
    n1442,
    n1704,
    n1355
  );


  or
  g2293
  (
    n2274,
    n1599,
    n1036,
    n912,
    n1286
  );


  nor
  g2294
  (
    n1943,
    n1252,
    n1288,
    n1163,
    n1310
  );


  and
  g2295
  (
    n2036,
    n1718,
    n1210,
    n1500,
    n1671
  );


  nor
  g2296
  (
    n1840,
    n1583,
    n1095,
    n1278,
    n1138
  );


  xor
  g2297
  (
    n2107,
    n531,
    n121,
    n523,
    n1481
  );


  xor
  g2298
  (
    n2322,
    n1722,
    n1659,
    n1618,
    n1444
  );


  xor
  g2299
  (
    n1933,
    n1154,
    n1316,
    n994,
    n968
  );


  or
  g2300
  (
    n2213,
    n1080,
    n1394,
    n476,
    n638
  );


  nor
  g2301
  (
    n2502,
    n1521,
    n1019,
    n601,
    n617
  );


  and
  g2302
  (
    n2156,
    n1582,
    n747,
    n1707,
    n613
  );


  xnor
  g2303
  (
    n2230,
    n907,
    n986,
    n1136,
    n1191
  );


  or
  g2304
  (
    n1993,
    n642,
    n637,
    n1281,
    n657
  );


  xor
  g2305
  (
    n2323,
    n935,
    n1314,
    n1186,
    n888
  );


  nand
  g2306
  (
    n2235,
    n753,
    n827,
    n855,
    n1606
  );


  and
  g2307
  (
    n2134,
    n1326,
    n1283,
    n1679,
    n1077
  );


  nor
  g2308
  (
    n1970,
    n1421,
    n845,
    n1022,
    n726
  );


  and
  g2309
  (
    n1893,
    n843,
    n1341,
    n1563,
    n1525
  );


  or
  g2310
  (
    n1929,
    n867,
    n580,
    n1586,
    n509
  );


  or
  g2311
  (
    n2196,
    n1645,
    n1038,
    n678,
    n1698
  );


  xor
  g2312
  (
    n2204,
    n895,
    n1005,
    n818,
    n967
  );


  or
  g2313
  (
    n2058,
    n1486,
    n1529,
    n1446,
    n961
  );


  xnor
  g2314
  (
    n2329,
    n1225,
    n727,
    n925,
    n1733
  );


  nor
  g2315
  (
    n2205,
    n1619,
    n123,
    n1124,
    n120
  );


  nand
  g2316
  (
    n2135,
    n915,
    n990,
    n1439,
    n538
  );


  nor
  g2317
  (
    n2207,
    n1472,
    n847,
    n1485,
    n1411
  );


  xnor
  g2318
  (
    n2356,
    n1683,
    n873,
    n1035,
    n1350
  );


  nor
  g2319
  (
    n2234,
    n925,
    n872,
    n1538,
    n582
  );


  xnor
  g2320
  (
    n1797,
    n1697,
    n1059,
    n1177,
    n1413
  );


  or
  g2321
  (
    n2468,
    n981,
    n958,
    n1676,
    n1137
  );


  xnor
  g2322
  (
    n1901,
    n561,
    n1568,
    n1517,
    n556
  );


  xnor
  g2323
  (
    n1812,
    n1654,
    n1260,
    n1363,
    n121
  );


  nand
  g2324
  (
    n2009,
    n1360,
    n960,
    n549,
    n930
  );


  nand
  g2325
  (
    n1957,
    n506,
    n1724,
    n1187,
    n742
  );


  xnor
  g2326
  (
    n1750,
    n543,
    n1097,
    n1140,
    n658
  );


  xor
  g2327
  (
    n2418,
    n1709,
    n1184,
    n1601,
    n1729
  );


  xnor
  g2328
  (
    n2007,
    n1622,
    n1489,
    n1227,
    n900
  );


  nand
  g2329
  (
    n2258,
    n1055,
    n1591,
    n1449,
    n125
  );


  and
  g2330
  (
    n2148,
    n1713,
    n1035,
    n1242,
    n1608
  );


  xor
  g2331
  (
    n1816,
    n1613,
    n1614,
    n797,
    n832
  );


  xor
  g2332
  (
    n1909,
    n789,
    n1484,
    n639,
    n1412
  );


  or
  g2333
  (
    n1921,
    n1046,
    n780,
    n1573,
    n1329
  );


  or
  g2334
  (
    n2095,
    n563,
    n1366,
    n1677,
    n493
  );


  nand
  g2335
  (
    n2154,
    n1475,
    n470,
    n658,
    n1631
  );


  and
  g2336
  (
    n1903,
    n1494,
    n1570,
    n1444,
    n588
  );


  xnor
  g2337
  (
    n1838,
    n1307,
    n1512,
    n1012,
    n643
  );


  and
  g2338
  (
    n2361,
    n576,
    n1694,
    n1227,
    n659
  );


  nand
  g2339
  (
    n1877,
    n1569,
    n1023,
    n1020,
    n1194
  );


  nor
  g2340
  (
    n1926,
    n1440,
    n809,
    n1524,
    n1550
  );


  nand
  g2341
  (
    n1968,
    n611,
    n1312,
    n786,
    n1433
  );


  xnor
  g2342
  (
    n1894,
    n1477,
    n1496,
    n1329,
    n1541
  );


  and
  g2343
  (
    n2313,
    n1268,
    n1389,
    n500,
    n1033
  );


  xnor
  g2344
  (
    n2240,
    n1591,
    n1720,
    n1678,
    n473
  );


  nor
  g2345
  (
    n2379,
    n1421,
    n1409,
    n832,
    n1438
  );


  xnor
  g2346
  (
    n2308,
    n874,
    n1064,
    n1689,
    n788
  );


  xnor
  g2347
  (
    n2139,
    n806,
    n817,
    n929,
    n585
  );


  nor
  g2348
  (
    n2492,
    n1291,
    n772,
    n955,
    n1517
  );


  nand
  g2349
  (
    n2112,
    n1322,
    n780,
    n1400,
    n1695
  );


  xnor
  g2350
  (
    n2040,
    n824,
    n1495,
    n1498,
    n1690
  );


  and
  g2351
  (
    n2446,
    n470,
    n1106,
    n676,
    n1437
  );


  and
  g2352
  (
    n1986,
    n1507,
    n1006,
    n884,
    n1029
  );


  and
  g2353
  (
    n2454,
    n1033,
    n913,
    n691,
    n841
  );


  or
  g2354
  (
    n1917,
    n563,
    n960,
    n1318,
    n1339
  );


  nand
  g2355
  (
    n2293,
    n1664,
    n1133,
    n116,
    n859
  );


  nor
  g2356
  (
    n1978,
    n1698,
    n534,
    n757,
    n980
  );


  or
  g2357
  (
    n1785,
    n1569,
    n1254,
    n1135,
    n858
  );


  and
  g2358
  (
    n1802,
    n1181,
    n872,
    n920,
    n1551
  );


  or
  g2359
  (
    n2394,
    n1473,
    n1207,
    n1487,
    n1678
  );


  nand
  g2360
  (
    n2076,
    n848,
    n850,
    n1321,
    n946
  );


  xor
  g2361
  (
    n2326,
    n512,
    n1489,
    n661,
    n1669
  );


  nand
  g2362
  (
    n2190,
    n1358,
    n984,
    n118,
    n829
  );


  and
  g2363
  (
    n1814,
    n594,
    n530,
    n1558,
    n1016
  );


  nand
  g2364
  (
    n1897,
    n1602,
    n981,
    n1523,
    n1297
  );


  nand
  g2365
  (
    n2357,
    n944,
    n1622,
    n1546,
    n1616
  );


  xor
  g2366
  (
    n2453,
    n489,
    n1461,
    n644,
    n1101
  );


  nand
  g2367
  (
    n2455,
    n961,
    n1379,
    n733,
    n1542
  );


  nor
  g2368
  (
    n2358,
    n1082,
    n675,
    n1637,
    n741
  );


  nor
  g2369
  (
    n2060,
    n546,
    n1574,
    n1328,
    n121
  );


  nor
  g2370
  (
    n2460,
    n1452,
    n125,
    n1382,
    n1717
  );


  xnor
  g2371
  (
    n2497,
    n990,
    n1498,
    n906,
    n1421
  );


  and
  g2372
  (
    n2498,
    n479,
    n1298,
    n1251,
    n1316
  );


  or
  g2373
  (
    n1976,
    n525,
    n908,
    n779,
    n1631
  );


  xor
  g2374
  (
    n2192,
    n1582,
    n904,
    n1298,
    n1289
  );


  or
  g2375
  (
    n2424,
    n828,
    n877,
    n1703,
    n1451
  );


  xor
  g2376
  (
    n1958,
    n1080,
    n1603,
    n1467,
    n1375
  );


  nand
  g2377
  (
    n2386,
    n1165,
    n1151,
    n1725,
    n1172
  );


  xor
  g2378
  (
    n2166,
    n965,
    n817,
    n550,
    n1283
  );


  and
  g2379
  (
    n1961,
    n822,
    n1666,
    n496,
    n1043
  );


  or
  g2380
  (
    n1975,
    n723,
    n699,
    n1722,
    n500
  );


  and
  g2381
  (
    n1856,
    n1719,
    n519,
    n1311,
    n715
  );


  and
  g2382
  (
    n2441,
    n1537,
    n783,
    n1417,
    n812
  );


  nor
  g2383
  (
    n1862,
    n664,
    n1053,
    n1405,
    n1535
  );


  nor
  g2384
  (
    n2085,
    n797,
    n1188,
    n1239,
    n1348
  );


  xnor
  g2385
  (
    n2220,
    n578,
    n1416,
    n1592,
    n1455
  );


  or
  g2386
  (
    n1918,
    n789,
    n1253,
    n616,
    n1090
  );


  or
  g2387
  (
    n1778,
    n565,
    n1431,
    n815,
    n1011
  );


  xor
  g2388
  (
    n2494,
    n1323,
    n1354,
    n1212,
    n1330
  );


  xnor
  g2389
  (
    n2225,
    n1713,
    n537,
    n597,
    n1448
  );


  and
  g2390
  (
    n1774,
    n1302,
    n1588,
    n1329,
    n1056
  );


  xnor
  g2391
  (
    n2402,
    n926,
    n714,
    n1401,
    n1617
  );


  xnor
  g2392
  (
    n2269,
    n1263,
    n1677,
    n1118,
    n540
  );


  nor
  g2393
  (
    n2404,
    n929,
    n1479,
    n1399,
    n1074
  );


  nor
  g2394
  (
    n1886,
    n1652,
    n1635,
    n1160,
    n724
  );


  and
  g2395
  (
    n2461,
    n1479,
    n1661,
    n1315,
    n680
  );


  xor
  g2396
  (
    n2452,
    n962,
    n1724,
    n1487,
    n1426
  );


  and
  g2397
  (
    n1757,
    n1552,
    n1167,
    n1029,
    n1185
  );


  xor
  g2398
  (
    n1902,
    n1649,
    n557,
    n1136,
    n1604
  );


  or
  g2399
  (
    n1916,
    n1730,
    n678,
    n1373,
    n631
  );


  nand
  g2400
  (
    n1890,
    n1259,
    n1443,
    n1008,
    n826
  );


  xor
  g2401
  (
    n2070,
    n1242,
    n1585,
    n1550,
    n1575
  );


  nand
  g2402
  (
    n2099,
    n702,
    n1601,
    n1228,
    n1548
  );


  xor
  g2403
  (
    n2064,
    n1372,
    n1410,
    n1551,
    n1597
  );


  xnor
  g2404
  (
    n1905,
    n613,
    n1180,
    n1313,
    n1117
  );


  and
  g2405
  (
    n2168,
    n1440,
    n932,
    n750,
    n1624
  );


  nor
  g2406
  (
    n1805,
    n673,
    n976,
    n1609,
    n852
  );


  or
  g2407
  (
    n1818,
    n1222,
    n1548,
    n782,
    n1681
  );


  nand
  g2408
  (
    n1988,
    n879,
    n1549,
    n510,
    n1049
  );


  nor
  g2409
  (
    n2215,
    n1684,
    n851,
    n706,
    n1042
  );


  xor
  g2410
  (
    n1896,
    n822,
    n1115,
    n1211,
    n1478
  );


  and
  g2411
  (
    n1907,
    n1480,
    n1535,
    n596,
    n774
  );


  or
  g2412
  (
    n2013,
    n1361,
    n1161,
    n892,
    n1547
  );


  xnor
  g2413
  (
    n1932,
    n1030,
    n1069,
    n708,
    n729
  );


  or
  g2414
  (
    n2464,
    n1220,
    n478,
    n1141,
    n880
  );


  nand
  g2415
  (
    n2153,
    n1476,
    n681,
    n1060,
    n951
  );


  xor
  g2416
  (
    n2202,
    n1361,
    n889,
    n792,
    n771
  );


  xnor
  g2417
  (
    n2177,
    n744,
    n754,
    n1717,
    n1316
  );


  nor
  g2418
  (
    n1980,
    n1123,
    n1376,
    n1615,
    n552
  );


  nor
  g2419
  (
    n1783,
    n656,
    n1471,
    n679,
    n612
  );


  or
  g2420
  (
    n2336,
    n1387,
    n744,
    n1197,
    n962
  );


  xnor
  g2421
  (
    n1766,
    n1060,
    n847,
    n1243,
    n1536
  );


  nor
  g2422
  (
    n2251,
    n1312,
    n1415,
    n1014,
    n650
  );


  or
  g2423
  (
    n2485,
    n1737,
    n1032,
    n1687,
    n1084
  );


  nor
  g2424
  (
    n1922,
    n689,
    n1718,
    n1064,
    n627
  );


  nand
  g2425
  (
    n2217,
    n555,
    n1374,
    n1139,
    n1216
  );


  xor
  g2426
  (
    n2051,
    n1173,
    n736,
    n739,
    n1266
  );


  xor
  g2427
  (
    n2382,
    n1501,
    n734,
    n1491,
    n1345
  );


  nor
  g2428
  (
    n1952,
    n525,
    n1190,
    n1330,
    n1044
  );


  xor
  g2429
  (
    n2025,
    n992,
    n1074,
    n938,
    n1166
  );


  nand
  g2430
  (
    n1801,
    n1219,
    n1669,
    n1386,
    n1040
  );


  nand
  g2431
  (
    n1887,
    n1201,
    n776,
    n1340,
    n1334
  );


  xor
  g2432
  (
    n2360,
    n1633,
    n820,
    n936,
    n1015
  );


  or
  g2433
  (
    n1949,
    n1287,
    n915,
    n1407,
    n1274
  );


  nand
  g2434
  (
    n1989,
    n932,
    n1208,
    n1692,
    n768
  );


  nand
  g2435
  (
    n2388,
    n1635,
    n1444,
    n700,
    n898
  );


  nor
  g2436
  (
    n2054,
    n1737,
    n1170,
    n1406,
    n116
  );


  and
  g2437
  (
    n2239,
    n1544,
    n1442,
    n1366,
    n1531
  );


  or
  g2438
  (
    n2305,
    n577,
    n1337,
    n1465,
    n1382
  );


  nor
  g2439
  (
    n1984,
    n1675,
    n1690,
    n1259,
    n1270
  );


  xnor
  g2440
  (
    n2362,
    n1020,
    n1586,
    n1204,
    n1471
  );


  xnor
  g2441
  (
    n2211,
    n1683,
    n1301,
    n1292,
    n1607
  );


  xor
  g2442
  (
    n2363,
    n1464,
    n1098,
    n1078,
    n1231
  );


  and
  g2443
  (
    n1844,
    n1646,
    n1384,
    n648,
    n1541
  );


  and
  g2444
  (
    n2324,
    n1378,
    n1114,
    n976,
    n701
  );


  or
  g2445
  (
    n2068,
    n1226,
    n600,
    n1298,
    n863
  );


  nand
  g2446
  (
    n2249,
    n1091,
    n1282,
    n119,
    n623
  );


  or
  g2447
  (
    n2457,
    n634,
    n1411,
    n1467,
    n1297
  );


  xor
  g2448
  (
    n2028,
    n1621,
    n1441,
    n1657,
    n1606
  );


  and
  g2449
  (
    n1913,
    n1221,
    n700,
    n554,
    n1544
  );


  xor
  g2450
  (
    n1940,
    n854,
    n1309,
    n1114,
    n787
  );


  nor
  g2451
  (
    n1843,
    n1301,
    n635,
    n1540,
    n1008
  );


  or
  g2452
  (
    n2061,
    n626,
    n1624,
    n712,
    n904
  );


  xnor
  g2453
  (
    n1931,
    n998,
    n1513,
    n1650,
    n1330
  );


  xor
  g2454
  (
    n2221,
    n1396,
    n773,
    n1133,
    n1538
  );


  and
  g2455
  (
    n1804,
    n1663,
    n530,
    n909,
    n1648
  );


  or
  g2456
  (
    n1923,
    n761,
    n1510,
    n635,
    n561
  );


  nor
  g2457
  (
    n1937,
    n1581,
    n1271,
    n1089,
    n498
  );


  nor
  g2458
  (
    n1751,
    n1608,
    n1492,
    n835,
    n1507
  );


  and
  g2459
  (
    n2152,
    n1356,
    n1548,
    n1331,
    n1584
  );


  xnor
  g2460
  (
    n2458,
    n875,
    n1366,
    n1459,
    n717
  );


  nand
  g2461
  (
    n1853,
    n1482,
    n1266,
    n1684,
    n1119
  );


  and
  g2462
  (
    n1841,
    n998,
    n1222,
    n620,
    n1521
  );


  and
  g2463
  (
    n2298,
    n1730,
    n1490,
    n1322,
    n1134
  );


  and
  g2464
  (
    n2466,
    n758,
    n1664,
    n1397,
    n1422
  );


  xnor
  g2465
  (
    n2262,
    n774,
    n1412,
    n746,
    n1247
  );


  xor
  g2466
  (
    n1852,
    n1657,
    n1736,
    n1327,
    n1012
  );


  nor
  g2467
  (
    n2160,
    n1527,
    n1353,
    n1231,
    n1453
  );


  or
  g2468
  (
    n2341,
    n864,
    n865,
    n686,
    n672
  );


  xor
  g2469
  (
    n2275,
    n1199,
    n1197,
    n1702,
    n577
  );


  nor
  g2470
  (
    n1928,
    n1666,
    n815,
    n773,
    n991
  );


  nand
  g2471
  (
    n2290,
    n930,
    n1072,
    n1590,
    n565
  );


  and
  g2472
  (
    n2410,
    n714,
    n1462,
    n1045,
    n1653
  );


  nor
  g2473
  (
    n1849,
    n1505,
    n954,
    n1295,
    n1390
  );


  xor
  g2474
  (
    n2641,
    n2130,
    n2146,
    n2268,
    n1835
  );


  or
  g2475
  (
    n2654,
    n2412,
    n2411,
    n2178,
    n2128
  );


  or
  g2476
  (
    n2648,
    n2282,
    n2242,
    n1772,
    n1892
  );


  xnor
  g2477
  (
    n2585,
    n2286,
    n2438,
    n1815,
    n2235
  );


  and
  g2478
  (
    n2650,
    n2001,
    n2254,
    n1863,
    n2238
  );


  xnor
  g2479
  (
    n2572,
    n1867,
    n1821,
    n1960,
    n2115
  );


  or
  g2480
  (
    n2550,
    n2252,
    n2353,
    n2005,
    n2047
  );


  or
  g2481
  (
    n2653,
    n2211,
    n1807,
    n2199,
    n2423
  );


  xnor
  g2482
  (
    n2674,
    n1830,
    n1857,
    n2000,
    n1843
  );


  nand
  g2483
  (
    n2633,
    n2150,
    n2088,
    n1864,
    n2320
  );


  xnor
  g2484
  (
    n2507,
    n1766,
    n2249,
    n2439,
    n1829
  );


  xor
  g2485
  (
    n2619,
    n1840,
    n2343,
    n2201,
    n2127
  );


  or
  g2486
  (
    n2598,
    n2229,
    n2148,
    n1812,
    n1986
  );


  nor
  g2487
  (
    n2651,
    n2061,
    n2010,
    n1968,
    n2259
  );


  xnor
  g2488
  (
    n2524,
    n2064,
    n2042,
    n2085,
    n1948
  );


  or
  g2489
  (
    n2593,
    n1873,
    n2195,
    n1854,
    n1832
  );


  or
  g2490
  (
    n2661,
    n1822,
    n2237,
    n2440,
    n2291
  );


  nor
  g2491
  (
    n2643,
    n1778,
    n2285,
    n2078,
    n1775
  );


  or
  g2492
  (
    n2520,
    n2153,
    n2395,
    n1824,
    n2212
  );


  and
  g2493
  (
    n2560,
    n2038,
    n1894,
    n1860,
    n2221
  );


  or
  g2494
  (
    n2611,
    n2069,
    n2176,
    n2145,
    n2327
  );


  nor
  g2495
  (
    n2536,
    n1844,
    n2113,
    n2244,
    n1862
  );


  and
  g2496
  (
    n2631,
    n1833,
    n1827,
    n2152,
    n2057
  );


  xnor
  g2497
  (
    n2531,
    n2151,
    n1810,
    n2086,
    n2335
  );


  xor
  g2498
  (
    n2665,
    n2016,
    n2154,
    n1871,
    n2453
  );


  and
  g2499
  (
    n2679,
    n2223,
    n2300,
    n2400,
    n2135
  );


  xnor
  g2500
  (
    n2618,
    n1970,
    n1790,
    n1918,
    n2364
  );


  xnor
  g2501
  (
    n2597,
    n2202,
    n1904,
    n2275,
    n1893
  );


  nor
  g2502
  (
    n2581,
    n1774,
    n1977,
    n1791,
    n2386
  );


  and
  g2503
  (
    n2594,
    n2448,
    n2402,
    n2206,
    n2339
  );


  and
  g2504
  (
    n2678,
    n1980,
    n2329,
    n1962,
    n1955
  );


  nand
  g2505
  (
    n2535,
    n2272,
    n1915,
    n2279,
    n2370
  );


  xnor
  g2506
  (
    n2655,
    n2375,
    n1811,
    n1999,
    n1911
  );


  nor
  g2507
  (
    n2533,
    n2014,
    n2326,
    n2276,
    n1965
  );


  xor
  g2508
  (
    n2517,
    n1912,
    n2156,
    n1878,
    n2295
  );


  nand
  g2509
  (
    n2578,
    n1966,
    n2186,
    n2379,
    n2445
  );


  and
  g2510
  (
    n2516,
    n2099,
    n2209,
    n2012,
    n2302
  );


  xor
  g2511
  (
    n2541,
    n2068,
    n2435,
    n2294,
    n2261
  );


  nor
  g2512
  (
    n2532,
    n2287,
    n2278,
    n2250,
    n2214
  );


  nor
  g2513
  (
    n2623,
    n2031,
    n2369,
    n1800,
    n2055
  );


  nor
  g2514
  (
    n2647,
    n1913,
    n2441,
    n1946,
    n2349
  );


  nand
  g2515
  (
    n2591,
    n2257,
    n1937,
    n2174,
    n2418
  );


  or
  g2516
  (
    n2577,
    n2305,
    n1759,
    n2399,
    n1785
  );


  or
  g2517
  (
    n2612,
    n1817,
    n2280,
    n2160,
    n1856
  );


  and
  g2518
  (
    n2630,
    n2110,
    n2104,
    n1853,
    n2389
  );


  xnor
  g2519
  (
    n2639,
    n2319,
    n2158,
    n1763,
    n2376
  );


  and
  g2520
  (
    n2660,
    n2427,
    n2454,
    n1909,
    n2312
  );


  and
  g2521
  (
    n2656,
    n2308,
    n2106,
    n2233,
    n2018
  );


  or
  g2522
  (
    n2556,
    n1865,
    n1819,
    n2098,
    n2290
  );


  nor
  g2523
  (
    n2610,
    n1839,
    n2301,
    n2415,
    n1938
  );


  and
  g2524
  (
    n2638,
    n2120,
    n2048,
    n1764,
    n2270
  );


  and
  g2525
  (
    n2571,
    n2125,
    n2071,
    n1927,
    n2367
  );


  and
  g2526
  (
    n2519,
    n2204,
    n1998,
    n1762,
    n2118
  );


  nand
  g2527
  (
    n2671,
    n2167,
    n2025,
    n2137,
    n2341
  );


  xnor
  g2528
  (
    n2545,
    n2215,
    n1761,
    n2283,
    n2333
  );


  and
  g2529
  (
    n2552,
    n2119,
    n1818,
    n1834,
    n2187
  );


  xnor
  g2530
  (
    n2505,
    n1795,
    n1877,
    n1969,
    n2245
  );


  and
  g2531
  (
    n2669,
    n2044,
    n2234,
    n2059,
    n2050
  );


  nand
  g2532
  (
    n2554,
    n2314,
    n2166,
    n2361,
    n2181
  );


  or
  g2533
  (
    n2549,
    n1950,
    n2103,
    n2109,
    n1934
  );


  and
  g2534
  (
    n2551,
    n2425,
    n1806,
    n2413,
    n2046
  );


  and
  g2535
  (
    n2543,
    n2112,
    n1984,
    n1942,
    n2424
  );


  nor
  g2536
  (
    n2670,
    n2419,
    n1768,
    n2348,
    n2208
  );


  and
  g2537
  (
    n2657,
    n2456,
    n2081,
    n2139,
    n2360
  );


  or
  g2538
  (
    n2646,
    n1801,
    n2321,
    n2019,
    n2105
  );


  nor
  g2539
  (
    n2642,
    n1976,
    n1826,
    n1972,
    n1845
  );


  and
  g2540
  (
    n2676,
    n1870,
    n2039,
    n2262,
    n1851
  );


  xnor
  g2541
  (
    n2652,
    n2188,
    n1978,
    n2102,
    n1951
  );


  and
  g2542
  (
    n2615,
    n2023,
    n1841,
    n1885,
    n2318
  );


  and
  g2543
  (
    n2609,
    n1947,
    n2449,
    n2388,
    n2062
  );


  nand
  g2544
  (
    n2625,
    n2365,
    n1989,
    n2008,
    n1985
  );


  xnor
  g2545
  (
    n2546,
    n1786,
    n1975,
    n2284,
    n2332
  );


  nor
  g2546
  (
    n2603,
    n2277,
    n2450,
    n2394,
    n2074
  );


  xor
  g2547
  (
    n2569,
    n2240,
    n1929,
    n1881,
    n2207
  );


  nand
  g2548
  (
    n2566,
    n1898,
    n1872,
    n2269,
    n2218
  );


  xor
  g2549
  (
    n2522,
    n2004,
    n2310,
    n2239,
    n1943
  );


  and
  g2550
  (
    n2530,
    n2385,
    n1794,
    n2434,
    n2095
  );


  and
  g2551
  (
    n2521,
    n2027,
    n2180,
    n2183,
    n2315
  );


  nor
  g2552
  (
    n2539,
    n2281,
    n1990,
    n1825,
    n2368
  );


  or
  g2553
  (
    n2605,
    n2003,
    n2011,
    n1941,
    n2253
  );


  nand
  g2554
  (
    n2664,
    n2219,
    n2403,
    n2296,
    n1804
  );


  xor
  g2555
  (
    n2514,
    n1883,
    n1930,
    n1887,
    n2304
  );


  xor
  g2556
  (
    n2547,
    n2354,
    n2271,
    n2442,
    n1789
  );


  nor
  g2557
  (
    n2600,
    n2210,
    n2136,
    n2017,
    n2013
  );


  and
  g2558
  (
    n2644,
    n2328,
    n1842,
    n2266,
    n1917
  );


  nor
  g2559
  (
    n2599,
    n2089,
    n1875,
    n2426,
    n1926
  );


  xor
  g2560
  (
    n2673,
    n1890,
    n2248,
    n2065,
    n2350
  );


  nand
  g2561
  (
    n2553,
    n2165,
    n2192,
    n1945,
    n2116
  );


  and
  g2562
  (
    n2645,
    n2124,
    n2397,
    n2224,
    n1808
  );


  or
  g2563
  (
    n2509,
    n1820,
    n1838,
    n1897,
    n1848
  );


  xnor
  g2564
  (
    n2621,
    n2138,
    n2100,
    n1953,
    n1855
  );


  or
  g2565
  (
    n2586,
    n2142,
    n1828,
    n2222,
    n2351
  );


  or
  g2566
  (
    n2662,
    n2052,
    n2063,
    n1900,
    n2322
  );


  xnor
  g2567
  (
    n2616,
    n1993,
    n1799,
    n2316,
    n2101
  );


  nand
  g2568
  (
    n2523,
    n1776,
    n1936,
    n1932,
    n2420
  );


  nor
  g2569
  (
    n2672,
    n2034,
    n1902,
    n1886,
    n2363
  );


  nand
  g2570
  (
    n2525,
    n1925,
    n2429,
    n1837,
    n2340
  );


  xnor
  g2571
  (
    n2629,
    n2227,
    n2359,
    n2433,
    n2182
  );


  and
  g2572
  (
    n2557,
    n2092,
    n1770,
    n1995,
    n2377
  );


  or
  g2573
  (
    n2518,
    n1796,
    n1798,
    n2225,
    n2372
  );


  xnor
  g2574
  (
    n2677,
    n2073,
    n2371,
    n1994,
    n1905
  );


  xor
  g2575
  (
    n2511,
    n2036,
    n2196,
    n1997,
    n2457
  );


  and
  g2576
  (
    n2659,
    n2177,
    n1831,
    n2094,
    n2410
  );


  nand
  g2577
  (
    n2555,
    n2256,
    n1852,
    n2396,
    n2049
  );


  xnor
  g2578
  (
    n2575,
    n1923,
    n1813,
    n2198,
    n2337
  );


  nor
  g2579
  (
    n2537,
    n1868,
    n1988,
    n2297,
    n1802
  );


  or
  g2580
  (
    n2587,
    n2409,
    n2444,
    n2338,
    n2140
  );


  xnor
  g2581
  (
    n2565,
    n2060,
    n2264,
    n2406,
    n1952
  );


  or
  g2582
  (
    n2624,
    n1916,
    n1793,
    n2431,
    n2197
  );


  or
  g2583
  (
    n2580,
    n1958,
    n2452,
    n2288,
    n1919
  );


  xnor
  g2584
  (
    n2540,
    n1760,
    n2355,
    n1792,
    n2390
  );


  and
  g2585
  (
    n2637,
    n2179,
    n2357,
    n2306,
    n2006
  );


  nor
  g2586
  (
    n2632,
    n2366,
    n2307,
    n2173,
    n1788
  );


  or
  g2587
  (
    n2576,
    n1781,
    n2077,
    n2067,
    n2163
  );


  xor
  g2588
  (
    n2513,
    n2381,
    n2053,
    n2324,
    n2026
  );


  nand
  g2589
  (
    n2595,
    n1859,
    n2289,
    n1928,
    n2387
  );


  nand
  g2590
  (
    n2626,
    n2122,
    n2162,
    n2323,
    n2216
  );


  xor
  g2591
  (
    n2564,
    n2293,
    n2408,
    n1992,
    n1982
  );


  xor
  g2592
  (
    n2640,
    n1884,
    n2093,
    n2455,
    n2309
  );


  xor
  g2593
  (
    n2675,
    n1771,
    n2203,
    n2380,
    n2084
  );


  and
  g2594
  (
    n2567,
    n2241,
    n1935,
    n2422,
    n1803
  );


  nand
  g2595
  (
    n2573,
    n2133,
    n1922,
    n2002,
    n1847
  );


  xor
  g2596
  (
    n2583,
    n2121,
    n1963,
    n1805,
    n1858
  );


  nand
  g2597
  (
    n2592,
    n2168,
    n2267,
    n2217,
    n2352
  );


  nor
  g2598
  (
    n2617,
    n2230,
    n2443,
    n1957,
    n2021
  );


  or
  g2599
  (
    n2606,
    n2255,
    n2416,
    n1880,
    n2149
  );


  xor
  g2600
  (
    n2589,
    n2129,
    n2330,
    n2417,
    n1939
  );


  and
  g2601
  (
    n2596,
    n2051,
    n2317,
    n2383,
    n1773
  );


  xor
  g2602
  (
    n2506,
    n2079,
    n2205,
    n2232,
    n2056
  );


  nor
  g2603
  (
    n2608,
    n1949,
    n2428,
    n2298,
    n2213
  );


  nor
  g2604
  (
    n2601,
    n2043,
    n2111,
    n2247,
    n1959
  );


  or
  g2605
  (
    n2542,
    n1823,
    n1861,
    n1809,
    n2347
  );


  nand
  g2606
  (
    n2613,
    n1906,
    n1780,
    n2131,
    n1891
  );


  xor
  g2607
  (
    n2527,
    n2260,
    n2083,
    n2345,
    n2382
  );


  xor
  g2608
  (
    n2620,
    n2299,
    n2391,
    n2144,
    n1846
  );


  xor
  g2609
  (
    n2579,
    n1971,
    n1895,
    n1869,
    n2108
  );


  nand
  g2610
  (
    n2666,
    n1816,
    n2458,
    n1866,
    n2058
  );


  and
  g2611
  (
    n2584,
    n1921,
    n1769,
    n2447,
    n1903
  );


  or
  g2612
  (
    n2563,
    n1967,
    n2313,
    n1991,
    n2407
  );


  xnor
  g2613
  (
    n2508,
    n2334,
    n1964,
    n1888,
    n2414
  );


  or
  g2614
  (
    n2512,
    n1777,
    n2029,
    n2421,
    n1908
  );


  or
  g2615
  (
    n2528,
    n1850,
    n2096,
    n2161,
    n2147
  );


  xnor
  g2616
  (
    n2627,
    n2032,
    n2273,
    n2446,
    n2020
  );


  xnor
  g2617
  (
    n2574,
    n2373,
    n2097,
    n1973,
    n2157
  );


  nand
  g2618
  (
    n2538,
    n2033,
    n2132,
    n2075,
    n2066
  );


  nand
  g2619
  (
    n2570,
    n2028,
    n2045,
    n1767,
    n2404
  );


  xnor
  g2620
  (
    n2668,
    n2384,
    n2040,
    n1874,
    n2170
  );


  nand
  g2621
  (
    n2559,
    n2303,
    n2193,
    n2022,
    n2331
  );


  and
  g2622
  (
    n2568,
    n1814,
    n2251,
    n1779,
    n2009
  );


  xnor
  g2623
  (
    n2602,
    n2030,
    n2175,
    n2430,
    n1996
  );


  nand
  g2624
  (
    n2526,
    n2200,
    n2076,
    n2405,
    n2346
  );


  xnor
  g2625
  (
    n2588,
    n1849,
    n2189,
    n2311,
    n1899
  );


  nor
  g2626
  (
    n2622,
    n2191,
    n1889,
    n2292,
    n2159
  );


  and
  g2627
  (
    n2544,
    n2185,
    n2356,
    n1765,
    n1931
  );


  xor
  g2628
  (
    n2510,
    n1914,
    n1901,
    n2451,
    n1924
  );


  nand
  g2629
  (
    n2663,
    n1979,
    n2114,
    n2190,
    n2091
  );


  xnor
  g2630
  (
    n2667,
    n2041,
    n2070,
    n2344,
    n2123
  );


  or
  g2631
  (
    n2590,
    n2325,
    n2265,
    n2107,
    n1961
  );


  xor
  g2632
  (
    n2548,
    n2228,
    n2090,
    n1940,
    n1954
  );


  or
  g2633
  (
    n2604,
    n2437,
    n2171,
    n2054,
    n2194
  );


  xnor
  g2634
  (
    n2515,
    n2392,
    n2024,
    n2274,
    n2243
  );


  xnor
  g2635
  (
    n2614,
    n2126,
    n2231,
    n1896,
    n1784
  );


  xor
  g2636
  (
    n2534,
    n1907,
    n2015,
    n2184,
    n1933
  );


  xnor
  g2637
  (
    n2636,
    n2258,
    n1836,
    n2358,
    n1882
  );


  nor
  g2638
  (
    n2649,
    n2141,
    n2143,
    n2362,
    n2155
  );


  xor
  g2639
  (
    n2562,
    n2432,
    n2374,
    n2378,
    n1782
  );


  nand
  g2640
  (
    n2658,
    n1879,
    n1983,
    n2263,
    n1944
  );


  xor
  g2641
  (
    n2558,
    n2436,
    n2117,
    n2080,
    n2393
  );


  xnor
  g2642
  (
    n2634,
    n2336,
    n1920,
    n2401,
    n2134
  );


  nor
  g2643
  (
    n2582,
    n1981,
    n2398,
    n2220,
    n2087
  );


  xnor
  g2644
  (
    n2607,
    n1876,
    n1910,
    n2226,
    n1787
  );


  nand
  g2645
  (
    n2529,
    n1797,
    n2169,
    n1783,
    n2007
  );


  and
  g2646
  (
    n2628,
    n1987,
    n2035,
    n2172,
    n2037
  );


  nor
  g2647
  (
    n2561,
    n2246,
    n2342,
    n2164,
    n1956
  );


  xnor
  g2648
  (
    n2635,
    n2082,
    n2236,
    n1974,
    n2072
  );


  xor
  g2649
  (
    n2688,
    n1737,
    n2508,
    n1738,
    n2511
  );


  or
  g2650
  (
    n2686,
    n1741,
    n1739,
    n2506,
    n1740
  );


  or
  g2651
  (
    n2687,
    n1746,
    n1743,
    n1742
  );


  and
  g2652
  (
    n2681,
    n1740,
    n1746,
    n1741,
    n1744
  );


  nand
  g2653
  (
    n2685,
    n2507,
    n1745,
    n1741,
    n1744
  );


  nor
  g2654
  (
    n2682,
    n2510,
    n1744,
    n1745,
    n1739
  );


  xor
  g2655
  (
    n2683,
    n1738,
    n2505,
    n1745,
    n2513
  );


  and
  g2656
  (
    n2680,
    n1743,
    n2509,
    n2512,
    n1739
  );


  xnor
  g2657
  (
    n2684,
    n1743,
    n1738,
    n1740,
    n1742
  );


  nand
  g2658
  (
    n2689,
    n2482,
    n2464,
    n2462,
    n2684
  );


  nand
  g2659
  (
    n2692,
    n2687,
    n2476,
    n2461,
    n2467
  );


  xor
  g2660
  (
    n2690,
    n2685,
    n2481,
    n2469,
    n2459
  );


  nand
  g2661
  (
    n2693,
    n2474,
    n2687,
    n2683,
    n2465
  );


  or
  g2662
  (
    n2691,
    n2463,
    n2477,
    n2681,
    n2470
  );


  and
  g2663
  (
    n2695,
    n2460,
    n2479,
    n2466,
    n2473
  );


  nor
  g2664
  (
    n2696,
    n2468,
    n2682,
    n2471,
    n2475
  );


  nand
  g2665
  (
    n2694,
    n2686,
    n2472,
    n2480,
    n2478
  );


  and
  g2666
  (
    n2713,
    n2526,
    n2691,
    n2542,
    n2690
  );


  nor
  g2667
  (
    n2708,
    n2690,
    n2693,
    n2522,
    n2519
  );


  or
  g2668
  (
    n2714,
    n2546,
    n2533,
    n2690,
    n2545
  );


  nand
  g2669
  (
    n2703,
    n2527,
    n2689,
    n2693
  );


  xnor
  g2670
  (
    n2705,
    n2534,
    n2515,
    n2555,
    n2548
  );


  nand
  g2671
  (
    n2712,
    n2531,
    n1747,
    n2553,
    n2530
  );


  nand
  g2672
  (
    n2698,
    n2543,
    n2528,
    n2551,
    n2547
  );


  xnor
  g2673
  (
    n2697,
    n2544,
    n2691,
    n2692,
    n2563
  );


  xor
  g2674
  (
    n2701,
    n2520,
    n2517,
    n2689,
    n2550
  );


  nor
  g2675
  (
    n2700,
    n2691,
    n2538,
    n1746,
    n2521
  );


  nor
  g2676
  (
    n2706,
    n2525,
    n2524,
    n1747,
    n2541
  );


  xor
  g2677
  (
    n2702,
    n2549,
    n2554,
    n2692,
    n2540
  );


  and
  g2678
  (
    n2710,
    n2690,
    n2561,
    n2689,
    n2516
  );


  and
  g2679
  (
    n2704,
    n2552,
    n2558,
    n2691,
    n2539
  );


  nand
  g2680
  (
    n2699,
    n2514,
    n2692,
    n2562,
    n2557
  );


  or
  g2681
  (
    n2709,
    n2523,
    n2529,
    n2556,
    n2536
  );


  or
  g2682
  (
    n2711,
    n2535,
    n2560,
    n2564,
    n2692
  );


  or
  g2683
  (
    n2707,
    n2532,
    n2559,
    n2518,
    n2537
  );


  buf
  g2684
  (
    n2720,
    n2702
  );


  not
  g2685
  (
    n2716,
    n2699
  );


  buf
  g2686
  (
    n2717,
    n2697
  );


  buf
  g2687
  (
    n2715,
    n2700
  );


  not
  g2688
  (
    n2719,
    n2698
  );


  not
  g2689
  (
    n2718,
    n2701
  );


  xnor
  g2690
  (
    n2736,
    n2580,
    n2614,
    n2716,
    n2577
  );


  nor
  g2691
  (
    n2737,
    n2715,
    n2581,
    n2607,
    n2628
  );


  or
  g2692
  (
    n2730,
    n2597,
    n2715,
    n2629,
    n2719
  );


  and
  g2693
  (
    n2743,
    n2589,
    n2575,
    n2693,
    n2579
  );


  nor
  g2694
  (
    n2738,
    n2585,
    n2591,
    n2605,
    n2718
  );


  nor
  g2695
  (
    n2726,
    n2587,
    n2588,
    n2717,
    n2566
  );


  or
  g2696
  (
    n2727,
    n2582,
    n2622,
    n2720,
    n2610
  );


  xnor
  g2697
  (
    n2744,
    n2584,
    n2693,
    n2578,
    n2717
  );


  xnor
  g2698
  (
    n2734,
    n2613,
    n2571,
    n2694,
    n2606
  );


  xor
  g2699
  (
    n2735,
    n2719,
    n2719,
    n2604,
    n2611
  );


  xor
  g2700
  (
    n2731,
    n2573,
    n2720,
    n2583
  );


  xnor
  g2701
  (
    n2728,
    n2596,
    n2603,
    n2568,
    n2616
  );


  xnor
  g2702
  (
    n2732,
    n2625,
    n2615,
    n2715,
    n2694
  );


  nand
  g2703
  (
    n2729,
    n2621,
    n2717,
    n2576,
    n2574
  );


  xnor
  g2704
  (
    n2722,
    n2608,
    n2609,
    n2715,
    n2617
  );


  xnor
  g2705
  (
    n2742,
    n2718,
    n2592,
    n2716,
    n2627
  );


  xor
  g2706
  (
    n2725,
    n2483,
    n2612,
    n2602,
    n2572
  );


  xnor
  g2707
  (
    n2740,
    n2569,
    n2720,
    n2719,
    n2590
  );


  or
  g2708
  (
    n2724,
    n2717,
    n2593,
    n2716,
    n2601
  );


  nand
  g2709
  (
    n2721,
    n2718,
    n2586,
    n2600,
    n2595
  );


  or
  g2710
  (
    n2723,
    n2694,
    n2618,
    n2624,
    n2619
  );


  and
  g2711
  (
    n2733,
    n2598,
    n2570,
    n2594,
    n2599
  );


  xor
  g2712
  (
    n2739,
    n2620,
    n2630,
    n2716,
    n2565
  );


  xor
  g2713
  (
    n2741,
    n2718,
    n2626,
    n2567,
    n2623
  );


  nand
  g2714
  (
    n2764,
    n2712,
    n2728,
    n2669,
    n2723
  );


  or
  g2715
  (
    n2762,
    n2729,
    n2709,
    n2631,
    n2666
  );


  xnor
  g2716
  (
    n2759,
    n2646,
    n2724,
    n2643,
    n2721
  );


  xor
  g2717
  (
    n2766,
    n2722,
    n2730,
    n2652,
    n2727
  );


  xnor
  g2718
  (
    n2751,
    n2495,
    n2703,
    n2491,
    n2639
  );


  or
  g2719
  (
    n2754,
    n2663,
    n2635,
    n2657,
    n2634
  );


  xnor
  g2720
  (
    n2749,
    n2726,
    n2727,
    n2642,
    n2658
  );


  xnor
  g2721
  (
    n2767,
    n2485,
    n2488,
    n2725
  );


  xor
  g2722
  (
    n2755,
    n2723,
    n2645,
    n2656,
    n2722
  );


  and
  g2723
  (
    n2745,
    n2724,
    n2484,
    n2638,
    n2661
  );


  and
  g2724
  (
    n2770,
    n2714,
    n2688,
    n2711,
    n2644
  );


  nor
  g2725
  (
    n2748,
    n2648,
    n2727,
    n2704,
    n2725
  );


  xnor
  g2726
  (
    n2752,
    n2489,
    n2659,
    n2727,
    n2492
  );


  nor
  g2727
  (
    n2768,
    n2664,
    n2726,
    n2710,
    n2662
  );


  nand
  g2728
  (
    n2758,
    n2723,
    n2708,
    n2649,
    n2725
  );


  nand
  g2729
  (
    n2753,
    n2487,
    n2655,
    n2726,
    n2641
  );


  xnor
  g2730
  (
    n2757,
    n2723,
    n2650,
    n2728,
    n2713
  );


  nor
  g2731
  (
    n2750,
    n2651,
    n2721,
    n2493,
    n2647
  );


  and
  g2732
  (
    n2756,
    n2486,
    n2494,
    n2640,
    n2729
  );


  xor
  g2733
  (
    n2761,
    n2636,
    n2722,
    n2654,
    n2706
  );


  xnor
  g2734
  (
    n2760,
    n2728,
    n2688,
    n2653,
    n2707
  );


  xor
  g2735
  (
    n2765,
    n2633,
    n2726,
    n2729,
    n2495
  );


  nand
  g2736
  (
    n2746,
    n2665,
    n2705,
    n2730,
    n2494
  );


  and
  g2737
  (
    n2769,
    n2722,
    n2724,
    n2660,
    n2637
  );


  or
  g2738
  (
    n2763,
    n2724,
    n2668,
    n2729,
    n2667
  );


  or
  g2739
  (
    n2747,
    n2721,
    n2632,
    n2728,
    n2490
  );


  not
  g2740
  (
    n2773,
    n2695
  );


  not
  g2741
  (
    n2771,
    n2695
  );


  and
  g2742
  (
    n2775,
    n2695,
    n2695,
    n2694,
    n2696
  );


  xnor
  g2743
  (
    n2774,
    n2745,
    n2696,
    n2746,
    n2747
  );


  xnor
  g2744
  (
    n2772,
    n2749,
    n2748,
    n2696
  );


  or
  g2745
  (
    n2786,
    n2739,
    n2732,
    n2773,
    n2737
  );


  nand
  g2746
  (
    n2790,
    n2738,
    n2773,
    n2737,
    n2774
  );


  and
  g2747
  (
    n2788,
    n2736,
    n2774,
    n2742,
    n2731
  );


  xor
  g2748
  (
    n2787,
    n2731,
    n2771,
    n2737,
    n2734
  );


  xor
  g2749
  (
    n2776,
    n2740,
    n2772,
    n2733,
    n2731
  );


  or
  g2750
  (
    n2785,
    n2731,
    n2734,
    n2732,
    n2736
  );


  nor
  g2751
  (
    n2780,
    n2735,
    n2741,
    n2736
  );


  xor
  g2752
  (
    n2792,
    n2740,
    n2742
  );


  and
  g2753
  (
    n2782,
    n2742,
    n2738,
    n2771,
    n2739
  );


  nor
  g2754
  (
    n2778,
    n2771,
    n2730,
    n2734,
    n2775
  );


  xnor
  g2755
  (
    n2781,
    n2738,
    n2730,
    n2732,
    n2773
  );


  nand
  g2756
  (
    n2784,
    n2740,
    n2772,
    n2743,
    n2736
  );


  or
  g2757
  (
    n2791,
    n2738,
    n2741,
    n2735,
    n2734
  );


  and
  g2758
  (
    n2783,
    n2741,
    n2739,
    n2774,
    n2733
  );


  xnor
  g2759
  (
    n2777,
    n2771,
    n2732,
    n2773,
    n2772
  );


  nor
  g2760
  (
    n2779,
    n2739,
    n2735,
    n2733
  );


  nand
  g2761
  (
    n2789,
    n2737,
    n2772,
    n2774,
    n2735
  );


  nand
  g2762
  (
    n2812,
    n2783,
    n2792
  );


  xor
  g2763
  (
    n2814,
    n2776,
    n2674,
    n2789,
    n2760
  );


  xor
  g2764
  (
    AntiSAT_key_wire,
    n2790,
    n458,
    n2767,
    n2787
  );


  and
  g2765
  (
    n2801,
    n2671,
    n2672,
    n2787,
    n2786
  );


  xor
  g2766
  (
    n2817,
    n2750,
    n2792,
    n2758,
    n2778
  );


  nand
  g2767
  (
    n2818,
    n459,
    n2778,
    n2777,
    n2776
  );


  nand
  g2768
  (
    n2796,
    n458,
    n2785,
    n2755
  );


  nand
  g2769
  (
    n2795,
    n460,
    n2790,
    n458,
    n459
  );


  or
  g2770
  (
    n2804,
    n2776,
    n2763,
    n2792
  );


  nand
  g2771
  (
    n2794,
    n2779,
    n2791,
    n2677,
    n2782
  );


  or
  g2772
  (
    n2805,
    n1747,
    n2670,
    n2791,
    n2786
  );


  nand
  g2773
  (
    n2808,
    n2765,
    n2766,
    n2790,
    n2786
  );


  and
  g2774
  (
    n2802,
    n2751,
    n2768,
    n2770,
    n2787
  );


  xor
  g2775
  (
    n2797,
    n2789,
    n459,
    n460,
    n2783
  );


  xnor
  g2776
  (
    n2811,
    n2753,
    n2791,
    n2784,
    n2790
  );


  and
  g2777
  (
    n2807,
    n2783,
    n2788,
    n2787
  );


  nand
  g2778
  (
    n2806,
    n2781,
    n2778,
    n460,
    n2779
  );


  nor
  g2779
  (
    n2799,
    n2788,
    n2782,
    n2754,
    n2780
  );


  and
  g2780
  (
    n2800,
    n2762,
    n2781,
    n2756,
    n2761
  );


  nor
  g2781
  (
    n2798,
    n2777,
    n2675,
    n2752,
    n2780
  );


  xnor
  g2782
  (
    n2810,
    n2788,
    n2676,
    n459,
    n2764
  );


  xor
  g2783
  (
    n2813,
    n2780,
    n2779,
    n2785
  );


  nand
  g2784
  (
    n2793,
    n2789,
    n457,
    n2784,
    n2769
  );


  nor
  g2785
  (
    n2816,
    n2789,
    n2784,
    n2777,
    n2781
  );


  nor
  g2786
  (
    n2803,
    n458,
    n2759,
    n2757,
    n2791
  );


  and
  g2787
  (
    n2809,
    n2782,
    n2786,
    n2673,
    n460
  );


  and
  g2788
  (
    n2822,
    n2799,
    n2800,
    n2743,
    n2814
  );


  nor
  g2789
  (
    n2820,
    n2815,
    n2807,
    n2805,
    n2802
  );


  nor
  g2790
  (
    n2825,
    n2796,
    n2811,
    n2800
  );


  xor
  g2791
  (
    n2827,
    n2817,
    n2744,
    n2798,
    n2775
  );


  xnor
  g2792
  (
    n2831,
    n2743,
    n2817,
    n2797,
    n2744
  );


  nand
  g2793
  (
    n2830,
    n2804,
    n2810,
    n2816,
    n2818
  );


  nand
  g2794
  (
    n2821,
    n2798,
    n2809,
    n2816,
    n2810
  );


  nand
  g2795
  (
    n2826,
    n2743,
    n2799,
    n2744,
    n2812
  );


  or
  g2796
  (
    n2828,
    n2812,
    n2807,
    n2804,
    n2818
  );


  nor
  g2797
  (
    n2824,
    n2803,
    n2775,
    n2802
  );


  xnor
  g2798
  (
    n2829,
    n2805,
    n2806,
    n2814,
    n2744
  );


  nand
  g2799
  (
    n2823,
    n2806,
    n2808,
    n2813
  );


  xnor
  g2800
  (
    n2819,
    n2813,
    n2801,
    n2809
  );


  and
  g2801
  (
    n2832,
    n2803,
    n2795,
    n2815,
    n2797
  );


  buf
  g2802
  (
    n2840,
    n2825
  );


  not
  g2803
  (
    n2839,
    n461
  );


  buf
  g2804
  (
    n2833,
    n2496
  );


  buf
  g2805
  (
    n2837,
    n2827
  );


  buf
  g2806
  (
    n2835,
    n2826
  );


  buf
  g2807
  (
    n2838,
    n2828
  );


  not
  g2808
  (
    n2841,
    n2824
  );


  nor
  g2809
  (
    n2836,
    n2831,
    n2829,
    n2832
  );


  nor
  g2810
  (
    n2834,
    n2496,
    n461,
    n2830
  );


  not
  g2811
  (
    n2844,
    n2833
  );


  buf
  g2812
  (
    n2845,
    n2834
  );


  buf
  g2813
  (
    n2843,
    n2833
  );


  buf
  g2814
  (
    n2842,
    n2833
  );


  xor
  g2815
  (
    n2847,
    n2837,
    n461,
    n2497,
    n2835
  );


  nor
  g2816
  (
    n2853,
    n2843,
    n2499,
    n25,
    n2836
  );


  nor
  g2817
  (
    n2852,
    n2500,
    n2497,
    n2498,
    n2844
  );


  and
  g2818
  (
    n2849,
    n2834,
    n462,
    n2845
  );


  and
  g2819
  (
    n2850,
    n2844,
    n2835,
    n2836
  );


  nor
  g2820
  (
    n2854,
    n2837,
    n2500,
    n2845,
    n2843
  );


  xnor
  g2821
  (
    n2851,
    n2835,
    n2499,
    n2844,
    n462
  );


  nor
  g2822
  (
    n2846,
    n2837,
    n2498,
    n2834,
    n2845
  );


  and
  g2823
  (
    n2848,
    n2843,
    n462,
    n2836,
    n25
  );


  not
  g2824
  (
    n2856,
    n2853
  );


  buf
  g2825
  (
    n2855,
    n2854
  );


  and
  g2826
  (
    n2859,
    n127,
    n128,
    n2856,
    n464
  );


  xor
  g2827
  (
    n2861,
    n126,
    n127,
    n2856,
    n463
  );


  and
  g2828
  (
    n2860,
    n2856,
    n2855,
    n128,
    n126
  );


  and
  g2829
  (
    n2858,
    n126,
    n127,
    n2856,
    n2855
  );


  and
  g2830
  (
    n2857,
    n127,
    n126,
    n463
  );


  xor
  g2831
  (
    n2862,
    n464,
    n463,
    n2855
  );


  xor
  g2832
  (
    n2864,
    n2840,
    n465,
    n466
  );


  nand
  g2833
  (
    n2866,
    n465,
    n2838,
    n2839,
    n2862
  );


  xnor
  g2834
  (
    n2869,
    n2861,
    n2839,
    n464,
    n2859
  );


  xnor
  g2835
  (
    n2870,
    n2840,
    n465,
    n2838,
    n2841
  );


  xor
  g2836
  (
    n2867,
    n2841,
    n2861,
    n2837,
    n2839
  );


  or
  g2837
  (
    n2865,
    n464,
    n2862,
    n2838,
    n2839
  );


  nand
  g2838
  (
    n2868,
    n2860,
    n2838,
    n2840,
    n2841
  );


  nor
  g2839
  (
    n2863,
    n2860,
    n2840,
    n2859,
    n2841
  );


  nor
  g2840
  (
    n2871,
    n2869,
    n2866,
    n29,
    n2870
  );


  and
  g2841
  (
    n2879,
    n2864,
    n27,
    n468
  );


  nor
  g2842
  (
    n2882,
    n29,
    n30,
    n27
  );


  nor
  g2843
  (
    n2873,
    n26,
    n26,
    n2868,
    n466
  );


  nor
  g2844
  (
    n2877,
    n26,
    n28,
    n2869,
    n2868
  );


  nor
  g2845
  (
    n2884,
    n466,
    n29,
    n2867,
    n2504
  );


  xor
  g2846
  (
    n2883,
    n2866,
    n2868,
    n2867,
    n30
  );


  xnor
  g2847
  (
    n2885,
    n2864,
    n2867,
    n2863,
    n128
  );


  xnor
  g2848
  (
    n2880,
    n467,
    n467,
    n2869,
    n2503
  );


  xnor
  g2849
  (
    n2881,
    n28,
    n28,
    n128,
    n2865
  );


  or
  g2850
  (
    n2872,
    n2866,
    n27,
    n30,
    n28
  );


  or
  g2851
  (
    n2878,
    n2863,
    n467,
    n2502
  );


  nand
  g2852
  (
    n2874,
    n2503,
    n2501,
    n2865,
    n2870
  );


  nor
  g2853
  (
    n2876,
    n466,
    n2870,
    n2501,
    n2865
  );


  nor
  g2854
  (
    n2875,
    n2864,
    n26,
    n29,
    n2502
  );


  not
  g2855
  (
    n2892,
    n2874
  );


  not
  g2856
  (
    n2896,
    n2875
  );


  buf
  g2857
  (
    n2895,
    n2871
  );


  not
  g2858
  (
    n2899,
    n2879
  );


  not
  g2859
  (
    n2886,
    n2877
  );


  buf
  g2860
  (
    n2900,
    n2876
  );


  buf
  g2861
  (
    n2891,
    n2880
  );


  buf
  g2862
  (
    n2893,
    n2878
  );


  not
  g2863
  (
    n2897,
    n2875
  );


  not
  g2864
  (
    n2890,
    n2873
  );


  not
  g2865
  (
    n2894,
    n2871
  );


  not
  g2866
  (
    n2888,
    n2878
  );


  xnor
  g2867
  (
    n2887,
    n2877,
    n2873,
    n2876
  );


  nand
  g2868
  (
    n2898,
    n2874,
    n2872,
    n2877,
    n2879
  );


  or
  g2869
  (
    n2901,
    n2875,
    n2876,
    n2872
  );


  nand
  g2870
  (
    n2889,
    n2879,
    n2871,
    n2874,
    n2878
  );


  buf
  g2871
  (
    n2907,
    n2887
  );


  not
  g2872
  (
    n2906,
    n2890
  );


  not
  g2873
  (
    n2913,
    n2886
  );


  buf
  g2874
  (
    n2912,
    n2887
  );


  buf
  g2875
  (
    n2905,
    n2891
  );


  buf
  g2876
  (
    n2908,
    n2889
  );


  not
  g2877
  (
    n2904,
    n2889
  );


  buf
  g2878
  (
    n2909,
    n2886
  );


  not
  g2879
  (
    n2910,
    n2891
  );


  not
  g2880
  (
    n2902,
    n2890
  );


  buf
  g2881
  (
    n2903,
    n2888
  );


  not
  g2882
  (
    n2911,
    n2888
  );


  buf
  g2883
  (
    n2914,
    n2902
  );


  not
  g2884
  (
    n2915,
    n2902
  );


  nor
  g2885
  (
    n2916,
    n2903,
    n2903,
    n2915,
    n2902
  );


  nand
  g2886
  (
    n2920,
    n2903,
    n2916,
    n2904
  );


  nand
  g2887
  (
    n2919,
    n2906,
    n2904,
    n2903
  );


  nand
  g2888
  (
    n2918,
    n2916,
    n2905,
    n2904
  );


  nand
  g2889
  (
    n2917,
    n2906,
    n2916,
    n2905
  );


  nand
  g2890
  (
    n2922,
    n2896,
    n2906,
    n2893,
    n2901
  );


  nor
  g2891
  (
    n2932,
    n2920,
    n2900,
    n2884,
    n2679
  );


  nor
  g2892
  (
    n2925,
    n2892,
    n2883,
    n2918,
    n2880
  );


  nand
  g2893
  (
    n2930,
    n2919,
    n2920,
    n2881,
    n2899
  );


  nand
  g2894
  (
    n2926,
    n2880,
    n468,
    n2918,
    n2899
  );


  and
  g2895
  (
    n2924,
    n2917,
    n2882,
    n2895,
    n2919
  );


  xnor
  g2896
  (
    n2923,
    n2917,
    n2883,
    n2894,
    n2885
  );


  nand
  g2897
  (
    n2929,
    n2897,
    n2895,
    n2918,
    n2917
  );


  xnor
  g2898
  (
    n2935,
    n2920,
    n2885,
    n2896,
    n2881
  );


  and
  g2899
  (
    n2934,
    n2884,
    n2919,
    n2901
  );


  xor
  g2900
  (
    n2933,
    n2504,
    n468,
    n2882
  );


  xnor
  g2901
  (
    n2928,
    n2918,
    n2882,
    n2897,
    n2881
  );


  nand
  g2902
  (
    n2927,
    n2893,
    n2901,
    n2885,
    n2898
  );


  xnor
  g2903
  (
    n2931,
    n2884,
    n2892,
    n2920,
    n2894
  );


  and
  g2904
  (
    n2921,
    n2900,
    n2898,
    n2678,
    n2883
  );


  nand
  g2905
  (
    n2946,
    n2913,
    n2912,
    n2909
  );


  and
  g2906
  (
    n2937,
    n2910,
    n2931,
    n2929,
    n2912
  );


  xnor
  g2907
  (
    n2939,
    n2933,
    n2930,
    n2928,
    n2912
  );


  and
  g2908
  (
    n2940,
    n2913,
    n2912,
    n2907,
    n2911
  );


  xnor
  g2909
  (
    n2945,
    n2907,
    n2907,
    n2932,
    n2910
  );


  nor
  g2910
  (
    n2942,
    n2909,
    n2906,
    n2907,
    n2934
  );


  xor
  g2911
  (
    n2936,
    n2910,
    n2929,
    n2932,
    n2911
  );


  xnor
  g2912
  (
    n2943,
    n2935,
    n2908,
    n2913,
    n2930
  );


  nor
  g2913
  (
    n2938,
    n2908,
    n2910,
    n2931,
    n2911
  );


  xor
  g2914
  (
    n2941,
    n2935,
    n2908,
    n2934
  );


  nor
  g2915
  (
    n2944,
    n2911,
    n2909,
    n2933,
    n2913
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_30
  (
    gbar_input_0_0,
    keyIn_0_30,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_31
  (
    gbar_input_0_1,
    keyIn_0_31,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_2,
    keyIn_0_32,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_3,
    keyIn_0_33,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_4,
    keyIn_0_34,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_5,
    keyIn_0_35,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_6,
    keyIn_0_36,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_7,
    keyIn_0_37,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_8,
    keyIn_0_38,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_9,
    keyIn_0_39,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_10,
    keyIn_0_40,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_11,
    keyIn_0_41,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_12,
    keyIn_0_42,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_13,
    keyIn_0_43,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_14,
    keyIn_0_44,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_15,
    keyIn_0_45,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_16,
    keyIn_0_46,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_17,
    keyIn_0_47,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_18,
    keyIn_0_48,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_19,
    keyIn_0_49,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_20,
    keyIn_0_50,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_21,
    keyIn_0_51,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_22,
    keyIn_0_52,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_23,
    keyIn_0_53,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_24,
    keyIn_0_54,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_25,
    keyIn_0_55,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_26,
    keyIn_0_56,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_27,
    keyIn_0_57,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_28,
    keyIn_0_58,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_29,
    keyIn_0_59,
    n30
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n2815,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

