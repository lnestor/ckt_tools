// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_205 written by SynthGen on 2021/04/05 11:08:36
module Stat_1000_205( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n174, n148, n179, n165, n178, n151, n168, n139,
 n194, n150, n186, n124, n181, n147, n135, n182,
 n601, n613, n610, n611, n598, n608, n623, n605,
 n621, n602, n620, n606, n617, n622, n1031, n1032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n174, n148, n179, n165, n178, n151, n168, n139,
 n194, n150, n186, n124, n181, n147, n135, n182,
 n601, n613, n610, n611, n598, n608, n623, n605,
 n621, n602, n620, n606, n617, n622, n1031, n1032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n136, n137, n138,
 n140, n141, n142, n143, n144, n145, n146, n149,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n166, n167, n169,
 n170, n171, n172, n173, n175, n176, n177, n180,
 n183, n184, n185, n187, n188, n189, n190, n191,
 n192, n193, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n599, n600, n603,
 n604, n607, n609, n612, n614, n615, n616, n618,
 n619, n624, n625, n626, n627, n628, n629, n630,
 n631, n632, n633, n634, n635, n636, n637, n638,
 n639, n640, n641, n642, n643, n644, n645, n646,
 n647, n648, n649, n650, n651, n652, n653, n654,
 n655, n656, n657, n658, n659, n660, n661, n662,
 n663, n664, n665, n666, n667, n668, n669, n670,
 n671, n672, n673, n674, n675, n676, n677, n678,
 n679, n680, n681, n682, n683, n684, n685, n686,
 n687, n688, n689, n690, n691, n692, n693, n694,
 n695, n696, n697, n698, n699, n700, n701, n702,
 n703, n704, n705, n706, n707, n708, n709, n710,
 n711, n712, n713, n714, n715, n716, n717, n718,
 n719, n720, n721, n722, n723, n724, n725, n726,
 n727, n728, n729, n730, n731, n732, n733, n734,
 n735, n736, n737, n738, n739, n740, n741, n742,
 n743, n744, n745, n746, n747, n748, n749, n750,
 n751, n752, n753, n754, n755, n756, n757, n758,
 n759, n760, n761, n762, n763, n764, n765, n766,
 n767, n768, n769, n770, n771, n772, n773, n774,
 n775, n776, n777, n778, n779, n780, n781, n782,
 n783, n784, n785, n786, n787, n788, n789, n790,
 n791, n792, n793, n794, n795, n796, n797, n798,
 n799, n800, n801, n802, n803, n804, n805, n806,
 n807, n808, n809, n810, n811, n812, n813, n814,
 n815, n816, n817, n818, n819, n820, n821, n822,
 n823, n824, n825, n826, n827, n828, n829, n830,
 n831, n832, n833, n834, n835, n836, n837, n838,
 n839, n840, n841, n842, n843, n844, n845, n846,
 n847, n848, n849, n850, n851, n852, n853, n854,
 n855, n856, n857, n858, n859, n860, n861, n862,
 n863, n864, n865, n866, n867, n868, n869, n870,
 n871, n872, n873, n874, n875, n876, n877, n878,
 n879, n880, n881, n882, n883, n884, n885, n886,
 n887, n888, n889, n890, n891, n892, n893, n894,
 n895, n896, n897, n898, n899, n900, n901, n902,
 n903, n904, n905, n906, n907, n908, n909, n910,
 n911, n912, n913, n914, n915, n916, n917, n918,
 n919, n920, n921, n922, n923, n924, n925, n926,
 n927, n928, n929, n930, n931, n932, n933, n934,
 n935, n936, n937, n938, n939, n940, n941, n942,
 n943, n944, n945, n946, n947, n948, n949, n950,
 n951, n952, n953, n954, n955, n956, n957, n958,
 n959, n960, n961, n962, n963, n964, n965, n966,
 n967, n968, n969, n970, n971, n972, n973, n974,
 n975, n976, n977, n978, n979, n980, n981, n982,
 n983, n984, n985, n986, n987, n988, n989, n990,
 n991, n992, n993, n994, n995, n996, n997, n998,
 n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
 n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
 n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
 n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030;

not  g0 (n87, n14);
buf  g1 (n68, n17);
not  g2 (n103, n14);
not  g3 (n62, n2);
not  g4 (n56, n21);
not  g5 (n34, n20);
buf  g6 (n49, n9);
not  g7 (n53, n20);
not  g8 (n72, n18);
not  g9 (n117, n16);
not  g10 (n40, n6);
buf  g11 (n79, n19);
not  g12 (n71, n21);
not  g13 (n108, n13);
buf  g14 (n69, n9);
buf  g15 (n102, n6);
buf  g16 (n74, n5);
buf  g17 (n38, n8);
buf  g18 (n80, n10);
buf  g19 (n43, n15);
buf  g20 (n41, n13);
buf  g21 (n110, n22);
buf  g22 (n46, n23);
buf  g23 (n115, n11);
not  g24 (n113, n4);
not  g25 (n70, n6);
buf  g26 (n47, n3);
buf  g27 (n109, n4);
not  g28 (n54, n23);
not  g29 (n86, n15);
buf  g30 (n84, n23);
not  g31 (n52, n6);
not  g32 (n101, n7);
not  g33 (n111, n7);
buf  g34 (n104, n21);
not  g35 (n78, n15);
buf  g36 (n100, n17);
not  g37 (n37, n11);
buf  g38 (n67, n8);
buf  g39 (n61, n15);
not  g40 (n94, n17);
not  g41 (n95, n9);
not  g42 (n96, n5);
not  g43 (n57, n12);
not  g44 (n90, n24);
not  g45 (n33, n9);
not  g46 (n58, n13);
buf  g47 (n98, n22);
buf  g48 (n83, n19);
not  g49 (n92, n20);
buf  g50 (n105, n5);
buf  g51 (n35, n10);
not  g52 (n114, n16);
not  g53 (n44, n10);
buf  g54 (n75, n23);
not  g55 (n89, n7);
buf  g56 (n76, n17);
buf  g57 (n106, n12);
not  g58 (n59, n14);
not  g59 (n107, n4);
not  g60 (n55, n11);
buf  g61 (n60, n18);
buf  g62 (n42, n18);
not  g63 (n77, n19);
not  g64 (n88, n1);
buf  g65 (n39, n21);
not  g66 (n66, n12);
not  g67 (n64, n14);
not  g68 (n48, n22);
not  g69 (n91, n11);
buf  g70 (n45, n4);
buf  g71 (n51, n8);
not  g72 (n85, n24);
not  g73 (n93, n8);
buf  g74 (n63, n13);
not  g75 (n116, n10);
not  g76 (n81, n16);
not  g77 (n73, n19);
not  g78 (n112, n20);
not  g79 (n65, n22);
buf  g80 (n36, n5);
buf  g81 (n97, n7);
buf  g82 (n82, n12);
buf  g83 (n99, n16);
not  g84 (n50, n18);
not  g85 (n168, n63);
not  g86 (n165, n75);
buf  g87 (n150, n73);
buf  g88 (n123, n72);
not  g89 (n185, n56);
buf  g90 (n162, n48);
buf  g91 (n158, n56);
buf  g92 (n147, n46);
not  g93 (n166, n53);
buf  g94 (n181, n56);
not  g95 (n132, n65);
not  g96 (n159, n68);
buf  g97 (n167, n54);
not  g98 (n155, n41);
buf  g99 (n153, n59);
not  g100 (n136, n75);
not  g101 (n143, n52);
not  g102 (n175, n63);
not  g103 (n188, n53);
buf  g104 (n193, n63);
not  g105 (n157, n74);
buf  g106 (n196, n62);
buf  g107 (n137, n53);
buf  g108 (n124, n75);
not  g109 (n141, n64);
not  g110 (n135, n70);
buf  g111 (n133, n61);
not  g112 (n118, n55);
not  g113 (n179, n67);
buf  g114 (n160, n68);
buf  g115 (n119, n42);
buf  g116 (n184, n50);
buf  g117 (n134, n74);
buf  g118 (n126, n35);
buf  g119 (n120, n53);
not  g120 (n163, n61);
not  g121 (n170, n77);
buf  g122 (n194, n67);
not  g123 (n145, n70);
not  g124 (n177, n45);
not  g125 (n142, n46);
buf  g126 (n169, n57);
not  g127 (n139, n57);
buf  g128 (n171, n50);
buf  g129 (n195, n36);
not  g130 (n154, n49);
buf  g131 (n122, n50);
buf  g132 (n149, n52);
not  g133 (n173, n61);
buf  g134 (n144, n76);
not  g135 (n176, n64);
buf  g136 (n183, n47);
buf  g137 (n131, n59);
buf  g138 (n191, n72);
not  g139 (n182, n59);
buf  g140 (n121, n60);
buf  g141 (n125, n50);
not  g142 (n129, n60);
buf  g143 (n128, n58);
nand g144 (n192, n58, n55, n76, n74);
nor  g145 (n146, n40, n62, n54, n77);
or   g146 (n127, n73, n72, n51, n54);
and  g147 (n172, n51, n65, n57, n70);
nor  g148 (n164, n62, n66, n67, n46);
or   g149 (n180, n65, n37, n69, n44);
and  g150 (n174, n70, n51, n72, n65);
nor  g151 (n189, n62, n49, n74, n46);
or   g152 (n156, n68, n68, n73, n33);
or   g153 (n148, n52, n55, n39, n48);
nand g154 (n151, n59, n71, n64, n38);
nor  g155 (n152, n49, n47, n76, n58);
xor  g156 (n161, n73, n71, n66, n43);
xnor g157 (n190, n48, n54, n60, n75);
or   g158 (n178, n48, n66, n58, n47);
nor  g159 (n187, n67, n76, n69, n60);
xor  g160 (n130, n57, n71, n56, n63);
or   g161 (n186, n49, n66, n69, n34);
nor  g162 (n138, n52, n69, n47, n61);
xor  g163 (n140, n55, n71, n64, n51);
not  g164 (n217, n162);
buf  g165 (n212, n28);
not  g166 (n221, n29);
buf  g167 (n199, n79);
not  g168 (n252, n158);
buf  g169 (n232, n25);
not  g170 (n234, n194);
buf  g171 (n229, n79);
not  g172 (n250, n177);
not  g173 (n254, n129);
not  g174 (n211, n182);
buf  g175 (n264, n178);
not  g176 (n244, n146);
buf  g177 (n240, n30);
buf  g178 (n262, n148);
not  g179 (n245, n77);
not  g180 (n243, n183);
not  g181 (n201, n153);
buf  g182 (n270, n125);
buf  g183 (n225, n144);
not  g184 (n215, n124);
not  g185 (n213, n136);
buf  g186 (n220, n163);
buf  g187 (n228, n152);
not  g188 (n236, n128);
not  g189 (n266, n195);
buf  g190 (n202, n137);
buf  g191 (n198, n150);
not  g192 (n257, n26);
buf  g193 (n261, n78);
buf  g194 (n248, n196);
not  g195 (n241, n142);
buf  g196 (n223, n30);
buf  g197 (n269, n191);
not  g198 (n230, n31);
not  g199 (n226, n186);
buf  g200 (n246, n30);
not  g201 (n216, n24);
buf  g202 (n203, n161);
buf  g203 (n222, n176);
buf  g204 (n204, n138);
buf  g205 (n206, n31);
buf  g206 (n259, n25);
buf  g207 (n210, n30);
buf  g208 (n209, n78);
not  g209 (n238, n193);
buf  g210 (n251, n132);
not  g211 (n258, n80);
not  g212 (n242, n31);
buf  g213 (n205, n164);
buf  g214 (n208, n160);
not  g215 (n255, n156);
or   g216 (n263, n174, n135, n143);
nor  g217 (n227, n26, n27, n79);
nand g218 (n197, n78, n175, n145);
or   g219 (n267, n187, n184, n181);
nor  g220 (n256, n170, n185, n31);
xnor g221 (n268, n192, n141, n28);
and  g222 (n249, n189, n126, n32);
nand g223 (n200, n127, n78, n80);
xor  g224 (n218, n26, n155, n168);
and  g225 (n207, n171, n29);
xnor g226 (n237, n159, n180, n147);
nor  g227 (n239, n134, n25, n139);
or   g228 (n224, n133, n77, n190);
xnor g229 (n253, n29, n28, n79);
xnor g230 (n260, n27, n130, n165);
nand g231 (n219, n26, n140, n172);
xnor g232 (n233, n166, n167, n27);
nor  g233 (n247, n157, n169, n173);
nand g234 (n235, n123, n28, n179);
xor  g235 (n231, n32, n131, n154);
nor  g236 (n265, n27, n149, n24);
nor  g237 (n214, n188, n151, n25);
not  g238 (n438, n99);
buf  g239 (n393, n253);
not  g240 (n428, n98);
buf  g241 (n374, n242);
not  g242 (n408, n236);
not  g243 (n354, n248);
buf  g244 (n353, n229);
not  g245 (n467, n84);
buf  g246 (n497, n90);
buf  g247 (n361, n234);
buf  g248 (n494, n101);
not  g249 (n462, n199);
not  g250 (n471, n94);
buf  g251 (n477, n222);
not  g252 (n420, n208);
buf  g253 (n454, n234);
not  g254 (n280, n235);
not  g255 (n401, n97);
not  g256 (n434, n86);
buf  g257 (n414, n109);
not  g258 (n271, n227);
buf  g259 (n491, n228);
buf  g260 (n440, n264);
buf  g261 (n368, n250);
buf  g262 (n415, n200);
not  g263 (n444, n242);
not  g264 (n395, n84);
not  g265 (n335, n253);
buf  g266 (n442, n95);
not  g267 (n389, n224);
not  g268 (n383, n229);
buf  g269 (n480, n102);
not  g270 (n476, n233);
buf  g271 (n326, n105);
not  g272 (n288, n81);
buf  g273 (n452, n198);
buf  g274 (n427, n202);
not  g275 (n329, n226);
not  g276 (n364, n82);
not  g277 (n313, n104);
buf  g278 (n423, n241);
not  g279 (n449, n262);
not  g280 (n277, n243);
buf  g281 (n330, n209);
not  g282 (n299, n242);
buf  g283 (n404, n245);
buf  g284 (n490, n99);
not  g285 (n387, n109);
buf  g286 (n338, n213);
not  g287 (n465, n262);
buf  g288 (n334, n241);
buf  g289 (n390, n99);
not  g290 (n314, n251);
not  g291 (n296, n239);
buf  g292 (n429, n231);
buf  g293 (n402, n259);
not  g294 (n397, n248);
not  g295 (n304, n207);
not  g296 (n370, n270);
not  g297 (n424, n106);
buf  g298 (n305, n256);
not  g299 (n486, n110);
not  g300 (n351, n239);
not  g301 (n275, n243);
buf  g302 (n413, n266);
buf  g303 (n483, n265);
not  g304 (n484, n255);
not  g305 (n380, n218);
not  g306 (n410, n101);
buf  g307 (n306, n85);
not  g308 (n436, n232);
not  g309 (n391, n211);
buf  g310 (n367, n230);
not  g311 (n324, n254);
not  g312 (n307, n265);
buf  g313 (n319, n232);
not  g314 (n336, n257);
not  g315 (n388, n219);
buf  g316 (n282, n103);
not  g317 (n355, n263);
not  g318 (n312, n233);
buf  g319 (n430, n264);
not  g320 (n488, n100);
not  g321 (n362, n237);
not  g322 (n448, n233);
buf  g323 (n371, n214);
buf  g324 (n341, n261);
buf  g325 (n495, n90);
buf  g326 (n392, n221);
not  g327 (n381, n258);
buf  g328 (n283, n93);
buf  g329 (n363, n252);
buf  g330 (n350, n241);
not  g331 (n375, n87);
not  g332 (n399, n208);
not  g333 (n287, n206);
buf  g334 (n366, n239);
not  g335 (n333, n260);
not  g336 (n411, n247);
not  g337 (n400, n228);
buf  g338 (n455, n110);
buf  g339 (n479, n244);
not  g340 (n281, n96);
buf  g341 (n446, n94);
not  g342 (n472, n265);
not  g343 (n365, n213);
buf  g344 (n290, n254);
not  g345 (n273, n204);
buf  g346 (n496, n224);
buf  g347 (n426, n106);
buf  g348 (n403, n204);
buf  g349 (n385, n86);
not  g350 (n372, n229);
buf  g351 (n318, n247);
not  g352 (n422, n249);
not  g353 (n456, n230);
buf  g354 (n379, n253);
not  g355 (n396, n102);
not  g356 (n492, n103);
buf  g357 (n487, n109);
buf  g358 (n441, n106);
not  g359 (n316, n205);
not  g360 (n382, n108);
not  g361 (n289, n92);
buf  g362 (n322, n232);
not  g363 (n278, n251);
buf  g364 (n466, n212);
buf  g365 (n356, n100);
not  g366 (n418, n261);
buf  g367 (n344, n97);
not  g368 (n447, n84);
buf  g369 (n272, n268);
not  g370 (n464, n265);
not  g371 (n274, n89);
buf  g372 (n310, n108);
buf  g373 (n470, n270);
buf  g374 (n332, n105);
not  g375 (n433, n223);
buf  g376 (n352, n215);
not  g377 (n419, n89);
buf  g378 (n405, n106);
not  g379 (n317, n227);
buf  g380 (n417, n215);
not  g381 (n302, n235);
not  g382 (n489, n97);
not  g383 (n345, n232);
buf  g384 (n359, n110);
buf  g385 (n386, n259);
buf  g386 (n327, n246);
not  g387 (n321, n95);
buf  g388 (n349, n255);
not  g389 (n279, n86);
not  g390 (n340, n268);
not  g391 (n298, n85);
buf  g392 (n377, n81);
not  g393 (n445, n91);
not  g394 (n308, n217);
not  g395 (n478, n248);
buf  g396 (n421, n235);
buf  g397 (n301, n107);
not  g398 (n431, n230);
not  g399 (n311, n269);
not  g400 (n407, n205);
buf  g401 (n451, n262);
buf  g402 (n343, n105);
buf  g403 (n463, n236);
buf  g404 (n291, n210);
buf  g405 (n346, n231);
not  g406 (n315, n266);
not  g407 (n384, n97);
not  g408 (n457, n212);
buf  g409 (n303, n258);
not  g410 (n460, n240);
not  g411 (n328, n85);
not  g412 (n453, n228);
not  g413 (n450, n92);
buf  g414 (n300, n95);
not  g415 (n323, n94);
buf  g416 (n295, n201);
buf  g417 (n376, n259);
not  g418 (n475, n237);
buf  g419 (n294, n256);
buf  g420 (n468, n216);
buf  g421 (n412, n245);
not  g422 (n276, n108);
buf  g423 (n409, n90);
and  g424 (n459, n84, n222);
nor  g425 (n439, n82, n98, n250, n260);
nand g426 (n432, n268, n236, n251, n233);
nand g427 (n284, n107, n259, n231, n267);
xor  g428 (n378, n255, n85, n80, n269);
nor  g429 (n360, n226, n254, n266);
and  g430 (n493, n100, n245, n257, n95);
and  g431 (n297, n83, n82, n87, n91);
and  g432 (n425, n255, n107, n240, n92);
nand g433 (n285, n98, n108, n238, n223);
nor  g434 (n416, n234, n96, n237, n264);
nor  g435 (n320, n104, n245, n218, n225);
xnor g436 (n481, n239, n241, n105, n92);
xnor g437 (n342, n96, n104, n263, n94);
or   g438 (n293, n261, n250, n257, n91);
or   g439 (n461, n98, n89, n263, n221);
xor  g440 (n325, n249, n269, n246, n253);
and  g441 (n485, n100, n83, n90, n88);
or   g442 (n443, n209, n99, n249, n88);
xor  g443 (n398, n268, n87, n235, n230);
and  g444 (n358, n263, n270, n81, n210);
or   g445 (n339, n219, n93, n91, n270);
or   g446 (n394, n248, n261, n211, n249);
nor  g447 (n406, n254, n238, n203, n243);
or   g448 (n482, n267, n225, n238, n103);
and  g449 (n458, n220, n247, n206, n229);
xor  g450 (n331, n246, n217, n260, n236);
or   g451 (n357, n247, n197, n82, n252);
nand g452 (n369, n101, n252, n244, n264);
and  g453 (n337, n81, n207, n258, n256);
and  g454 (n435, n267, n214, n252, n107);
nor  g455 (n473, n267, n251, n87, n88);
nor  g456 (n347, n240, n101, n244, n109);
or   g457 (n437, n220, n244, n269, n93);
nand g458 (n292, n256, n83, n250, n231);
or   g459 (n373, n243, n88, n102, n260);
nor  g460 (n309, n103, n89, n83, n234);
or   g461 (n474, n262, n104, n240, n228);
nand g462 (n469, n242, n216, n96, n257);
xor  g463 (n348, n238, n93, n80, n237);
and  g464 (n286, n246, n258, n86, n102);
buf  g465 (n527, n275);
not  g466 (n511, n291);
buf  g467 (n528, n285);
not  g468 (n522, n283);
buf  g469 (n512, n300);
not  g470 (n521, n279);
buf  g471 (n506, n293);
buf  g472 (n513, n276);
buf  g473 (n504, n278);
not  g474 (n499, n286);
not  g475 (n516, n296);
buf  g476 (n503, n290);
not  g477 (n523, n284);
not  g478 (n520, n274);
buf  g479 (n517, n271);
not  g480 (n500, n280);
not  g481 (n507, n287);
not  g482 (n501, n298);
buf  g483 (n519, n282);
not  g484 (n518, n277);
not  g485 (n505, n288);
buf  g486 (n515, n289);
buf  g487 (n526, n302);
buf  g488 (n508, n297);
not  g489 (n525, n281);
not  g490 (n498, n292);
buf  g491 (n509, n272);
buf  g492 (n524, n294);
buf  g493 (n502, n273);
not  g494 (n514, n299);
buf  g495 (n529, n301);
buf  g496 (n510, n295);
not  g497 (n566, n501);
not  g498 (n558, n514);
buf  g499 (n559, n506);
buf  g500 (n544, n505);
not  g501 (n569, n499);
buf  g502 (n568, n498);
not  g503 (n563, n508);
not  g504 (n545, n508);
buf  g505 (n553, n511);
not  g506 (n530, n498);
not  g507 (n540, n512);
not  g508 (n531, n506);
not  g509 (n535, n502);
not  g510 (n561, n506);
buf  g511 (n549, n111);
buf  g512 (n552, n499);
buf  g513 (n536, n512);
buf  g514 (n541, n510);
not  g515 (n548, n506);
not  g516 (n550, n511);
buf  g517 (n538, n505);
buf  g518 (n537, n510);
buf  g519 (n560, n503);
not  g520 (n554, n498);
buf  g521 (n567, n503);
not  g522 (n562, n500);
nand g523 (n556, n513, n503);
xor  g524 (n557, n515, n513);
and  g525 (n555, n511, n514, n508, n515);
or   g526 (n534, n515, n507, n511, n508);
or   g527 (n547, n502, n507, n110, n505);
nor  g528 (n533, n500, n509, n502, n501);
nor  g529 (n564, n516, n498, n510, n505);
or   g530 (n546, n507, n509, n514, n512);
or   g531 (n565, n510, n507, n499, n512);
or   g532 (n551, n509, n500, n504);
nand g533 (n539, n501, n502, n516, n513);
nand g534 (n543, n509, n504, n499, n501);
nand g535 (n542, n513, n111, n516, n500);
nand g536 (n532, n514, n515, n503, n504);
not  g537 (n570, n542);
buf  g538 (n578, n532);
buf  g539 (n583, n531);
not  g540 (n575, n535);
not  g541 (n572, n530);
not  g542 (n584, n536);
not  g543 (n574, n541);
not  g544 (n571, n537);
buf  g545 (n573, n543);
not  g546 (n576, n533);
not  g547 (n585, n534);
buf  g548 (n579, n539);
buf  g549 (n581, n545);
buf  g550 (n582, n544);
not  g551 (n580, n540);
not  g552 (n577, n538);
buf  g553 (n587, n304);
buf  g554 (n594, n576);
buf  g555 (n595, n305);
not  g556 (n588, n578);
nor  g557 (n591, n573, n303);
xor  g558 (n589, n306, n570);
and  g559 (n593, n571, n572);
and  g560 (n586, n575, n579);
xnor g561 (n592, n577, n111);
nor  g562 (n590, n574, n111);
not  g563 (n608, n516);
not  g564 (n599, n590);
not  g565 (n613, n592);
not  g566 (n612, n588);
not  g567 (n601, n587);
not  g568 (n606, n590);
buf  g569 (n609, n587);
not  g570 (n617, n590);
buf  g571 (n623, n593);
not  g572 (n596, n591);
not  g573 (n610, n589);
buf  g574 (n598, n588);
buf  g575 (n614, n589);
not  g576 (n615, n586);
buf  g577 (n604, n586);
not  g578 (n616, n591);
not  g579 (n620, n592);
buf  g580 (n619, n589);
not  g581 (n602, n593);
buf  g582 (n618, n587);
buf  g583 (n605, n587);
not  g584 (n622, n588);
buf  g585 (n624, n517);
buf  g586 (n625, n591);
not  g587 (n597, n590);
buf  g588 (n621, n588);
buf  g589 (n603, n586);
buf  g590 (n607, n586);
buf  g591 (n600, n592);
nor  g592 (n611, n591, n592, n589);
buf  g593 (n631, n313);
buf  g594 (n637, n551);
buf  g595 (n629, n552);
buf  g596 (n636, n563);
or   g597 (n630, n564, n615, n549, n613);
and  g598 (n627, n311, n557, n610, n618);
or   g599 (n632, n619, n585, n622, n546);
xor  g600 (n634, n556, n555, n580, n560);
nand g601 (n638, n620, n582, n307, n616);
xor  g602 (n628, n553, n562, n315, n581);
or   g603 (n635, n617, n312, n316, n317);
and  g604 (n633, n314, n561, n548, n624);
nor  g605 (n626, n583, n547, n612, n310);
xnor g606 (n640, n614, n584, n550, n621);
nor  g607 (n639, n309, n559, n623, n554);
nand g608 (n641, n611, n308, n558, n625);
not  g609 (n644, n631);
buf  g610 (n647, n630);
buf  g611 (n643, n629);
buf  g612 (n650, n628);
buf  g613 (n649, n323);
buf  g614 (n646, n632);
not  g615 (n651, n320);
not  g616 (n642, n322);
and  g617 (n645, n319, n626, n318, n629);
or   g618 (n648, n630, n627, n631, n321);
not  g619 (n661, n648);
buf  g620 (n654, n646);
nor  g621 (n653, n645, n326, n651, n334);
xnor g622 (n656, n333, n642, n644, n518);
and  g623 (n657, n332, n325, n517);
nor  g624 (n655, n335, n329, n520, n519);
nand g625 (n652, n328, n519, n518, n651);
and  g626 (n658, n647, n643, n650, n519);
or   g627 (n660, n518, n518, n331, n520);
xor  g628 (n662, n520, n519, n324, n327);
nand g629 (n659, n517, n520, n330, n649);
buf  g630 (n667, n638);
buf  g631 (n673, n568);
buf  g632 (n702, n633);
not  g633 (n697, n659);
not  g634 (n703, n344);
not  g635 (n688, n566);
not  g636 (n704, n639);
buf  g637 (n666, n113);
buf  g638 (n680, n657);
buf  g639 (n699, n662);
buf  g640 (n692, n656);
buf  g641 (n690, n653);
not  g642 (n681, n654);
not  g643 (n685, n112);
buf  g644 (n686, n112);
buf  g645 (n678, n654);
not  g646 (n689, n652);
not  g647 (n705, n658);
buf  g648 (n693, n660);
buf  g649 (n683, n640);
buf  g650 (n675, n113);
not  g651 (n665, n637);
buf  g652 (n677, n660);
buf  g653 (n701, n635);
not  g654 (n679, n634);
buf  g655 (n663, n636);
and  g656 (n695, n658, n347, n661, n345);
nand g657 (n698, n338, n343, n662);
nor  g658 (n694, n112, n653, n641);
xor  g659 (n669, n639, n661, n635, n640);
or   g660 (n691, n636, n348, n653, n654);
nand g661 (n706, n652, n354, n353, n340);
nand g662 (n676, n656, n652, n339, n352);
nor  g663 (n664, n641, n351, n652, n569);
xnor g664 (n671, n341, n659, n655, n657);
and  g665 (n672, n656, n634, n655);
and  g666 (n682, n637, n114, n342, n349);
nor  g667 (n696, n337, n657, n658);
and  g668 (n670, n350, n654, n632, n656);
or   g669 (n668, n638, n355, n659, n567);
nor  g670 (n674, n346, n662, n565, n660);
xor  g671 (n700, n336, n655, n661, n113);
nor  g672 (n684, n113, n660, n114, n633);
and  g673 (n687, n657, n661, n659, n112);
nor  g674 (n747, n464, n436, n473, n684);
and  g675 (n744, n474, n454, n448, n463);
xnor g676 (n746, n389, n481, n356, n415);
and  g677 (n728, n467, n685, n452, n381);
and  g678 (n709, n453, n481, n458, n444);
and  g679 (n754, n479, n663, n373, n482);
xor  g680 (n712, n486, n694, n469, n693);
and  g681 (n742, n363, n691, n382, n686);
xor  g682 (n768, n688, n455, n458, n478);
nor  g683 (n745, n457, n476, n695, n452);
nand g684 (n753, n481, n685, n466, n693);
and  g685 (n740, n372, n683, n692, n481);
nor  g686 (n785, n446, n687, n406, n423);
or   g687 (n711, n429, n681, n689, n470);
nor  g688 (n765, n485, n487, n455, n365);
and  g689 (n735, n433, n469, n487, n402);
xor  g690 (n770, n439, n370, n443, n690);
xnor g691 (n707, n412, n692, n394, n671);
or   g692 (n763, n366, n479, n453, n386);
xor  g693 (n760, n692, n420, n427, n694);
nand g694 (n714, n688, n404, n418, n486);
and  g695 (n773, n459, n688, n457, n484);
and  g696 (n741, n424, n673, n685, n475);
or   g697 (n776, n422, n395, n474, n469);
or   g698 (n772, n466, n689, n442, n683);
or   g699 (n736, n425, n387, n460, n691);
xor  g700 (n748, n447, n693, n465, n455);
xnor g701 (n771, n397, n441, n377, n446);
and  g702 (n758, n362, n456, n470, n467);
nor  g703 (n780, n693, n694, n376, n477);
or   g704 (n775, n449, n476, n459, n695);
xnor g705 (n731, n385, n676, n691, n480);
xor  g706 (n730, n485, n692, n465, n411);
or   g707 (n749, n465, n485, n471, n478);
xor  g708 (n743, n468, n456, n681, n460);
nand g709 (n764, n407, n694, n487, n484);
xor  g710 (n724, n431, n450, n674, n413);
and  g711 (n729, n438, n446, n368, n448);
xor  g712 (n738, n393, n419, n483, n461);
xor  g713 (n786, n375, n447, n474, n484);
xor  g714 (n727, n401, n690, n450, n379);
nand g715 (n719, n471, n687, n417, n400);
or   g716 (n721, n440, n677, n408, n484);
xnor g717 (n722, n460, n468, n388, n467);
nand g718 (n732, n466, n472, n688);
xnor g719 (n781, n434, n696, n390, n462);
nand g720 (n774, n474, n432, n680, n687);
xnor g721 (n710, n462, n684, n454, n686);
and  g722 (n769, n384, n480, n478, n471);
nor  g723 (n756, n466, n683, n396, n691);
or   g724 (n761, n416, n695, n479, n469);
xnor g725 (n708, n409, n430, n684, n453);
xor  g726 (n767, n398, n482, n463, n451);
xnor g727 (n726, n454, n451, n445, n480);
xnor g728 (n750, n449, n479, n360, n472);
nor  g729 (n762, n477, n374, n681, n403);
or   g730 (n725, n696, n392, n668, n447);
and  g731 (n733, n486, n686, n359, n480);
xor  g732 (n766, n378, n468, n391, n690);
xnor g733 (n720, n421, n670, n483, n459);
or   g734 (n734, n426, n364, n461, n678);
nand g735 (n784, n399, n369, n477, n682);
xor  g736 (n715, n451, n471, n665, n683);
xnor g737 (n752, n465, n666, n357, n695);
and  g738 (n723, n667, n468, n470, n696);
nand g739 (n779, n669, n358, n482, n684);
nor  g740 (n759, n690, n682, n475);
xnor g741 (n777, n414, n467, n696, n470);
xor  g742 (n782, n458, n380, n435, n685);
or   g743 (n718, n371, n475, n473, n449);
xor  g744 (n755, n672, n452, n461, n457);
xor  g745 (n713, n463, n464, n478, n361);
and  g746 (n739, n448, n689, n383);
and  g747 (n737, n456, n428, n487, n686);
xnor g748 (n716, n473, n477, n464, n367);
or   g749 (n751, n405, n464, n664, n462);
and  g750 (n783, n482, n483, n472, n675);
xor  g751 (n717, n679, n476, n485, n450);
and  g752 (n778, n437, n473, n483, n410);
nand g753 (n757, n486, n475, n687, n476);
buf  g754 (n842, n758);
not  g755 (n906, n114);
not  g756 (n797, n723);
not  g757 (n942, n728);
buf  g758 (n795, n747);
buf  g759 (n863, n725);
not  g760 (n798, n785);
not  g761 (n843, n523);
not  g762 (n883, n117);
not  g763 (n933, n715);
not  g764 (n849, n716);
not  g765 (n817, n521);
buf  g766 (n917, n527);
buf  g767 (n877, n769);
buf  g768 (n929, n741);
not  g769 (n836, n731);
not  g770 (n846, n784);
not  g771 (n810, n732);
not  g772 (n901, n720);
not  g773 (n946, n528);
not  g774 (n805, n762);
not  g775 (n879, n521);
not  g776 (n923, n773);
not  g777 (n804, n710);
not  g778 (n918, n595);
not  g779 (n889, n528);
buf  g780 (n848, n760);
buf  g781 (n945, n753);
not  g782 (n893, n525);
not  g783 (n847, n758);
not  g784 (n818, n748);
not  g785 (n807, n723);
buf  g786 (n854, n785);
not  g787 (n834, n756);
buf  g788 (n788, n770);
not  g789 (n868, n765);
not  g790 (n808, n116);
buf  g791 (n799, n761);
not  g792 (n900, n734);
buf  g793 (n855, n724);
buf  g794 (n878, n709);
buf  g795 (n902, n718);
not  g796 (n895, n780);
not  g797 (n794, n751);
buf  g798 (n914, n752);
not  g799 (n845, n736);
not  g800 (n894, n742);
buf  g801 (n857, n743);
not  g802 (n821, n709);
buf  g803 (n884, n755);
buf  g804 (n861, n526);
nor  g805 (n856, n766, n724, n593);
nand g806 (n882, n747, n730, n710);
xnor g807 (n787, n736, n525, n732);
nor  g808 (n947, n766, n744, n738);
nor  g809 (n791, n708, n722, n733);
nor  g810 (n892, n748, n765, n784);
xor  g811 (n824, n779, n755, n708);
xnor g812 (n871, n786, n526, n726);
xor  g813 (n819, n786, n782, n719);
xnor g814 (n922, n716, n734, n743);
nor  g815 (n872, n748, n529, n751);
and  g816 (n812, n712, n771, n707);
and  g817 (n909, n711, n783, n772);
nand g818 (n809, n774, n767, n735);
nor  g819 (n875, n714, n716, n776);
and  g820 (n865, n594, n726, n773);
xnor g821 (n858, n768, n780, n734);
xnor g822 (n935, n725, n764, n752);
xor  g823 (n938, n715, n594, n523);
nand g824 (n862, n760, n719, n529);
and  g825 (n851, n786, n779, n526);
nand g826 (n801, n738, n737, n707);
and  g827 (n860, n763, n757, n713);
nor  g828 (n832, n778, n116, n763);
and  g829 (n925, n729, n524, n750);
xor  g830 (n880, n780, n767, n521);
xnor g831 (n859, n739, n748, n728);
xnor g832 (n790, n718, n713, n759);
or   g833 (n850, n766, n781, n711);
xnor g834 (n939, n735, n762, n754);
or   g835 (n853, n744, n773, n761);
or   g836 (n913, n711, n732, n766);
xnor g837 (n800, n115, n729, n720);
nand g838 (n873, n746, n744, n736);
and  g839 (n911, n708, n733, n709);
and  g840 (n813, n741, n528, n746);
and  g841 (n910, n727, n742, n751);
nor  g842 (n874, n750, n32, n761);
or   g843 (n932, n760, n749, n719);
xor  g844 (n915, n117, n728, n716);
nor  g845 (n830, n764, n755);
nand g846 (n891, n771, n739, n707);
or   g847 (n931, n731, n753, n757);
xnor g848 (n890, n722, n115, n727);
nor  g849 (n886, n115, n739, n754);
and  g850 (n927, n594, n752, n730);
xor  g851 (n803, n743, n774, n778);
xor  g852 (n814, n785, n723, n777);
and  g853 (n820, n721, n525, n723);
or   g854 (n904, n775, n529, n759);
xor  g855 (n796, n763, n773, n751);
and  g856 (n816, n749, n772, n725);
nand g857 (n869, n744, n522, n732);
or   g858 (n907, n117, n762, n743);
xor  g859 (n888, n730, n754, n722);
xor  g860 (n827, n756, n772, n738);
xor  g861 (n792, n786, n781, n718);
xnor g862 (n941, n726, n775, n720);
nor  g863 (n898, n775, n729, n745);
or   g864 (n839, n771, n774, n772);
nand g865 (n815, n720, n721, n768);
xnor g866 (n885, n767, n746, n770);
and  g867 (n934, n595, n760, n741);
nor  g868 (n829, n717, n759, n710);
xor  g869 (n823, n768, n745, n737);
nor  g870 (n926, n528, n724, n524);
nand g871 (n806, n781, n777, n769);
nand g872 (n930, n776, n737, n750);
xor  g873 (n887, n758, n594, n721);
or   g874 (n905, n764, n742, n747);
nor  g875 (n825, n741, n115, n725);
and  g876 (n896, n527, n783, n522);
nor  g877 (n940, n708, n521, n117);
and  g878 (n936, n722, n759, n526);
and  g879 (n833, n761, n775, n770);
nand g880 (n919, n595, n739, n782);
xnor g881 (n944, n758, n713, n523);
nand g882 (n831, n740, n769, n733);
and  g883 (n876, n745, n779, n774);
nand g884 (n864, n756, n529, n731);
xnor g885 (n943, n746, n740, n724);
xor  g886 (n826, n707, n714, n522);
and  g887 (n822, n765, n735, n727);
or   g888 (n881, n777, n778, n769);
and  g889 (n852, n733, n753, n757);
xnor g890 (n921, n771, n765, n747);
xor  g891 (n899, n784, n735, n742);
nor  g892 (n866, n523, n712);
nand g893 (n903, n736, n715, n721);
and  g894 (n924, n776, n731, n734);
xor  g895 (n916, n726, n527, n714);
nand g896 (n912, n525, n776, n768);
and  g897 (n908, n709, n756, n752);
xnor g898 (n867, n737, n717, n783);
xnor g899 (n841, n712, n782, n717);
xor  g900 (n837, n116, n715, n714);
xnor g901 (n838, n729, n749, n753);
nor  g902 (n811, n719, n767, n717);
and  g903 (n793, n738, n764, n749);
xnor g904 (n840, n711, n740, n763);
xor  g905 (n802, n783, n730, n785);
or   g906 (n844, n116, n778, n524);
nand g907 (n789, n114, n784, n728);
nand g908 (n828, n757, n740, n782);
nor  g909 (n835, n595, n780, n754);
nor  g910 (n937, n524, n777, n522);
nand g911 (n928, n593, n781, n718);
or   g912 (n897, n762, n770, n779);
and  g913 (n920, n727, n710, n750);
xor  g914 (n870, n527, n713, n745);
xor  g915 (n953, n808, n832, n793, n799);
or   g916 (n950, n792, n787, n813, n836);
xnor g917 (n960, n830, n820, n842, n841);
xor  g918 (n965, n816, n851, n814, n803);
nor  g919 (n952, n806, n801, n800, n797);
xnor g920 (n956, n837, n789, n818, n809);
or   g921 (n961, n810, n858, n833, n825);
xor  g922 (n964, n850, n848, n802, n839);
xnor g923 (n963, n791, n828, n854, n855);
xnor g924 (n949, n852, n788, n821, n815);
and  g925 (n957, n845, n838, n844, n847);
xnor g926 (n951, n846, n811, n795, n831);
and  g927 (n959, n840, n857, n796, n849);
and  g928 (n955, n819, n804, n817, n843);
or   g929 (n958, n822, n790, n835, n827);
xor  g930 (n962, n829, n826, n853, n834);
and  g931 (n954, n824, n807, n805, n856);
or   g932 (n948, n812, n798, n823, n794);
nor  g933 (n979, n698, n965, n699, n701);
or   g934 (n980, n948, n701, n495, n489);
nor  g935 (n975, n497, n492, n704, n960);
or   g936 (n976, n953, n488, n961, n702);
or   g937 (n972, n699, n964, n493, n494);
xnor g938 (n984, n698, n496, n963, n700);
xor  g939 (n966, n491, n495, n961, n706);
and  g940 (n991, n697, n963, n706, n960);
nand g941 (n978, n706, n495, n700, n704);
xor  g942 (n967, n698, n702, n959, n496);
nor  g943 (n987, n494, n703, n962, n497);
nor  g944 (n992, n699, n962, n955, n704);
xnor g945 (n989, n700, n702, n494, n705);
nand g946 (n970, n957, n490, n962, n956);
nor  g947 (n974, n490, n697, n965);
nand g948 (n983, n706, n491, n959, n497);
xnor g949 (n993, n494, n949, n488, n493);
nor  g950 (n977, n951, n497, n963, n699);
xnor g951 (n985, n493, n952, n964, n488);
nand g952 (n986, n492, n496, n488, n701);
xnor g953 (n988, n950, n961, n489, n700);
or   g954 (n982, n964, n965, n489, n490);
xnor g955 (n969, n492, n958, n705, n703);
nand g956 (n968, n960, n954, n701, n496);
and  g957 (n973, n493, n703, n705, n698);
or   g958 (n981, n704, n492, n702, n958);
nand g959 (n971, n697, n703, n490, n495);
xor  g960 (n990, n489, n705, n491);
nand g961 (n1000, n922, n897, n918, n875);
nand g962 (n1010, n990, n879, n930, n914);
nand g963 (n1003, n873, n887, n920, n933);
or   g964 (n999, n970, n945, n984, n971);
nand g965 (n1017, n862, n924, n928, n888);
or   g966 (n996, n934, n940, n869, n890);
or   g967 (n998, n884, n892, n880, n923);
xnor g968 (n1012, n909, n885, n966, n896);
or   g969 (n1021, n878, n931, n944, n900);
or   g970 (n1005, n993, n906, n988, n893);
xnor g971 (n1008, n883, n886, n937, n908);
nand g972 (n1016, n912, n904, n927, n972);
or   g973 (n1014, n867, n877, n868, n973);
and  g974 (n1022, n982, n943, n939, n986);
nand g975 (n1006, n874, n974, n917, n864);
or   g976 (n1004, n872, n921, n975, n901);
xnor g977 (n1009, n915, n905, n898, n895);
xor  g978 (n1001, n891, n882, n976, n938);
xnor g979 (n1015, n910, n981, n870, n942);
nand g980 (n1013, n993, n983, n935, n916);
and  g981 (n997, n936, n866, n894, n978);
or   g982 (n1007, n989, n863, n871, n926);
and  g983 (n1002, n987, n903, n876, n977);
xor  g984 (n1020, n985, n980, n865, n899);
xnor g985 (n995, n979, n889, n992, n907);
nor  g986 (n1011, n991, n929, n859, n860);
or   g987 (n1019, n881, n969, n941, n919);
nor  g988 (n1018, n967, n913, n932, n968);
nor  g989 (n994, n911, n902, n861, n925);
nor  g990 (n1028, n1019, n1013, n1006, n1002);
nor  g991 (n1026, n1001, n1014, n999, n1015);
or   g992 (n1024, n998, n996, n1022, n1000);
xnor g993 (n1029, n1008, n1021, n995, n1017);
nor  g994 (n1023, n1007, n1003, n1018, n997);
or   g995 (n1027, n1005, n32, n994, n1010);
and  g996 (n1030, n1016, n1012, n947, n1009);
xor  g997 (n1025, n1020, n946, n1004, n1011);
nor  g998 (n1032, n1030, n1027, n1028, n1024);
xnor g999 (n1031, n1029, n1025, n1026, n1023);
endmodule
