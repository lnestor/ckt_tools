

module Stat_100_57
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n83,
  n102,
  n88,
  n70,
  n77,
  n92,
  n95,
  n115,
  n94,
  n99,
  n71,
  n106,
  n104,
  n78,
  n100,
  n87,
  n75,
  n98,
  n103,
  n127,
  n124,
  n121,
  n128,
  n129,
  n126,
  n130,
  n120,
  n123,
  n122,
  n125,
  n132,
  n131,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n83;
  output n102;
  output n88;
  output n70;
  output n77;
  output n92;
  output n95;
  output n115;
  output n94;
  output n99;
  output n71;
  output n106;
  output n104;
  output n78;
  output n100;
  output n87;
  output n75;
  output n98;
  output n103;
  output n127;
  output n124;
  output n121;
  output n128;
  output n129;
  output n126;
  output n130;
  output n120;
  output n123;
  output n122;
  output n125;
  output n132;
  output n131;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n72;
  wire n73;
  wire n74;
  wire n76;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n84;
  wire n85;
  wire n86;
  wire n89;
  wire n90;
  wire n91;
  wire n93;
  wire n96;
  wire n97;
  wire n101;
  wire n105;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n35,
    n2
  );


  buf
  g1
  (
    n41,
    n3
  );


  buf
  g2
  (
    KeyWire_0_42,
    n1
  );


  not
  g3
  (
    KeyWire_0_15,
    n1
  );


  not
  g4
  (
    n37,
    n3
  );


  buf
  g5
  (
    n36,
    n1
  );


  not
  g6
  (
    KeyWire_0_16,
    n2
  );


  buf
  g7
  (
    KeyWire_0_28,
    n2
  );


  not
  g8
  (
    KeyWire_0_59,
    n2
  );


  buf
  g9
  (
    n38,
    n1
  );


  not
  g10
  (
    KeyWire_0_35,
    n33
  );


  not
  g11
  (
    KeyWire_0_34,
    n34
  );


  buf
  g12
  (
    KeyWire_0_26,
    n35
  );


  buf
  g13
  (
    n44,
    n37
  );


  buf
  g14
  (
    n49,
    n34
  );


  not
  g15
  (
    n55,
    n36
  );


  buf
  g16
  (
    n43,
    n35
  );


  buf
  g17
  (
    KeyWire_0_58,
    n36
  );


  buf
  g18
  (
    KeyWire_0_36,
    n34
  );


  buf
  g19
  (
    KeyWire_0_5,
    n36
  );


  buf
  g20
  (
    n47,
    n35
  );


  and
  g21
  (
    KeyWire_0_25,
    n37,
    n33
  );


  or
  g22
  (
    KeyWire_0_38,
    n33,
    n35,
    n34,
    n36
  );


  not
  g23
  (
    KeyWire_0_17,
    n45
  );


  not
  g24
  (
    KeyWire_0_7,
    n45
  );


  buf
  g25
  (
    KeyWire_0_19,
    n47
  );


  not
  g26
  (
    n69,
    n46
  );


  not
  g27
  (
    KeyWire_0_56,
    n49
  );


  not
  g28
  (
    n58,
    n46
  );


  not
  g29
  (
    KeyWire_0_4,
    n44
  );


  not
  g30
  (
    n57,
    n45
  );


  not
  g31
  (
    n60,
    n48
  );


  not
  g32
  (
    n67,
    n43
  );


  buf
  g33
  (
    KeyWire_0_13,
    n45
  );


  nor
  g34
  (
    n56,
    n46,
    n47,
    n49,
    n44
  );


  and
  g35
  (
    KeyWire_0_60,
    n44,
    n48,
    n47
  );


  xnor
  g36
  (
    KeyWire_0_43,
    n46,
    n44,
    n48
  );


  xnor
  g37
  (
    n118,
    n4,
    n27,
    n29,
    n62
  );


  nand
  g38
  (
    KeyWire_0_41,
    n61,
    n20,
    n17
  );


  and
  g39
  (
    KeyWire_0_33,
    n65,
    n22,
    n31,
    n56
  );


  nand
  g40
  (
    n77,
    n61,
    n28,
    n51,
    n63
  );


  nor
  g41
  (
    KeyWire_0_55,
    n11,
    n17,
    n14,
    n64
  );


  or
  g42
  (
    KeyWire_0_62,
    n54,
    n14,
    n24,
    n28
  );


  nand
  g43
  (
    n93,
    n30,
    n65,
    n26,
    n66
  );


  xnor
  g44
  (
    n117,
    n61,
    n5,
    n32,
    n13
  );


  nand
  g45
  (
    n105,
    n64,
    n16,
    n3,
    n25
  );


  and
  g46
  (
    n81,
    n60,
    n13,
    n55,
    n20
  );


  and
  g47
  (
    KeyWire_0_24,
    n9,
    n3,
    n63,
    n15
  );


  xnor
  g48
  (
    KeyWire_0_18,
    n64,
    n50,
    n8,
    n21
  );


  nor
  g49
  (
    KeyWire_0_30,
    n55,
    n30,
    n49,
    n23
  );


  nand
  g50
  (
    KeyWire_0_37,
    n6,
    n19,
    n27,
    n53
  );


  nand
  g51
  (
    KeyWire_0_12,
    n65,
    n18,
    n31,
    n9
  );


  nor
  g52
  (
    KeyWire_0_29,
    n53,
    n5,
    n8,
    n18
  );


  and
  g53
  (
    KeyWire_0_45,
    n67,
    n7,
    n58,
    n11
  );


  xnor
  g54
  (
    n71,
    n66,
    n25,
    n22
  );


  xnor
  g55
  (
    n114,
    n69,
    n10,
    n9
  );


  or
  g56
  (
    KeyWire_0_46,
    n62,
    n51,
    n12,
    n58
  );


  and
  g57
  (
    KeyWire_0_54,
    n69,
    n57,
    n13,
    n54
  );


  or
  g58
  (
    KeyWire_0_31,
    n4,
    n30,
    n29,
    n27
  );


  nor
  g59
  (
    KeyWire_0_9,
    n27,
    n56,
    n19,
    n23
  );


  xor
  g60
  (
    KeyWire_0_48,
    n59,
    n23,
    n16,
    n14
  );


  xor
  g61
  (
    KeyWire_0_50,
    n58,
    n10,
    n24,
    n6
  );


  xnor
  g62
  (
    KeyWire_0_0,
    n18,
    n32,
    n57,
    n28
  );


  or
  g63
  (
    KeyWire_0_47,
    n32,
    n16,
    n13,
    n56
  );


  nand
  g64
  (
    n86,
    n49,
    n67,
    n31
  );


  xor
  g65
  (
    KeyWire_0_49,
    n21,
    n16,
    n30,
    n22
  );


  and
  g66
  (
    KeyWire_0_40,
    n21,
    n59,
    n69,
    n29
  );


  and
  g67
  (
    KeyWire_0_23,
    n63,
    n65,
    n50,
    n68
  );


  and
  g68
  (
    n91,
    n29,
    n7,
    n17,
    n61
  );


  xnor
  g69
  (
    n96,
    n60,
    n57,
    n7,
    n24
  );


  nor
  g70
  (
    KeyWire_0_1,
    n68,
    n19,
    n26,
    n53
  );


  xnor
  g71
  (
    KeyWire_0_10,
    n24,
    n56,
    n17,
    n55
  );


  nor
  g72
  (
    n89,
    n60,
    n14,
    n28,
    n15
  );


  and
  g73
  (
    KeyWire_0_39,
    n5,
    n12,
    n52,
    n15
  );


  nor
  g74
  (
    KeyWire_0_27,
    n9,
    n51,
    n62,
    n21
  );


  nor
  g75
  (
    n103,
    n58,
    n55,
    n5,
    n12
  );


  xnor
  g76
  (
    KeyWire_0_51,
    n66,
    n4,
    n51,
    n60
  );


  xor
  g77
  (
    KeyWire_0_2,
    n57,
    n4,
    n8,
    n20
  );


  or
  g78
  (
    KeyWire_0_22,
    n32,
    n25,
    n10,
    n23
  );


  nor
  g79
  (
    n88,
    n62,
    n50,
    n53,
    n11
  );


  nand
  g80
  (
    KeyWire_0_21,
    n68,
    n52,
    n15,
    n54
  );


  and
  g81
  (
    KeyWire_0_61,
    n66,
    n26,
    n6,
    n19
  );


  nand
  g82
  (
    KeyWire_0_11,
    n54,
    n59,
    n26,
    n31
  );


  and
  g83
  (
    KeyWire_0_53,
    n59,
    n18,
    n67,
    n7
  );


  xor
  g84
  (
    KeyWire_0_63,
    n63,
    n22,
    n11,
    n12
  );


  or
  g85
  (
    n83,
    n64,
    n8,
    n68,
    n69
  );


  nand
  g86
  (
    KeyWire_0_57,
    n50,
    n52,
    n6
  );


  nand
  g87
  (
    KeyWire_0_32,
    n89,
    n103,
    n96,
    n92
  );


  or
  g88
  (
    KeyWire_0_6,
    n114,
    n111,
    n42,
    n41
  );


  or
  g89
  (
    KeyWire_0_52,
    n108,
    n107,
    n38,
    n116
  );


  nand
  g90
  (
    KeyWire_0_8,
    n112,
    n40,
    n109
  );


  nand
  g91
  (
    n126,
    n39,
    n98,
    n118,
    n42
  );


  nor
  g92
  (
    n127,
    n38,
    n106,
    n95,
    n97
  );


  or
  g93
  (
    KeyWire_0_3,
    n113,
    n41,
    n93,
    n101
  );


  xor
  g94
  (
    n132,
    n102,
    n105,
    n40,
    n91
  );


  nand
  g95
  (
    KeyWire_0_14,
    n117,
    n110,
    n119,
    n94
  );


  nand
  g96
  (
    n130,
    n39,
    n39,
    n40,
    n104
  );


  xor
  g97
  (
    KeyWire_0_20,
    n99,
    n37,
    n42,
    n38
  );


  and
  g98
  (
    n128,
    n100,
    n41,
    n38
  );


  nor
  g99
  (
    KeyWire_0_44,
    n115,
    n39,
    n90,
    n42
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n119,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n73,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n112,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n121,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n61,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n51,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n125,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n59,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n122,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n94,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n74,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n107,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n104,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n63,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n120,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n33,
    KeyNOTWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n42,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n64,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n101,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n66,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n129,
    KeyNOTWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n80,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n76,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n70,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n95,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n54,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n46,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n111,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n34,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n85,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n92,
    KeyNOTWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n97,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n131,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n82,
    KeyNOTWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n50,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n53,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    n52,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n90,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n48,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n98,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n72,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n106,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n40,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n65,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n124,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n79,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n113,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n116,
    keyIn_0_47,
    KeyWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n75,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n110,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n102,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n115,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n123,
    keyIn_0_52,
    KeyWire_0_52
  );


  xnor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n84,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n109,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n100,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n62,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n108,
    KeyNOTWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    n45,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n39,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n68,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n78,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n87,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n99,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

