

module Stat_100_41
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n112,
  n131,
  n117,
  n108,
  n125,
  n121,
  n130,
  n118,
  n102,
  n116,
  n110,
  n124,
  n128,
  n122,
  n114,
  n104,
  n109,
  n113,
  n123,
  n101,
  n127,
  n105,
  n119,
  n103,
  n120,
  n106,
  n132,
  n129,
  n107,
  n126,
  n111,
  n115,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n112;
  output n131;
  output n117;
  output n108;
  output n125;
  output n121;
  output n130;
  output n118;
  output n102;
  output n116;
  output n110;
  output n124;
  output n128;
  output n122;
  output n114;
  output n104;
  output n109;
  output n113;
  output n123;
  output n101;
  output n127;
  output n105;
  output n119;
  output n103;
  output n120;
  output n106;
  output n132;
  output n129;
  output n107;
  output n126;
  output n111;
  output n115;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyNOTWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyNOTWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    KeyWire_0_16,
    n4
  );


  not
  g1
  (
    KeyWire_0_32,
    n2
  );


  not
  g2
  (
    KeyWire_0_29,
    n3
  );


  buf
  g3
  (
    n42,
    n3
  );


  buf
  g4
  (
    KeyWire_0_51,
    n2
  );


  not
  g5
  (
    KeyWire_0_26,
    n1
  );


  buf
  g6
  (
    n37,
    n3
  );


  not
  g7
  (
    n38,
    n4
  );


  buf
  g8
  (
    n36,
    n1
  );


  not
  g9
  (
    KeyWire_0_38,
    n1
  );


  buf
  g10
  (
    n33,
    n2
  );


  not
  g11
  (
    n44,
    n4
  );


  not
  g12
  (
    KeyWire_0_60,
    n13
  );


  buf
  g13
  (
    KeyWire_0_6,
    n15
  );


  buf
  g14
  (
    KeyWire_0_50,
    n27
  );


  not
  g15
  (
    KeyWire_0_24,
    n8
  );


  not
  g16
  (
    n51,
    n31
  );


  not
  g17
  (
    n73,
    n33
  );


  buf
  g18
  (
    KeyWire_0_12,
    n31
  );


  not
  g19
  (
    n75,
    n19
  );


  or
  g20
  (
    KeyWire_0_17,
    n11,
    n21,
    n18,
    n42
  );


  nor
  g21
  (
    KeyWire_0_31,
    n22,
    n41,
    n36,
    n18
  );


  nand
  g22
  (
    n78,
    n35,
    n17,
    n25,
    n20
  );


  nand
  g23
  (
    KeyWire_0_18,
    n37,
    n39,
    n42,
    n43
  );


  nor
  g24
  (
    KeyWire_0_1,
    n22,
    n19,
    n35,
    n44
  );


  or
  g25
  (
    KeyWire_0_23,
    n18,
    n13,
    n7,
    n28
  );


  xor
  g26
  (
    KeyWire_0_30,
    n43,
    n30,
    n39,
    n38
  );


  xor
  g27
  (
    KeyWire_0_14,
    n29,
    n24,
    n6,
    n26
  );


  nor
  g28
  (
    KeyWire_0_11,
    n40,
    n14,
    n9,
    n11
  );


  and
  g29
  (
    KeyWire_0_55,
    n7,
    n16,
    n10,
    n19
  );


  or
  g30
  (
    KeyWire_0_42,
    n9,
    n35,
    n16,
    n42
  );


  and
  g31
  (
    KeyWire_0_19,
    n29,
    n41,
    n37,
    n20
  );


  and
  g32
  (
    KeyWire_0_15,
    n37,
    n44,
    n23,
    n27
  );


  nand
  g33
  (
    n63,
    n32,
    n25,
    n34,
    n5
  );


  and
  g34
  (
    n52,
    n14,
    n38,
    n44,
    n8
  );


  xor
  g35
  (
    KeyWire_0_59,
    n9,
    n23,
    n22,
    n15
  );


  and
  g36
  (
    n70,
    n17,
    n6,
    n33,
    n43
  );


  nand
  g37
  (
    KeyWire_0_8,
    n12,
    n24,
    n5,
    n26
  );


  or
  g38
  (
    KeyWire_0_45,
    n24,
    n16,
    n32,
    n13
  );


  and
  g39
  (
    KeyWire_0_4,
    n29,
    n11,
    n7,
    n26
  );


  nand
  g40
  (
    KeyWire_0_47,
    n30,
    n36,
    n40,
    n6
  );


  nor
  g41
  (
    KeyWire_0_63,
    n30,
    n39,
    n21,
    n10
  );


  nand
  g42
  (
    KeyWire_0_52,
    n25,
    n10,
    n41,
    n31
  );


  nand
  g43
  (
    KeyWire_0_7,
    n14,
    n15,
    n5,
    n8
  );


  nor
  g44
  (
    KeyWire_0_0,
    n38,
    n27,
    n36,
    n32
  );


  and
  g45
  (
    n68,
    n17,
    n34,
    n33,
    n20
  );


  xor
  g46
  (
    n77,
    n28,
    n23,
    n12,
    n40
  );


  xor
  g47
  (
    KeyWire_0_21,
    n34,
    n21,
    n12,
    n28
  );


  buf
  g48
  (
    KeyWire_0_2,
    n45
  );


  not
  g49
  (
    KeyWire_0_5,
    n49
  );


  buf
  g50
  (
    KeyWire_0_9,
    n48
  );


  buf
  g51
  (
    n92,
    n45
  );


  buf
  g52
  (
    KeyWire_0_40,
    n46
  );


  buf
  g53
  (
    n91,
    n48
  );


  buf
  g54
  (
    KeyWire_0_13,
    n46
  );


  not
  g55
  (
    n90,
    n50
  );


  buf
  g56
  (
    KeyWire_0_44,
    n50
  );


  buf
  g57
  (
    n89,
    n49
  );


  buf
  g58
  (
    KeyWire_0_48,
    n51
  );


  not
  g59
  (
    n88,
    n51
  );


  buf
  g60
  (
    KeyWire_0_10,
    n48
  );


  buf
  g61
  (
    n100,
    n50
  );


  not
  g62
  (
    KeyWire_0_46,
    n46
  );


  buf
  g63
  (
    KeyWire_0_61,
    n45
  );


  buf
  g64
  (
    KeyWire_0_43,
    n47
  );


  not
  g65
  (
    n97,
    n47
  );


  not
  g66
  (
    n99,
    n47
  );


  not
  g67
  (
    KeyWire_0_53,
    n49
  );


  or
  g68
  (
    n120,
    n97,
    n64,
    n98,
    n70
  );


  xnor
  g69
  (
    KeyWire_0_33,
    n60,
    n80,
    n95
  );


  or
  g70
  (
    KeyWire_0_62,
    n78,
    n74,
    n71,
    n77
  );


  or
  g71
  (
    n130,
    n57,
    n63,
    n69,
    n99
  );


  xnor
  g72
  (
    KeyWire_0_25,
    n88,
    n56,
    n72,
    n58
  );


  or
  g73
  (
    n128,
    n70,
    n91,
    n94,
    n60
  );


  or
  g74
  (
    n113,
    n71,
    n54,
    n51,
    n59
  );


  nand
  g75
  (
    KeyWire_0_20,
    n86,
    n94,
    n62
  );


  nand
  g76
  (
    n129,
    n82,
    n75,
    n52,
    n61
  );


  and
  g77
  (
    KeyWire_0_3,
    n62,
    n85,
    n54,
    n75
  );


  xor
  g78
  (
    n108,
    n59,
    n79,
    n68,
    n91
  );


  xor
  g79
  (
    n114,
    n69,
    n92,
    n53,
    n65
  );


  xor
  g80
  (
    KeyWire_0_36,
    n83,
    n91,
    n60,
    n68
  );


  nand
  g81
  (
    KeyWire_0_22,
    n74,
    n72,
    n89,
    n65
  );


  xor
  g82
  (
    KeyWire_0_41,
    n68,
    n64,
    n81,
    n92
  );


  xnor
  g83
  (
    KeyWire_0_28,
    n53,
    n92,
    n99,
    n98
  );


  or
  g84
  (
    KeyWire_0_35,
    n56,
    n56,
    n61,
    n66
  );


  nand
  g85
  (
    n106,
    n65,
    n99,
    n93,
    n74
  );


  nand
  g86
  (
    n118,
    n73,
    n55,
    n78,
    n76
  );


  xnor
  g87
  (
    KeyWire_0_49,
    n95,
    n87,
    n71,
    n55
  );


  nor
  g88
  (
    n107,
    n97,
    n70,
    n84,
    n79
  );


  nor
  g89
  (
    KeyWire_0_54,
    n58,
    n77,
    n66,
    n52
  );


  nand
  g90
  (
    KeyWire_0_27,
    n63,
    n80,
    n59,
    n93
  );


  nand
  g91
  (
    n109,
    n64,
    n72,
    n100,
    n57
  );


  nor
  g92
  (
    KeyWire_0_56,
    n58,
    n67,
    n73,
    n66
  );


  xor
  g93
  (
    n117,
    n100,
    n73,
    n80,
    n96
  );


  and
  g94
  (
    KeyWire_0_39,
    n54,
    n67,
    n90,
    n61
  );


  xnor
  g95
  (
    KeyWire_0_37,
    n76,
    n75,
    n52,
    n53
  );


  or
  g96
  (
    KeyWire_0_34,
    n67,
    n93,
    n96,
    n78
  );


  or
  g97
  (
    n131,
    n98,
    n96,
    n94,
    n79
  );


  nor
  g98
  (
    KeyWire_0_57,
    n69,
    n97,
    n57,
    n100
  );


  or
  g99
  (
    KeyWire_0_58,
    n55,
    n76,
    n63,
    n77
  );


  xnor
  KeyGate_0_0
  (
    n57,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n80,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n96,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n112,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n48,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n84,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n66,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n67,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n47,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n81,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n86,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n65,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n71,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n85,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n49,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n53,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n40,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n61,
    KeyNOTWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n45,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n69,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n115,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n62,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n104,
    KeyNOTWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n74,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n72,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n121,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n41,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n122,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n110,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n34,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n60,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n64,
    KeyNOTWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n39,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    n102,
    keyIn_0_33,
    KeyWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n132,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n101,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n119,
    keyIn_0_36,
    KeyWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n111,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n43,
    KeyNOTWire_0_38
  );


  xnor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n124,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n83,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n105,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n58,
    keyIn_0_42,
    KeyWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n87,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    n82,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n79,
    KeyNOTWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n98,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n46,
    KeyNOTWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n94,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    KeyNOTWire_0_49,
    keyIn_0_49,
    KeyWire_0_49
  );


  not
  KeyNOTGate_0_49
  (
    n123,
    KeyNOTWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n76,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n35,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n54,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n95,
    keyIn_0_53,
    KeyWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n103,
    KeyNOTWire_0_54
  );


  xor
  KeyGate_0_55
  (
    n50,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n126,
    keyIn_0_56,
    KeyWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n116,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n127,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    n55,
    keyIn_0_59,
    KeyWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n59,
    KeyNOTWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n93,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n125,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n56,
    KeyNOTWire_0_63
  );


endmodule

