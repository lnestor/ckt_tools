

module Stat_1000_204
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n968,
  n967,
  n957,
  n984,
  n953,
  n962,
  n979,
  n976,
  n969,
  n960,
  n981,
  n977,
  n974,
  n956,
  n985,
  n952,
  n973,
  n971,
  n1031,
  n1023,
  n1025,
  n1030,
  n1032,
  n1027,
  n1021,
  n1026,
  n1019,
  n1020,
  n1029,
  n1024,
  n1028,
  n1022,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n968;output n967;output n957;output n984;output n953;output n962;output n979;output n976;output n969;output n960;output n981;output n977;output n974;output n956;output n985;output n952;output n973;output n971;output n1031;output n1023;output n1025;output n1030;output n1032;output n1027;output n1021;output n1026;output n1019;output n1020;output n1029;output n1024;output n1028;output n1022;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n954;wire n955;wire n958;wire n959;wire n961;wire n963;wire n964;wire n965;wire n966;wire n970;wire n972;wire n975;wire n978;wire n980;wire n982;wire n983;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyNOTWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyNOTWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyNOTWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyNOTWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyNOTWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyNOTWire_0_21;wire KeyWire_0_22;wire KeyNOTWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyNOTWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyNOTWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;wire KeyNOTWire_0_31;

  buf
  g0
  (
    n69,
    n8
  );


  not
  g1
  (
    n53,
    n27
  );


  buf
  g2
  (
    n79,
    n25
  );


  buf
  g3
  (
    n61,
    n28
  );


  not
  g4
  (
    n33,
    n18
  );


  buf
  g5
  (
    n91,
    n11
  );


  not
  g6
  (
    n87,
    n24
  );


  not
  g7
  (
    KeyWire_0_4,
    n16
  );


  not
  g8
  (
    n77,
    n21
  );


  not
  g9
  (
    n94,
    n27
  );


  not
  g10
  (
    n82,
    n20
  );


  buf
  g11
  (
    n65,
    n4
  );


  not
  g12
  (
    n66,
    n24
  );


  not
  g13
  (
    n72,
    n11
  );


  not
  g14
  (
    n38,
    n12
  );


  buf
  g15
  (
    n60,
    n7
  );


  buf
  g16
  (
    n49,
    n15
  );


  not
  g17
  (
    n56,
    n17
  );


  buf
  g18
  (
    n46,
    n22
  );


  buf
  g19
  (
    n55,
    n27
  );


  buf
  g20
  (
    n85,
    n20
  );


  not
  g21
  (
    n58,
    n18
  );


  buf
  g22
  (
    n89,
    n23
  );


  buf
  g23
  (
    n39,
    n13
  );


  not
  g24
  (
    n48,
    n8
  );


  not
  g25
  (
    n81,
    n10
  );


  not
  g26
  (
    n40,
    n3
  );


  not
  g27
  (
    n68,
    n23
  );


  buf
  g28
  (
    n73,
    n17
  );


  not
  g29
  (
    n34,
    n16
  );


  buf
  g30
  (
    n63,
    n2
  );


  not
  g31
  (
    n57,
    n2
  );


  buf
  g32
  (
    n59,
    n20
  );


  not
  g33
  (
    n92,
    n28
  );


  not
  g34
  (
    n36,
    n15
  );


  not
  g35
  (
    n35,
    n1
  );


  not
  g36
  (
    n52,
    n23
  );


  not
  g37
  (
    n64,
    n25
  );


  buf
  g38
  (
    n41,
    n19
  );


  not
  g39
  (
    n78,
    n21
  );


  not
  g40
  (
    n42,
    n19
  );


  not
  g41
  (
    n54,
    n26
  );


  buf
  g42
  (
    n37,
    n3
  );


  not
  g43
  (
    n84,
    n19
  );


  not
  g44
  (
    n43,
    n25
  );


  not
  g45
  (
    n47,
    n17
  );


  not
  g46
  (
    n44,
    n22
  );


  buf
  g47
  (
    n90,
    n24
  );


  buf
  g48
  (
    n74,
    n7
  );


  buf
  g49
  (
    n86,
    n18
  );


  buf
  g50
  (
    n71,
    n21
  );


  buf
  g51
  (
    n80,
    n21
  );


  not
  g52
  (
    n93,
    n6
  );


  not
  g53
  (
    n70,
    n14
  );


  buf
  g54
  (
    n88,
    n22
  );


  buf
  g55
  (
    n45,
    n6
  );


  xor
  g56
  (
    n83,
    n26,
    n19
  );


  nor
  g57
  (
    n51,
    n5,
    n22,
    n14,
    n9
  );


  or
  g58
  (
    n76,
    n1,
    n20,
    n10,
    n18
  );


  xor
  g59
  (
    n67,
    n5,
    n23,
    n26,
    n17
  );


  xnor
  g60
  (
    n50,
    n12,
    n9,
    n4,
    n24
  );


  xnor
  g61
  (
    n75,
    n26,
    n13,
    n25,
    n27
  );


  buf
  g62
  (
    n244,
    n45
  );


  buf
  g63
  (
    n233,
    n71
  );


  buf
  g64
  (
    n259,
    n41
  );


  buf
  g65
  (
    n274,
    n78
  );


  not
  g66
  (
    n310,
    n60
  );


  not
  g67
  (
    n278,
    n59
  );


  buf
  g68
  (
    n247,
    n39
  );


  buf
  g69
  (
    n116,
    n70
  );


  buf
  g70
  (
    KeyWire_0_8,
    n40
  );


  not
  g71
  (
    n163,
    n68
  );


  not
  g72
  (
    n301,
    n44
  );


  buf
  g73
  (
    n238,
    n42
  );


  buf
  g74
  (
    n192,
    n65
  );


  not
  g75
  (
    KeyWire_0_7,
    n63
  );


  buf
  g76
  (
    n161,
    n79
  );


  not
  g77
  (
    n281,
    n58
  );


  buf
  g78
  (
    n280,
    n33
  );


  not
  g79
  (
    n196,
    n36
  );


  not
  g80
  (
    n118,
    n50
  );


  not
  g81
  (
    n139,
    n47
  );


  not
  g82
  (
    n124,
    n84
  );


  buf
  g83
  (
    n100,
    n56
  );


  not
  g84
  (
    n154,
    n81
  );


  buf
  g85
  (
    n112,
    n87
  );


  not
  g86
  (
    n242,
    n58
  );


  not
  g87
  (
    n143,
    n86
  );


  not
  g88
  (
    n252,
    n45
  );


  not
  g89
  (
    n240,
    n56
  );


  not
  g90
  (
    n202,
    n42
  );


  buf
  g91
  (
    n129,
    n83
  );


  buf
  g92
  (
    KeyWire_0_23,
    n76
  );


  not
  g93
  (
    n146,
    n48
  );


  buf
  g94
  (
    n212,
    n62
  );


  buf
  g95
  (
    n268,
    n64
  );


  buf
  g96
  (
    n302,
    n66
  );


  not
  g97
  (
    n209,
    n50
  );


  buf
  g98
  (
    n219,
    n71
  );


  not
  g99
  (
    n251,
    n86
  );


  not
  g100
  (
    n113,
    n81
  );


  buf
  g101
  (
    n234,
    n73
  );


  not
  g102
  (
    n117,
    n37
  );


  not
  g103
  (
    n164,
    n70
  );


  not
  g104
  (
    n204,
    n50
  );


  not
  g105
  (
    n134,
    n82
  );


  not
  g106
  (
    n241,
    n85
  );


  buf
  g107
  (
    n109,
    n79
  );


  not
  g108
  (
    n131,
    n78
  );


  buf
  g109
  (
    KeyWire_0_26,
    n37
  );


  not
  g110
  (
    n261,
    n39
  );


  not
  g111
  (
    n144,
    n66
  );


  buf
  g112
  (
    n174,
    n78
  );


  buf
  g113
  (
    n288,
    n83
  );


  not
  g114
  (
    n218,
    n77
  );


  not
  g115
  (
    n176,
    n63
  );


  buf
  g116
  (
    n297,
    n69
  );


  not
  g117
  (
    n215,
    n77
  );


  not
  g118
  (
    n184,
    n46
  );


  not
  g119
  (
    n152,
    n46
  );


  not
  g120
  (
    n142,
    n60
  );


  not
  g121
  (
    n160,
    n64
  );


  buf
  g122
  (
    n305,
    n85
  );


  buf
  g123
  (
    n275,
    n59
  );


  buf
  g124
  (
    n248,
    n71
  );


  not
  g125
  (
    n193,
    n44
  );


  buf
  g126
  (
    n208,
    n44
  );


  not
  g127
  (
    n226,
    n72
  );


  not
  g128
  (
    n220,
    n42
  );


  buf
  g129
  (
    n236,
    n77
  );


  buf
  g130
  (
    n148,
    n69
  );


  not
  g131
  (
    n270,
    n67
  );


  not
  g132
  (
    n158,
    n33
  );


  not
  g133
  (
    n262,
    n73
  );


  buf
  g134
  (
    n243,
    n87
  );


  buf
  g135
  (
    n290,
    n64
  );


  not
  g136
  (
    n298,
    n86
  );


  not
  g137
  (
    n216,
    n69
  );


  buf
  g138
  (
    n291,
    n41
  );


  buf
  g139
  (
    n180,
    n46
  );


  buf
  g140
  (
    n185,
    n63
  );


  not
  g141
  (
    n159,
    n82
  );


  not
  g142
  (
    n165,
    n52
  );


  buf
  g143
  (
    n155,
    n38
  );


  not
  g144
  (
    n122,
    n81
  );


  not
  g145
  (
    n266,
    n36
  );


  buf
  g146
  (
    n171,
    n75
  );


  not
  g147
  (
    n287,
    n78
  );


  buf
  g148
  (
    n145,
    n87
  );


  not
  g149
  (
    n293,
    n57
  );


  not
  g150
  (
    n211,
    n67
  );


  buf
  g151
  (
    n181,
    n79
  );


  buf
  g152
  (
    n115,
    n85
  );


  not
  g153
  (
    n311,
    n43
  );


  not
  g154
  (
    n175,
    n40
  );


  buf
  g155
  (
    n182,
    n48
  );


  not
  g156
  (
    n141,
    n65
  );


  buf
  g157
  (
    n303,
    n33
  );


  not
  g158
  (
    n230,
    n39
  );


  not
  g159
  (
    n173,
    n85
  );


  buf
  g160
  (
    n150,
    n75
  );


  not
  g161
  (
    n272,
    n49
  );


  not
  g162
  (
    KeyWire_0_17,
    n76
  );


  not
  g163
  (
    n224,
    n38
  );


  not
  g164
  (
    KeyWire_0_27,
    n44
  );


  buf
  g165
  (
    n156,
    n54
  );


  buf
  g166
  (
    n225,
    n55
  );


  buf
  g167
  (
    n231,
    n36
  );


  buf
  g168
  (
    n166,
    n58
  );


  buf
  g169
  (
    n101,
    n51
  );


  not
  g170
  (
    n235,
    n72
  );


  not
  g171
  (
    n294,
    n59
  );


  buf
  g172
  (
    n123,
    n82
  );


  not
  g173
  (
    n135,
    n71
  );


  buf
  g174
  (
    n108,
    n64
  );


  not
  g175
  (
    n308,
    n43
  );


  buf
  g176
  (
    n210,
    n37
  );


  buf
  g177
  (
    n203,
    n42
  );


  not
  g178
  (
    n125,
    n76
  );


  not
  g179
  (
    n140,
    n75
  );


  not
  g180
  (
    n277,
    n76
  );


  buf
  g181
  (
    n197,
    n34
  );


  buf
  g182
  (
    n273,
    n33
  );


  not
  g183
  (
    n98,
    n57
  );


  not
  g184
  (
    n102,
    n52
  );


  not
  g185
  (
    n172,
    n80
  );


  not
  g186
  (
    n130,
    n86
  );


  not
  g187
  (
    n201,
    n73
  );


  not
  g188
  (
    n151,
    n80
  );


  buf
  g189
  (
    n205,
    n52
  );


  buf
  g190
  (
    n217,
    n43
  );


  not
  g191
  (
    n147,
    n53
  );


  not
  g192
  (
    n195,
    n61
  );


  buf
  g193
  (
    n284,
    n62
  );


  buf
  g194
  (
    n126,
    n72
  );


  not
  g195
  (
    n312,
    n74
  );


  not
  g196
  (
    n198,
    n55
  );


  buf
  g197
  (
    n190,
    n48
  );


  buf
  g198
  (
    n96,
    n35
  );


  buf
  g199
  (
    n120,
    n48
  );


  not
  g200
  (
    n286,
    n70
  );


  buf
  g201
  (
    n255,
    n56
  );


  not
  g202
  (
    n228,
    n35
  );


  buf
  g203
  (
    n128,
    n68
  );


  buf
  g204
  (
    n296,
    n54
  );


  not
  g205
  (
    n95,
    n43
  );


  not
  g206
  (
    n221,
    n87
  );


  not
  g207
  (
    n199,
    n54
  );


  buf
  g208
  (
    n183,
    n40
  );


  buf
  g209
  (
    n295,
    n53
  );


  buf
  g210
  (
    KeyWire_0_15,
    n51
  );


  not
  g211
  (
    n137,
    n58
  );


  buf
  g212
  (
    n194,
    n69
  );


  buf
  g213
  (
    n257,
    n45
  );


  not
  g214
  (
    n207,
    n74
  );


  not
  g215
  (
    n97,
    n60
  );


  not
  g216
  (
    n267,
    n79
  );


  not
  g217
  (
    n200,
    n62
  );


  buf
  g218
  (
    n168,
    n61
  );


  buf
  g219
  (
    n133,
    n63
  );


  buf
  g220
  (
    n229,
    n49
  );


  not
  g221
  (
    n214,
    n65
  );


  buf
  g222
  (
    n179,
    n41
  );


  not
  g223
  (
    n239,
    n34
  );


  not
  g224
  (
    n114,
    n80
  );


  not
  g225
  (
    n162,
    n55
  );


  buf
  g226
  (
    n232,
    n80
  );


  buf
  g227
  (
    n304,
    n68
  );


  buf
  g228
  (
    n264,
    n49
  );


  buf
  g229
  (
    n223,
    n61
  );


  not
  g230
  (
    n249,
    n74
  );


  not
  g231
  (
    n177,
    n66
  );


  not
  g232
  (
    n99,
    n53
  );


  buf
  g233
  (
    n253,
    n66
  );


  not
  g234
  (
    n121,
    n82
  );


  buf
  g235
  (
    n153,
    n84
  );


  buf
  g236
  (
    n246,
    n36
  );


  not
  g237
  (
    n178,
    n54
  );


  not
  g238
  (
    n300,
    n65
  );


  buf
  g239
  (
    n282,
    n72
  );


  buf
  g240
  (
    n213,
    n47
  );


  buf
  g241
  (
    n299,
    n53
  );


  not
  g242
  (
    n191,
    n46
  );


  not
  g243
  (
    n170,
    n75
  );


  not
  g244
  (
    n260,
    n83
  );


  buf
  g245
  (
    n106,
    n35
  );


  buf
  g246
  (
    n206,
    n70
  );


  not
  g247
  (
    n105,
    n38
  );


  buf
  g248
  (
    n127,
    n52
  );


  not
  g249
  (
    n271,
    n51
  );


  not
  g250
  (
    n289,
    n51
  );


  not
  g251
  (
    n157,
    n34
  );


  not
  g252
  (
    n265,
    n62
  );


  not
  g253
  (
    n307,
    n55
  );


  not
  g254
  (
    n186,
    n74
  );


  buf
  g255
  (
    KeyWire_0_12,
    n81
  );


  not
  g256
  (
    n279,
    n73
  );


  not
  g257
  (
    n258,
    n35
  );


  not
  g258
  (
    n250,
    n38
  );


  buf
  g259
  (
    n188,
    n47
  );


  not
  g260
  (
    n227,
    n45
  );


  buf
  g261
  (
    n138,
    n61
  );


  buf
  g262
  (
    n292,
    n41
  );


  buf
  g263
  (
    n276,
    n47
  );


  not
  g264
  (
    n169,
    n56
  );


  not
  g265
  (
    n306,
    n57
  );


  buf
  g266
  (
    n104,
    n83
  );


  buf
  g267
  (
    n119,
    n50
  );


  not
  g268
  (
    n254,
    n67
  );


  buf
  g269
  (
    n309,
    n39
  );


  not
  g270
  (
    n149,
    n59
  );


  not
  g271
  (
    n245,
    n67
  );


  not
  g272
  (
    n269,
    n57
  );


  not
  g273
  (
    n103,
    n77
  );


  buf
  g274
  (
    n132,
    n68
  );


  not
  g275
  (
    n263,
    n37
  );


  not
  g276
  (
    KeyWire_0_21,
    n60
  );


  not
  g277
  (
    n189,
    n84
  );


  nand
  g278
  (
    n136,
    n40,
    n49
  );


  xnor
  g279
  (
    n283,
    n34,
    n84
  );


  not
  g280
  (
    n422,
    n115
  );


  buf
  g281
  (
    n515,
    n252
  );


  not
  g282
  (
    n506,
    n274
  );


  buf
  g283
  (
    n320,
    n306
  );


  not
  g284
  (
    n380,
    n275
  );


  not
  g285
  (
    n488,
    n222
  );


  buf
  g286
  (
    n465,
    n302
  );


  buf
  g287
  (
    n388,
    n194
  );


  not
  g288
  (
    n360,
    n209
  );


  buf
  g289
  (
    n348,
    n241
  );


  not
  g290
  (
    n385,
    n281
  );


  buf
  g291
  (
    n510,
    n284
  );


  not
  g292
  (
    n521,
    n148
  );


  buf
  g293
  (
    n502,
    n233
  );


  buf
  g294
  (
    n410,
    n153
  );


  buf
  g295
  (
    n436,
    n131
  );


  not
  g296
  (
    n389,
    n246
  );


  not
  g297
  (
    n492,
    n192
  );


  buf
  g298
  (
    n413,
    n244
  );


  not
  g299
  (
    n401,
    n295
  );


  buf
  g300
  (
    n334,
    n95
  );


  buf
  g301
  (
    n325,
    n194
  );


  buf
  g302
  (
    n359,
    n179
  );


  not
  g303
  (
    n527,
    n279
  );


  buf
  g304
  (
    n343,
    n237
  );


  or
  g305
  (
    n407,
    n120,
    n107,
    n238
  );


  nor
  g306
  (
    n368,
    n204,
    n119,
    n146,
    n122
  );


  nand
  g307
  (
    n361,
    n234,
    n244,
    n209,
    n205
  );


  nand
  g308
  (
    n322,
    n189,
    n162,
    n194,
    n143
  );


  and
  g309
  (
    n376,
    n232,
    n132,
    n256,
    n240
  );


  xor
  g310
  (
    n524,
    n197,
    n129,
    n227,
    n154
  );


  nand
  g311
  (
    KeyWire_0_0,
    n98,
    n303,
    n122,
    n123
  );


  nand
  g312
  (
    n347,
    n131,
    n243,
    n197,
    n114
  );


  or
  g313
  (
    n326,
    n250,
    n200,
    n180,
    n214
  );


  nor
  g314
  (
    n365,
    n149,
    n252,
    n120,
    n248
  );


  nand
  g315
  (
    n481,
    n222,
    n227,
    n183,
    n198
  );


  xnor
  g316
  (
    n315,
    n287,
    n273,
    n305,
    n111
  );


  or
  g317
  (
    n509,
    n190,
    n256,
    n192,
    n201
  );


  xor
  g318
  (
    n471,
    n221,
    n218,
    n157,
    n300
  );


  nor
  g319
  (
    KeyWire_0_18,
    n113,
    n126,
    n160,
    n198
  );


  xor
  g320
  (
    n335,
    n152,
    n304,
    n291,
    n230
  );


  nand
  g321
  (
    n454,
    n303,
    n137,
    n197,
    n225
  );


  or
  g322
  (
    n406,
    n265,
    n285,
    n261,
    n166
  );


  nor
  g323
  (
    n450,
    n263,
    n258,
    n140,
    n186
  );


  nand
  g324
  (
    n369,
    n132,
    n188,
    n281,
    n161
  );


  xor
  g325
  (
    n329,
    n287,
    n224,
    n213,
    n272
  );


  or
  g326
  (
    n372,
    n182,
    n167,
    n96,
    n186
  );


  and
  g327
  (
    n351,
    n257,
    n126,
    n169,
    n155
  );


  or
  g328
  (
    n392,
    n292,
    n311,
    n163,
    n180
  );


  xnor
  g329
  (
    n536,
    n211,
    n114,
    n226,
    n204
  );


  xnor
  g330
  (
    n434,
    n181,
    n261,
    n262,
    n172
  );


  nand
  g331
  (
    n513,
    n297,
    n259,
    n156
  );


  xnor
  g332
  (
    n331,
    n217,
    n280,
    n235,
    n267
  );


  xor
  g333
  (
    n512,
    n187,
    n212,
    n191,
    n160
  );


  and
  g334
  (
    n340,
    n133,
    n293,
    n147,
    n260
  );


  and
  g335
  (
    n328,
    n264,
    n275,
    n212,
    n127
  );


  nor
  g336
  (
    n519,
    n110,
    n215,
    n254,
    n284
  );


  xor
  g337
  (
    n429,
    n302,
    n228,
    n220,
    n117
  );


  xor
  g338
  (
    n445,
    n311,
    n301,
    n156
  );


  and
  g339
  (
    n461,
    n269,
    n118,
    n250,
    n248
  );


  xnor
  g340
  (
    n474,
    n208,
    n161,
    n298,
    n300
  );


  and
  g341
  (
    n458,
    n285,
    n189,
    n283,
    n133
  );


  xnor
  g342
  (
    KeyWire_0_19,
    n132,
    n281,
    n307,
    n187
  );


  xor
  g343
  (
    n336,
    n242,
    n143,
    n192,
    n247
  );


  and
  g344
  (
    n396,
    n182,
    n292,
    n307,
    n240
  );


  xnor
  g345
  (
    n468,
    n115,
    n230,
    n271,
    n268
  );


  and
  g346
  (
    n467,
    n215,
    n207,
    n276,
    n231
  );


  xnor
  g347
  (
    n425,
    n176,
    n185,
    n239,
    n291
  );


  and
  g348
  (
    n428,
    n186,
    n274,
    n262,
    n256
  );


  and
  g349
  (
    n377,
    n128,
    n243,
    n105,
    n312
  );


  and
  g350
  (
    n456,
    n128,
    n112,
    n174,
    n251
  );


  xnor
  g351
  (
    n324,
    n257,
    n293,
    n116,
    n136
  );


  or
  g352
  (
    n400,
    n240,
    n137,
    n229,
    n290
  );


  nor
  g353
  (
    n391,
    n195,
    n151,
    n207,
    n310
  );


  and
  g354
  (
    n432,
    n119,
    n254,
    n150,
    n249
  );


  nor
  g355
  (
    n424,
    n190,
    n209,
    n267,
    n126
  );


  nand
  g356
  (
    n350,
    n145,
    n287,
    n129,
    n264
  );


  xnor
  g357
  (
    n316,
    n247,
    n142,
    n284,
    n299
  );


  or
  g358
  (
    n358,
    n221,
    n308,
    n268,
    n302
  );


  xor
  g359
  (
    n490,
    n179,
    n251,
    n295,
    n289
  );


  nand
  g360
  (
    n382,
    n238,
    n248,
    n149,
    n121
  );


  or
  g361
  (
    n446,
    n177,
    n118,
    n131,
    n191
  );


  nand
  g362
  (
    n356,
    n290,
    n232,
    n231,
    n223
  );


  nand
  g363
  (
    n491,
    n261,
    n282,
    n127,
    n300
  );


  or
  g364
  (
    n375,
    n130,
    n152,
    n211,
    n164
  );


  or
  g365
  (
    n395,
    n193,
    n147,
    n108,
    n245
  );


  nand
  g366
  (
    n397,
    n183,
    n310,
    n168,
    n180
  );


  nand
  g367
  (
    n405,
    n151,
    n224,
    n102,
    n110
  );


  and
  g368
  (
    n433,
    n295,
    n303,
    n164,
    n130
  );


  nor
  g369
  (
    n473,
    n203,
    n188,
    n182,
    n197
  );


  nor
  g370
  (
    n323,
    n192,
    n127,
    n170,
    n157
  );


  xnor
  g371
  (
    n470,
    n280,
    n148,
    n237,
    n135
  );


  nand
  g372
  (
    n330,
    n123,
    n161,
    n239,
    n133
  );


  nand
  g373
  (
    n440,
    n119,
    n114,
    n175,
    n117
  );


  xnor
  g374
  (
    n525,
    n157,
    n171,
    n238
  );


  nand
  g375
  (
    n399,
    n205,
    n174,
    n182,
    n200
  );


  nand
  g376
  (
    n487,
    n208,
    n276,
    n181,
    n202
  );


  nand
  g377
  (
    n498,
    n198,
    n181,
    n231,
    n210
  );


  or
  g378
  (
    n416,
    n116,
    n275,
    n273,
    n124
  );


  xnor
  g379
  (
    n507,
    n135,
    n282,
    n144,
    n226
  );


  xor
  g380
  (
    KeyWire_0_16,
    n232,
    n195,
    n201,
    n306
  );


  nor
  g381
  (
    n533,
    n113,
    n139,
    n162,
    n178
  );


  or
  g382
  (
    n370,
    n199,
    n278,
    n220,
    n134
  );


  xnor
  g383
  (
    n530,
    n269,
    n159,
    n257,
    n264
  );


  nor
  g384
  (
    n535,
    n153,
    n134,
    n196,
    n117
  );


  xnor
  g385
  (
    n408,
    n220,
    n289,
    n183,
    n247
  );


  nor
  g386
  (
    n520,
    n97,
    n199,
    n311,
    n125
  );


  or
  g387
  (
    n341,
    n218,
    n246,
    n127,
    n233
  );


  nand
  g388
  (
    n353,
    n233,
    n170,
    n139,
    n158
  );


  nor
  g389
  (
    n415,
    n125,
    n265,
    n169,
    n189
  );


  xnor
  g390
  (
    n384,
    n159,
    n160,
    n219,
    n106
  );


  xnor
  g391
  (
    n466,
    n250,
    n301,
    n270,
    n132
  );


  nor
  g392
  (
    n534,
    n137,
    n277,
    n164,
    n138
  );


  and
  g393
  (
    n398,
    n238,
    n174,
    n186,
    n206
  );


  xnor
  g394
  (
    n532,
    n220,
    n288,
    n279,
    n225
  );


  or
  g395
  (
    n459,
    n241,
    n138,
    n297,
    n150
  );


  xor
  g396
  (
    n478,
    n158,
    n228,
    n149,
    n237
  );


  or
  g397
  (
    n448,
    n258,
    n154,
    n202,
    n204
  );


  nor
  g398
  (
    n414,
    n296,
    n130,
    n185,
    n274
  );


  and
  g399
  (
    n318,
    n263,
    n249,
    n286,
    n142
  );


  nor
  g400
  (
    n503,
    n114,
    n279,
    n294,
    n283
  );


  xnor
  g401
  (
    n486,
    n266,
    n190,
    n234,
    n163
  );


  xor
  g402
  (
    n423,
    n184,
    n118,
    n155,
    n295
  );


  and
  g403
  (
    n362,
    n212,
    n140,
    n223,
    n281
  );


  xor
  g404
  (
    KeyWire_0_9,
    n144,
    n128,
    n206,
    n293
  );


  nor
  g405
  (
    n420,
    n239,
    n250,
    n310,
    n252
  );


  or
  g406
  (
    n319,
    n294,
    n162,
    n235,
    n213
  );


  nor
  g407
  (
    n390,
    n247,
    n145,
    n169,
    n305
  );


  nor
  g408
  (
    n526,
    n101,
    n171,
    n143,
    n312
  );


  or
  g409
  (
    n497,
    n149,
    n183,
    n305,
    n165
  );


  xor
  g410
  (
    n484,
    n206,
    n218,
    n151,
    n139
  );


  nor
  g411
  (
    n374,
    n249,
    n268,
    n272,
    n211
  );


  xor
  g412
  (
    n452,
    n194,
    n161,
    n258,
    n239
  );


  nor
  g413
  (
    n495,
    n271,
    n152,
    n138,
    n270
  );


  and
  g414
  (
    n494,
    n156,
    n291,
    n171,
    n308
  );


  or
  g415
  (
    n313,
    n141,
    n120,
    n255
  );


  nor
  g416
  (
    n485,
    n282,
    n229,
    n178,
    n145
  );


  nor
  g417
  (
    n505,
    n219,
    n244,
    n307,
    n170
  );


  xor
  g418
  (
    n443,
    n211,
    n209,
    n305,
    n283
  );


  xor
  g419
  (
    n455,
    n241,
    n109,
    n168,
    n262
  );


  or
  g420
  (
    n508,
    n189,
    n306,
    n245,
    n289
  );


  or
  g421
  (
    n531,
    n286,
    n205,
    n258,
    n228
  );


  xnor
  g422
  (
    n516,
    n107,
    n289,
    n144,
    n270
  );


  nand
  g423
  (
    n381,
    n278,
    n147,
    n185,
    n304
  );


  xnor
  g424
  (
    n537,
    n263,
    n172,
    n103,
    n205
  );


  xor
  g425
  (
    n480,
    n184,
    n301,
    n179,
    n146
  );


  and
  g426
  (
    n464,
    n175,
    n196,
    n141,
    n165
  );


  and
  g427
  (
    n349,
    n219,
    n300,
    n296,
    n199
  );


  xor
  g428
  (
    n449,
    n290,
    n292,
    n135,
    n166
  );


  xnor
  g429
  (
    n344,
    n100,
    n168,
    n298,
    n142
  );


  xor
  g430
  (
    n462,
    n187,
    n165,
    n271,
    n210
  );


  and
  g431
  (
    n373,
    n108,
    n140,
    n285,
    n272
  );


  xor
  g432
  (
    n418,
    n118,
    n309,
    n163,
    n282
  );


  xor
  g433
  (
    n421,
    n273,
    n213,
    n280,
    n166
  );


  nor
  g434
  (
    n511,
    n252,
    n165,
    n116,
    n288
  );


  nor
  g435
  (
    n447,
    n271,
    n279,
    n302,
    n122
  );


  and
  g436
  (
    n489,
    n117,
    n259,
    n301,
    n123
  );


  nand
  g437
  (
    n430,
    n172,
    n218,
    n99,
    n260
  );


  nor
  g438
  (
    n327,
    n277,
    n172,
    n265,
    n125
  );


  nor
  g439
  (
    n332,
    n254,
    n249,
    n124,
    n164
  );


  xor
  g440
  (
    n366,
    n276,
    n200,
    n236,
    n126
  );


  xnor
  g441
  (
    n517,
    n213,
    n157,
    n122,
    n221
  );


  and
  g442
  (
    n475,
    n241,
    n216,
    n296,
    n178
  );


  xor
  g443
  (
    n367,
    n141,
    n115,
    n112,
    n296
  );


  xnor
  g444
  (
    n460,
    n150,
    n173,
    n188,
    n266
  );


  xor
  g445
  (
    n442,
    n145,
    n304,
    n288,
    n203
  );


  or
  g446
  (
    n393,
    n169,
    n146,
    n261,
    n124
  );


  nor
  g447
  (
    KeyWire_0_14,
    n217,
    n173,
    n308,
    n159
  );


  xor
  g448
  (
    n499,
    n160,
    n297,
    n193,
    n128
  );


  xor
  g449
  (
    n501,
    n229,
    n185,
    n280,
    n225
  );


  and
  g450
  (
    n402,
    n224,
    n299,
    n210
  );


  nor
  g451
  (
    n518,
    n177,
    n304,
    n204,
    n215
  );


  nand
  g452
  (
    n379,
    n106,
    n294,
    n167,
    n153
  );


  and
  g453
  (
    n522,
    n248,
    n269,
    n255,
    n188
  );


  xnor
  g454
  (
    n476,
    n216,
    n176,
    n170,
    n299
  );


  or
  g455
  (
    n317,
    n309,
    n264,
    n255,
    n175
  );


  xnor
  g456
  (
    n411,
    n286,
    n227,
    n195,
    n236
  );


  and
  g457
  (
    n528,
    n141,
    n235,
    n263,
    n129
  );


  xor
  g458
  (
    n453,
    n148,
    n253,
    n243,
    n153
  );


  xor
  g459
  (
    n472,
    n136,
    n173,
    n278,
    n276
  );


  nor
  g460
  (
    n469,
    n159,
    n303,
    n190,
    n312
  );


  and
  g461
  (
    n431,
    n288,
    n253,
    n196,
    n232
  );


  and
  g462
  (
    KeyWire_0_29,
    n137,
    n158,
    n176,
    n140
  );


  and
  g463
  (
    n387,
    n207,
    n254,
    n155,
    n146
  );


  xor
  g464
  (
    n479,
    n119,
    n163,
    n272,
    n166
  );


  or
  g465
  (
    n403,
    n135,
    n230,
    n222,
    n291
  );


  or
  g466
  (
    n483,
    n262,
    n150,
    n202,
    n310
  );


  or
  g467
  (
    n339,
    n139,
    n177,
    n290,
    n234
  );


  xor
  g468
  (
    n457,
    n246,
    n116,
    n113,
    n215
  );


  nor
  g469
  (
    n493,
    n200,
    n268,
    n226,
    n158
  );


  and
  g470
  (
    n412,
    n193,
    n222,
    n226,
    n143
  );


  nor
  g471
  (
    n378,
    n277,
    n267,
    n307,
    n191
  );


  or
  g472
  (
    n417,
    n246,
    n308,
    n179,
    n242
  );


  xnor
  g473
  (
    n363,
    n278,
    n242,
    n124,
    n233
  );


  xor
  g474
  (
    KeyWire_0_30,
    n236,
    n136,
    n256,
    n123
  );


  xnor
  g475
  (
    n371,
    n230,
    n113,
    n287,
    n275
  );


  xnor
  g476
  (
    n345,
    n109,
    n237,
    n298,
    n144
  );


  or
  g477
  (
    n314,
    n214,
    n184,
    n235,
    n298
  );


  nor
  g478
  (
    n477,
    n236,
    n216,
    n181,
    n136
  );


  xnor
  g479
  (
    n441,
    n231,
    n177,
    n253,
    n104
  );


  xnor
  g480
  (
    n427,
    n178,
    n286,
    n221,
    n196
  );


  nand
  g481
  (
    n496,
    n125,
    n223,
    n111,
    n133
  );


  xor
  g482
  (
    n409,
    n201,
    n212,
    n203,
    n245
  );


  nor
  g483
  (
    n386,
    n174,
    n147,
    n306,
    n217
  );


  xor
  g484
  (
    n383,
    n175,
    n223,
    n167,
    n115
  );


  nor
  g485
  (
    n529,
    n208,
    n270,
    n201,
    n199
  );


  xor
  g486
  (
    n364,
    n267,
    n195,
    n173,
    n180
  );


  xor
  g487
  (
    n500,
    n152,
    n142,
    n202,
    n121
  );


  xor
  g488
  (
    n482,
    n216,
    n155,
    n255,
    n154
  );


  or
  g489
  (
    n463,
    n251,
    n198,
    n134,
    n227
  );


  xor
  g490
  (
    n333,
    n121,
    n176,
    n269,
    n130
  );


  or
  g491
  (
    n523,
    n265,
    n266,
    n309
  );


  or
  g492
  (
    n357,
    n240,
    n129,
    n228,
    n225
  );


  or
  g493
  (
    n394,
    n284,
    n259,
    n138,
    n121
  );


  nand
  g494
  (
    n426,
    n277,
    n214,
    n208,
    n229
  );


  and
  g495
  (
    n342,
    n253,
    n266,
    n219,
    n191
  );


  and
  g496
  (
    n321,
    n207,
    n154,
    n260,
    n151
  );


  nor
  g497
  (
    KeyWire_0_2,
    n206,
    n243,
    n162,
    n242
  );


  and
  g498
  (
    n514,
    n299,
    n184,
    n260,
    n134
  );


  xnor
  g499
  (
    n346,
    n294,
    n203,
    n187,
    n148
  );


  or
  g500
  (
    n451,
    n168,
    n257,
    n217,
    n167
  );


  xnor
  g501
  (
    n404,
    n293,
    n273,
    n224,
    n274
  );


  nor
  g502
  (
    n355,
    n131,
    n292,
    n214,
    n285
  );


  and
  g503
  (
    n435,
    n245,
    n283,
    n234,
    n244
  );


  xnor
  g504
  (
    n338,
    n193,
    n311,
    n297,
    n251
  );


  not
  g505
  (
    KeyWire_0_28,
    n324
  );


  not
  g506
  (
    n565,
    n341
  );


  buf
  g507
  (
    n559,
    n343
  );


  buf
  g508
  (
    n567,
    n332
  );


  buf
  g509
  (
    n539,
    n318
  );


  buf
  g510
  (
    n553,
    n333
  );


  not
  g511
  (
    n560,
    n336
  );


  not
  g512
  (
    n556,
    n321
  );


  buf
  g513
  (
    n543,
    n313
  );


  not
  g514
  (
    n549,
    n337
  );


  not
  g515
  (
    n545,
    n329
  );


  not
  g516
  (
    n554,
    n315
  );


  buf
  g517
  (
    n551,
    n330
  );


  buf
  g518
  (
    n561,
    n331
  );


  not
  g519
  (
    n542,
    n326
  );


  buf
  g520
  (
    n558,
    n328
  );


  buf
  g521
  (
    n541,
    n325
  );


  buf
  g522
  (
    n562,
    n340
  );


  not
  g523
  (
    n546,
    n316
  );


  buf
  g524
  (
    n538,
    n323
  );


  buf
  g525
  (
    n566,
    n320
  );


  not
  g526
  (
    n552,
    n319
  );


  buf
  g527
  (
    n555,
    n342
  );


  not
  g528
  (
    n547,
    n322
  );


  not
  g529
  (
    n564,
    n314
  );


  buf
  g530
  (
    n550,
    n338
  );


  buf
  g531
  (
    n540,
    n339
  );


  buf
  g532
  (
    n557,
    n334
  );


  buf
  g533
  (
    n568,
    n344
  );


  buf
  g534
  (
    n544,
    n327
  );


  buf
  g535
  (
    n563,
    n317
  );


  not
  g536
  (
    n548,
    n335
  );


  xor
  g537
  (
    n587,
    n389,
    n555,
    n350,
    n538
  );


  or
  g538
  (
    n609,
    n397,
    n560,
    n379,
    n551
  );


  nor
  g539
  (
    n593,
    n544,
    n548,
    n557,
    n550
  );


  nand
  g540
  (
    n573,
    n552,
    n358,
    n538,
    n558
  );


  xor
  g541
  (
    n608,
    n346,
    n382,
    n391,
    n556
  );


  xnor
  g542
  (
    n588,
    n549,
    n540,
    n557,
    n548
  );


  xor
  g543
  (
    n605,
    n558,
    n551,
    n542
  );


  or
  g544
  (
    n610,
    n549,
    n405,
    n406,
    n556
  );


  or
  g545
  (
    n581,
    n543,
    n407,
    n357,
    n551
  );


  nand
  g546
  (
    n604,
    n553,
    n549,
    n403,
    n547
  );


  xnor
  g547
  (
    n599,
    n553,
    n559,
    n372,
    n366
  );


  xor
  g548
  (
    n592,
    n562,
    n400,
    n553,
    n549
  );


  xnor
  g549
  (
    n584,
    n556,
    n557,
    n560,
    n351
  );


  xor
  g550
  (
    n611,
    n396,
    n393,
    n392,
    n561
  );


  nand
  g551
  (
    n574,
    n557,
    n378,
    n554,
    n547
  );


  xnor
  g552
  (
    n591,
    n552,
    n545,
    n558,
    n561
  );


  nand
  g553
  (
    n606,
    n563,
    n362,
    n556,
    n545
  );


  xnor
  g554
  (
    n579,
    n552,
    n554,
    n348,
    n386
  );


  xor
  g555
  (
    n603,
    n543,
    n373,
    n552,
    n560
  );


  xor
  g556
  (
    n595,
    n558,
    n365,
    n539,
    n554
  );


  or
  g557
  (
    n576,
    n371,
    n561,
    n548,
    n559
  );


  and
  g558
  (
    n597,
    n395,
    n555,
    n375,
    n547
  );


  nor
  g559
  (
    n596,
    n347,
    n541,
    n367,
    n399
  );


  nand
  g560
  (
    n572,
    n388,
    n540,
    n368,
    n408
  );


  nor
  g561
  (
    n589,
    n561,
    n555,
    n398,
    n544
  );


  nor
  g562
  (
    n577,
    n550,
    n359,
    n410,
    n544
  );


  nor
  g563
  (
    n594,
    n364,
    n550,
    n354,
    n562
  );


  xor
  g564
  (
    KeyWire_0_20,
    n548,
    n562,
    n352,
    n546
  );


  and
  g565
  (
    n600,
    n394,
    n380,
    n550,
    n401
  );


  xnor
  g566
  (
    n570,
    n559,
    n541,
    n387
  );


  xor
  g567
  (
    n583,
    n545,
    n374,
    n377,
    n543
  );


  and
  g568
  (
    n578,
    n538,
    n546,
    n360,
    n361
  );


  nand
  g569
  (
    n571,
    n562,
    n538,
    n543,
    n404
  );


  xor
  g570
  (
    n598,
    n409,
    n411,
    n560,
    n355
  );


  nor
  g571
  (
    n602,
    n540,
    n544,
    n356,
    n376
  );


  or
  g572
  (
    n601,
    n369,
    n546,
    n349
  );


  xor
  g573
  (
    n575,
    n545,
    n381,
    n363,
    n390
  );


  nor
  g574
  (
    n586,
    n383,
    n402,
    n547,
    n555
  );


  nand
  g575
  (
    n607,
    n559,
    n551,
    n353,
    n385
  );


  nor
  g576
  (
    n590,
    n370,
    n384,
    n541,
    n539
  );


  or
  g577
  (
    n580,
    n539,
    n345,
    n542,
    n554
  );


  or
  g578
  (
    n585,
    n539,
    n540,
    n542,
    n553
  );


  buf
  g579
  (
    n710,
    n425
  );


  not
  g580
  (
    n704,
    n423
  );


  buf
  g581
  (
    n616,
    n526
  );


  buf
  g582
  (
    n663,
    n519
  );


  not
  g583
  (
    n639,
    n457
  );


  buf
  g584
  (
    n671,
    n518
  );


  buf
  g585
  (
    n674,
    n452
  );


  not
  g586
  (
    n656,
    n494
  );


  not
  g587
  (
    n638,
    n604
  );


  buf
  g588
  (
    n682,
    n414
  );


  buf
  g589
  (
    n654,
    n418
  );


  buf
  g590
  (
    n633,
    n480
  );


  not
  g591
  (
    n643,
    n590
  );


  buf
  g592
  (
    n667,
    n495
  );


  not
  g593
  (
    n673,
    n570
  );


  not
  g594
  (
    n650,
    n571
  );


  not
  g595
  (
    n689,
    n492
  );


  buf
  g596
  (
    n670,
    n601
  );


  not
  g597
  (
    n620,
    n578
  );


  buf
  g598
  (
    n641,
    n606
  );


  not
  g599
  (
    n653,
    n599
  );


  not
  g600
  (
    n617,
    n474
  );


  buf
  g601
  (
    n632,
    n594
  );


  not
  g602
  (
    n694,
    n586
  );


  buf
  g603
  (
    n708,
    n588
  );


  buf
  g604
  (
    n651,
    n600
  );


  not
  g605
  (
    n669,
    n609
  );


  buf
  g606
  (
    n627,
    n603
  );


  not
  g607
  (
    n705,
    n580
  );


  buf
  g608
  (
    n649,
    n517
  );


  not
  g609
  (
    n677,
    n597
  );


  buf
  g610
  (
    n692,
    n606
  );


  buf
  g611
  (
    n672,
    n593
  );


  buf
  g612
  (
    n644,
    n603
  );


  and
  g613
  (
    n681,
    n584,
    n466
  );


  nand
  g614
  (
    n684,
    n522,
    n500,
    n472
  );


  xor
  g615
  (
    n648,
    n590,
    n481,
    n593
  );


  nor
  g616
  (
    n629,
    n523,
    n522,
    n484
  );


  or
  g617
  (
    n699,
    n470,
    n415,
    n525
  );


  nor
  g618
  (
    n647,
    n434,
    n601,
    n485
  );


  xnor
  g619
  (
    n675,
    n525,
    n511,
    n476
  );


  xnor
  g620
  (
    n614,
    n413,
    n486,
    n591
  );


  nand
  g621
  (
    n652,
    n607,
    n438,
    n462
  );


  and
  g622
  (
    n662,
    n579,
    n589,
    n524
  );


  xor
  g623
  (
    n626,
    n589,
    n468,
    n600
  );


  nor
  g624
  (
    n621,
    n488,
    n611,
    n513
  );


  xor
  g625
  (
    n623,
    n524,
    n523,
    n499
  );


  or
  g626
  (
    n660,
    n464,
    n602,
    n465
  );


  xor
  g627
  (
    n707,
    n510,
    n508,
    n603
  );


  or
  g628
  (
    n695,
    n574,
    n427,
    n599
  );


  xor
  g629
  (
    n679,
    n442,
    n420,
    n514
  );


  xnor
  g630
  (
    n655,
    n597,
    n610,
    n606
  );


  xnor
  g631
  (
    n622,
    n595,
    n610,
    n523
  );


  xor
  g632
  (
    n698,
    n597,
    n525,
    n512
  );


  nor
  g633
  (
    n657,
    n455,
    n603,
    n460
  );


  or
  g634
  (
    n640,
    n467,
    n443,
    n421
  );


  or
  g635
  (
    n624,
    n497,
    n596,
    n608
  );


  nand
  g636
  (
    n618,
    n521,
    n439,
    n482
  );


  xor
  g637
  (
    n666,
    n597,
    n610,
    n430
  );


  or
  g638
  (
    n680,
    n431,
    n602,
    n594
  );


  xor
  g639
  (
    n625,
    n473,
    n582,
    n605
  );


  nand
  g640
  (
    n615,
    n609,
    n489,
    n422
  );


  xnor
  g641
  (
    n645,
    n583,
    n501,
    n461
  );


  or
  g642
  (
    n612,
    n446,
    n428,
    n594
  );


  nor
  g643
  (
    n696,
    n502,
    n504,
    n475
  );


  xor
  g644
  (
    n700,
    n604,
    n520,
    n445
  );


  xor
  g645
  (
    n637,
    n424,
    n435,
    n451
  );


  nor
  g646
  (
    n676,
    n471,
    n606,
    n515
  );


  nand
  g647
  (
    n697,
    n605,
    n595,
    n449
  );


  nor
  g648
  (
    n646,
    n441,
    n573,
    n608
  );


  and
  g649
  (
    n613,
    n509,
    n526,
    n609
  );


  xor
  g650
  (
    KeyWire_0_5,
    n607,
    n516,
    n600
  );


  and
  g651
  (
    n693,
    n506,
    n604,
    n575
  );


  xor
  g652
  (
    n659,
    n598,
    n444,
    n607
  );


  nor
  g653
  (
    n642,
    n602,
    n432,
    n426
  );


  xnor
  g654
  (
    n668,
    n604,
    n463,
    n599
  );


  nand
  g655
  (
    n701,
    n587,
    n601,
    n577
  );


  and
  g656
  (
    n709,
    n419,
    n483,
    n412
  );


  nand
  g657
  (
    n702,
    n598,
    n505,
    n576
  );


  nor
  g658
  (
    n635,
    n596,
    n507,
    n477
  );


  or
  g659
  (
    n687,
    n503,
    n456,
    n522
  );


  nand
  g660
  (
    n683,
    n498,
    n608,
    n600
  );


  nand
  g661
  (
    n630,
    n610,
    n609,
    n491
  );


  or
  g662
  (
    n690,
    n524,
    n522,
    n440
  );


  xor
  g663
  (
    n686,
    n416,
    n453,
    n469
  );


  xnor
  g664
  (
    n661,
    n447,
    n601,
    n433
  );


  or
  g665
  (
    n678,
    n496,
    n596,
    n525
  );


  and
  g666
  (
    n665,
    n607,
    n436,
    n478
  );


  or
  g667
  (
    n685,
    n602,
    n605,
    n585
  );


  xor
  g668
  (
    n691,
    n611,
    n448,
    n458
  );


  nand
  g669
  (
    n664,
    n591,
    n595,
    n487
  );


  and
  g670
  (
    n703,
    n524,
    n479,
    n596
  );


  nor
  g671
  (
    n628,
    n490,
    n526,
    n599
  );


  or
  g672
  (
    n658,
    n572,
    n595,
    n598
  );


  and
  g673
  (
    n634,
    n592,
    n581,
    n523
  );


  nand
  g674
  (
    n688,
    n598,
    n592,
    n493
  );


  or
  g675
  (
    n619,
    n454,
    n459,
    n605
  );


  xor
  g676
  (
    n706,
    n450,
    n608,
    n594
  );


  nor
  g677
  (
    n631,
    n429,
    n417,
    n437
  );


  not
  g678
  (
    n789,
    n698
  );


  not
  g679
  (
    n712,
    n701
  );


  buf
  g680
  (
    n716,
    n689
  );


  buf
  g681
  (
    n794,
    n681
  );


  not
  g682
  (
    n719,
    n657
  );


  buf
  g683
  (
    n726,
    n694
  );


  not
  g684
  (
    n742,
    n696
  );


  buf
  g685
  (
    n715,
    n652
  );


  not
  g686
  (
    n782,
    n699
  );


  buf
  g687
  (
    n778,
    n685
  );


  not
  g688
  (
    n786,
    n648
  );


  buf
  g689
  (
    n757,
    n612
  );


  not
  g690
  (
    n725,
    n618
  );


  xnor
  g691
  (
    n779,
    n687,
    n683,
    n644
  );


  and
  g692
  (
    n720,
    n671,
    n628,
    n657
  );


  and
  g693
  (
    n740,
    n663,
    n563,
    n692,
    n665
  );


  xor
  g694
  (
    n746,
    n673,
    n635,
    n678,
    n669
  );


  or
  g695
  (
    n792,
    n699,
    n704,
    n675,
    n686
  );


  nor
  g696
  (
    n753,
    n566,
    n687,
    n565,
    n677
  );


  nand
  g697
  (
    n744,
    n693,
    n690,
    n661,
    n678
  );


  and
  g698
  (
    n751,
    n696,
    n621,
    n654,
    n564
  );


  and
  g699
  (
    n769,
    n690,
    n692,
    n630,
    n685
  );


  and
  g700
  (
    n730,
    n658,
    n658,
    n662,
    n689
  );


  and
  g701
  (
    n721,
    n681,
    n667,
    n657,
    n666
  );


  nand
  g702
  (
    n729,
    n659,
    n675,
    n702,
    n697
  );


  nand
  g703
  (
    n745,
    n659,
    n653,
    n636,
    n686
  );


  nor
  g704
  (
    n758,
    n663,
    n633,
    n680,
    n614
  );


  or
  g705
  (
    n766,
    n705,
    n673,
    n653,
    n649
  );


  xor
  g706
  (
    n755,
    n564,
    n702,
    n674,
    n566
  );


  xor
  g707
  (
    n761,
    n684,
    n653,
    n689,
    n691
  );


  xor
  g708
  (
    n734,
    n674,
    n656,
    n700,
    n704
  );


  or
  g709
  (
    n732,
    n620,
    n649,
    n683,
    n703
  );


  or
  g710
  (
    n723,
    n706,
    n694,
    n651,
    n674
  );


  xor
  g711
  (
    n780,
    n691,
    n646,
    n656
  );


  xor
  g712
  (
    n773,
    n658,
    n659,
    n563,
    n691
  );


  and
  g713
  (
    n722,
    n648,
    n650,
    n669,
    n660
  );


  and
  g714
  (
    n748,
    n646,
    n651,
    n687,
    n670
  );


  or
  g715
  (
    n763,
    n676,
    n655,
    n688,
    n654
  );


  nand
  g716
  (
    n733,
    n658,
    n703,
    n672,
    n662
  );


  xor
  g717
  (
    n777,
    n627,
    n647,
    n694,
    n684
  );


  nand
  g718
  (
    n776,
    n702,
    n674,
    n654,
    n678
  );


  nor
  g719
  (
    n790,
    n654,
    n647,
    n698,
    n677
  );


  xnor
  g720
  (
    n727,
    n697,
    n672,
    n565,
    n649
  );


  or
  g721
  (
    n767,
    n661,
    n671,
    n664,
    n701
  );


  or
  g722
  (
    KeyWire_0_13,
    n677,
    n655,
    n704,
    n637
  );


  and
  g723
  (
    n749,
    n666,
    n653,
    n697,
    n706
  );


  and
  g724
  (
    n775,
    n672,
    n705,
    n615,
    n565
  );


  xnor
  g725
  (
    n717,
    n703,
    n657,
    n699,
    n704
  );


  and
  g726
  (
    n735,
    n663,
    n659,
    n632,
    n644
  );


  xor
  g727
  (
    n738,
    n675,
    n660,
    n631,
    n626
  );


  and
  g728
  (
    n714,
    n690,
    n639,
    n649,
    n695
  );


  or
  g729
  (
    n768,
    n640,
    n701,
    n695,
    n670
  );


  or
  g730
  (
    KeyWire_0_6,
    n651,
    n655,
    n648,
    n669
  );


  xor
  g731
  (
    n765,
    n680,
    n617,
    n673,
    n645
  );


  xor
  g732
  (
    n756,
    n676,
    n702,
    n651,
    n667
  );


  nor
  g733
  (
    n760,
    n696,
    n689,
    n661,
    n685
  );


  xnor
  g734
  (
    n784,
    n641,
    n650,
    n670,
    n625
  );


  or
  g735
  (
    n741,
    n701,
    n700,
    n566,
    n675
  );


  nor
  g736
  (
    n739,
    n693,
    n661,
    n662,
    n668
  );


  and
  g737
  (
    n752,
    n706,
    n652,
    n664,
    n662
  );


  nand
  g738
  (
    n788,
    n699,
    n698,
    n679,
    n673
  );


  xor
  g739
  (
    n754,
    n685,
    n665,
    n613,
    n681
  );


  and
  g740
  (
    n737,
    n677,
    n694,
    n648,
    n664
  );


  nand
  g741
  (
    n762,
    n697,
    n693,
    n688,
    n686
  );


  and
  g742
  (
    n736,
    n681,
    n668,
    n705
  );


  nor
  g743
  (
    n791,
    n684,
    n676,
    n705,
    n683
  );


  xnor
  g744
  (
    n781,
    n688,
    n666,
    n668
  );


  and
  g745
  (
    n759,
    n691,
    n682,
    n652,
    n643
  );


  nand
  g746
  (
    n728,
    n682,
    n700,
    n678,
    n564
  );


  and
  g747
  (
    KeyWire_0_24,
    n700,
    n680,
    n687,
    n698
  );


  nor
  g748
  (
    n793,
    n619,
    n652,
    n660,
    n703
  );


  xor
  g749
  (
    n743,
    n690,
    n622,
    n566,
    n671
  );


  xor
  g750
  (
    n783,
    n671,
    n623,
    n638,
    n672
  );


  or
  g751
  (
    n774,
    n629,
    n684,
    n656,
    n647
  );


  xnor
  g752
  (
    n772,
    n692,
    n683,
    n634,
    n706
  );


  nor
  g753
  (
    n731,
    n563,
    n616,
    n696,
    n624
  );


  nor
  g754
  (
    n770,
    n656,
    n660,
    n679,
    n665
  );


  nor
  g755
  (
    n785,
    n650,
    n667,
    n647,
    n679
  );


  nor
  g756
  (
    n713,
    n676,
    n669,
    n650,
    n655
  );


  and
  g757
  (
    n711,
    n693,
    n679,
    n695,
    n645
  );


  nand
  g758
  (
    n787,
    n695,
    n670,
    n564,
    n664
  );


  or
  g759
  (
    n771,
    n665,
    n682,
    n646
  );


  xnor
  g760
  (
    n750,
    n663,
    n692,
    n680,
    n667
  );


  and
  g761
  (
    n724,
    n688,
    n565,
    n642,
    n686
  );


  buf
  g762
  (
    n808,
    n713
  );


  not
  g763
  (
    n804,
    n716
  );


  buf
  g764
  (
    n800,
    n718
  );


  buf
  g765
  (
    n802,
    n722
  );


  buf
  g766
  (
    n798,
    n715
  );


  not
  g767
  (
    n803,
    n721
  );


  buf
  g768
  (
    n801,
    n711
  );


  not
  g769
  (
    n805,
    n717
  );


  not
  g770
  (
    n796,
    n719
  );


  not
  g771
  (
    n806,
    n724
  );


  buf
  g772
  (
    n799,
    n714
  );


  not
  g773
  (
    n797,
    n720
  );


  not
  g774
  (
    n795,
    n723
  );


  not
  g775
  (
    n807,
    n712
  );


  buf
  g776
  (
    n823,
    n798
  );


  nand
  g777
  (
    n818,
    n526,
    n802,
    n803
  );


  nor
  g778
  (
    n809,
    n808,
    n799,
    n800,
    n806
  );


  xnor
  g779
  (
    KeyWire_0_3,
    n807,
    n796,
    n312,
    n795
  );


  xnor
  g780
  (
    n811,
    n800,
    n798,
    n805,
    n796
  );


  xnor
  g781
  (
    n822,
    n806,
    n804
  );


  nand
  g782
  (
    n816,
    n805,
    n804,
    n799
  );


  or
  g783
  (
    n821,
    n807,
    n795,
    n800,
    n806
  );


  and
  g784
  (
    n810,
    n801,
    n808,
    n800,
    n798
  );


  nor
  g785
  (
    n824,
    n796,
    n802,
    n805,
    n795
  );


  or
  g786
  (
    n813,
    n799,
    n797,
    n802
  );


  nor
  g787
  (
    n815,
    n798,
    n801,
    n795,
    n88
  );


  nand
  g788
  (
    KeyWire_0_1,
    n801,
    n803
  );


  nor
  g789
  (
    n812,
    n807,
    n802,
    n801,
    n808
  );


  xor
  g790
  (
    n819,
    n807,
    n804,
    n805,
    n797
  );


  xnor
  g791
  (
    n820,
    n797,
    n796,
    n707,
    n808
  );


  not
  g792
  (
    n827,
    n725
  );


  not
  g793
  (
    n830,
    n726
  );


  xnor
  g794
  (
    n829,
    n813,
    n809
  );


  xor
  g795
  (
    n825,
    n729,
    n810,
    n728,
    n816
  );


  and
  g796
  (
    n826,
    n811,
    n814,
    n815,
    n731
  );


  nor
  g797
  (
    n828,
    n817,
    n727,
    n730,
    n812
  );


  not
  g798
  (
    n835,
    n826
  );


  and
  g799
  (
    n831,
    n527,
    n830
  );


  or
  g800
  (
    n832,
    n826,
    n826,
    n827,
    n829
  );


  nand
  g801
  (
    n836,
    n830,
    n830,
    n828,
    n827
  );


  and
  g802
  (
    n833,
    n828,
    n527,
    n827
  );


  nor
  g803
  (
    n834,
    n826,
    n829,
    n527
  );


  and
  g804
  (
    n837,
    n828,
    n828,
    n825,
    n829
  );


  or
  g805
  (
    n841,
    n819,
    n824,
    n529,
    n532
  );


  xnor
  g806
  (
    n838,
    n837,
    n832,
    n530,
    n531
  );


  xor
  g807
  (
    n840,
    n529,
    n822,
    n528,
    n818
  );


  nor
  g808
  (
    n839,
    n532,
    n836,
    n531,
    n821
  );


  xnor
  g809
  (
    n843,
    n831,
    n834,
    n529,
    n835
  );


  nand
  g810
  (
    n842,
    n531,
    n528,
    n527,
    n532
  );


  xnor
  g811
  (
    n845,
    n531,
    n529,
    n530
  );


  nor
  g812
  (
    n846,
    n837,
    n836,
    n528,
    n820
  );


  nand
  g813
  (
    n844,
    n530,
    n833,
    n528,
    n823
  );


  buf
  g814
  (
    n851,
    n841
  );


  not
  g815
  (
    n859,
    n843
  );


  buf
  g816
  (
    n857,
    n843
  );


  not
  g817
  (
    n861,
    n843
  );


  not
  g818
  (
    n860,
    n844
  );


  not
  g819
  (
    n848,
    n842
  );


  buf
  g820
  (
    n858,
    n843
  );


  not
  g821
  (
    n862,
    n842
  );


  buf
  g822
  (
    n847,
    n841
  );


  buf
  g823
  (
    n850,
    n838
  );


  buf
  g824
  (
    n852,
    n840
  );


  buf
  g825
  (
    n849,
    n841
  );


  not
  g826
  (
    n853,
    n842
  );


  not
  g827
  (
    n856,
    n841
  );


  buf
  g828
  (
    n854,
    n842
  );


  buf
  g829
  (
    n855,
    n839
  );


  and
  g830
  (
    n914,
    n92,
    n785,
    n28,
    n780
  );


  nor
  g831
  (
    n874,
    n782,
    n861,
    n846,
    n794
  );


  nand
  g832
  (
    KeyWire_0_10,
    n786,
    n738,
    n92,
    n568
  );


  and
  g833
  (
    n912,
    n783,
    n848,
    n769,
    n747
  );


  nand
  g834
  (
    n876,
    n707,
    n30,
    n788,
    n779
  );


  xnor
  g835
  (
    n894,
    n774,
    n88,
    n567,
    n850
  );


  nand
  g836
  (
    n868,
    n784,
    n854,
    n789,
    n772
  );


  nor
  g837
  (
    n884,
    n848,
    n754,
    n859,
    n771
  );


  nand
  g838
  (
    n864,
    n790,
    n764,
    n776,
    n775
  );


  nor
  g839
  (
    n905,
    n791,
    n777,
    n762,
    n742
  );


  nand
  g840
  (
    n902,
    n847,
    n854,
    n768,
    n855
  );


  nand
  g841
  (
    n911,
    n786,
    n784,
    n790,
    n765
  );


  or
  g842
  (
    n925,
    n756,
    n91,
    n29
  );


  and
  g843
  (
    n901,
    n778,
    n851,
    n739,
    n844
  );


  nand
  g844
  (
    n879,
    n852,
    n788,
    n778,
    n862
  );


  nand
  g845
  (
    n872,
    n734,
    n788,
    n760,
    n708
  );


  xor
  g846
  (
    n906,
    n736,
    n763,
    n785,
    n567
  );


  and
  g847
  (
    n923,
    n785,
    n783,
    n856,
    n740
  );


  and
  g848
  (
    n887,
    n853,
    n861,
    n89,
    n93
  );


  xor
  g849
  (
    n885,
    n751,
    n776,
    n782,
    n791
  );


  xor
  g850
  (
    n866,
    n792,
    n775,
    n791,
    n781
  );


  nand
  g851
  (
    n908,
    n793,
    n859,
    n787,
    n853
  );


  nor
  g852
  (
    n869,
    n845,
    n732,
    n857,
    n794
  );


  xnor
  g853
  (
    n924,
    n852,
    n860,
    n849,
    n848
  );


  nor
  g854
  (
    n903,
    n752,
    n761,
    n94,
    n776
  );


  xnor
  g855
  (
    n873,
    n793,
    n88,
    n780,
    n746
  );


  and
  g856
  (
    n870,
    n779,
    n567,
    n93,
    n847
  );


  xnor
  g857
  (
    n922,
    n854,
    n743,
    n844,
    n852
  );


  xnor
  g858
  (
    n881,
    n90,
    n785,
    n789,
    n757
  );


  and
  g859
  (
    n895,
    n856,
    n775,
    n94,
    n787
  );


  nor
  g860
  (
    n871,
    n847,
    n846,
    n784,
    n855
  );


  and
  g861
  (
    n863,
    n845,
    n758,
    n776,
    n790
  );


  nand
  g862
  (
    n882,
    n846,
    n774,
    n852,
    n791
  );


  xnor
  g863
  (
    n891,
    n769,
    n860,
    n778,
    n90
  );


  nand
  g864
  (
    n875,
    n777,
    n848,
    n91,
    n778
  );


  xor
  g865
  (
    n888,
    n568,
    n789,
    n781
  );


  xor
  g866
  (
    n877,
    n858,
    n845,
    n749,
    n568
  );


  nand
  g867
  (
    n892,
    n857,
    n29,
    n783,
    n766
  );


  nor
  g868
  (
    n899,
    n779,
    n708,
    n794,
    n782
  );


  nor
  g869
  (
    n867,
    n781,
    n768,
    n862,
    n780
  );


  xnor
  g870
  (
    n893,
    n745,
    n790,
    n767,
    n773
  );


  xor
  g871
  (
    n919,
    n759,
    n847,
    n857,
    n861
  );


  xnor
  g872
  (
    n910,
    n767,
    n786,
    n92,
    n770
  );


  nor
  g873
  (
    n886,
    n568,
    n856,
    n748,
    n792
  );


  xnor
  g874
  (
    n897,
    n858,
    n845,
    n862,
    n708
  );


  nand
  g875
  (
    n917,
    n707,
    n851,
    n709,
    n855
  );


  nor
  g876
  (
    n907,
    n88,
    n787,
    n792,
    n753
  );


  nand
  g877
  (
    n909,
    n772,
    n771,
    n28,
    n851
  );


  xnor
  g878
  (
    n896,
    n89,
    n787,
    n780,
    n854
  );


  xor
  g879
  (
    n926,
    n855,
    n777,
    n90,
    n858
  );


  xor
  g880
  (
    n889,
    n708,
    n735,
    n846,
    n773
  );


  nand
  g881
  (
    n900,
    n770,
    n92,
    n850,
    n707
  );


  and
  g882
  (
    n880,
    n793,
    n567,
    n89,
    n856
  );


  nand
  g883
  (
    n878,
    n792,
    n750,
    n744,
    n788
  );


  and
  g884
  (
    n921,
    n29,
    n849,
    n90,
    n858
  );


  xnor
  g885
  (
    n918,
    n777,
    n782,
    n849,
    n844
  );


  or
  g886
  (
    n916,
    n861,
    n794,
    n779,
    n853
  );


  xor
  g887
  (
    n913,
    n781,
    n860,
    n853,
    n775
  );


  nor
  g888
  (
    n915,
    n29,
    n859,
    n793,
    n783
  );


  and
  g889
  (
    n920,
    n94,
    n737,
    n733,
    n849
  );


  xor
  g890
  (
    n883,
    n851,
    n786,
    n93
  );


  nor
  g891
  (
    n904,
    n862,
    n850,
    n755,
    n741
  );


  xor
  g892
  (
    n890,
    n860,
    n94,
    n89,
    n857
  );


  xnor
  g893
  (
    n898,
    n91,
    n859,
    n850,
    n784
  );


  buf
  g894
  (
    n930,
    n864
  );


  not
  g895
  (
    n931,
    n865
  );


  not
  g896
  (
    n927,
    n865
  );


  buf
  g897
  (
    n929,
    n863
  );


  and
  g898
  (
    n928,
    n863,
    n864,
    n866
  );


  or
  g899
  (
    n947,
    n927,
    n879,
    n867,
    n876
  );


  or
  g900
  (
    n950,
    n873,
    n874,
    n929,
    n881
  );


  and
  g901
  (
    n932,
    n868,
    n876,
    n928,
    n869
  );


  xnor
  g902
  (
    n944,
    n878,
    n874,
    n931
  );


  xnor
  g903
  (
    n941,
    n880,
    n930,
    n929,
    n873
  );


  xnor
  g904
  (
    KeyWire_0_25,
    n875,
    n881,
    n879,
    n930
  );


  nand
  g905
  (
    n951,
    n872,
    n881,
    n930,
    n931
  );


  xnor
  g906
  (
    n939,
    n873,
    n928,
    n868
  );


  nand
  g907
  (
    n938,
    n870,
    n871,
    n929
  );


  nand
  g908
  (
    n934,
    n872,
    n878,
    n879,
    n927
  );


  nor
  g909
  (
    n946,
    n880,
    n870,
    n872,
    n931
  );


  xnor
  g910
  (
    n936,
    n880,
    n867,
    n878,
    n877
  );


  xor
  g911
  (
    n940,
    n930,
    n869,
    n874,
    n875
  );


  xor
  g912
  (
    n945,
    n867,
    n871,
    n870,
    n931
  );


  xor
  g913
  (
    n933,
    n871,
    n927,
    n879,
    n868
  );


  nor
  g914
  (
    n948,
    n927,
    n877,
    n867,
    n928
  );


  xor
  g915
  (
    n949,
    n878,
    n881,
    n877,
    n871
  );


  xnor
  g916
  (
    n942,
    n873,
    n870,
    n875,
    n869
  );


  nor
  g917
  (
    n943,
    n872,
    n876,
    n877
  );


  and
  g918
  (
    n937,
    n869,
    n928,
    n880,
    n875
  );


  nand
  g919
  (
    n958,
    n908,
    n886,
    n884
  );


  nand
  g920
  (
    n955,
    n883,
    n898,
    n891,
    n901
  );


  nor
  g921
  (
    n982,
    n951,
    n947,
    n900,
    n945
  );


  xnor
  g922
  (
    n976,
    n948,
    n900,
    n949
  );


  and
  g923
  (
    n983,
    n887,
    n892,
    n889,
    n907
  );


  nand
  g924
  (
    n961,
    n896,
    n905,
    n894
  );


  and
  g925
  (
    n953,
    n893,
    n887,
    n946,
    n897
  );


  xnor
  g926
  (
    n964,
    n896,
    n947,
    n949,
    n883
  );


  xor
  g927
  (
    n975,
    n883,
    n904,
    n951,
    n897
  );


  xnor
  g928
  (
    n956,
    n903,
    n892,
    n950,
    n882
  );


  nand
  g929
  (
    n984,
    n888,
    n902,
    n905,
    n951
  );


  nor
  g930
  (
    n970,
    n900,
    n890,
    n939,
    n949
  );


  nand
  g931
  (
    n962,
    n889,
    n897,
    n940,
    n903
  );


  or
  g932
  (
    n957,
    n898,
    n906,
    n947,
    n944
  );


  and
  g933
  (
    n969,
    n896,
    n943,
    n895,
    n907
  );


  xnor
  g934
  (
    n952,
    n935,
    n906,
    n901,
    n897
  );


  nand
  g935
  (
    n968,
    n882,
    n892,
    n883,
    n950
  );


  xnor
  g936
  (
    n974,
    n887,
    n891,
    n884,
    n893
  );


  nor
  g937
  (
    KeyWire_0_22,
    n946,
    n882,
    n893,
    n894
  );


  xnor
  g938
  (
    n981,
    n895,
    n888,
    n886,
    n907
  );


  and
  g939
  (
    n973,
    n885,
    n890,
    n905,
    n902
  );


  nand
  g940
  (
    n966,
    n891,
    n894,
    n902,
    n948
  );


  xor
  g941
  (
    n986,
    n889,
    n936,
    n891,
    n932
  );


  and
  g942
  (
    n980,
    n890,
    n901,
    n902,
    n884
  );


  nand
  g943
  (
    n959,
    n941,
    n890,
    n899,
    n904
  );


  or
  g944
  (
    n978,
    n947,
    n899,
    n903,
    n889
  );


  or
  g945
  (
    n977,
    n885,
    n892,
    n895,
    n901
  );


  nand
  g946
  (
    n985,
    n900,
    n887,
    n906,
    n934
  );


  nand
  g947
  (
    n954,
    n907,
    n904,
    n938,
    n942
  );


  nand
  g948
  (
    n979,
    n904,
    n899,
    n888,
    n948
  );


  xnor
  g949
  (
    n967,
    n898,
    n896,
    n886,
    n882
  );


  xnor
  g950
  (
    n960,
    n933,
    n893,
    n899,
    n950
  );


  xor
  g951
  (
    n963,
    n885,
    n885,
    n950,
    n903
  );


  and
  g952
  (
    n971,
    n898,
    n888,
    n906,
    n894
  );


  nor
  g953
  (
    n965,
    n884,
    n895,
    n937,
    n948
  );


  xnor
  g954
  (
    n992,
    n910,
    n974,
    n975,
    n971
  );


  or
  g955
  (
    n987,
    n535,
    n970,
    n973,
    n533
  );


  xnor
  g956
  (
    n990,
    n908,
    n533,
    n972,
    n534
  );


  and
  g957
  (
    n989,
    n911,
    n534,
    n977
  );


  and
  g958
  (
    n991,
    n533,
    n533,
    n908,
    n910
  );


  or
  g959
  (
    n993,
    n911,
    n909,
    n910
  );


  or
  g960
  (
    n994,
    n912,
    n976,
    n909,
    n532
  );


  xor
  g961
  (
    KeyWire_0_31,
    n908,
    n911,
    n910,
    n909
  );


  or
  g962
  (
    n988,
    n911,
    n534,
    n535,
    n978
  );


  or
  g963
  (
    n1010,
    n536,
    n913
  );


  nand
  g964
  (
    n1014,
    n986,
    n915,
    n994
  );


  or
  g965
  (
    n1002,
    n710,
    n912,
    n536,
    n918
  );


  xor
  g966
  (
    n1001,
    n984,
    n993,
    n912,
    n569
  );


  nand
  g967
  (
    n997,
    n537,
    n32,
    n981,
    n995
  );


  xnor
  g968
  (
    n1009,
    n915,
    n985,
    n916,
    n32
  );


  and
  g969
  (
    n1004,
    n917,
    n30,
    n611,
    n979
  );


  nand
  g970
  (
    n1005,
    n32,
    n30,
    n917
  );


  or
  g971
  (
    n1013,
    n989,
    n914,
    n710,
    n994
  );


  nand
  g972
  (
    n996,
    n991,
    n995,
    n914,
    n913
  );


  and
  g973
  (
    n1006,
    n992,
    n32,
    n537,
    n987
  );


  xnor
  g974
  (
    n998,
    n535,
    n918,
    n995,
    n537
  );


  xor
  g975
  (
    n1018,
    n536,
    n569,
    n915,
    n917
  );


  xnor
  g976
  (
    n1008,
    n709,
    n535,
    n991,
    n913
  );


  or
  g977
  (
    n1015,
    n31,
    n537,
    n993,
    n914
  );


  or
  g978
  (
    n1000,
    n914,
    n709,
    n990,
    n31
  );


  and
  g979
  (
    n1003,
    n918,
    n993,
    n31,
    n710
  );


  xnor
  g980
  (
    n1016,
    n912,
    n951,
    n988,
    n916
  );


  nand
  g981
  (
    n1011,
    n569,
    n983,
    n31,
    n989
  );


  nor
  g982
  (
    n1012,
    n916,
    n988,
    n982,
    n569
  );


  and
  g983
  (
    n1017,
    n992,
    n710,
    n709,
    n917
  );


  nor
  g984
  (
    KeyWire_0_11,
    n611,
    n915,
    n993,
    n995
  );


  xor
  g985
  (
    n999,
    n990,
    n994,
    n916,
    n980
  );


  or
  g986
  (
    n1029,
    n1005,
    n923,
    n1004,
    n1002
  );


  nand
  g987
  (
    n1024,
    n922,
    n998,
    n925,
    n1006
  );


  xor
  g988
  (
    n1019,
    n996,
    n920,
    n925
  );


  xnor
  g989
  (
    n1032,
    n1000,
    n1016,
    n926,
    n1010
  );


  nand
  g990
  (
    n1022,
    n919,
    n921,
    n925
  );


  nand
  g991
  (
    n1020,
    n920,
    n923,
    n922,
    n1001
  );


  or
  g992
  (
    n1021,
    n920,
    n1011,
    n1018,
    n1007
  );


  xnor
  g993
  (
    n1030,
    n920,
    n923,
    n921,
    n997
  );


  and
  g994
  (
    n1023,
    n924,
    n918,
    n1009,
    n1017
  );


  nor
  g995
  (
    n1028,
    n923,
    n924,
    n926
  );


  nand
  g996
  (
    n1031,
    n1014,
    n919,
    n921,
    n924
  );


  xor
  g997
  (
    n1027,
    n1012,
    n1013,
    n924,
    n922
  );


  or
  g998
  (
    n1026,
    n919,
    n1008,
    n922,
    n999
  );


  or
  g999
  (
    n1025,
    n1015,
    n919,
    n926,
    n1003
  );


  xor
  KeyGate_0_0
  (
    n352,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n817,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n337,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n814,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n62,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n636,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n718,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n285,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n187,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n437,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n865,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n1007,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n110,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n764,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n419,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n111,
    KeyNOTWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n354,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n167,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n439,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n444,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n582,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n222,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    KeyNOTWire_0_22,
    keyIn_0_22,
    KeyWire_0_22
  );


  not
  KeyNOTGate_0_22
  (
    n972,
    KeyNOTWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n107,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n747,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n935,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n256,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n237,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n569,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n504,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n438,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n995,
    KeyNOTWire_0_31
  );


endmodule

