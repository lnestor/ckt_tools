

module Stat_4000_401
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n3772,
  n3769,
  n3786,
  n3787,
  n3783,
  n3784,
  n3792,
  n3793,
  n3790,
  n3989,
  n4000,
  n3998,
  n3987,
  n3996,
  n3995,
  n3997,
  n3986,
  n3999,
  n3993,
  n3991,
  n3994,
  n3985,
  n4002,
  n3988,
  n4023,
  n4025,
  n4021,
  n4024,
  n4022,
  n4018,
  n4020,
  n4032,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n3772;
  output n3769;
  output n3786;
  output n3787;
  output n3783;
  output n3784;
  output n3792;
  output n3793;
  output n3790;
  output n3989;
  output n4000;
  output n3998;
  output n3987;
  output n3996;
  output n3995;
  output n3997;
  output n3986;
  output n3999;
  output n3993;
  output n3991;
  output n3994;
  output n3985;
  output n4002;
  output n3988;
  output n4023;
  output n4025;
  output n4021;
  output n4024;
  output n4022;
  output n4018;
  output n4020;
  output n4032;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2453;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2482;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2521;
  wire n2522;
  wire n2523;
  wire n2524;
  wire n2525;
  wire n2526;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire n2553;
  wire n2554;
  wire n2555;
  wire n2556;
  wire n2557;
  wire n2558;
  wire n2559;
  wire n2560;
  wire n2561;
  wire n2562;
  wire n2563;
  wire n2564;
  wire n2565;
  wire n2566;
  wire n2567;
  wire n2568;
  wire n2569;
  wire n2570;
  wire n2571;
  wire n2572;
  wire n2573;
  wire n2574;
  wire n2575;
  wire n2576;
  wire n2577;
  wire n2578;
  wire n2579;
  wire n2580;
  wire n2581;
  wire n2582;
  wire n2583;
  wire n2584;
  wire n2585;
  wire n2586;
  wire n2587;
  wire n2588;
  wire n2589;
  wire n2590;
  wire n2591;
  wire n2592;
  wire n2593;
  wire n2594;
  wire n2595;
  wire n2596;
  wire n2597;
  wire n2598;
  wire n2599;
  wire n2600;
  wire n2601;
  wire n2602;
  wire n2603;
  wire n2604;
  wire n2605;
  wire n2606;
  wire n2607;
  wire n2608;
  wire n2609;
  wire n2610;
  wire n2611;
  wire n2612;
  wire n2613;
  wire n2614;
  wire n2615;
  wire n2616;
  wire n2617;
  wire n2618;
  wire n2619;
  wire n2620;
  wire n2621;
  wire n2622;
  wire n2623;
  wire n2624;
  wire n2625;
  wire n2626;
  wire n2627;
  wire n2628;
  wire n2629;
  wire n2630;
  wire n2631;
  wire n2632;
  wire n2633;
  wire n2634;
  wire n2635;
  wire n2636;
  wire n2637;
  wire n2638;
  wire n2639;
  wire n2640;
  wire n2641;
  wire n2642;
  wire n2643;
  wire n2644;
  wire n2645;
  wire n2646;
  wire n2647;
  wire n2648;
  wire n2649;
  wire n2650;
  wire n2651;
  wire n2652;
  wire n2653;
  wire n2654;
  wire n2655;
  wire n2656;
  wire n2657;
  wire n2658;
  wire n2659;
  wire n2660;
  wire n2661;
  wire n2662;
  wire n2663;
  wire n2664;
  wire n2665;
  wire n2666;
  wire n2667;
  wire n2668;
  wire n2669;
  wire n2670;
  wire n2671;
  wire n2672;
  wire n2673;
  wire n2674;
  wire n2675;
  wire n2676;
  wire n2677;
  wire n2678;
  wire n2679;
  wire n2680;
  wire n2681;
  wire n2682;
  wire n2683;
  wire n2684;
  wire n2685;
  wire n2686;
  wire n2687;
  wire n2688;
  wire n2689;
  wire n2690;
  wire n2691;
  wire n2692;
  wire n2693;
  wire n2694;
  wire n2695;
  wire n2696;
  wire n2697;
  wire n2698;
  wire n2699;
  wire n2700;
  wire n2701;
  wire n2702;
  wire n2703;
  wire n2704;
  wire n2705;
  wire n2706;
  wire n2707;
  wire n2708;
  wire n2709;
  wire n2710;
  wire n2711;
  wire n2712;
  wire n2713;
  wire n2714;
  wire n2715;
  wire n2716;
  wire n2717;
  wire n2718;
  wire n2719;
  wire n2720;
  wire n2721;
  wire n2722;
  wire n2723;
  wire n2724;
  wire n2725;
  wire n2726;
  wire n2727;
  wire n2728;
  wire n2729;
  wire n2730;
  wire n2731;
  wire n2732;
  wire n2733;
  wire n2734;
  wire n2735;
  wire n2736;
  wire n2737;
  wire n2738;
  wire n2739;
  wire n2740;
  wire n2741;
  wire n2742;
  wire n2743;
  wire n2744;
  wire n2745;
  wire n2746;
  wire n2747;
  wire n2748;
  wire n2749;
  wire n2750;
  wire n2751;
  wire n2752;
  wire n2753;
  wire n2754;
  wire n2755;
  wire n2756;
  wire n2757;
  wire n2758;
  wire n2759;
  wire n2760;
  wire n2761;
  wire n2762;
  wire n2763;
  wire n2764;
  wire n2765;
  wire n2766;
  wire n2767;
  wire n2768;
  wire n2769;
  wire n2770;
  wire n2771;
  wire n2772;
  wire n2773;
  wire n2774;
  wire n2775;
  wire n2776;
  wire n2777;
  wire n2778;
  wire n2779;
  wire n2780;
  wire n2781;
  wire n2782;
  wire n2783;
  wire n2784;
  wire n2785;
  wire n2786;
  wire n2787;
  wire n2788;
  wire n2789;
  wire n2790;
  wire n2791;
  wire n2792;
  wire n2793;
  wire n2794;
  wire n2795;
  wire n2796;
  wire n2797;
  wire n2798;
  wire n2799;
  wire n2800;
  wire n2801;
  wire n2802;
  wire n2803;
  wire n2804;
  wire n2805;
  wire n2806;
  wire n2807;
  wire n2808;
  wire n2809;
  wire n2810;
  wire n2811;
  wire n2812;
  wire n2813;
  wire n2814;
  wire n2815;
  wire n2816;
  wire n2817;
  wire n2818;
  wire n2819;
  wire n2820;
  wire n2821;
  wire n2822;
  wire n2823;
  wire n2824;
  wire n2825;
  wire n2826;
  wire n2827;
  wire n2828;
  wire n2829;
  wire n2830;
  wire n2831;
  wire n2832;
  wire n2833;
  wire n2834;
  wire n2835;
  wire n2836;
  wire n2837;
  wire n2838;
  wire n2839;
  wire n2840;
  wire n2841;
  wire n2842;
  wire n2843;
  wire n2844;
  wire n2845;
  wire n2846;
  wire n2847;
  wire n2848;
  wire n2849;
  wire n2850;
  wire n2851;
  wire n2852;
  wire n2853;
  wire n2854;
  wire n2855;
  wire n2856;
  wire n2857;
  wire n2858;
  wire n2859;
  wire n2860;
  wire n2861;
  wire n2862;
  wire n2863;
  wire n2864;
  wire n2865;
  wire n2866;
  wire n2867;
  wire n2868;
  wire n2869;
  wire n2870;
  wire n2871;
  wire n2872;
  wire n2873;
  wire n2874;
  wire n2875;
  wire n2876;
  wire n2877;
  wire n2878;
  wire n2879;
  wire n2880;
  wire n2881;
  wire n2882;
  wire n2883;
  wire n2884;
  wire n2885;
  wire n2886;
  wire n2887;
  wire n2888;
  wire n2889;
  wire n2890;
  wire n2891;
  wire n2892;
  wire n2893;
  wire n2894;
  wire n2895;
  wire n2896;
  wire n2897;
  wire n2898;
  wire n2899;
  wire n2900;
  wire n2901;
  wire n2902;
  wire n2903;
  wire n2904;
  wire n2905;
  wire n2906;
  wire n2907;
  wire n2908;
  wire n2909;
  wire n2910;
  wire n2911;
  wire n2912;
  wire n2913;
  wire n2914;
  wire n2915;
  wire n2916;
  wire n2917;
  wire n2918;
  wire n2919;
  wire n2920;
  wire n2921;
  wire n2922;
  wire n2923;
  wire n2924;
  wire n2925;
  wire n2926;
  wire n2927;
  wire n2928;
  wire n2929;
  wire n2930;
  wire n2931;
  wire n2932;
  wire n2933;
  wire n2934;
  wire n2935;
  wire n2936;
  wire n2937;
  wire n2938;
  wire n2939;
  wire n2940;
  wire n2941;
  wire n2942;
  wire n2943;
  wire n2944;
  wire n2945;
  wire n2946;
  wire n2947;
  wire n2948;
  wire n2949;
  wire n2950;
  wire n2951;
  wire n2952;
  wire n2953;
  wire n2954;
  wire n2955;
  wire n2956;
  wire n2957;
  wire n2958;
  wire n2959;
  wire n2960;
  wire n2961;
  wire n2962;
  wire n2963;
  wire n2964;
  wire n2965;
  wire n2966;
  wire n2967;
  wire n2968;
  wire n2969;
  wire n2970;
  wire n2971;
  wire n2972;
  wire n2973;
  wire n2974;
  wire n2975;
  wire n2976;
  wire n2977;
  wire n2978;
  wire n2979;
  wire n2980;
  wire n2981;
  wire n2982;
  wire n2983;
  wire n2984;
  wire n2985;
  wire n2986;
  wire n2987;
  wire n2988;
  wire n2989;
  wire n2990;
  wire n2991;
  wire n2992;
  wire n2993;
  wire n2994;
  wire n2995;
  wire n2996;
  wire n2997;
  wire n2998;
  wire n2999;
  wire n3000;
  wire n3001;
  wire n3002;
  wire n3003;
  wire n3004;
  wire n3005;
  wire n3006;
  wire n3007;
  wire n3008;
  wire n3009;
  wire n3010;
  wire n3011;
  wire n3012;
  wire n3013;
  wire n3014;
  wire n3015;
  wire n3016;
  wire n3017;
  wire n3018;
  wire n3019;
  wire n3020;
  wire n3021;
  wire n3022;
  wire n3023;
  wire n3024;
  wire n3025;
  wire n3026;
  wire n3027;
  wire n3028;
  wire n3029;
  wire n3030;
  wire n3031;
  wire n3032;
  wire n3033;
  wire n3034;
  wire n3035;
  wire n3036;
  wire n3037;
  wire n3038;
  wire n3039;
  wire n3040;
  wire n3041;
  wire n3042;
  wire n3043;
  wire n3044;
  wire n3045;
  wire n3046;
  wire n3047;
  wire n3048;
  wire n3049;
  wire n3050;
  wire n3051;
  wire n3052;
  wire n3053;
  wire n3054;
  wire n3055;
  wire n3056;
  wire n3057;
  wire n3058;
  wire n3059;
  wire n3060;
  wire n3061;
  wire n3062;
  wire n3063;
  wire n3064;
  wire n3065;
  wire n3066;
  wire n3067;
  wire n3068;
  wire n3069;
  wire n3070;
  wire n3071;
  wire n3072;
  wire n3073;
  wire n3074;
  wire n3075;
  wire n3076;
  wire n3077;
  wire n3078;
  wire n3079;
  wire n3080;
  wire n3081;
  wire n3082;
  wire n3083;
  wire n3084;
  wire n3085;
  wire n3086;
  wire n3087;
  wire n3088;
  wire n3089;
  wire n3090;
  wire n3091;
  wire n3092;
  wire n3093;
  wire n3094;
  wire n3095;
  wire n3096;
  wire n3097;
  wire n3098;
  wire n3099;
  wire n3100;
  wire n3101;
  wire n3102;
  wire n3103;
  wire n3104;
  wire n3105;
  wire n3106;
  wire n3107;
  wire n3108;
  wire n3109;
  wire n3110;
  wire n3111;
  wire n3112;
  wire n3113;
  wire n3114;
  wire n3115;
  wire n3116;
  wire n3117;
  wire n3118;
  wire n3119;
  wire n3120;
  wire n3121;
  wire n3122;
  wire n3123;
  wire n3124;
  wire n3125;
  wire n3126;
  wire n3127;
  wire n3128;
  wire n3129;
  wire n3130;
  wire n3131;
  wire n3132;
  wire n3133;
  wire n3134;
  wire n3135;
  wire n3136;
  wire n3137;
  wire n3138;
  wire n3139;
  wire n3140;
  wire n3141;
  wire n3142;
  wire n3143;
  wire n3144;
  wire n3145;
  wire n3146;
  wire n3147;
  wire n3148;
  wire n3149;
  wire n3150;
  wire n3151;
  wire n3152;
  wire n3153;
  wire n3154;
  wire n3155;
  wire n3156;
  wire n3157;
  wire n3158;
  wire n3159;
  wire n3160;
  wire n3161;
  wire n3162;
  wire n3163;
  wire n3164;
  wire n3165;
  wire n3166;
  wire n3167;
  wire n3168;
  wire n3169;
  wire n3170;
  wire n3171;
  wire n3172;
  wire n3173;
  wire n3174;
  wire n3175;
  wire n3176;
  wire n3177;
  wire n3178;
  wire n3179;
  wire n3180;
  wire n3181;
  wire n3182;
  wire n3183;
  wire n3184;
  wire n3185;
  wire n3186;
  wire n3187;
  wire n3188;
  wire n3189;
  wire n3190;
  wire n3191;
  wire n3192;
  wire n3193;
  wire n3194;
  wire n3195;
  wire n3196;
  wire n3197;
  wire n3198;
  wire n3199;
  wire n3200;
  wire n3201;
  wire n3202;
  wire n3203;
  wire n3204;
  wire n3205;
  wire n3206;
  wire n3207;
  wire n3208;
  wire n3209;
  wire n3210;
  wire n3211;
  wire n3212;
  wire n3213;
  wire n3214;
  wire n3215;
  wire n3216;
  wire n3217;
  wire n3218;
  wire n3219;
  wire n3220;
  wire n3221;
  wire n3222;
  wire n3223;
  wire n3224;
  wire n3225;
  wire n3226;
  wire n3227;
  wire n3228;
  wire n3229;
  wire n3230;
  wire n3231;
  wire n3232;
  wire n3233;
  wire n3234;
  wire n3235;
  wire n3236;
  wire n3237;
  wire n3238;
  wire n3239;
  wire n3240;
  wire n3241;
  wire n3242;
  wire n3243;
  wire n3244;
  wire n3245;
  wire n3246;
  wire n3247;
  wire n3248;
  wire n3249;
  wire n3250;
  wire n3251;
  wire n3252;
  wire n3253;
  wire n3254;
  wire n3255;
  wire n3256;
  wire n3257;
  wire n3258;
  wire n3259;
  wire n3260;
  wire n3261;
  wire n3262;
  wire n3263;
  wire n3264;
  wire n3265;
  wire n3266;
  wire n3267;
  wire n3268;
  wire n3269;
  wire n3270;
  wire n3271;
  wire n3272;
  wire n3273;
  wire n3274;
  wire n3275;
  wire n3276;
  wire n3277;
  wire n3278;
  wire n3279;
  wire n3280;
  wire n3281;
  wire n3282;
  wire n3283;
  wire n3284;
  wire n3285;
  wire n3286;
  wire n3287;
  wire n3288;
  wire n3289;
  wire n3290;
  wire n3291;
  wire n3292;
  wire n3293;
  wire n3294;
  wire n3295;
  wire n3296;
  wire n3297;
  wire n3298;
  wire n3299;
  wire n3300;
  wire n3301;
  wire n3302;
  wire n3303;
  wire n3304;
  wire n3305;
  wire n3306;
  wire n3307;
  wire n3308;
  wire n3309;
  wire n3310;
  wire n3311;
  wire n3312;
  wire n3313;
  wire n3314;
  wire n3315;
  wire n3316;
  wire n3317;
  wire n3318;
  wire n3319;
  wire n3320;
  wire n3321;
  wire n3322;
  wire n3323;
  wire n3324;
  wire n3325;
  wire n3326;
  wire n3327;
  wire n3328;
  wire n3329;
  wire n3330;
  wire n3331;
  wire n3332;
  wire n3333;
  wire n3334;
  wire n3335;
  wire n3336;
  wire n3337;
  wire n3338;
  wire n3339;
  wire n3340;
  wire n3341;
  wire n3342;
  wire n3343;
  wire n3344;
  wire n3345;
  wire n3346;
  wire n3347;
  wire n3348;
  wire n3349;
  wire n3350;
  wire n3351;
  wire n3352;
  wire n3353;
  wire n3354;
  wire n3355;
  wire n3356;
  wire n3357;
  wire n3358;
  wire n3359;
  wire n3360;
  wire n3361;
  wire n3362;
  wire n3363;
  wire n3364;
  wire n3365;
  wire n3366;
  wire n3367;
  wire n3368;
  wire n3369;
  wire n3370;
  wire n3371;
  wire n3372;
  wire n3373;
  wire n3374;
  wire n3375;
  wire n3376;
  wire n3377;
  wire n3378;
  wire n3379;
  wire n3380;
  wire n3381;
  wire n3382;
  wire n3383;
  wire n3384;
  wire n3385;
  wire n3386;
  wire n3387;
  wire n3388;
  wire n3389;
  wire n3390;
  wire n3391;
  wire n3392;
  wire n3393;
  wire n3394;
  wire n3395;
  wire n3396;
  wire n3397;
  wire n3398;
  wire n3399;
  wire n3400;
  wire n3401;
  wire n3402;
  wire n3403;
  wire n3404;
  wire n3405;
  wire n3406;
  wire n3407;
  wire n3408;
  wire n3409;
  wire n3410;
  wire n3411;
  wire n3412;
  wire n3413;
  wire n3414;
  wire n3415;
  wire n3416;
  wire n3417;
  wire n3418;
  wire n3419;
  wire n3420;
  wire n3421;
  wire n3422;
  wire n3423;
  wire n3424;
  wire n3425;
  wire n3426;
  wire n3427;
  wire n3428;
  wire n3429;
  wire n3430;
  wire n3431;
  wire n3432;
  wire n3433;
  wire n3434;
  wire n3435;
  wire n3436;
  wire n3437;
  wire n3438;
  wire n3439;
  wire n3440;
  wire n3441;
  wire n3442;
  wire n3443;
  wire n3444;
  wire n3445;
  wire n3446;
  wire n3447;
  wire n3448;
  wire n3449;
  wire n3450;
  wire n3451;
  wire n3452;
  wire n3453;
  wire n3454;
  wire n3455;
  wire n3456;
  wire n3457;
  wire n3458;
  wire n3459;
  wire n3460;
  wire n3461;
  wire n3462;
  wire n3463;
  wire n3464;
  wire n3465;
  wire n3466;
  wire n3467;
  wire n3468;
  wire n3469;
  wire n3470;
  wire n3471;
  wire n3472;
  wire n3473;
  wire n3474;
  wire n3475;
  wire n3476;
  wire n3477;
  wire n3478;
  wire n3479;
  wire n3480;
  wire n3481;
  wire n3482;
  wire n3483;
  wire n3484;
  wire n3485;
  wire n3486;
  wire n3487;
  wire n3488;
  wire n3489;
  wire n3490;
  wire n3491;
  wire n3492;
  wire n3493;
  wire n3494;
  wire n3495;
  wire n3496;
  wire n3497;
  wire n3498;
  wire n3499;
  wire n3500;
  wire n3501;
  wire n3502;
  wire n3503;
  wire n3504;
  wire n3505;
  wire n3506;
  wire n3507;
  wire n3508;
  wire n3509;
  wire n3510;
  wire n3511;
  wire n3512;
  wire n3513;
  wire n3514;
  wire n3515;
  wire n3516;
  wire n3517;
  wire n3518;
  wire n3519;
  wire n3520;
  wire n3521;
  wire n3522;
  wire n3523;
  wire n3524;
  wire n3525;
  wire n3526;
  wire n3527;
  wire n3528;
  wire n3529;
  wire n3530;
  wire n3531;
  wire n3532;
  wire n3533;
  wire n3534;
  wire n3535;
  wire n3536;
  wire n3537;
  wire n3538;
  wire n3539;
  wire n3540;
  wire n3541;
  wire n3542;
  wire n3543;
  wire n3544;
  wire n3545;
  wire n3546;
  wire n3547;
  wire n3548;
  wire n3549;
  wire n3550;
  wire n3551;
  wire n3552;
  wire n3553;
  wire n3554;
  wire n3555;
  wire n3556;
  wire n3557;
  wire n3558;
  wire n3559;
  wire n3560;
  wire n3561;
  wire n3562;
  wire n3563;
  wire n3564;
  wire n3565;
  wire n3566;
  wire n3567;
  wire n3568;
  wire n3569;
  wire n3570;
  wire n3571;
  wire n3572;
  wire n3573;
  wire n3574;
  wire n3575;
  wire n3576;
  wire n3577;
  wire n3578;
  wire n3579;
  wire n3580;
  wire n3581;
  wire n3582;
  wire n3583;
  wire n3584;
  wire n3585;
  wire n3586;
  wire n3587;
  wire n3588;
  wire n3589;
  wire n3590;
  wire n3591;
  wire n3592;
  wire n3593;
  wire n3594;
  wire n3595;
  wire n3596;
  wire n3597;
  wire n3598;
  wire n3599;
  wire n3600;
  wire n3601;
  wire n3602;
  wire n3603;
  wire n3604;
  wire n3605;
  wire n3606;
  wire n3607;
  wire n3608;
  wire n3609;
  wire n3610;
  wire n3611;
  wire n3612;
  wire n3613;
  wire n3614;
  wire n3615;
  wire n3616;
  wire n3617;
  wire n3618;
  wire n3619;
  wire n3620;
  wire n3621;
  wire n3622;
  wire n3623;
  wire n3624;
  wire n3625;
  wire n3626;
  wire n3627;
  wire n3628;
  wire n3629;
  wire n3630;
  wire n3631;
  wire n3632;
  wire n3633;
  wire n3634;
  wire n3635;
  wire n3636;
  wire n3637;
  wire n3638;
  wire n3639;
  wire n3640;
  wire n3641;
  wire n3642;
  wire n3643;
  wire n3644;
  wire n3645;
  wire n3646;
  wire n3647;
  wire n3648;
  wire n3649;
  wire n3650;
  wire n3651;
  wire n3652;
  wire n3653;
  wire n3654;
  wire n3655;
  wire n3656;
  wire n3657;
  wire n3658;
  wire n3659;
  wire n3660;
  wire n3661;
  wire n3662;
  wire n3663;
  wire n3664;
  wire n3665;
  wire n3666;
  wire n3667;
  wire n3668;
  wire n3669;
  wire n3670;
  wire n3671;
  wire n3672;
  wire n3673;
  wire n3674;
  wire n3675;
  wire n3676;
  wire n3677;
  wire n3678;
  wire n3679;
  wire n3680;
  wire n3681;
  wire n3682;
  wire n3683;
  wire n3684;
  wire n3685;
  wire n3686;
  wire n3687;
  wire n3688;
  wire n3689;
  wire n3690;
  wire n3691;
  wire n3692;
  wire n3693;
  wire n3694;
  wire n3695;
  wire n3696;
  wire n3697;
  wire n3698;
  wire n3699;
  wire n3700;
  wire n3701;
  wire n3702;
  wire n3703;
  wire n3704;
  wire n3705;
  wire n3706;
  wire n3707;
  wire n3708;
  wire n3709;
  wire n3710;
  wire n3711;
  wire n3712;
  wire n3713;
  wire n3714;
  wire n3715;
  wire n3716;
  wire n3717;
  wire n3718;
  wire n3719;
  wire n3720;
  wire n3721;
  wire n3722;
  wire n3723;
  wire n3724;
  wire n3725;
  wire n3726;
  wire n3727;
  wire n3728;
  wire n3729;
  wire n3730;
  wire n3731;
  wire n3732;
  wire n3733;
  wire n3734;
  wire n3735;
  wire n3736;
  wire n3737;
  wire n3738;
  wire n3739;
  wire n3740;
  wire n3741;
  wire n3742;
  wire n3743;
  wire n3744;
  wire n3745;
  wire n3746;
  wire n3747;
  wire n3748;
  wire n3749;
  wire n3750;
  wire n3751;
  wire n3752;
  wire n3753;
  wire n3754;
  wire n3755;
  wire n3756;
  wire n3757;
  wire n3758;
  wire n3759;
  wire n3760;
  wire n3761;
  wire n3762;
  wire n3763;
  wire n3764;
  wire n3765;
  wire n3766;
  wire n3767;
  wire n3768;
  wire n3770;
  wire n3771;
  wire n3773;
  wire n3774;
  wire n3775;
  wire n3776;
  wire n3777;
  wire n3778;
  wire n3779;
  wire n3780;
  wire n3781;
  wire n3782;
  wire n3785;
  wire n3788;
  wire n3789;
  wire n3791;
  wire n3794;
  wire n3795;
  wire n3796;
  wire n3797;
  wire n3798;
  wire n3799;
  wire n3800;
  wire n3801;
  wire n3802;
  wire n3803;
  wire n3804;
  wire n3805;
  wire n3806;
  wire n3807;
  wire n3808;
  wire n3809;
  wire n3810;
  wire n3811;
  wire n3812;
  wire n3813;
  wire n3814;
  wire n3815;
  wire n3816;
  wire n3817;
  wire n3818;
  wire n3819;
  wire n3820;
  wire n3821;
  wire n3822;
  wire n3823;
  wire n3824;
  wire n3825;
  wire n3826;
  wire n3827;
  wire n3828;
  wire n3829;
  wire n3830;
  wire n3831;
  wire n3832;
  wire n3833;
  wire n3834;
  wire n3835;
  wire n3836;
  wire n3837;
  wire n3838;
  wire n3839;
  wire n3840;
  wire n3841;
  wire n3842;
  wire n3843;
  wire n3844;
  wire n3845;
  wire n3846;
  wire n3847;
  wire n3848;
  wire n3849;
  wire n3850;
  wire n3851;
  wire n3852;
  wire n3853;
  wire n3854;
  wire n3855;
  wire n3856;
  wire n3857;
  wire n3858;
  wire n3859;
  wire n3860;
  wire n3861;
  wire n3862;
  wire n3863;
  wire n3864;
  wire n3865;
  wire n3866;
  wire n3867;
  wire n3868;
  wire n3869;
  wire n3870;
  wire n3871;
  wire n3872;
  wire n3873;
  wire n3874;
  wire n3875;
  wire n3876;
  wire n3877;
  wire n3878;
  wire n3879;
  wire n3880;
  wire n3881;
  wire n3882;
  wire n3883;
  wire n3884;
  wire n3885;
  wire n3886;
  wire n3887;
  wire n3888;
  wire n3889;
  wire n3890;
  wire n3891;
  wire n3892;
  wire n3893;
  wire n3894;
  wire n3895;
  wire n3896;
  wire n3897;
  wire n3898;
  wire n3899;
  wire n3900;
  wire n3901;
  wire n3902;
  wire n3903;
  wire n3904;
  wire n3905;
  wire n3906;
  wire n3907;
  wire n3908;
  wire n3909;
  wire n3910;
  wire n3911;
  wire n3912;
  wire n3913;
  wire n3914;
  wire n3915;
  wire n3916;
  wire n3917;
  wire n3918;
  wire n3919;
  wire n3920;
  wire n3921;
  wire n3922;
  wire n3923;
  wire n3924;
  wire n3925;
  wire n3926;
  wire n3927;
  wire n3928;
  wire n3929;
  wire n3930;
  wire n3931;
  wire n3932;
  wire n3933;
  wire n3934;
  wire n3935;
  wire n3936;
  wire n3937;
  wire n3938;
  wire n3939;
  wire n3940;
  wire n3941;
  wire n3942;
  wire n3943;
  wire n3944;
  wire n3945;
  wire n3946;
  wire n3947;
  wire n3948;
  wire n3949;
  wire n3950;
  wire n3951;
  wire n3952;
  wire n3953;
  wire n3954;
  wire n3955;
  wire n3956;
  wire n3957;
  wire n3958;
  wire n3959;
  wire n3960;
  wire n3961;
  wire n3962;
  wire n3963;
  wire n3964;
  wire n3965;
  wire n3966;
  wire n3967;
  wire n3968;
  wire n3969;
  wire n3970;
  wire n3971;
  wire n3972;
  wire n3973;
  wire n3974;
  wire n3975;
  wire n3976;
  wire n3977;
  wire n3978;
  wire n3979;
  wire n3980;
  wire n3981;
  wire n3982;
  wire n3983;
  wire n3984;
  wire n3990;
  wire n3992;
  wire n4001;
  wire n4003;
  wire n4004;
  wire n4005;
  wire n4006;
  wire n4007;
  wire n4008;
  wire n4009;
  wire n4010;
  wire n4011;
  wire n4012;
  wire n4013;
  wire n4014;
  wire n4015;
  wire n4016;
  wire n4017;
  wire n4019;
  wire n4026;
  wire n4027;
  wire n4028;
  wire n4029;
  wire n4030;
  wire n4031;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyNOTWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;
  wire KeyNOTWire_0_63;

  not
  g0
  (
    n145,
    n28
  );


  not
  g1
  (
    n56,
    n19
  );


  buf
  g2
  (
    n152,
    n21
  );


  buf
  g3
  (
    n114,
    n24
  );


  not
  g4
  (
    n99,
    n23
  );


  not
  g5
  (
    n50,
    n24
  );


  not
  g6
  (
    n143,
    n32
  );


  buf
  g7
  (
    n85,
    n17
  );


  not
  g8
  (
    n103,
    n7
  );


  not
  g9
  (
    n151,
    n27
  );


  buf
  g10
  (
    n111,
    n2
  );


  buf
  g11
  (
    n157,
    n10
  );


  buf
  g12
  (
    n130,
    n26
  );


  not
  g13
  (
    n106,
    n6
  );


  not
  g14
  (
    n34,
    n28
  );


  not
  g15
  (
    n69,
    n12
  );


  buf
  g16
  (
    n41,
    n20
  );


  not
  g17
  (
    n107,
    n32
  );


  buf
  g18
  (
    n135,
    n23
  );


  buf
  g19
  (
    n46,
    n8
  );


  buf
  g20
  (
    n131,
    n2
  );


  buf
  g21
  (
    n73,
    n14
  );


  buf
  g22
  (
    n90,
    n11
  );


  buf
  g23
  (
    n77,
    n18
  );


  buf
  g24
  (
    n39,
    n19
  );


  buf
  g25
  (
    n160,
    n2
  );


  not
  g26
  (
    n96,
    n26
  );


  not
  g27
  (
    n52,
    n4
  );


  buf
  g28
  (
    n53,
    n14
  );


  not
  g29
  (
    n89,
    n32
  );


  buf
  g30
  (
    n158,
    n31
  );


  not
  g31
  (
    n81,
    n17
  );


  buf
  g32
  (
    n139,
    n16
  );


  not
  g33
  (
    n51,
    n29
  );


  not
  g34
  (
    n155,
    n31
  );


  not
  g35
  (
    n154,
    n29
  );


  not
  g36
  (
    n86,
    n4
  );


  buf
  g37
  (
    n66,
    n11
  );


  buf
  g38
  (
    n55,
    n17
  );


  not
  g39
  (
    n118,
    n8
  );


  not
  g40
  (
    n92,
    n1
  );


  buf
  g41
  (
    n138,
    n15
  );


  buf
  g42
  (
    n100,
    n4
  );


  not
  g43
  (
    n110,
    n32
  );


  not
  g44
  (
    n97,
    n9
  );


  not
  g45
  (
    n95,
    n1
  );


  not
  g46
  (
    n68,
    n28
  );


  not
  g47
  (
    n128,
    n10
  );


  not
  g48
  (
    n105,
    n6
  );


  buf
  g49
  (
    n43,
    n22
  );


  not
  g50
  (
    n104,
    n23
  );


  not
  g51
  (
    n36,
    n20
  );


  not
  g52
  (
    n59,
    n22
  );


  buf
  g53
  (
    n91,
    n24
  );


  not
  g54
  (
    n148,
    n8
  );


  not
  g55
  (
    n122,
    n9
  );


  not
  g56
  (
    n146,
    n29
  );


  not
  g57
  (
    n74,
    n16
  );


  not
  g58
  (
    n108,
    n3
  );


  buf
  g59
  (
    n102,
    n16
  );


  buf
  g60
  (
    n58,
    n12
  );


  buf
  g61
  (
    n127,
    n20
  );


  buf
  g62
  (
    n40,
    n9
  );


  not
  g63
  (
    n48,
    n27
  );


  buf
  g64
  (
    n75,
    n15
  );


  not
  g65
  (
    KeyWire_0_11,
    n20
  );


  buf
  g66
  (
    n149,
    n21
  );


  not
  g67
  (
    n144,
    n13
  );


  buf
  g68
  (
    n125,
    n18
  );


  buf
  g69
  (
    n136,
    n12
  );


  not
  g70
  (
    n83,
    n25
  );


  buf
  g71
  (
    n93,
    n13
  );


  buf
  g72
  (
    n129,
    n18
  );


  buf
  g73
  (
    n113,
    n28
  );


  buf
  g74
  (
    n120,
    n3
  );


  not
  g75
  (
    n38,
    n30
  );


  not
  g76
  (
    n101,
    n7
  );


  buf
  g77
  (
    n159,
    n11
  );


  not
  g78
  (
    n79,
    n15
  );


  not
  g79
  (
    n112,
    n6
  );


  buf
  g80
  (
    n72,
    n14
  );


  not
  g81
  (
    n132,
    n2
  );


  buf
  g82
  (
    n49,
    n12
  );


  not
  g83
  (
    n88,
    n27
  );


  not
  g84
  (
    KeyWire_0_56,
    n23
  );


  not
  g85
  (
    n78,
    n10
  );


  not
  g86
  (
    n67,
    n21
  );


  buf
  g87
  (
    n150,
    n7
  );


  not
  g88
  (
    n115,
    n19
  );


  buf
  g89
  (
    n153,
    n27
  );


  buf
  g90
  (
    n147,
    n11
  );


  buf
  g91
  (
    n71,
    n17
  );


  not
  g92
  (
    n44,
    n31
  );


  buf
  g93
  (
    n80,
    n25
  );


  not
  g94
  (
    n121,
    n9
  );


  not
  g95
  (
    n134,
    n3
  );


  not
  g96
  (
    n62,
    n30
  );


  not
  g97
  (
    n119,
    n22
  );


  buf
  g98
  (
    n64,
    n24
  );


  buf
  g99
  (
    n82,
    n15
  );


  not
  g100
  (
    n116,
    n30
  );


  buf
  g101
  (
    n109,
    n1
  );


  not
  g102
  (
    n65,
    n19
  );


  buf
  g103
  (
    n142,
    n3
  );


  not
  g104
  (
    n61,
    n29
  );


  not
  g105
  (
    n126,
    n13
  );


  buf
  g106
  (
    n57,
    n1
  );


  buf
  g107
  (
    n47,
    n16
  );


  not
  g108
  (
    n137,
    n21
  );


  not
  g109
  (
    n45,
    n18
  );


  not
  g110
  (
    n156,
    n14
  );


  buf
  g111
  (
    n60,
    n5
  );


  not
  g112
  (
    n54,
    n26
  );


  buf
  g113
  (
    n141,
    n8
  );


  buf
  g114
  (
    n94,
    n7
  );


  not
  g115
  (
    KeyWire_0_8,
    n6
  );


  buf
  g116
  (
    n33,
    n4
  );


  not
  g117
  (
    n84,
    n5
  );


  buf
  g118
  (
    n124,
    n13
  );


  buf
  g119
  (
    n117,
    n30
  );


  buf
  g120
  (
    n87,
    n10
  );


  buf
  g121
  (
    n140,
    n22
  );


  not
  g122
  (
    n123,
    n5
  );


  buf
  g123
  (
    n70,
    n31
  );


  not
  g124
  (
    n42,
    n25
  );


  not
  g125
  (
    n98,
    n26
  );


  not
  g126
  (
    n37,
    n25
  );


  buf
  g127
  (
    n63,
    n5
  );


  not
  g128
  (
    n493,
    n127
  );


  not
  g129
  (
    n174,
    n55
  );


  not
  g130
  (
    n560,
    n138
  );


  not
  g131
  (
    n639,
    n40
  );


  buf
  g132
  (
    n229,
    n76
  );


  not
  g133
  (
    n491,
    n69
  );


  buf
  g134
  (
    n531,
    n143
  );


  buf
  g135
  (
    n330,
    n61
  );


  not
  g136
  (
    n588,
    n64
  );


  buf
  g137
  (
    n280,
    n70
  );


  not
  g138
  (
    n234,
    n58
  );


  not
  g139
  (
    n420,
    n79
  );


  not
  g140
  (
    n215,
    n86
  );


  buf
  g141
  (
    n323,
    n33
  );


  buf
  g142
  (
    n545,
    n114
  );


  not
  g143
  (
    n263,
    n123
  );


  not
  g144
  (
    n395,
    n39
  );


  not
  g145
  (
    n437,
    n79
  );


  buf
  g146
  (
    n208,
    n141
  );


  buf
  g147
  (
    n196,
    n150
  );


  not
  g148
  (
    n412,
    n97
  );


  buf
  g149
  (
    n165,
    n100
  );


  buf
  g150
  (
    n222,
    n51
  );


  buf
  g151
  (
    n522,
    n118
  );


  buf
  g152
  (
    n385,
    n160
  );


  not
  g153
  (
    n613,
    n126
  );


  not
  g154
  (
    n163,
    n134
  );


  not
  g155
  (
    n576,
    n95
  );


  not
  g156
  (
    n509,
    n80
  );


  buf
  g157
  (
    n529,
    n127
  );


  not
  g158
  (
    n181,
    n72
  );


  not
  g159
  (
    n466,
    n55
  );


  not
  g160
  (
    n518,
    n86
  );


  not
  g161
  (
    n306,
    n124
  );


  not
  g162
  (
    n625,
    n126
  );


  buf
  g163
  (
    n177,
    n80
  );


  buf
  g164
  (
    n533,
    n107
  );


  buf
  g165
  (
    n379,
    n53
  );


  buf
  g166
  (
    n450,
    n40
  );


  buf
  g167
  (
    n464,
    n71
  );


  not
  g168
  (
    n328,
    n136
  );


  buf
  g169
  (
    n508,
    n152
  );


  not
  g170
  (
    KeyWire_0_13,
    n112
  );


  not
  g171
  (
    n349,
    n153
  );


  buf
  g172
  (
    n394,
    n104
  );


  buf
  g173
  (
    n569,
    n119
  );


  buf
  g174
  (
    n305,
    n131
  );


  not
  g175
  (
    n340,
    n82
  );


  buf
  g176
  (
    n178,
    n154
  );


  buf
  g177
  (
    n352,
    n119
  );


  buf
  g178
  (
    n503,
    n126
  );


  not
  g179
  (
    n247,
    n99
  );


  buf
  g180
  (
    n188,
    n156
  );


  buf
  g181
  (
    n570,
    n130
  );


  buf
  g182
  (
    n510,
    n92
  );


  not
  g183
  (
    n413,
    n68
  );


  not
  g184
  (
    n392,
    n108
  );


  not
  g185
  (
    n374,
    n118
  );


  not
  g186
  (
    n337,
    n73
  );


  buf
  g187
  (
    n494,
    n105
  );


  buf
  g188
  (
    n512,
    n151
  );


  not
  g189
  (
    n598,
    n46
  );


  not
  g190
  (
    n168,
    n78
  );


  not
  g191
  (
    n276,
    n140
  );


  not
  g192
  (
    n206,
    n92
  );


  not
  g193
  (
    n281,
    n51
  );


  buf
  g194
  (
    n219,
    n81
  );


  buf
  g195
  (
    n517,
    n45
  );


  not
  g196
  (
    n182,
    n44
  );


  not
  g197
  (
    n389,
    n70
  );


  not
  g198
  (
    n393,
    n102
  );


  buf
  g199
  (
    n442,
    n44
  );


  buf
  g200
  (
    n422,
    n104
  );


  buf
  g201
  (
    n506,
    n37
  );


  not
  g202
  (
    n478,
    n107
  );


  buf
  g203
  (
    n479,
    n93
  );


  buf
  g204
  (
    n590,
    n66
  );


  not
  g205
  (
    n405,
    n56
  );


  not
  g206
  (
    n254,
    n54
  );


  buf
  g207
  (
    n179,
    n58
  );


  not
  g208
  (
    n652,
    n42
  );


  not
  g209
  (
    n628,
    n69
  );


  buf
  g210
  (
    n198,
    n145
  );


  not
  g211
  (
    n513,
    n44
  );


  buf
  g212
  (
    n191,
    n52
  );


  buf
  g213
  (
    n398,
    n43
  );


  not
  g214
  (
    n217,
    n112
  );


  not
  g215
  (
    n342,
    n122
  );


  not
  g216
  (
    n551,
    n111
  );


  buf
  g217
  (
    n425,
    n103
  );


  buf
  g218
  (
    n614,
    n77
  );


  not
  g219
  (
    n262,
    n102
  );


  buf
  g220
  (
    n242,
    n96
  );


  buf
  g221
  (
    n583,
    n34
  );


  buf
  g222
  (
    n331,
    n128
  );


  buf
  g223
  (
    n482,
    n52
  );


  buf
  g224
  (
    n492,
    n89
  );


  buf
  g225
  (
    n444,
    n153
  );


  buf
  g226
  (
    n472,
    n157
  );


  not
  g227
  (
    n351,
    n77
  );


  not
  g228
  (
    n357,
    n90
  );


  buf
  g229
  (
    n654,
    n159
  );


  not
  g230
  (
    n212,
    n159
  );


  buf
  g231
  (
    n363,
    n123
  );


  not
  g232
  (
    n429,
    n57
  );


  not
  g233
  (
    n456,
    n93
  );


  not
  g234
  (
    n205,
    n112
  );


  not
  g235
  (
    n186,
    n108
  );


  not
  g236
  (
    n660,
    n139
  );


  buf
  g237
  (
    n621,
    n78
  );


  buf
  g238
  (
    n426,
    n35
  );


  buf
  g239
  (
    n346,
    n142
  );


  not
  g240
  (
    n431,
    n81
  );


  not
  g241
  (
    n534,
    n88
  );


  not
  g242
  (
    n582,
    n153
  );


  buf
  g243
  (
    n228,
    n140
  );


  not
  g244
  (
    n599,
    n105
  );


  not
  g245
  (
    n185,
    n57
  );


  buf
  g246
  (
    n428,
    n150
  );


  not
  g247
  (
    n348,
    n115
  );


  not
  g248
  (
    n370,
    n140
  );


  not
  g249
  (
    n383,
    n124
  );


  not
  g250
  (
    n611,
    n135
  );


  not
  g251
  (
    n375,
    n146
  );


  buf
  g252
  (
    n221,
    n71
  );


  not
  g253
  (
    n463,
    n137
  );


  buf
  g254
  (
    n310,
    n149
  );


  buf
  g255
  (
    n287,
    n83
  );


  buf
  g256
  (
    n211,
    n145
  );


  buf
  g257
  (
    KeyWire_0_22,
    n63
  );


  not
  g258
  (
    n246,
    n144
  );


  buf
  g259
  (
    n487,
    n41
  );


  not
  g260
  (
    n344,
    n96
  );


  buf
  g261
  (
    n194,
    n123
  );


  buf
  g262
  (
    n409,
    n106
  );


  buf
  g263
  (
    n244,
    n122
  );


  buf
  g264
  (
    n581,
    n105
  );


  buf
  g265
  (
    n270,
    n66
  );


  buf
  g266
  (
    n641,
    n135
  );


  not
  g267
  (
    n334,
    n92
  );


  buf
  g268
  (
    n557,
    n103
  );


  not
  g269
  (
    n433,
    n50
  );


  buf
  g270
  (
    n336,
    n88
  );


  buf
  g271
  (
    n252,
    n35
  );


  not
  g272
  (
    n586,
    n85
  );


  buf
  g273
  (
    n476,
    n156
  );


  buf
  g274
  (
    n171,
    n128
  );


  not
  g275
  (
    n397,
    n144
  );


  buf
  g276
  (
    n249,
    n141
  );


  buf
  g277
  (
    n238,
    n90
  );


  not
  g278
  (
    n258,
    n125
  );


  buf
  g279
  (
    n519,
    n61
  );


  buf
  g280
  (
    n668,
    n121
  );


  not
  g281
  (
    n653,
    n155
  );


  not
  g282
  (
    n218,
    n100
  );


  not
  g283
  (
    n274,
    n153
  );


  buf
  g284
  (
    n484,
    n131
  );


  buf
  g285
  (
    n233,
    n144
  );


  buf
  g286
  (
    n189,
    n83
  );


  buf
  g287
  (
    n364,
    n129
  );


  buf
  g288
  (
    n322,
    n85
  );


  not
  g289
  (
    n631,
    n118
  );


  not
  g290
  (
    n587,
    n36
  );


  buf
  g291
  (
    n605,
    n98
  );


  not
  g292
  (
    n530,
    n76
  );


  buf
  g293
  (
    n571,
    n136
  );


  not
  g294
  (
    n485,
    n158
  );


  not
  g295
  (
    n255,
    n117
  );


  buf
  g296
  (
    KeyWire_0_21,
    n70
  );


  buf
  g297
  (
    n457,
    n94
  );


  not
  g298
  (
    n608,
    n67
  );


  buf
  g299
  (
    n407,
    n150
  );


  not
  g300
  (
    n269,
    n107
  );


  buf
  g301
  (
    n319,
    n109
  );


  buf
  g302
  (
    n293,
    n110
  );


  not
  g303
  (
    n547,
    n38
  );


  buf
  g304
  (
    n486,
    n143
  );


  buf
  g305
  (
    n176,
    n70
  );


  not
  g306
  (
    n289,
    n125
  );


  buf
  g307
  (
    n642,
    n48
  );


  not
  g308
  (
    n505,
    n83
  );


  not
  g309
  (
    n200,
    n57
  );


  buf
  g310
  (
    n523,
    n69
  );


  not
  g311
  (
    n559,
    n62
  );


  buf
  g312
  (
    n589,
    n87
  );


  not
  g313
  (
    n562,
    n137
  );


  buf
  g314
  (
    n376,
    n146
  );


  buf
  g315
  (
    n489,
    n73
  );


  not
  g316
  (
    n520,
    n102
  );


  not
  g317
  (
    n665,
    n140
  );


  buf
  g318
  (
    n175,
    n102
  );


  buf
  g319
  (
    n532,
    n47
  );


  not
  g320
  (
    n295,
    n49
  );


  not
  g321
  (
    n514,
    n65
  );


  not
  g322
  (
    n292,
    n127
  );


  not
  g323
  (
    n169,
    n72
  );


  buf
  g324
  (
    n419,
    n76
  );


  buf
  g325
  (
    n193,
    n34
  );


  buf
  g326
  (
    n646,
    n122
  );


  not
  g327
  (
    n459,
    n65
  );


  buf
  g328
  (
    n256,
    n67
  );


  not
  g329
  (
    n602,
    n37
  );


  buf
  g330
  (
    n648,
    n111
  );


  buf
  g331
  (
    n481,
    n91
  );


  not
  g332
  (
    n378,
    n95
  );


  not
  g333
  (
    n390,
    n50
  );


  not
  g334
  (
    n417,
    n146
  );


  buf
  g335
  (
    n273,
    n157
  );


  buf
  g336
  (
    n438,
    n100
  );


  not
  g337
  (
    n275,
    n71
  );


  not
  g338
  (
    n657,
    n154
  );


  buf
  g339
  (
    n316,
    n152
  );


  buf
  g340
  (
    n544,
    n135
  );


  buf
  g341
  (
    n307,
    n132
  );


  not
  g342
  (
    n561,
    n146
  );


  buf
  g343
  (
    n638,
    n61
  );


  not
  g344
  (
    n241,
    n101
  );


  buf
  g345
  (
    n345,
    n101
  );


  not
  g346
  (
    n488,
    n99
  );


  buf
  g347
  (
    n315,
    n36
  );


  buf
  g348
  (
    n377,
    n73
  );


  buf
  g349
  (
    KeyWire_0_19,
    n120
  );


  buf
  g350
  (
    n593,
    n48
  );


  not
  g351
  (
    n524,
    n56
  );


  not
  g352
  (
    n272,
    n64
  );


  not
  g353
  (
    n591,
    n111
  );


  not
  g354
  (
    n670,
    n59
  );


  not
  g355
  (
    n525,
    n119
  );


  not
  g356
  (
    n257,
    n141
  );


  buf
  g357
  (
    n286,
    n60
  );


  buf
  g358
  (
    n396,
    n115
  );


  buf
  g359
  (
    n332,
    n41
  );


  not
  g360
  (
    n502,
    n117
  );


  not
  g361
  (
    n616,
    n122
  );


  buf
  g362
  (
    n304,
    n109
  );


  buf
  g363
  (
    n515,
    n106
  );


  buf
  g364
  (
    n403,
    n87
  );


  not
  g365
  (
    n355,
    n66
  );


  not
  g366
  (
    n659,
    n115
  );


  buf
  g367
  (
    n308,
    n117
  );


  buf
  g368
  (
    n265,
    n55
  );


  not
  g369
  (
    n354,
    n154
  );


  not
  g370
  (
    n404,
    n95
  );


  not
  g371
  (
    n656,
    n56
  );


  not
  g372
  (
    n297,
    n45
  );


  not
  g373
  (
    n227,
    n84
  );


  buf
  g374
  (
    n384,
    n131
  );


  buf
  g375
  (
    n239,
    n42
  );


  not
  g376
  (
    n435,
    n103
  );


  buf
  g377
  (
    n620,
    n138
  );


  buf
  g378
  (
    n264,
    n46
  );


  buf
  g379
  (
    n573,
    n128
  );


  buf
  g380
  (
    n356,
    n99
  );


  not
  g381
  (
    n467,
    n128
  );


  buf
  g382
  (
    n285,
    n38
  );


  buf
  g383
  (
    n418,
    n80
  );


  buf
  g384
  (
    n387,
    n110
  );


  not
  g385
  (
    n296,
    n65
  );


  not
  g386
  (
    n359,
    n130
  );


  buf
  g387
  (
    n578,
    n120
  );


  buf
  g388
  (
    n458,
    n152
  );


  not
  g389
  (
    n555,
    n125
  );


  not
  g390
  (
    n298,
    n82
  );


  buf
  g391
  (
    n441,
    n135
  );


  not
  g392
  (
    n402,
    n117
  );


  buf
  g393
  (
    n213,
    n160
  );


  buf
  g394
  (
    n204,
    n40
  );


  not
  g395
  (
    n454,
    n84
  );


  buf
  g396
  (
    n617,
    n127
  );


  not
  g397
  (
    n367,
    n157
  );


  buf
  g398
  (
    n552,
    n74
  );


  buf
  g399
  (
    n526,
    n96
  );


  not
  g400
  (
    n596,
    n56
  );


  not
  g401
  (
    n325,
    n90
  );


  not
  g402
  (
    n432,
    n98
  );


  buf
  g403
  (
    n268,
    n148
  );


  not
  g404
  (
    n666,
    n69
  );


  buf
  g405
  (
    n225,
    n62
  );


  buf
  g406
  (
    n282,
    n36
  );


  buf
  g407
  (
    n650,
    n94
  );


  not
  g408
  (
    n311,
    n82
  );


  not
  g409
  (
    n671,
    n110
  );


  buf
  g410
  (
    n399,
    n79
  );


  not
  g411
  (
    n439,
    n75
  );


  buf
  g412
  (
    n471,
    n60
  );


  buf
  g413
  (
    n300,
    n91
  );


  not
  g414
  (
    n283,
    n91
  );


  not
  g415
  (
    n302,
    n53
  );


  not
  g416
  (
    n366,
    n47
  );


  not
  g417
  (
    n511,
    n72
  );


  buf
  g418
  (
    n347,
    n78
  );


  buf
  g419
  (
    n243,
    n86
  );


  buf
  g420
  (
    n266,
    n133
  );


  buf
  g421
  (
    n538,
    n97
  );


  not
  g422
  (
    n209,
    n104
  );


  buf
  g423
  (
    n658,
    n44
  );


  not
  g424
  (
    n423,
    n160
  );


  buf
  g425
  (
    KeyWire_0_4,
    n98
  );


  not
  g426
  (
    n600,
    n151
  );


  not
  g427
  (
    n232,
    n149
  );


  buf
  g428
  (
    n259,
    n38
  );


  buf
  g429
  (
    n495,
    n62
  );


  not
  g430
  (
    n564,
    n68
  );


  buf
  g431
  (
    n549,
    n54
  );


  buf
  g432
  (
    n187,
    n113
  );


  not
  g433
  (
    n664,
    n105
  );


  not
  g434
  (
    n195,
    n35
  );


  buf
  g435
  (
    n542,
    n68
  );


  not
  g436
  (
    n368,
    n39
  );


  buf
  g437
  (
    n214,
    n36
  );


  buf
  g438
  (
    n382,
    n54
  );


  not
  g439
  (
    n543,
    n63
  );


  not
  g440
  (
    n635,
    n124
  );


  not
  g441
  (
    n572,
    n100
  );


  buf
  g442
  (
    n320,
    n71
  );


  buf
  g443
  (
    n386,
    n158
  );


  buf
  g444
  (
    n164,
    n75
  );


  buf
  g445
  (
    n301,
    n38
  );


  buf
  g446
  (
    n645,
    n156
  );


  not
  g447
  (
    n362,
    n54
  );


  not
  g448
  (
    n504,
    n152
  );


  buf
  g449
  (
    n446,
    n109
  );


  buf
  g450
  (
    n465,
    n88
  );


  not
  g451
  (
    n408,
    n159
  );


  not
  g452
  (
    n190,
    n52
  );


  buf
  g453
  (
    n558,
    n138
  );


  not
  g454
  (
    n226,
    n42
  );


  buf
  g455
  (
    n371,
    n80
  );


  buf
  g456
  (
    n566,
    n136
  );


  buf
  g457
  (
    n312,
    n130
  );


  not
  g458
  (
    n601,
    n33
  );


  not
  g459
  (
    n180,
    n83
  );


  buf
  g460
  (
    n350,
    n55
  );


  not
  g461
  (
    KeyWire_0_18,
    n126
  );


  not
  g462
  (
    n460,
    n75
  );


  buf
  g463
  (
    n480,
    n57
  );


  not
  g464
  (
    n612,
    n87
  );


  not
  g465
  (
    n475,
    n41
  );


  not
  g466
  (
    n406,
    n113
  );


  buf
  g467
  (
    n197,
    n79
  );


  buf
  g468
  (
    n416,
    n147
  );


  buf
  g469
  (
    n563,
    n40
  );


  buf
  g470
  (
    n455,
    n134
  );


  not
  g471
  (
    n575,
    n111
  );


  buf
  g472
  (
    n585,
    n52
  );


  not
  g473
  (
    n649,
    n49
  );


  not
  g474
  (
    n303,
    n103
  );


  not
  g475
  (
    n235,
    n33
  );


  not
  g476
  (
    n615,
    n156
  );


  not
  g477
  (
    n445,
    n132
  );


  not
  g478
  (
    n647,
    n50
  );


  buf
  g479
  (
    n318,
    n139
  );


  not
  g480
  (
    n643,
    n137
  );


  buf
  g481
  (
    n216,
    n114
  );


  buf
  g482
  (
    n284,
    n104
  );


  not
  g483
  (
    n470,
    n133
  );


  buf
  g484
  (
    n497,
    n81
  );


  buf
  g485
  (
    n231,
    n85
  );


  not
  g486
  (
    n541,
    n157
  );


  buf
  g487
  (
    n498,
    n129
  );


  buf
  g488
  (
    n521,
    n51
  );


  not
  g489
  (
    n546,
    n109
  );


  buf
  g490
  (
    n577,
    n78
  );


  not
  g491
  (
    n373,
    n49
  );


  buf
  g492
  (
    n167,
    n74
  );


  not
  g493
  (
    n622,
    n97
  );


  not
  g494
  (
    n536,
    n77
  );


  not
  g495
  (
    n592,
    n39
  );


  not
  g496
  (
    n388,
    n116
  );


  not
  g497
  (
    n627,
    n114
  );


  buf
  g498
  (
    n170,
    n98
  );


  buf
  g499
  (
    n410,
    n34
  );


  buf
  g500
  (
    n597,
    n143
  );


  not
  g501
  (
    n637,
    n64
  );


  buf
  g502
  (
    n414,
    n84
  );


  buf
  g503
  (
    n291,
    n150
  );


  not
  g504
  (
    n427,
    n139
  );


  buf
  g505
  (
    n606,
    n142
  );


  not
  g506
  (
    n661,
    n60
  );


  buf
  g507
  (
    n313,
    n96
  );


  buf
  g508
  (
    n636,
    n49
  );


  not
  g509
  (
    n447,
    n159
  );


  not
  g510
  (
    n499,
    n50
  );


  buf
  g511
  (
    n327,
    n158
  );


  not
  g512
  (
    n443,
    n129
  );


  buf
  g513
  (
    n183,
    n62
  );


  not
  g514
  (
    n224,
    n114
  );


  not
  g515
  (
    n619,
    n75
  );


  buf
  g516
  (
    n338,
    n124
  );


  not
  g517
  (
    n288,
    n120
  );


  not
  g518
  (
    n250,
    n47
  );


  buf
  g519
  (
    n424,
    n93
  );


  not
  g520
  (
    n309,
    n106
  );


  not
  g521
  (
    n236,
    n132
  );


  buf
  g522
  (
    n230,
    n93
  );


  buf
  g523
  (
    n299,
    n88
  );


  not
  g524
  (
    n240,
    n147
  );


  buf
  g525
  (
    n430,
    n142
  );


  buf
  g526
  (
    n251,
    n108
  );


  buf
  g527
  (
    n626,
    n48
  );


  buf
  g528
  (
    n550,
    n41
  );


  buf
  g529
  (
    n329,
    n148
  );


  not
  g530
  (
    n411,
    n120
  );


  buf
  g531
  (
    n343,
    n113
  );


  not
  g532
  (
    n609,
    n116
  );


  buf
  g533
  (
    n326,
    n118
  );


  not
  g534
  (
    n161,
    n141
  );


  not
  g535
  (
    n260,
    n119
  );


  not
  g536
  (
    n314,
    n137
  );


  buf
  g537
  (
    n669,
    n106
  );


  buf
  g538
  (
    n483,
    n139
  );


  buf
  g539
  (
    n192,
    n133
  );


  not
  g540
  (
    n535,
    n133
  );


  not
  g541
  (
    n474,
    n74
  );


  not
  g542
  (
    n341,
    n33
  );


  buf
  g543
  (
    n527,
    n64
  );


  not
  g544
  (
    n436,
    n53
  );


  not
  g545
  (
    n358,
    n129
  );


  buf
  g546
  (
    n162,
    n48
  );


  not
  g547
  (
    n434,
    n63
  );


  buf
  g548
  (
    n633,
    n89
  );


  not
  g549
  (
    n468,
    n58
  );


  not
  g550
  (
    n369,
    n73
  );


  buf
  g551
  (
    n278,
    n65
  );


  buf
  g552
  (
    n603,
    n155
  );


  not
  g553
  (
    n223,
    n86
  );


  buf
  g554
  (
    n473,
    n158
  );


  buf
  g555
  (
    n539,
    n145
  );


  buf
  g556
  (
    n663,
    n76
  );


  buf
  g557
  (
    n199,
    n89
  );


  not
  g558
  (
    n496,
    n66
  );


  buf
  g559
  (
    n540,
    n134
  );


  not
  g560
  (
    n248,
    n151
  );


  buf
  g561
  (
    n271,
    n143
  );


  buf
  g562
  (
    n610,
    n95
  );


  buf
  g563
  (
    n261,
    n154
  );


  buf
  g564
  (
    n237,
    n116
  );


  buf
  g565
  (
    n365,
    n37
  );


  not
  g566
  (
    n644,
    n34
  );


  not
  g567
  (
    n317,
    n89
  );


  buf
  g568
  (
    n184,
    n151
  );


  buf
  g569
  (
    n290,
    n101
  );


  buf
  g570
  (
    n537,
    n94
  );


  not
  g571
  (
    n220,
    n134
  );


  buf
  g572
  (
    n440,
    n67
  );


  buf
  g573
  (
    n380,
    n123
  );


  buf
  g574
  (
    n210,
    n37
  );


  buf
  g575
  (
    n360,
    n142
  );


  not
  g576
  (
    n554,
    n58
  );


  buf
  g577
  (
    n579,
    n145
  );


  buf
  g578
  (
    n490,
    n148
  );


  buf
  g579
  (
    n401,
    n131
  );


  not
  g580
  (
    n166,
    n51
  );


  not
  g581
  (
    n632,
    n125
  );


  buf
  g582
  (
    KeyWire_0_14,
    n53
  );


  not
  g583
  (
    n574,
    n87
  );


  buf
  g584
  (
    n516,
    n115
  );


  not
  g585
  (
    n630,
    n101
  );


  buf
  g586
  (
    n651,
    n90
  );


  not
  g587
  (
    n201,
    n82
  );


  not
  g588
  (
    n335,
    n148
  );


  buf
  g589
  (
    n607,
    n60
  );


  not
  g590
  (
    n500,
    n121
  );


  not
  g591
  (
    n203,
    n97
  );


  not
  g592
  (
    n324,
    n132
  );


  buf
  g593
  (
    n567,
    n45
  );


  buf
  g594
  (
    n333,
    n85
  );


  not
  g595
  (
    n580,
    n59
  );


  not
  g596
  (
    n451,
    n42
  );


  buf
  g597
  (
    n584,
    n74
  );


  buf
  g598
  (
    n640,
    n136
  );


  buf
  g599
  (
    n553,
    n121
  );


  buf
  g600
  (
    n568,
    n112
  );


  not
  g601
  (
    n400,
    n92
  );


  not
  g602
  (
    n462,
    n155
  );


  buf
  g603
  (
    n501,
    n43
  );


  not
  g604
  (
    n361,
    n155
  );


  not
  g605
  (
    n604,
    n130
  );


  not
  g606
  (
    n202,
    n138
  );


  buf
  g607
  (
    n449,
    n121
  );


  buf
  g608
  (
    n321,
    n113
  );


  buf
  g609
  (
    n372,
    n47
  );


  not
  g610
  (
    n172,
    n63
  );


  not
  g611
  (
    n339,
    n68
  );


  not
  g612
  (
    n565,
    n147
  );


  not
  g613
  (
    n507,
    n59
  );


  not
  g614
  (
    n391,
    n84
  );


  not
  g615
  (
    n353,
    n46
  );


  not
  g616
  (
    n624,
    n45
  );


  not
  g617
  (
    n267,
    n144
  );


  buf
  g618
  (
    n477,
    n149
  );


  not
  g619
  (
    n662,
    n39
  );


  buf
  g620
  (
    n629,
    n147
  );


  not
  g621
  (
    n173,
    n35
  );


  buf
  g622
  (
    n245,
    n67
  );


  buf
  g623
  (
    n253,
    n110
  );


  buf
  g624
  (
    n618,
    n77
  );


  buf
  g625
  (
    n594,
    n99
  );


  buf
  g626
  (
    n294,
    n149
  );


  not
  g627
  (
    n279,
    n46
  );


  not
  g628
  (
    n548,
    n59
  );


  buf
  g629
  (
    n556,
    n43
  );


  not
  g630
  (
    n528,
    n81
  );


  not
  g631
  (
    n623,
    n116
  );


  not
  g632
  (
    n415,
    n72
  );


  buf
  g633
  (
    n667,
    n94
  );


  not
  g634
  (
    n277,
    n107
  );


  buf
  g635
  (
    n448,
    n91
  );


  not
  g636
  (
    n453,
    n108
  );


  buf
  g637
  (
    n207,
    n43
  );


  not
  g638
  (
    n381,
    n61
  );


  not
  g639
  (
    n1148,
    n580
  );


  not
  g640
  (
    n1336,
    n246
  );


  not
  g641
  (
    n1036,
    n376
  );


  not
  g642
  (
    n2116,
    n509
  );


  buf
  g643
  (
    n1476,
    n264
  );


  buf
  g644
  (
    n1326,
    n306
  );


  not
  g645
  (
    n1070,
    n312
  );


  not
  g646
  (
    n795,
    n669
  );


  buf
  g647
  (
    n1628,
    n463
  );


  not
  g648
  (
    n1657,
    n576
  );


  buf
  g649
  (
    n1842,
    n581
  );


  buf
  g650
  (
    n1631,
    n439
  );


  buf
  g651
  (
    n1923,
    n279
  );


  buf
  g652
  (
    n1032,
    n625
  );


  not
  g653
  (
    n1684,
    n633
  );


  not
  g654
  (
    n1038,
    n238
  );


  not
  g655
  (
    n1682,
    n229
  );


  not
  g656
  (
    n1022,
    n640
  );


  not
  g657
  (
    n1922,
    n455
  );


  not
  g658
  (
    n2048,
    n388
  );


  not
  g659
  (
    n813,
    n602
  );


  buf
  g660
  (
    n2059,
    n642
  );


  not
  g661
  (
    n1150,
    n539
  );


  buf
  g662
  (
    n1529,
    n665
  );


  not
  g663
  (
    n1174,
    n657
  );


  buf
  g664
  (
    n828,
    n618
  );


  buf
  g665
  (
    n1295,
    n167
  );


  not
  g666
  (
    n1074,
    n373
  );


  buf
  g667
  (
    n826,
    n581
  );


  buf
  g668
  (
    n2133,
    n570
  );


  not
  g669
  (
    n1055,
    n428
  );


  not
  g670
  (
    n1392,
    n301
  );


  buf
  g671
  (
    n1508,
    n441
  );


  not
  g672
  (
    n1368,
    n534
  );


  buf
  g673
  (
    n1729,
    n329
  );


  buf
  g674
  (
    n768,
    n392
  );


  not
  g675
  (
    n1548,
    n309
  );


  not
  g676
  (
    n846,
    n411
  );


  buf
  g677
  (
    n872,
    n321
  );


  not
  g678
  (
    n1283,
    n414
  );


  buf
  g679
  (
    n1945,
    n255
  );


  not
  g680
  (
    n1512,
    n453
  );


  buf
  g681
  (
    n1853,
    n343
  );


  not
  g682
  (
    n1086,
    n202
  );


  buf
  g683
  (
    n776,
    n409
  );


  buf
  g684
  (
    n1457,
    n443
  );


  buf
  g685
  (
    n1267,
    n407
  );


  not
  g686
  (
    n2070,
    n195
  );


  not
  g687
  (
    n1388,
    n351
  );


  buf
  g688
  (
    n1469,
    n635
  );


  not
  g689
  (
    n1587,
    n403
  );


  not
  g690
  (
    n2054,
    n297
  );


  not
  g691
  (
    n1535,
    n172
  );


  not
  g692
  (
    n1409,
    n303
  );


  buf
  g693
  (
    n2147,
    n527
  );


  buf
  g694
  (
    n1594,
    n333
  );


  buf
  g695
  (
    n1390,
    n522
  );


  not
  g696
  (
    n2140,
    n201
  );


  not
  g697
  (
    n1484,
    n329
  );


  not
  g698
  (
    n1081,
    n478
  );


  buf
  g699
  (
    n1609,
    n197
  );


  not
  g700
  (
    n704,
    n633
  );


  not
  g701
  (
    n1536,
    n376
  );


  buf
  g702
  (
    n1565,
    n404
  );


  buf
  g703
  (
    n2055,
    n663
  );


  buf
  g704
  (
    n2023,
    n205
  );


  not
  g705
  (
    n1758,
    n208
  );


  buf
  g706
  (
    n1818,
    n276
  );


  not
  g707
  (
    n889,
    n531
  );


  not
  g708
  (
    n1692,
    n336
  );


  buf
  g709
  (
    n1488,
    n402
  );


  not
  g710
  (
    n1870,
    n339
  );


  buf
  g711
  (
    n2016,
    n402
  );


  not
  g712
  (
    n1239,
    n161
  );


  not
  g713
  (
    n1294,
    n570
  );


  not
  g714
  (
    n1837,
    n385
  );


  not
  g715
  (
    n1685,
    n573
  );


  not
  g716
  (
    n1761,
    n424
  );


  not
  g717
  (
    n944,
    n408
  );


  buf
  g718
  (
    n733,
    n347
  );


  buf
  g719
  (
    n1528,
    n203
  );


  not
  g720
  (
    n1834,
    n313
  );


  not
  g721
  (
    n843,
    n197
  );


  not
  g722
  (
    KeyWire_0_59,
    n266
  );


  buf
  g723
  (
    n2076,
    n586
  );


  not
  g724
  (
    n1963,
    n613
  );


  not
  g725
  (
    n1816,
    n530
  );


  not
  g726
  (
    n1266,
    n343
  );


  buf
  g727
  (
    n760,
    n363
  );


  not
  g728
  (
    n1677,
    n161
  );


  not
  g729
  (
    KeyWire_0_34,
    n498
  );


  not
  g730
  (
    n1595,
    n370
  );


  not
  g731
  (
    n1701,
    n583
  );


  buf
  g732
  (
    n1833,
    n257
  );


  not
  g733
  (
    n1333,
    n515
  );


  buf
  g734
  (
    n1563,
    n495
  );


  buf
  g735
  (
    n1598,
    n287
  );


  buf
  g736
  (
    n1747,
    n517
  );


  buf
  g737
  (
    n1307,
    n477
  );


  buf
  g738
  (
    n1557,
    n368
  );


  not
  g739
  (
    n1315,
    n189
  );


  not
  g740
  (
    n1427,
    n629
  );


  buf
  g741
  (
    n1664,
    n433
  );


  buf
  g742
  (
    KeyWire_0_29,
    n248
  );


  not
  g743
  (
    n2075,
    n241
  );


  buf
  g744
  (
    n2000,
    n335
  );


  not
  g745
  (
    n2158,
    n430
  );


  buf
  g746
  (
    n1224,
    n518
  );


  not
  g747
  (
    n1982,
    n270
  );


  buf
  g748
  (
    n2060,
    n382
  );


  not
  g749
  (
    n787,
    n410
  );


  buf
  g750
  (
    n1337,
    n389
  );


  not
  g751
  (
    n945,
    n230
  );


  not
  g752
  (
    n685,
    n428
  );


  buf
  g753
  (
    n873,
    n586
  );


  buf
  g754
  (
    n1065,
    n599
  );


  buf
  g755
  (
    n745,
    n660
  );


  not
  g756
  (
    n1033,
    n497
  );


  not
  g757
  (
    n1796,
    n590
  );


  buf
  g758
  (
    KeyWire_0_26,
    n242
  );


  not
  g759
  (
    n792,
    n585
  );


  buf
  g760
  (
    n1251,
    n246
  );


  buf
  g761
  (
    n1447,
    n173
  );


  not
  g762
  (
    n1568,
    n444
  );


  not
  g763
  (
    n862,
    n285
  );


  buf
  g764
  (
    n984,
    n425
  );


  buf
  g765
  (
    n1054,
    n256
  );


  not
  g766
  (
    n988,
    n278
  );


  not
  g767
  (
    n848,
    n309
  );


  not
  g768
  (
    n1600,
    n491
  );


  not
  g769
  (
    n1420,
    n593
  );


  buf
  g770
  (
    n1031,
    n401
  );


  buf
  g771
  (
    n913,
    n532
  );


  not
  g772
  (
    n1357,
    n378
  );


  buf
  g773
  (
    n1791,
    n636
  );


  buf
  g774
  (
    n1769,
    n394
  );


  not
  g775
  (
    n1592,
    n614
  );


  not
  g776
  (
    n2160,
    n379
  );


  buf
  g777
  (
    n983,
    n320
  );


  buf
  g778
  (
    n800,
    n287
  );


  not
  g779
  (
    n1793,
    n606
  );


  not
  g780
  (
    n2028,
    n516
  );


  not
  g781
  (
    n751,
    n560
  );


  buf
  g782
  (
    n2139,
    n232
  );


  buf
  g783
  (
    n706,
    n642
  );


  buf
  g784
  (
    n1200,
    n250
  );


  not
  g785
  (
    n1317,
    n321
  );


  not
  g786
  (
    n2115,
    n329
  );


  not
  g787
  (
    n1374,
    n350
  );


  not
  g788
  (
    n1010,
    n181
  );


  not
  g789
  (
    n1708,
    n162
  );


  buf
  g790
  (
    n1013,
    n598
  );


  buf
  g791
  (
    n1415,
    n665
  );


  not
  g792
  (
    n2117,
    n407
  );


  buf
  g793
  (
    n918,
    n312
  );


  buf
  g794
  (
    n1716,
    n394
  );


  buf
  g795
  (
    n1369,
    n625
  );


  not
  g796
  (
    n1124,
    n559
  );


  not
  g797
  (
    n1932,
    n242
  );


  buf
  g798
  (
    n1840,
    n459
  );


  not
  g799
  (
    n1971,
    n440
  );


  buf
  g800
  (
    n747,
    n249
  );


  buf
  g801
  (
    n1218,
    n436
  );


  buf
  g802
  (
    n1160,
    n276
  );


  not
  g803
  (
    n1057,
    n225
  );


  not
  g804
  (
    n1211,
    n325
  );


  not
  g805
  (
    n1553,
    n656
  );


  not
  g806
  (
    n1227,
    n196
  );


  buf
  g807
  (
    n875,
    n328
  );


  not
  g808
  (
    n708,
    n638
  );


  buf
  g809
  (
    n995,
    n521
  );


  buf
  g810
  (
    n2134,
    n227
  );


  buf
  g811
  (
    n1001,
    n357
  );


  buf
  g812
  (
    n1698,
    n297
  );


  buf
  g813
  (
    n1771,
    n261
  );


  not
  g814
  (
    n1979,
    n206
  );


  not
  g815
  (
    n816,
    n570
  );


  not
  g816
  (
    n992,
    n431
  );


  buf
  g817
  (
    n1705,
    n640
  );


  buf
  g818
  (
    n772,
    n333
  );


  not
  g819
  (
    n1524,
    n200
  );


  not
  g820
  (
    n1353,
    n177
  );


  buf
  g821
  (
    n1459,
    n480
  );


  not
  g822
  (
    n2077,
    n609
  );


  not
  g823
  (
    n1732,
    n274
  );


  buf
  g824
  (
    n1398,
    n291
  );


  buf
  g825
  (
    n785,
    n391
  );


  buf
  g826
  (
    n1672,
    n507
  );


  buf
  g827
  (
    KeyWire_0_62,
    n241
  );


  buf
  g828
  (
    n1984,
    n233
  );


  not
  g829
  (
    n1396,
    n296
  );


  not
  g830
  (
    n1966,
    n470
  );


  buf
  g831
  (
    n1994,
    n624
  );


  buf
  g832
  (
    n1702,
    n204
  );


  buf
  g833
  (
    n2154,
    n632
  );


  buf
  g834
  (
    n2022,
    n605
  );


  not
  g835
  (
    n1309,
    n548
  );


  buf
  g836
  (
    n783,
    n576
  );


  not
  g837
  (
    n1175,
    n662
  );


  buf
  g838
  (
    n1428,
    n520
  );


  not
  g839
  (
    n1821,
    n231
  );


  buf
  g840
  (
    n842,
    n429
  );


  buf
  g841
  (
    n1872,
    n463
  );


  buf
  g842
  (
    n1412,
    n431
  );


  not
  g843
  (
    n1958,
    n634
  );


  buf
  g844
  (
    n749,
    n584
  );


  not
  g845
  (
    n1259,
    n231
  );


  not
  g846
  (
    n1318,
    n652
  );


  not
  g847
  (
    n1106,
    n521
  );


  not
  g848
  (
    n1989,
    n331
  );


  not
  g849
  (
    n1083,
    n481
  );


  buf
  g850
  (
    n2142,
    n532
  );


  buf
  g851
  (
    n1015,
    n400
  );


  buf
  g852
  (
    n1851,
    n198
  );


  buf
  g853
  (
    n895,
    n535
  );


  buf
  g854
  (
    n1522,
    n616
  );


  not
  g855
  (
    n1615,
    n604
  );


  buf
  g856
  (
    n1939,
    n223
  );


  buf
  g857
  (
    n2017,
    n393
  );


  buf
  g858
  (
    n936,
    n525
  );


  not
  g859
  (
    n993,
    n316
  );


  not
  g860
  (
    n1744,
    n343
  );


  not
  g861
  (
    n938,
    n283
  );


  buf
  g862
  (
    n1772,
    n613
  );


  buf
  g863
  (
    n2067,
    n507
  );


  buf
  g864
  (
    n709,
    n439
  );


  buf
  g865
  (
    n1449,
    n187
  );


  not
  g866
  (
    n2081,
    n614
  );


  not
  g867
  (
    n1216,
    n608
  );


  not
  g868
  (
    n683,
    n630
  );


  buf
  g869
  (
    n971,
    n409
  );


  buf
  g870
  (
    n1496,
    n564
  );


  not
  g871
  (
    n1857,
    n389
  );


  buf
  g872
  (
    n2145,
    n489
  );


  not
  g873
  (
    n1072,
    n415
  );


  buf
  g874
  (
    n1873,
    n437
  );


  not
  g875
  (
    n1110,
    n413
  );


  buf
  g876
  (
    n1815,
    n297
  );


  buf
  g877
  (
    n1859,
    n567
  );


  not
  g878
  (
    n1091,
    n607
  );


  buf
  g879
  (
    n2103,
    n378
  );


  not
  g880
  (
    n933,
    n172
  );


  buf
  g881
  (
    n1380,
    n386
  );


  not
  g882
  (
    n998,
    n198
  );


  buf
  g883
  (
    n2144,
    n221
  );


  not
  g884
  (
    n2121,
    n302
  );


  not
  g885
  (
    n1338,
    n277
  );


  buf
  g886
  (
    n824,
    n268
  );


  not
  g887
  (
    n1464,
    n165
  );


  buf
  g888
  (
    n2074,
    n437
  );


  buf
  g889
  (
    n950,
    n533
  );


  buf
  g890
  (
    n1432,
    n258
  );


  not
  g891
  (
    n1865,
    n312
  );


  not
  g892
  (
    n1136,
    n435
  );


  buf
  g893
  (
    n1654,
    n403
  );


  not
  g894
  (
    n915,
    n377
  );


  not
  g895
  (
    n1511,
    n206
  );


  not
  g896
  (
    n871,
    n504
  );


  not
  g897
  (
    n844,
    n164
  );


  buf
  g898
  (
    n851,
    n162
  );


  not
  g899
  (
    n1276,
    n344
  );


  buf
  g900
  (
    n2063,
    n257
  );


  buf
  g901
  (
    n2112,
    n621
  );


  buf
  g902
  (
    n754,
    n632
  );


  buf
  g903
  (
    n694,
    n188
  );


  buf
  g904
  (
    n1825,
    n190
  );


  buf
  g905
  (
    n791,
    n382
  );


  buf
  g906
  (
    n825,
    n626
  );


  buf
  g907
  (
    n1823,
    n668
  );


  buf
  g908
  (
    n876,
    n613
  );


  not
  g909
  (
    n1981,
    n238
  );


  not
  g910
  (
    n1650,
    n488
  );


  buf
  g911
  (
    n1225,
    n383
  );


  buf
  g912
  (
    n1446,
    n623
  );


  not
  g913
  (
    n2053,
    n243
  );


  not
  g914
  (
    n1108,
    n460
  );


  buf
  g915
  (
    n1552,
    n429
  );


  not
  g916
  (
    n1205,
    n354
  );


  buf
  g917
  (
    n1079,
    n298
  );


  not
  g918
  (
    n1652,
    n267
  );


  buf
  g919
  (
    n1713,
    n498
  );


  not
  g920
  (
    n1454,
    n310
  );


  buf
  g921
  (
    n1616,
    n453
  );


  not
  g922
  (
    n1084,
    n656
  );


  buf
  g923
  (
    n2105,
    n502
  );


  buf
  g924
  (
    KeyWire_0_38,
    n554
  );


  buf
  g925
  (
    n1804,
    n487
  );


  not
  g926
  (
    n1406,
    n395
  );


  not
  g927
  (
    n1864,
    n204
  );


  not
  g928
  (
    n1291,
    n196
  );


  buf
  g929
  (
    n1786,
    n182
  );


  not
  g930
  (
    n1012,
    n384
  );


  not
  g931
  (
    n1005,
    n562
  );


  buf
  g932
  (
    n1444,
    n556
  );


  buf
  g933
  (
    n829,
    n396
  );


  buf
  g934
  (
    n1169,
    n348
  );


  not
  g935
  (
    n2004,
    n647
  );


  buf
  g936
  (
    n974,
    n260
  );


  buf
  g937
  (
    n2079,
    n375
  );


  buf
  g938
  (
    n1410,
    n506
  );


  not
  g939
  (
    n1092,
    n251
  );


  not
  g940
  (
    n1139,
    n651
  );


  buf
  g941
  (
    n2141,
    n494
  );


  not
  g942
  (
    n1688,
    n216
  );


  buf
  g943
  (
    n898,
    n496
  );


  not
  g944
  (
    n1877,
    n298
  );


  buf
  g945
  (
    n1610,
    n594
  );


  buf
  g946
  (
    n1117,
    n375
  );


  not
  g947
  (
    n1897,
    n331
  );


  buf
  g948
  (
    n1479,
    n410
  );


  not
  g949
  (
    n966,
    n500
  );


  not
  g950
  (
    n2162,
    n193
  );


  not
  g951
  (
    n1088,
    n544
  );


  not
  g952
  (
    n1782,
    n469
  );


  not
  g953
  (
    n967,
    n663
  );


  buf
  g954
  (
    n2156,
    n412
  );


  buf
  g955
  (
    n1644,
    n426
  );


  buf
  g956
  (
    n1413,
    n333
  );


  not
  g957
  (
    n1753,
    n226
  );


  buf
  g958
  (
    n1292,
    n554
  );


  buf
  g959
  (
    n1222,
    n240
  );


  not
  g960
  (
    n2064,
    n382
  );


  buf
  g961
  (
    n1120,
    n413
  );


  not
  g962
  (
    n827,
    n413
  );


  not
  g963
  (
    n1215,
    n324
  );


  buf
  g964
  (
    n817,
    n488
  );


  not
  g965
  (
    n734,
    n604
  );


  not
  g966
  (
    n1745,
    n493
  );


  not
  g967
  (
    n1442,
    n179
  );


  buf
  g968
  (
    n762,
    n486
  );


  buf
  g969
  (
    n1861,
    n510
  );


  buf
  g970
  (
    n1350,
    n449
  );


  buf
  g971
  (
    n2021,
    n619
  );


  buf
  g972
  (
    n1860,
    n630
  );


  not
  g973
  (
    n2088,
    n589
  );


  buf
  g974
  (
    n1187,
    n304
  );


  buf
  g975
  (
    n1911,
    n405
  );


  buf
  g976
  (
    n883,
    n572
  );


  not
  g977
  (
    n1576,
    n339
  );


  not
  g978
  (
    n2014,
    n575
  );


  not
  g979
  (
    n884,
    n269
  );


  not
  g980
  (
    n1930,
    n431
  );


  buf
  g981
  (
    n758,
    n418
  );


  not
  g982
  (
    n830,
    n508
  );


  buf
  g983
  (
    n820,
    n435
  );


  not
  g984
  (
    n1384,
    n426
  );


  not
  g985
  (
    n2157,
    n654
  );


  not
  g986
  (
    n1504,
    n282
  );


  not
  g987
  (
    n865,
    n241
  );


  buf
  g988
  (
    n1525,
    n390
  );


  not
  g989
  (
    n2082,
    n495
  );


  buf
  g990
  (
    n1327,
    n359
  );


  not
  g991
  (
    n1613,
    n216
  );


  buf
  g992
  (
    n1017,
    n401
  );


  not
  g993
  (
    n1142,
    n646
  );


  not
  g994
  (
    n1927,
    n175
  );


  buf
  g995
  (
    n1645,
    n380
  );


  not
  g996
  (
    n1289,
    n620
  );


  not
  g997
  (
    n859,
    n595
  );


  not
  g998
  (
    n2107,
    n295
  );


  not
  g999
  (
    n1992,
    n609
  );


  not
  g1000
  (
    n2015,
    n200
  );


  buf
  g1001
  (
    n986,
    n652
  );


  buf
  g1002
  (
    n1340,
    n463
  );


  buf
  g1003
  (
    n1736,
    n616
  );


  not
  g1004
  (
    n1207,
    n193
  );


  buf
  g1005
  (
    n1983,
    n508
  );


  buf
  g1006
  (
    n1405,
    n395
  );


  buf
  g1007
  (
    n1482,
    n443
  );


  not
  g1008
  (
    n1928,
    n653
  );


  not
  g1009
  (
    n1640,
    n410
  );


  buf
  g1010
  (
    n1544,
    n390
  );


  not
  g1011
  (
    KeyWire_0_61,
    n382
  );


  not
  g1012
  (
    n2032,
    n261
  );


  buf
  g1013
  (
    n1689,
    n162
  );


  buf
  g1014
  (
    n724,
    n617
  );


  buf
  g1015
  (
    n748,
    n399
  );


  buf
  g1016
  (
    n1501,
    n370
  );


  buf
  g1017
  (
    n1714,
    n179
  );


  buf
  g1018
  (
    n1310,
    n633
  );


  not
  g1019
  (
    KeyWire_0_41,
    n311
  );


  not
  g1020
  (
    n1844,
    n445
  );


  not
  g1021
  (
    n1324,
    n284
  );


  not
  g1022
  (
    n885,
    n453
  );


  buf
  g1023
  (
    n994,
    n163
  );


  not
  g1024
  (
    n839,
    n359
  );


  not
  g1025
  (
    n2106,
    n247
  );


  not
  g1026
  (
    n901,
    n234
  );


  buf
  g1027
  (
    n1248,
    n289
  );


  not
  g1028
  (
    n790,
    n236
  );


  buf
  g1029
  (
    n1313,
    n464
  );


  not
  g1030
  (
    n836,
    n233
  );


  buf
  g1031
  (
    n1836,
    n402
  );


  buf
  g1032
  (
    n1393,
    n466
  );


  buf
  g1033
  (
    n781,
    n615
  );


  not
  g1034
  (
    n1245,
    n529
  );


  buf
  g1035
  (
    n1591,
    n287
  );


  buf
  g1036
  (
    n1489,
    n175
  );


  buf
  g1037
  (
    n1797,
    n428
  );


  not
  g1038
  (
    n1290,
    n520
  );


  not
  g1039
  (
    n1360,
    n668
  );


  not
  g1040
  (
    n1542,
    n381
  );


  buf
  g1041
  (
    n1867,
    n338
  );


  not
  g1042
  (
    n1238,
    n594
  );


  buf
  g1043
  (
    n1530,
    n647
  );


  buf
  g1044
  (
    n799,
    n406
  );


  buf
  g1045
  (
    n1016,
    n217
  );


  not
  g1046
  (
    n1138,
    n663
  );


  buf
  g1047
  (
    n845,
    n364
  );


  not
  g1048
  (
    n963,
    n394
  );


  buf
  g1049
  (
    n1145,
    n654
  );


  buf
  g1050
  (
    n1909,
    n601
  );


  not
  g1051
  (
    n686,
    n314
  );


  buf
  g1052
  (
    n1363,
    n192
  );


  buf
  g1053
  (
    n1961,
    n649
  );


  buf
  g1054
  (
    n1739,
    n595
  );


  not
  g1055
  (
    n1445,
    n351
  );


  not
  g1056
  (
    KeyWire_0_28,
    n365
  );


  buf
  g1057
  (
    n1258,
    n638
  );


  not
  g1058
  (
    n1152,
    n161
  );


  not
  g1059
  (
    n674,
    n595
  );


  not
  g1060
  (
    n1474,
    n243
  );


  buf
  g1061
  (
    n1779,
    n438
  );


  not
  g1062
  (
    n1918,
    n562
  );


  buf
  g1063
  (
    n1402,
    n452
  );


  buf
  g1064
  (
    n1095,
    n164
  );


  buf
  g1065
  (
    n1165,
    n644
  );


  buf
  g1066
  (
    n1622,
    n298
  );


  buf
  g1067
  (
    n1249,
    n452
  );


  buf
  g1068
  (
    n1597,
    n171
  );


  buf
  g1069
  (
    n2013,
    n494
  );


  buf
  g1070
  (
    n921,
    n499
  );


  not
  g1071
  (
    n1726,
    n596
  );


  buf
  g1072
  (
    n1342,
    n511
  );


  not
  g1073
  (
    n904,
    n618
  );


  buf
  g1074
  (
    n717,
    n175
  );


  buf
  g1075
  (
    n1623,
    n550
  );


  not
  g1076
  (
    n1507,
    n432
  );


  not
  g1077
  (
    n1403,
    n505
  );


  buf
  g1078
  (
    n775,
    n481
  );


  not
  g1079
  (
    n1505,
    n430
  );


  buf
  g1080
  (
    n1451,
    n503
  );


  buf
  g1081
  (
    n1495,
    n587
  );


  buf
  g1082
  (
    n1467,
    n316
  );


  buf
  g1083
  (
    n1957,
    n441
  );


  not
  g1084
  (
    n2056,
    n555
  );


  not
  g1085
  (
    n2020,
    n275
  );


  buf
  g1086
  (
    n882,
    n559
  );


  not
  g1087
  (
    n1306,
    n369
  );


  buf
  g1088
  (
    n1471,
    n278
  );


  not
  g1089
  (
    n1781,
    n247
  );


  buf
  g1090
  (
    n1727,
    n341
  );


  not
  g1091
  (
    n1694,
    n500
  );


  buf
  g1092
  (
    n722,
    n176
  );


  not
  g1093
  (
    n2033,
    n214
  );


  not
  g1094
  (
    n2166,
    n467
  );


  buf
  g1095
  (
    n1988,
    n421
  );


  not
  g1096
  (
    n1443,
    n442
  );


  not
  g1097
  (
    n1641,
    n251
  );


  not
  g1098
  (
    n929,
    n562
  );


  not
  g1099
  (
    n1367,
    n653
  );


  buf
  g1100
  (
    n849,
    n222
  );


  buf
  g1101
  (
    n1183,
    n294
  );


  buf
  g1102
  (
    n1908,
    n233
  );


  not
  g1103
  (
    n922,
    n624
  );


  not
  g1104
  (
    n1257,
    n206
  );


  buf
  g1105
  (
    n2165,
    n286
  );


  not
  g1106
  (
    n1618,
    n305
  );


  not
  g1107
  (
    n1914,
    n368
  );


  not
  g1108
  (
    n1828,
    n263
  );


  not
  g1109
  (
    n2108,
    n289
  );


  not
  g1110
  (
    n739,
    n346
  );


  buf
  g1111
  (
    n999,
    n425
  );


  buf
  g1112
  (
    n1486,
    n632
  );


  buf
  g1113
  (
    n985,
    n226
  );


  not
  g1114
  (
    n1355,
    n543
  );


  buf
  g1115
  (
    n1087,
    n508
  );


  buf
  g1116
  (
    n1868,
    n221
  );


  buf
  g1117
  (
    n1075,
    n401
  );


  buf
  g1118
  (
    n1305,
    n587
  );


  buf
  g1119
  (
    n2031,
    n479
  );


  not
  g1120
  (
    n1284,
    n168
  );


  not
  g1121
  (
    n2071,
    n248
  );


  buf
  g1122
  (
    n982,
    n239
  );


  not
  g1123
  (
    n2096,
    n497
  );


  not
  g1124
  (
    n1855,
    n338
  );


  buf
  g1125
  (
    n1993,
    n631
  );


  buf
  g1126
  (
    n1558,
    n472
  );


  buf
  g1127
  (
    n1666,
    n285
  );


  not
  g1128
  (
    KeyWire_0_46,
    n628
  );


  not
  g1129
  (
    n2094,
    n409
  );


  buf
  g1130
  (
    n2002,
    n166
  );


  buf
  g1131
  (
    KeyWire_0_20,
    n476
  );


  not
  g1132
  (
    n1349,
    n179
  );


  buf
  g1133
  (
    n2090,
    n379
  );


  not
  g1134
  (
    n1460,
    n568
  );


  not
  g1135
  (
    n723,
    n460
  );


  not
  g1136
  (
    n1933,
    n260
  );


  buf
  g1137
  (
    n756,
    n521
  );


  buf
  g1138
  (
    n2043,
    n219
  );


  buf
  g1139
  (
    n1812,
    n190
  );


  not
  g1140
  (
    n1921,
    n488
  );


  buf
  g1141
  (
    n1049,
    n432
  );


  buf
  g1142
  (
    n928,
    n660
  );


  buf
  g1143
  (
    n1438,
    n443
  );


  buf
  g1144
  (
    n1206,
    n416
  );


  buf
  g1145
  (
    n1599,
    n255
  );


  not
  g1146
  (
    n1299,
    n473
  );


  buf
  g1147
  (
    n887,
    n205
  );


  buf
  g1148
  (
    n1977,
    n190
  );


  buf
  g1149
  (
    n1068,
    n457
  );


  buf
  g1150
  (
    n1630,
    n550
  );


  buf
  g1151
  (
    n1119,
    n322
  );


  buf
  g1152
  (
    n1439,
    n279
  );


  not
  g1153
  (
    n1627,
    n186
  );


  not
  g1154
  (
    n1827,
    n519
  );


  buf
  g1155
  (
    n2122,
    n602
  );


  buf
  g1156
  (
    n1556,
    n212
  );


  buf
  g1157
  (
    n1741,
    n484
  );


  buf
  g1158
  (
    n1004,
    n345
  );


  buf
  g1159
  (
    n1007,
    n474
  );


  buf
  g1160
  (
    n1112,
    n512
  );


  buf
  g1161
  (
    n855,
    n468
  );


  buf
  g1162
  (
    n1233,
    n173
  );


  buf
  g1163
  (
    n1456,
    n557
  );


  not
  g1164
  (
    n1799,
    n371
  );


  not
  g1165
  (
    n1899,
    n422
  );


  buf
  g1166
  (
    n713,
    n418
  );


  not
  g1167
  (
    n1064,
    n361
  );


  buf
  g1168
  (
    n1240,
    n445
  );


  not
  g1169
  (
    n805,
    n594
  );


  not
  g1170
  (
    n1843,
    n197
  );


  not
  g1171
  (
    n1792,
    n475
  );


  not
  g1172
  (
    n1241,
    n169
  );


  buf
  g1173
  (
    n682,
    n542
  );


  not
  g1174
  (
    n750,
    n262
  );


  buf
  g1175
  (
    n1925,
    n594
  );


  not
  g1176
  (
    n2050,
    n626
  );


  not
  g1177
  (
    n1356,
    n665
  );


  buf
  g1178
  (
    n919,
    n249
  );


  not
  g1179
  (
    n1231,
    n307
  );


  buf
  g1180
  (
    n1743,
    n343
  );


  buf
  g1181
  (
    n906,
    n536
  );


  not
  g1182
  (
    n1281,
    n213
  );


  buf
  g1183
  (
    n2025,
    n363
  );


  not
  g1184
  (
    n818,
    n543
  );


  buf
  g1185
  (
    n767,
    n425
  );


  not
  g1186
  (
    n1237,
    n485
  );


  not
  g1187
  (
    n1431,
    n412
  );


  buf
  g1188
  (
    n1775,
    n394
  );


  buf
  g1189
  (
    n1951,
    n319
  );


  buf
  g1190
  (
    n1102,
    n219
  );


  buf
  g1191
  (
    n779,
    n228
  );


  buf
  g1192
  (
    n1962,
    n191
  );


  buf
  g1193
  (
    n1730,
    n484
  );


  not
  g1194
  (
    n1904,
    n613
  );


  buf
  g1195
  (
    n1419,
    n520
  );


  buf
  g1196
  (
    n1990,
    n575
  );


  not
  g1197
  (
    n1819,
    n406
  );


  buf
  g1198
  (
    n953,
    n311
  );


  buf
  g1199
  (
    n2009,
    n471
  );


  buf
  g1200
  (
    n1649,
    n652
  );


  not
  g1201
  (
    n1448,
    n317
  );


  buf
  g1202
  (
    n675,
    n335
  );


  not
  g1203
  (
    n1056,
    n194
  );


  buf
  g1204
  (
    n912,
    n483
  );


  not
  g1205
  (
    n1098,
    n371
  );


  buf
  g1206
  (
    n1386,
    n615
  );


  not
  g1207
  (
    n1720,
    n496
  );


  buf
  g1208
  (
    n1892,
    n189
  );


  not
  g1209
  (
    n1361,
    n549
  );


  not
  g1210
  (
    n947,
    n395
  );


  buf
  g1211
  (
    n2011,
    n165
  );


  buf
  g1212
  (
    n1626,
    n250
  );


  not
  g1213
  (
    n2136,
    n487
  );


  buf
  g1214
  (
    n2080,
    n372
  );


  not
  g1215
  (
    n1637,
    n397
  );


  not
  g1216
  (
    n1133,
    n199
  );


  not
  g1217
  (
    n766,
    n662
  );


  not
  g1218
  (
    n1230,
    n170
  );


  not
  g1219
  (
    n905,
    n619
  );


  buf
  g1220
  (
    n1039,
    n307
  );


  not
  g1221
  (
    n2085,
    n188
  );


  buf
  g1222
  (
    n1734,
    n186
  );


  not
  g1223
  (
    n1541,
    n448
  );


  buf
  g1224
  (
    n1164,
    n482
  );


  not
  g1225
  (
    n1123,
    n483
  );


  not
  g1226
  (
    n1676,
    n350
  );


  not
  g1227
  (
    n1316,
    n454
  );


  buf
  g1228
  (
    n880,
    n631
  );


  not
  g1229
  (
    n1416,
    n294
  );


  buf
  g1230
  (
    n1906,
    n176
  );


  not
  g1231
  (
    n1566,
    n553
  );


  not
  g1232
  (
    n1399,
    n663
  );


  not
  g1233
  (
    n1322,
    n540
  );


  buf
  g1234
  (
    n1303,
    n448
  );


  buf
  g1235
  (
    n1748,
    n295
  );


  buf
  g1236
  (
    n1585,
    n559
  );


  buf
  g1237
  (
    n1509,
    n511
  );


  buf
  g1238
  (
    n1441,
    n574
  );


  not
  g1239
  (
    n1320,
    n554
  );


  not
  g1240
  (
    n1625,
    n345
  );


  not
  g1241
  (
    n1182,
    n531
  );


  buf
  g1242
  (
    n1076,
    n604
  );


  not
  g1243
  (
    n1875,
    n377
  );


  buf
  g1244
  (
    n2104,
    n466
  );


  buf
  g1245
  (
    n1339,
    n482
  );


  not
  g1246
  (
    n1767,
    n575
  );


  not
  g1247
  (
    n977,
    n617
  );


  not
  g1248
  (
    n2163,
    n220
  );


  not
  g1249
  (
    n688,
    n523
  );


  buf
  g1250
  (
    n1903,
    n478
  );


  not
  g1251
  (
    n958,
    n253
  );


  buf
  g1252
  (
    n1999,
    n556
  );


  not
  g1253
  (
    n2111,
    n337
  );


  not
  g1254
  (
    n1277,
    n508
  );


  not
  g1255
  (
    n1204,
    n522
  );


  buf
  g1256
  (
    n1293,
    n231
  );


  not
  g1257
  (
    n1662,
    n563
  );


  not
  g1258
  (
    n949,
    n641
  );


  buf
  g1259
  (
    n1040,
    n658
  );


  buf
  g1260
  (
    n1704,
    n424
  );


  buf
  g1261
  (
    n2114,
    n566
  );


  buf
  g1262
  (
    n1247,
    n534
  );


  not
  g1263
  (
    n1733,
    n175
  );


  buf
  g1264
  (
    n976,
    n670
  );


  not
  g1265
  (
    n925,
    n397
  );


  not
  g1266
  (
    n877,
    n302
  );


  buf
  g1267
  (
    n1463,
    n237
  );


  buf
  g1268
  (
    n2030,
    n364
  );


  buf
  g1269
  (
    n1547,
    n412
  );


  buf
  g1270
  (
    n1395,
    n373
  );


  not
  g1271
  (
    n1126,
    n276
  );


  not
  g1272
  (
    n1611,
    n199
  );


  buf
  g1273
  (
    n1890,
    n505
  );


  not
  g1274
  (
    n1659,
    n592
  );


  not
  g1275
  (
    n797,
    n291
  );


  not
  g1276
  (
    n911,
    n271
  );


  not
  g1277
  (
    n1208,
    n556
  );


  not
  g1278
  (
    n908,
    n317
  );


  not
  g1279
  (
    n1784,
    n587
  );


  buf
  g1280
  (
    n2036,
    n619
  );


  buf
  g1281
  (
    n1341,
    n272
  );


  not
  g1282
  (
    n899,
    n524
  );


  not
  g1283
  (
    n1731,
    n384
  );


  not
  g1284
  (
    n1468,
    n596
  );


  not
  g1285
  (
    n903,
    n627
  );


  buf
  g1286
  (
    n1069,
    n318
  );


  not
  g1287
  (
    n1605,
    n398
  );


  not
  g1288
  (
    n2095,
    n240
  );


  buf
  g1289
  (
    n1477,
    n355
  );


  not
  g1290
  (
    n1681,
    n440
  );


  buf
  g1291
  (
    n770,
    n185
  );


  not
  g1292
  (
    n2167,
    n352
  );


  not
  g1293
  (
    n1564,
    n191
  );


  buf
  g1294
  (
    n1889,
    n638
  );


  buf
  g1295
  (
    n1633,
    n509
  );


  not
  g1296
  (
    n1255,
    n399
  );


  buf
  g1297
  (
    n1268,
    n261
  );


  buf
  g1298
  (
    n847,
    n549
  );


  not
  g1299
  (
    n757,
    n551
  );


  buf
  g1300
  (
    n1862,
    n336
  );


  not
  g1301
  (
    n1061,
    n171
  );


  buf
  g1302
  (
    n1571,
    n606
  );


  buf
  g1303
  (
    n939,
    n191
  );


  buf
  g1304
  (
    n1185,
    n655
  );


  buf
  g1305
  (
    n1693,
    n427
  );


  not
  g1306
  (
    n1869,
    n446
  );


  not
  g1307
  (
    n832,
    n408
  );


  buf
  g1308
  (
    n721,
    n273
  );


  buf
  g1309
  (
    n1777,
    n420
  );


  buf
  g1310
  (
    n1304,
    n373
  );


  not
  g1311
  (
    n1429,
    n546
  );


  not
  g1312
  (
    n1789,
    n407
  );


  buf
  g1313
  (
    n1329,
    n588
  );


  not
  g1314
  (
    n1876,
    n537
  );


  buf
  g1315
  (
    n1936,
    n670
  );


  not
  g1316
  (
    n951,
    n580
  );


  not
  g1317
  (
    n1638,
    n486
  );


  not
  g1318
  (
    n1912,
    n296
  );


  not
  g1319
  (
    n1082,
    n187
  );


  buf
  g1320
  (
    n968,
    n655
  );


  buf
  g1321
  (
    n2137,
    n275
  );


  buf
  g1322
  (
    n1274,
    n607
  );


  not
  g1323
  (
    n1590,
    n427
  );


  buf
  g1324
  (
    n2120,
    n557
  );


  buf
  g1325
  (
    n1440,
    n589
  );


  buf
  g1326
  (
    n1179,
    n538
  );


  not
  g1327
  (
    n2034,
    n469
  );


  not
  g1328
  (
    n1394,
    n166
  );


  not
  g1329
  (
    n1213,
    n558
  );


  not
  g1330
  (
    n1668,
    n245
  );


  not
  g1331
  (
    n838,
    n492
  );


  not
  g1332
  (
    n1915,
    n526
  );


  not
  g1333
  (
    n1273,
    n388
  );


  buf
  g1334
  (
    n1243,
    n334
  );


  not
  g1335
  (
    n1115,
    n439
  );


  not
  g1336
  (
    n1674,
    n583
  );


  not
  g1337
  (
    n1973,
    n448
  );


  not
  g1338
  (
    n1724,
    n254
  );


  not
  g1339
  (
    n1871,
    n596
  );


  not
  g1340
  (
    n2078,
    n328
  );


  buf
  g1341
  (
    n926,
    n432
  );


  buf
  g1342
  (
    n696,
    n269
  );


  not
  g1343
  (
    n1109,
    n332
  );


  not
  g1344
  (
    n1907,
    n203
  );


  buf
  g1345
  (
    n1332,
    n462
  );


  not
  g1346
  (
    n755,
    n362
  );


  not
  g1347
  (
    n784,
    n592
  );


  not
  g1348
  (
    n1824,
    n316
  );


  not
  g1349
  (
    n1596,
    n360
  );


  buf
  g1350
  (
    n823,
    n464
  );


  buf
  g1351
  (
    n1354,
    n528
  );


  not
  g1352
  (
    n2164,
    n269
  );


  not
  g1353
  (
    n1312,
    n396
  );


  not
  g1354
  (
    n2143,
    n667
  );


  buf
  g1355
  (
    n2068,
    n301
  );


  buf
  g1356
  (
    n1382,
    n348
  );


  not
  g1357
  (
    n856,
    n583
  );


  buf
  g1358
  (
    n1144,
    n538
  );


  buf
  g1359
  (
    n809,
    n321
  );


  not
  g1360
  (
    n1172,
    n221
  );


  buf
  g1361
  (
    n1044,
    n544
  );


  buf
  g1362
  (
    n1146,
    n168
  );


  buf
  g1363
  (
    n1265,
    n356
  );


  not
  g1364
  (
    n1766,
    n501
  );


  buf
  g1365
  (
    n1620,
    n299
  );


  buf
  g1366
  (
    n1707,
    n315
  );


  buf
  g1367
  (
    n1838,
    n515
  );


  buf
  g1368
  (
    n1543,
    n277
  );


  not
  g1369
  (
    n1129,
    n368
  );


  not
  g1370
  (
    n1905,
    n646
  );


  not
  g1371
  (
    n1499,
    n612
  );


  buf
  g1372
  (
    n2007,
    n375
  );


  buf
  g1373
  (
    n1002,
    n568
  );


  not
  g1374
  (
    n729,
    n266
  );


  buf
  g1375
  (
    n1201,
    n471
  );


  not
  g1376
  (
    n1937,
    n326
  );


  not
  g1377
  (
    n1421,
    n216
  );


  buf
  g1378
  (
    n1286,
    n511
  );


  buf
  g1379
  (
    n1602,
    n232
  );


  not
  g1380
  (
    n2069,
    n193
  );


  buf
  g1381
  (
    n774,
    n590
  );


  not
  g1382
  (
    n1253,
    n629
  );


  buf
  g1383
  (
    n1391,
    n261
  );


  buf
  g1384
  (
    n1756,
    n251
  );


  buf
  g1385
  (
    n2041,
    n661
  );


  buf
  g1386
  (
    n1893,
    n610
  );


  not
  g1387
  (
    n1331,
    n174
  );


  buf
  g1388
  (
    n1573,
    n530
  );


  not
  g1389
  (
    n1695,
    n392
  );


  not
  g1390
  (
    n1549,
    n218
  );


  not
  g1391
  (
    n2146,
    n499
  );


  not
  g1392
  (
    n2046,
    n269
  );


  buf
  g1393
  (
    n1166,
    n195
  );


  not
  g1394
  (
    n1913,
    n661
  );


  not
  g1395
  (
    n1256,
    n191
  );


  not
  g1396
  (
    n1178,
    n577
  );


  buf
  g1397
  (
    n2151,
    n270
  );


  not
  g1398
  (
    n940,
    n509
  );


  not
  g1399
  (
    n1848,
    n239
  );


  not
  g1400
  (
    n1634,
    n312
  );


  not
  g1401
  (
    n712,
    n359
  );


  not
  g1402
  (
    n1883,
    n530
  );


  not
  g1403
  (
    n1521,
    n275
  );


  not
  g1404
  (
    n1527,
    n468
  );


  buf
  g1405
  (
    n730,
    n254
  );


  buf
  g1406
  (
    n1686,
    n550
  );


  not
  g1407
  (
    n1520,
    n368
  );


  buf
  g1408
  (
    KeyWire_0_0,
    n489
  );


  not
  g1409
  (
    n1790,
    n324
  );


  not
  g1410
  (
    n1715,
    n523
  );


  not
  g1411
  (
    n1581,
    n283
  );


  not
  g1412
  (
    n941,
    n535
  );


  not
  g1413
  (
    n853,
    n466
  );


  buf
  g1414
  (
    n2001,
    n367
  );


  buf
  g1415
  (
    n886,
    n457
  );


  not
  g1416
  (
    n1011,
    n178
  );


  not
  g1417
  (
    n1188,
    n245
  );


  not
  g1418
  (
    n1972,
    n299
  );


  buf
  g1419
  (
    n1328,
    n199
  );


  buf
  g1420
  (
    n1492,
    n335
  );


  not
  g1421
  (
    n1635,
    n217
  );


  buf
  g1422
  (
    n1619,
    n296
  );


  not
  g1423
  (
    n990,
    n344
  );


  buf
  g1424
  (
    n1722,
    n487
  );


  not
  g1425
  (
    n1643,
    n367
  );


  buf
  g1426
  (
    n2161,
    n418
  );


  buf
  g1427
  (
    n2008,
    n441
  );


  not
  g1428
  (
    n1728,
    n221
  );


  buf
  g1429
  (
    n1362,
    n283
  );


  buf
  g1430
  (
    n978,
    n377
  );


  buf
  g1431
  (
    KeyWire_0_44,
    n533
  );


  not
  g1432
  (
    n1603,
    n263
  );


  buf
  g1433
  (
    n1234,
    n655
  );


  not
  g1434
  (
    n1746,
    n615
  );


  not
  g1435
  (
    n1950,
    n161
  );


  not
  g1436
  (
    n1646,
    n281
  );


  buf
  g1437
  (
    n902,
    n497
  );


  buf
  g1438
  (
    n744,
    n516
  );


  not
  g1439
  (
    n1181,
    n539
  );


  buf
  g1440
  (
    n796,
    n284
  );


  buf
  g1441
  (
    n1929,
    n625
  );


  buf
  g1442
  (
    n673,
    n477
  );


  buf
  g1443
  (
    n2123,
    n366
  );


  not
  g1444
  (
    n2131,
    n650
  );


  buf
  g1445
  (
    n879,
    n235
  );


  buf
  g1446
  (
    n1768,
    n336
  );


  buf
  g1447
  (
    n1028,
    n281
  );


  not
  g1448
  (
    n1534,
    n569
  );


  not
  g1449
  (
    n1433,
    n582
  );


  buf
  g1450
  (
    KeyWire_0_10,
    n276
  );


  not
  g1451
  (
    n1161,
    n320
  );


  not
  g1452
  (
    n1503,
    n351
  );


  buf
  g1453
  (
    n1158,
    n491
  );


  not
  g1454
  (
    n1584,
    n271
  );


  buf
  g1455
  (
    n1121,
    n220
  );


  not
  g1456
  (
    n2058,
    n589
  );


  not
  g1457
  (
    n909,
    n531
  );


  not
  g1458
  (
    n1712,
    n549
  );


  buf
  g1459
  (
    n1986,
    n225
  );


  buf
  g1460
  (
    n1583,
    n425
  );


  buf
  g1461
  (
    n1621,
    n512
  );


  buf
  g1462
  (
    n727,
    n208
  );


  buf
  g1463
  (
    n1478,
    n513
  );


  not
  g1464
  (
    n1194,
    n415
  );


  not
  g1465
  (
    n1806,
    n183
  );


  not
  g1466
  (
    n1898,
    n537
  );


  buf
  g1467
  (
    n1458,
    n467
  );


  not
  g1468
  (
    n684,
    n199
  );


  buf
  g1469
  (
    n1037,
    n503
  );


  buf
  g1470
  (
    n1588,
    n222
  );


  not
  g1471
  (
    KeyWire_0_43,
    n177
  );


  not
  g1472
  (
    n914,
    n364
  );


  buf
  g1473
  (
    n1466,
    n282
  );


  buf
  g1474
  (
    n1046,
    n501
  );


  not
  g1475
  (
    n1203,
    n323
  );


  buf
  g1476
  (
    n1691,
    n473
  );


  buf
  g1477
  (
    n741,
    n581
  );


  buf
  g1478
  (
    n1567,
    n409
  );


  not
  g1479
  (
    n1533,
    n380
  );


  buf
  g1480
  (
    n878,
    n408
  );


  buf
  g1481
  (
    n735,
    n345
  );


  buf
  g1482
  (
    n860,
    n202
  );


  not
  g1483
  (
    n937,
    n366
  );


  buf
  g1484
  (
    n1757,
    n504
  );


  not
  g1485
  (
    n1487,
    n669
  );


  not
  g1486
  (
    n1586,
    n515
  );


  not
  g1487
  (
    n1943,
    n480
  );


  not
  g1488
  (
    n1254,
    n291
  );


  not
  g1489
  (
    n1809,
    n520
  );


  buf
  g1490
  (
    n1518,
    n450
  );


  buf
  g1491
  (
    n1180,
    n501
  );


  not
  g1492
  (
    n1058,
    n237
  );


  not
  g1493
  (
    n798,
    n430
  );


  buf
  g1494
  (
    n1795,
    n624
  );


  not
  g1495
  (
    n1651,
    n528
  );


  buf
  g1496
  (
    n746,
    n407
  );


  not
  g1497
  (
    n819,
    n358
  );


  not
  g1498
  (
    n1025,
    n436
  );


  buf
  g1499
  (
    n965,
    n651
  );


  not
  g1500
  (
    n1801,
    n209
  );


  buf
  g1501
  (
    KeyWire_0_52,
    n232
  );


  not
  g1502
  (
    n2006,
    n600
  );


  buf
  g1503
  (
    n2039,
    n423
  );


  buf
  g1504
  (
    n1719,
    n385
  );


  buf
  g1505
  (
    n987,
    n277
  );


  not
  g1506
  (
    n1236,
    n288
  );


  not
  g1507
  (
    n1157,
    n203
  );


  buf
  g1508
  (
    n1811,
    n426
  );


  buf
  g1509
  (
    n1047,
    n399
  );


  not
  g1510
  (
    n1073,
    n196
  );


  not
  g1511
  (
    KeyWire_0_32,
    n370
  );


  not
  g1512
  (
    n1264,
    n439
  );


  buf
  g1513
  (
    n2038,
    n422
  );


  buf
  g1514
  (
    n761,
    n624
  );


  not
  g1515
  (
    n957,
    n174
  );


  buf
  g1516
  (
    n1854,
    n229
  );


  not
  g1517
  (
    n788,
    n506
  );


  buf
  g1518
  (
    n2010,
    n323
  );


  buf
  g1519
  (
    n833,
    n602
  );


  not
  g1520
  (
    n1131,
    n554
  );


  not
  g1521
  (
    n1516,
    n661
  );


  buf
  g1522
  (
    n2148,
    n561
  );


  not
  g1523
  (
    n1364,
    n524
  );


  buf
  g1524
  (
    n1948,
    n249
  );


  not
  g1525
  (
    n1260,
    n196
  );


  buf
  g1526
  (
    n1829,
    n171
  );


  not
  g1527
  (
    n1545,
    n669
  );


  not
  g1528
  (
    n1697,
    n517
  );


  buf
  g1529
  (
    n742,
    n274
  );


  not
  g1530
  (
    n1358,
    n603
  );


  not
  g1531
  (
    n1279,
    n609
  );


  buf
  g1532
  (
    n858,
    n553
  );


  not
  g1533
  (
    n1149,
    n330
  );


  buf
  g1534
  (
    n1009,
    n419
  );


  not
  g1535
  (
    n948,
    n347
  );


  not
  g1536
  (
    n1385,
    n256
  );


  not
  g1537
  (
    n814,
    n184
  );


  buf
  g1538
  (
    n1593,
    n560
  );


  buf
  g1539
  (
    n1764,
    n400
  );


  buf
  g1540
  (
    n1680,
    n207
  );


  buf
  g1541
  (
    n1675,
    n389
  );


  buf
  g1542
  (
    n1252,
    n501
  );


  not
  g1543
  (
    n1938,
    n635
  );


  buf
  g1544
  (
    n2049,
    n369
  );


  buf
  g1545
  (
    n1228,
    n617
  );


  buf
  g1546
  (
    n935,
    n623
  );


  not
  g1547
  (
    n1882,
    n571
  );


  buf
  g1548
  (
    n1699,
    n599
  );


  buf
  g1549
  (
    n1917,
    n452
  );


  buf
  g1550
  (
    n1220,
    n182
  );


  not
  g1551
  (
    n1794,
    n574
  );


  not
  g1552
  (
    n1246,
    n183
  );


  not
  g1553
  (
    n1810,
    n423
  );


  buf
  g1554
  (
    n1116,
    n329
  );


  buf
  g1555
  (
    n1696,
    n446
  );


  buf
  g1556
  (
    n1352,
    n290
  );


  buf
  g1557
  (
    n1655,
    n416
  );


  not
  g1558
  (
    n1856,
    n545
  );


  buf
  g1559
  (
    n2101,
    n450
  );


  not
  g1560
  (
    n1717,
    n209
  );


  buf
  g1561
  (
    n2098,
    n178
  );


  not
  g1562
  (
    n769,
    n383
  );


  buf
  g1563
  (
    n841,
    n541
  );


  buf
  g1564
  (
    n2044,
    n490
  );


  not
  g1565
  (
    n975,
    n327
  );


  buf
  g1566
  (
    n1670,
    n258
  );


  buf
  g1567
  (
    n1805,
    n319
  );


  not
  g1568
  (
    n1219,
    n659
  );


  buf
  g1569
  (
    n1401,
    n591
  );


  buf
  g1570
  (
    n907,
    n327
  );


  buf
  g1571
  (
    n1498,
    n352
  );


  not
  g1572
  (
    n1430,
    n541
  );


  not
  g1573
  (
    n1330,
    n403
  );


  not
  g1574
  (
    n736,
    n525
  );


  not
  g1575
  (
    n1678,
    n560
  );


  not
  g1576
  (
    n2128,
    n626
  );


  buf
  g1577
  (
    n1043,
    n645
  );


  not
  g1578
  (
    n1952,
    n293
  );


  buf
  g1579
  (
    n1539,
    n229
  );


  not
  g1580
  (
    n1035,
    n412
  );


  buf
  g1581
  (
    n2012,
    n437
  );


  not
  g1582
  (
    n1387,
    n442
  );


  not
  g1583
  (
    n1849,
    n493
  );


  buf
  g1584
  (
    n1803,
    n567
  );


  not
  g1585
  (
    n1847,
    n557
  );


  buf
  g1586
  (
    n1721,
    n614
  );


  buf
  g1587
  (
    n1263,
    n565
  );


  not
  g1588
  (
    n854,
    n556
  );


  not
  g1589
  (
    n1308,
    n390
  );


  not
  g1590
  (
    n752,
    n601
  );


  buf
  g1591
  (
    n881,
    n391
  );


  not
  g1592
  (
    n1089,
    n167
  );


  buf
  g1593
  (
    n1019,
    n393
  );


  not
  g1594
  (
    n1969,
    n485
  );


  buf
  g1595
  (
    n1947,
    n349
  );


  not
  g1596
  (
    n1381,
    n585
  );


  buf
  g1597
  (
    n1090,
    n284
  );


  not
  g1598
  (
    n857,
    n308
  );


  not
  g1599
  (
    n1026,
    n225
  );


  buf
  g1600
  (
    n1629,
    n235
  );


  not
  g1601
  (
    n2026,
    n213
  );


  not
  g1602
  (
    n1742,
    n618
  );


  buf
  g1603
  (
    n1050,
    n376
  );


  not
  g1604
  (
    n2152,
    n642
  );


  buf
  g1605
  (
    n1538,
    n324
  );


  not
  g1606
  (
    n1041,
    n461
  );


  buf
  g1607
  (
    n910,
    n574
  );


  buf
  g1608
  (
    n1574,
    n292
  );


  buf
  g1609
  (
    n1377,
    n369
  );


  not
  g1610
  (
    n1546,
    n319
  );


  buf
  g1611
  (
    n1559,
    n252
  );


  not
  g1612
  (
    n1526,
    n582
  );


  buf
  g1613
  (
    n1472,
    n318
  );


  buf
  g1614
  (
    n1190,
    n229
  );


  not
  g1615
  (
    n1878,
    n527
  );


  buf
  g1616
  (
    n893,
    n478
  );


  not
  g1617
  (
    n1018,
    n212
  );


  not
  g1618
  (
    n1344,
    n262
  );


  not
  g1619
  (
    n681,
    n167
  );


  buf
  g1620
  (
    n1919,
    n168
  );


  not
  g1621
  (
    n1278,
    n337
  );


  buf
  g1622
  (
    n1155,
    n416
  );


  not
  g1623
  (
    n1663,
    n177
  );


  buf
  g1624
  (
    n1418,
    n644
  );


  buf
  g1625
  (
    n764,
    n172
  );


  buf
  g1626
  (
    n1151,
    n563
  );


  buf
  g1627
  (
    n1956,
    n476
  );


  not
  g1628
  (
    n1788,
    n300
  );


  not
  g1629
  (
    n991,
    n233
  );


  buf
  g1630
  (
    n1118,
    n315
  );


  buf
  g1631
  (
    n1198,
    n224
  );


  not
  g1632
  (
    n894,
    n278
  );


  buf
  g1633
  (
    n1537,
    n232
  );


  buf
  g1634
  (
    n1617,
    n330
  );


  not
  g1635
  (
    n1579,
    n194
  );


  not
  g1636
  (
    n1130,
    n410
  );


  buf
  g1637
  (
    n1197,
    n286
  );


  buf
  g1638
  (
    n1221,
    n516
  );


  buf
  g1639
  (
    n1506,
    n273
  );


  buf
  g1640
  (
    n1814,
    n495
  );


  not
  g1641
  (
    n1884,
    n616
  );


  not
  g1642
  (
    n1978,
    n256
  );


  buf
  g1643
  (
    n1934,
    n342
  );


  buf
  g1644
  (
    n1113,
    n542
  );


  not
  g1645
  (
    n1946,
    n598
  );


  not
  g1646
  (
    n765,
    n178
  );


  buf
  g1647
  (
    n1760,
    n169
  );


  buf
  g1648
  (
    n2124,
    n228
  );


  not
  g1649
  (
    n1515,
    n265
  );


  buf
  g1650
  (
    n822,
    n189
  );


  not
  g1651
  (
    n1096,
    n364
  );


  not
  g1652
  (
    n1280,
    n247
  );


  not
  g1653
  (
    n1817,
    n644
  );


  buf
  g1654
  (
    n1891,
    n585
  );


  not
  g1655
  (
    n869,
    n319
  );


  buf
  g1656
  (
    n700,
    n339
  );


  buf
  g1657
  (
    n2159,
    n513
  );


  buf
  g1658
  (
    n1270,
    n234
  );


  not
  g1659
  (
    n679,
    n396
  );


  buf
  g1660
  (
    n740,
    n509
  );


  buf
  g1661
  (
    n1998,
    n467
  );


  not
  g1662
  (
    n868,
    n578
  );


  not
  g1663
  (
    n2127,
    n219
  );


  not
  g1664
  (
    n864,
    n519
  );


  buf
  g1665
  (
    n695,
    n588
  );


  buf
  g1666
  (
    n1931,
    n332
  );


  buf
  g1667
  (
    n1671,
    n457
  );


  buf
  g1668
  (
    n1483,
    n300
  );


  not
  g1669
  (
    n1832,
    n522
  );


  not
  g1670
  (
    n1400,
    n498
  );


  not
  g1671
  (
    n1209,
    n218
  );


  buf
  g1672
  (
    n2037,
    n622
  );


  buf
  g1673
  (
    n1424,
    n546
  );


  buf
  g1674
  (
    n1711,
    n228
  );


  not
  g1675
  (
    n716,
    n422
  );


  buf
  g1676
  (
    n1125,
    n434
  );


  not
  g1677
  (
    n960,
    n178
  );


  not
  g1678
  (
    n2091,
    n497
  );


  not
  g1679
  (
    n1008,
    n608
  );


  buf
  g1680
  (
    n1195,
    n574
  );


  buf
  g1681
  (
    n1942,
    n634
  );


  not
  g1682
  (
    n1034,
    n317
  );


  not
  g1683
  (
    n804,
    n568
  );


  buf
  g1684
  (
    n1601,
    n496
  );


  buf
  g1685
  (
    n1606,
    n356
  );


  not
  g1686
  (
    n1359,
    n428
  );


  not
  g1687
  (
    n1314,
    n559
  );


  buf
  g1688
  (
    n916,
    n565
  );


  buf
  g1689
  (
    n1000,
    n215
  );


  not
  g1690
  (
    n1059,
    n263
  );


  not
  g1691
  (
    n955,
    n526
  );


  buf
  g1692
  (
    n1612,
    n610
  );


  not
  g1693
  (
    n1300,
    n637
  );


  not
  g1694
  (
    n1006,
    n460
  );


  buf
  g1695
  (
    n1540,
    n341
  );


  not
  g1696
  (
    n1661,
    n266
  );


  buf
  g1697
  (
    n1723,
    n543
  );


  buf
  g1698
  (
    n1555,
    n206
  );


  buf
  g1699
  (
    n2003,
    n421
  );


  buf
  g1700
  (
    n1062,
    n293
  );


  not
  g1701
  (
    n1926,
    n539
  );


  buf
  g1702
  (
    KeyWire_0_33,
    n513
  );


  not
  g1703
  (
    n874,
    n205
  );


  buf
  g1704
  (
    n1134,
    n567
  );


  not
  g1705
  (
    n1171,
    n584
  );


  buf
  g1706
  (
    n959,
    n587
  );


  not
  g1707
  (
    n1137,
    n519
  );


  not
  g1708
  (
    n1122,
    n641
  );


  not
  g1709
  (
    n1475,
    n449
  );


  not
  g1710
  (
    n2066,
    n641
  );


  not
  g1711
  (
    n1189,
    n297
  );


  buf
  g1712
  (
    n1184,
    n492
  );


  not
  g1713
  (
    n1024,
    n271
  );


  buf
  g1714
  (
    n678,
    n334
  );


  buf
  g1715
  (
    n1101,
    n643
  );


  not
  g1716
  (
    n1709,
    n601
  );


  buf
  g1717
  (
    n1301,
    n489
  );


  not
  g1718
  (
    n1575,
    n306
  );


  buf
  g1719
  (
    n810,
    n417
  );


  not
  g1720
  (
    n1080,
    n367
  );


  buf
  g1721
  (
    n1154,
    n631
  );


  buf
  g1722
  (
    n1029,
    n419
  );


  buf
  g1723
  (
    n956,
    n608
  );


  not
  g1724
  (
    n1170,
    n296
  );


  not
  g1725
  (
    n1335,
    n260
  );


  not
  g1726
  (
    n969,
    n659
  );


  not
  g1727
  (
    n1774,
    n547
  );


  buf
  g1728
  (
    n2087,
    n558
  );


  buf
  g1729
  (
    n942,
    n475
  );


  buf
  g1730
  (
    n1750,
    n607
  );


  buf
  g1731
  (
    n1569,
    n638
  );


  not
  g1732
  (
    n1497,
    n209
  );


  buf
  g1733
  (
    n1673,
    n643
  );


  not
  g1734
  (
    n870,
    n621
  );


  buf
  g1735
  (
    n863,
    n262
  );


  not
  g1736
  (
    n1656,
    n168
  );


  buf
  g1737
  (
    n693,
    n459
  );


  not
  g1738
  (
    n692,
    n664
  );


  not
  g1739
  (
    n1959,
    n387
  );


  not
  g1740
  (
    n1953,
    n363
  );


  not
  g1741
  (
    n1895,
    n493
  );


  buf
  g1742
  (
    n1223,
    n631
  );


  not
  g1743
  (
    n1935,
    n633
  );


  buf
  g1744
  (
    n720,
    n643
  );


  buf
  g1745
  (
    n1269,
    n265
  );


  buf
  g1746
  (
    n1480,
    n480
  );


  buf
  g1747
  (
    n1153,
    n169
  );


  not
  g1748
  (
    n1099,
    n355
  );


  buf
  g1749
  (
    n1718,
    n204
  );


  buf
  g1750
  (
    n1639,
    n454
  );


  buf
  g1751
  (
    n1881,
    n411
  );


  not
  g1752
  (
    n1737,
    n499
  );


  not
  g1753
  (
    n1288,
    n301
  );


  not
  g1754
  (
    n1014,
    n210
  );


  buf
  g1755
  (
    n808,
    n470
  );


  not
  g1756
  (
    n980,
    n414
  );


  not
  g1757
  (
    n931,
    n485
  );


  not
  g1758
  (
    n1111,
    n307
  );


  not
  g1759
  (
    n1885,
    n218
  );


  not
  g1760
  (
    n1852,
    n318
  );


  not
  g1761
  (
    n1052,
    n506
  );


  not
  g1762
  (
    n1192,
    n610
  );


  not
  g1763
  (
    n1491,
    n524
  );


  buf
  g1764
  (
    n1901,
    n380
  );


  not
  g1765
  (
    n1282,
    n403
  );


  buf
  g1766
  (
    n1048,
    n284
  );


  buf
  g1767
  (
    n1383,
    n272
  );


  buf
  g1768
  (
    n1578,
    n550
  );


  buf
  g1769
  (
    n1242,
    n208
  );


  buf
  g1770
  (
    n1143,
    n648
  );


  not
  g1771
  (
    n1755,
    n484
  );


  not
  g1772
  (
    n773,
    n324
  );


  not
  g1773
  (
    n1389,
    n330
  );


  not
  g1774
  (
    n1955,
    n582
  );


  buf
  g1775
  (
    n1964,
    n481
  );


  buf
  g1776
  (
    n1186,
    n254
  );


  buf
  g1777
  (
    n1485,
    n381
  );


  buf
  g1778
  (
    n1078,
    n185
  );


  buf
  g1779
  (
    n970,
    n361
  );


  not
  g1780
  (
    n2052,
    n522
  );


  buf
  g1781
  (
    n973,
    n465
  );


  not
  g1782
  (
    n2110,
    n478
  );


  buf
  g1783
  (
    n946,
    n468
  );


  buf
  g1784
  (
    n1191,
    n430
  );


  not
  g1785
  (
    n892,
    n479
  );


  not
  g1786
  (
    n1725,
    n406
  );


  buf
  g1787
  (
    n1490,
    n491
  );


  not
  g1788
  (
    n1071,
    n231
  );


  not
  g1789
  (
    n1196,
    n250
  );


  buf
  g1790
  (
    n1665,
    n292
  );


  not
  g1791
  (
    n1494,
    n181
  );


  not
  g1792
  (
    n2153,
    n585
  );


  buf
  g1793
  (
    n1193,
    n667
  );


  buf
  g1794
  (
    n1214,
    n300
  );


  buf
  g1795
  (
    KeyWire_0_7,
    n180
  );


  not
  g1796
  (
    n1826,
    n358
  );


  not
  g1797
  (
    n1896,
    n593
  );


  buf
  g1798
  (
    n1159,
    n200
  );


  buf
  g1799
  (
    n1970,
    n195
  );


  buf
  g1800
  (
    n676,
    n474
  );


  not
  g1801
  (
    n707,
    n304
  );


  not
  g1802
  (
    n1513,
    n444
  );


  buf
  g1803
  (
    n1163,
    n286
  );


  not
  g1804
  (
    n981,
    n405
  );


  buf
  g1805
  (
    n1683,
    n310
  );


  buf
  g1806
  (
    n2138,
    n365
  );


  buf
  g1807
  (
    n1841,
    n234
  );


  not
  g1808
  (
    n834,
    n455
  );


  buf
  g1809
  (
    n1319,
    n548
  );


  not
  g1810
  (
    n927,
    n429
  );


  not
  g1811
  (
    n1916,
    n236
  );


  buf
  g1812
  (
    n1173,
    n652
  );


  buf
  g1813
  (
    n1749,
    n405
  );


  buf
  g1814
  (
    n1285,
    n545
  );


  buf
  g1815
  (
    n1845,
    n591
  );


  buf
  g1816
  (
    n703,
    n448
  );


  buf
  g1817
  (
    n1275,
    n222
  );


  buf
  g1818
  (
    n1250,
    n447
  );


  not
  g1819
  (
    n2018,
    n201
  );


  not
  g1820
  (
    n1426,
    n386
  );


  buf
  g1821
  (
    n743,
    n236
  );


  buf
  g1822
  (
    n1261,
    n538
  );


  not
  g1823
  (
    n2024,
    n290
  );


  not
  g1824
  (
    n1297,
    n378
  );


  not
  g1825
  (
    n1636,
    n211
  );


  not
  g1826
  (
    n1097,
    n454
  );


  buf
  g1827
  (
    KeyWire_0_30,
    n226
  );


  buf
  g1828
  (
    n1785,
    n476
  );


  not
  g1829
  (
    n687,
    n452
  );


  not
  g1830
  (
    n1135,
    n250
  );


  not
  g1831
  (
    n1370,
    n646
  );


  buf
  g1832
  (
    n1376,
    n235
  );


  buf
  g1833
  (
    n1334,
    n331
  );


  buf
  g1834
  (
    n1831,
    n584
  );


  buf
  g1835
  (
    n1212,
    n560
  );


  buf
  g1836
  (
    n1103,
    n607
  );


  not
  g1837
  (
    n1778,
    n536
  );


  not
  g1838
  (
    n866,
    n174
  );


  buf
  g1839
  (
    n1453,
    n299
  );


  not
  g1840
  (
    n1262,
    n255
  );


  buf
  g1841
  (
    n753,
    n462
  );


  buf
  g1842
  (
    n1700,
    n552
  );


  not
  g1843
  (
    n2005,
    n424
  );


  not
  g1844
  (
    n1107,
    n540
  );


  buf
  g1845
  (
    n1132,
    n566
  );


  not
  g1846
  (
    n1321,
    n187
  );


  buf
  g1847
  (
    n1437,
    n166
  );


  buf
  g1848
  (
    n989,
    n252
  );


  buf
  g1849
  (
    n897,
    n502
  );


  buf
  g1850
  (
    n1455,
    n164
  );


  buf
  g1851
  (
    n2062,
    n174
  );


  not
  g1852
  (
    n1177,
    n657
  );


  buf
  g1853
  (
    n1604,
    n627
  );


  not
  g1854
  (
    n1105,
    n254
  );


  buf
  g1855
  (
    n701,
    n267
  );


  buf
  g1856
  (
    n1532,
    n637
  );


  buf
  g1857
  (
    n1287,
    n552
  );


  buf
  g1858
  (
    n1991,
    n436
  );


  buf
  g1859
  (
    n1822,
    n318
  );


  not
  g1860
  (
    n1807,
    n259
  );


  not
  g1861
  (
    n1679,
    n611
  );


  not
  g1862
  (
    n2102,
    n200
  );


  not
  g1863
  (
    n979,
    n447
  );


  buf
  g1864
  (
    n2125,
    n225
  );


  buf
  g1865
  (
    n1020,
    n354
  );


  not
  g1866
  (
    n1703,
    n385
  );


  buf
  g1867
  (
    n2065,
    n528
  );


  not
  g1868
  (
    n711,
    n391
  );


  buf
  g1869
  (
    n996,
    n598
  );


  buf
  g1870
  (
    n1347,
    n188
  );


  not
  g1871
  (
    n806,
    n290
  );


  buf
  g1872
  (
    n1562,
    n227
  );


  buf
  g1873
  (
    n1765,
    n544
  );


  not
  g1874
  (
    n699,
    n326
  );


  buf
  g1875
  (
    n1987,
    n223
  );


  buf
  g1876
  (
    n1980,
    n666
  );


  not
  g1877
  (
    n1975,
    n592
  );


  not
  g1878
  (
    n1229,
    n486
  );


  not
  g1879
  (
    n1104,
    n270
  );


  not
  g1880
  (
    n1759,
    n565
  );


  not
  g1881
  (
    n1302,
    n660
  );


  buf
  g1882
  (
    n728,
    n180
  );


  not
  g1883
  (
    n1967,
    n167
  );


  buf
  g1884
  (
    n1296,
    n264
  );


  buf
  g1885
  (
    n2035,
    n346
  );


  buf
  g1886
  (
    n1217,
    n230
  );


  not
  g1887
  (
    n896,
    n295
  );


  not
  g1888
  (
    n1093,
    n611
  );


  buf
  g1889
  (
    n1176,
    n537
  );


  not
  g1890
  (
    n1378,
    n561
  );


  buf
  g1891
  (
    n1996,
    n563
  );


  not
  g1892
  (
    n718,
    n336
  );


  not
  g1893
  (
    n1839,
    n586
  );


  not
  g1894
  (
    n2130,
    n184
  );


  buf
  g1895
  (
    n1435,
    n298
  );


  buf
  g1896
  (
    n1365,
    n259
  );


  not
  g1897
  (
    n1830,
    n456
  );


  buf
  g1898
  (
    n1434,
    n316
  );


  not
  g1899
  (
    n1298,
    n374
  );


  not
  g1900
  (
    KeyWire_0_17,
    n256
  );


  not
  g1901
  (
    n715,
    n437
  );


  buf
  g1902
  (
    n2093,
    n372
  );


  not
  g1903
  (
    n837,
    n564
  );


  buf
  g1904
  (
    n1667,
    n670
  );


  buf
  g1905
  (
    n737,
    n623
  );


  buf
  g1906
  (
    n1094,
    n361
  );


  buf
  g1907
  (
    n997,
    n571
  );


  buf
  g1908
  (
    n2040,
    n566
  );


  not
  g1909
  (
    n1417,
    n634
  );


  buf
  g1910
  (
    n2132,
    n479
  );


  not
  g1911
  (
    n1077,
    n471
  );


  not
  g1912
  (
    n2109,
    n305
  );


  not
  g1913
  (
    n1800,
    n227
  );


  not
  g1914
  (
    n1589,
    n622
  );


  buf
  g1915
  (
    n710,
    n214
  );


  not
  g1916
  (
    n2150,
    n627
  );


  buf
  g1917
  (
    n821,
    n473
  );


  buf
  g1918
  (
    n815,
    n355
  );


  buf
  g1919
  (
    n1808,
    n315
  );


  not
  g1920
  (
    n794,
    n639
  );


  buf
  g1921
  (
    n1465,
    n515
  );


  buf
  g1922
  (
    n934,
    n456
  );


  buf
  g1923
  (
    n1147,
    n442
  );


  not
  g1924
  (
    n1346,
    n259
  );


  not
  g1925
  (
    n1027,
    n391
  );


  buf
  g1926
  (
    n680,
    n347
  );


  buf
  g1927
  (
    n1960,
    n384
  );


  not
  g1928
  (
    n2118,
    n651
  );


  not
  g1929
  (
    n2129,
    n423
  );


  buf
  g1930
  (
    n850,
    n338
  );


  not
  g1931
  (
    n1411,
    n671
  );


  not
  g1932
  (
    n2027,
    n482
  );


  not
  g1933
  (
    n2092,
    n162
  );


  not
  g1934
  (
    n1470,
    n317
  );


  buf
  g1935
  (
    n1642,
    n588
  );


  not
  g1936
  (
    n1886,
    n383
  );


  not
  g1937
  (
    n861,
    n620
  );


  not
  g1938
  (
    n1066,
    n192
  );


  buf
  g1939
  (
    n1551,
    n626
  );


  not
  g1940
  (
    n1944,
    n304
  );


  buf
  g1941
  (
    n1941,
    n603
  );


  buf
  g1942
  (
    n714,
    n217
  );


  buf
  g1943
  (
    n1880,
    n547
  );


  not
  g1944
  (
    n1780,
    n649
  );


  not
  g1945
  (
    n1023,
    n491
  );


  buf
  g1946
  (
    n917,
    n605
  );


  not
  g1947
  (
    n1452,
    n173
  );


  buf
  g1948
  (
    n1311,
    n590
  );


  not
  g1949
  (
    n1902,
    n612
  );


  not
  g1950
  (
    n1199,
    n639
  );


  buf
  g1951
  (
    n1653,
    n332
  );


  not
  g1952
  (
    n2073,
    n505
  );


  xnor
  g1953
  (
    n1738,
    n252,
    n207,
    n466,
    n442
  );


  nand
  g1954
  (
    n1436,
    n341,
    n487,
    n377,
    n405
  );


  nor
  g1955
  (
    n782,
    n353,
    n237,
    n246,
    n367
  );


  xor
  g1956
  (
    n1706,
    n214,
    n623,
    n362,
    n657
  );


  and
  g1957
  (
    n807,
    n381,
    n396,
    n666,
    n434
  );


  or
  g1958
  (
    n1879,
    n313,
    n397,
    n224,
    n346
  );


  and
  g1959
  (
    n1404,
    n352,
    n619,
    n583,
    n463
  );


  nor
  g1960
  (
    n1976,
    n566,
    n664,
    n454,
    n305
  );


  nand
  g1961
  (
    n1607,
    n462,
    n310,
    n274,
    n472
  );


  xor
  g1962
  (
    n890,
    n414,
    n360,
    n622,
    n330
  );


  nand
  g1963
  (
    n812,
    n477,
    n635,
    n563,
    n421
  );


  and
  g1964
  (
    n1910,
    n265,
    n483,
    n577,
    n569
  );


  xnor
  g1965
  (
    n2089,
    n514,
    n198,
    n163,
    n611
  );


  nand
  g1966
  (
    n2113,
    n592,
    n362,
    n242,
    n629
  );


  and
  g1967
  (
    n1021,
    n293,
    n243,
    n608,
    n237
  );


  xnor
  g1968
  (
    n1156,
    n572,
    n547,
    n273,
    n288
  );


  xnor
  g1969
  (
    n1140,
    n597,
    n395,
    n662,
    n534
  );


  or
  g1970
  (
    n801,
    n511,
    n527,
    n286,
    n516
  );


  nand
  g1971
  (
    n1798,
    n386,
    n315,
    n282,
    n244
  );


  or
  g1972
  (
    n1450,
    n266,
    n288,
    n488,
    n194
  );


  xor
  g1973
  (
    n803,
    n213,
    n411,
    n660,
    n558
  );


  and
  g1974
  (
    n2045,
    n667,
    n379,
    n451,
    n558
  );


  or
  g1975
  (
    n1053,
    n309,
    n461,
    n614,
    n502
  );


  nand
  g1976
  (
    n705,
    n662,
    n450,
    n325,
    n356
  );


  nand
  g1977
  (
    n802,
    n640,
    n667,
    n518,
    n584
  );


  xnor
  g1978
  (
    n771,
    n649,
    n302,
    n340,
    n192
  );


  xor
  g1979
  (
    n2019,
    n402,
    n529,
    n541,
    n456
  );


  and
  g1980
  (
    n1554,
    n576,
    n581,
    n387,
    n253
  );


  nand
  g1981
  (
    n1461,
    n551,
    n622,
    n656,
    n455
  );


  nor
  g1982
  (
    n1379,
    n427,
    n597,
    n601,
    n650
  );


  xor
  g1983
  (
    n1371,
    n415,
    n440,
    n504,
    n605
  );


  nand
  g1984
  (
    n1647,
    n635,
    n169,
    n201,
    n617
  );


  or
  g1985
  (
    n835,
    n606,
    n182,
    n278,
    n534
  );


  nor
  g1986
  (
    n1888,
    n370,
    n289,
    n170,
    n365
  );


  xor
  g1987
  (
    n1375,
    n438,
    n246,
    n449,
    n387
  );


  nand
  g1988
  (
    n2086,
    n418,
    n311,
    n392,
    n519
  );


  xor
  g1989
  (
    n1063,
    n469,
    n240,
    n646,
    n304
  );


  xor
  g1990
  (
    n1271,
    n280,
    n458,
    n636,
    n630
  );


  nand
  g1991
  (
    n2083,
    n579,
    n536,
    n373,
    n657
  );


  and
  g1992
  (
    n1874,
    n475,
    n518,
    n181,
    n434
  );


  and
  g1993
  (
    n840,
    n280,
    n313,
    n435,
    n649
  );


  xor
  g1994
  (
    n1965,
    n541,
    n570,
    n490,
    n342
  );


  nor
  g1995
  (
    n1235,
    n634,
    n340,
    n283,
    n348
  );


  or
  g1996
  (
    n1687,
    n387,
    n458,
    n525,
    n181
  );


  or
  g1997
  (
    n961,
    n325,
    n287,
    n419,
    n620
  );


  xor
  g1998
  (
    n1473,
    n294,
    n533,
    n398,
    n227
  );


  nor
  g1999
  (
    n900,
    n658,
    n580,
    n490,
    n327
  );


  nand
  g2000
  (
    n725,
    n664,
    n306,
    n469,
    n465
  );


  xnor
  g2001
  (
    n1754,
    n354,
    n455,
    n504,
    n424
  );


  nand
  g2002
  (
    n2042,
    n380,
    n416,
    n184,
    n628
  );


  nor
  g2003
  (
    n1502,
    n285,
    n621,
    n505,
    n372
  );


  and
  g2004
  (
    n1210,
    n459,
    n470,
    n186,
    n514
  );


  nor
  g2005
  (
    KeyWire_0_47,
    n446,
    n512,
    n289,
    n422
  );


  or
  g2006
  (
    n1560,
    n357,
    n503,
    n639,
    n479
  );


  or
  g2007
  (
    n759,
    n482,
    n173,
    n645,
    n593
  );


  and
  g2008
  (
    n1085,
    n483,
    n664,
    n166,
    n282
  );


  nand
  g2009
  (
    n852,
    n322,
    n257,
    n618,
    n513
  );


  or
  g2010
  (
    n1202,
    n651,
    n445,
    n230,
    n611
  );


  or
  g2011
  (
    n691,
    n421,
    n578,
    n555,
    n599
  );


  nor
  g2012
  (
    n1740,
    n248,
    n600,
    n530,
    n186
  );


  nand
  g2013
  (
    n1735,
    n596,
    n575,
    n303,
    n426
  );


  nor
  g2014
  (
    n867,
    n244,
    n211,
    n224,
    n240
  );


  xor
  g2015
  (
    n1940,
    n441,
    n536,
    n375,
    n472
  );


  nor
  g2016
  (
    n1577,
    n369,
    n567,
    n238,
    n334
  );


  and
  g2017
  (
    n2149,
    n307,
    n252,
    n561,
    n323
  );


  or
  g2018
  (
    n954,
    n576,
    n320,
    n393,
    n241
  );


  and
  g2019
  (
    n1669,
    n347,
    n215,
    n310,
    n245
  );


  or
  g2020
  (
    n1481,
    n393,
    n457,
    n645,
    n494
  );


  xnor
  g2021
  (
    n1572,
    n419,
    n549,
    n268,
    n514
  );


  and
  g2022
  (
    n738,
    n208,
    n313,
    n456,
    n659
  );


  xnor
  g2023
  (
    KeyWire_0_63,
    n188,
    n420,
    n340,
    n374
  );


  nand
  g2024
  (
    n1523,
    n292,
    n475,
    n593,
    n198
  );


  nor
  g2025
  (
    n1514,
    n540,
    n285,
    n235,
    n432
  );


  xor
  g2026
  (
    n1232,
    n642,
    n397,
    n223,
    n401
  );


  xnor
  g2027
  (
    n2084,
    n648,
    n603,
    n510,
    n539
  );


  xor
  g2028
  (
    n1127,
    n510,
    n303,
    n573,
    n621
  );


  xor
  g2029
  (
    n1995,
    n242,
    n527,
    n230,
    n183
  );


  xnor
  g2030
  (
    n1751,
    n279,
    n665,
    n172,
    n579
  );


  nand
  g2031
  (
    n1162,
    n507,
    n653,
    n465,
    n348
  );


  and
  g2032
  (
    n2135,
    n185,
    n350,
    n204,
    n477
  );


  and
  g2033
  (
    n677,
    n213,
    n436,
    n639,
    n495
  );


  and
  g2034
  (
    n962,
    n384,
    n542,
    n540,
    n400
  );


  xor
  g2035
  (
    n1787,
    n163,
    n526,
    n288,
    n569
  );


  nor
  g2036
  (
    n1632,
    n417,
    n565,
    n218,
    n360
  );


  nor
  g2037
  (
    n1366,
    n668,
    n564,
    n238,
    n591
  );


  or
  g2038
  (
    n2100,
    n176,
    n510,
    n471,
    n190
  );


  xnor
  g2039
  (
    n2155,
    n308,
    n518,
    n243,
    n546
  );


  nand
  g2040
  (
    n811,
    n322,
    n440,
    n308,
    n413
  );


  or
  g2041
  (
    n920,
    n163,
    n568,
    n644,
    n668
  );


  or
  g2042
  (
    n1100,
    n643,
    n434,
    n353,
    n236
  );


  nor
  g2043
  (
    n1323,
    n274,
    n398,
    n212,
    n572
  );


  and
  g2044
  (
    n952,
    n294,
    n349,
    n661,
    n598
  );


  or
  g2045
  (
    n1974,
    n171,
    n378,
    n655,
    n308
  );


  or
  g2046
  (
    n1846,
    n228,
    n353,
    n358,
    n577
  );


  and
  g2047
  (
    n702,
    n612,
    n535,
    n429,
    n262
  );


  xor
  g2048
  (
    n1408,
    n202,
    n326,
    n197,
    n503
  );


  xnor
  g2049
  (
    n1325,
    n480,
    n411,
    n561,
    n211
  );


  nor
  g2050
  (
    n1550,
    n630,
    n219,
    n578,
    n620
  );


  and
  g2051
  (
    n1051,
    n326,
    n372,
    n571,
    n353
  );


  nand
  g2052
  (
    KeyWire_0_40,
    n481,
    n220,
    n264,
    n281
  );


  or
  g2053
  (
    n1042,
    n263,
    n337,
    n360,
    n216
  );


  nand
  g2054
  (
    n763,
    n195,
    n365,
    n461,
    n349
  );


  and
  g2055
  (
    n1763,
    n164,
    n647,
    n528,
    n547
  );


  or
  g2056
  (
    n1820,
    n277,
    n323,
    n573,
    n542
  );


  and
  g2057
  (
    n1517,
    n275,
    n340,
    n215,
    n366
  );


  or
  g2058
  (
    n1582,
    n352,
    n444,
    n320,
    n357
  );


  nand
  g2059
  (
    n1624,
    n220,
    n484,
    n453,
    n388
  );


  or
  g2060
  (
    n1414,
    n493,
    n325,
    n383,
    n647
  );


  xor
  g2061
  (
    n1762,
    n371,
    n363,
    n582,
    n356
  );


  xnor
  g2062
  (
    n1614,
    n648,
    n562,
    n603,
    n248
  );


  and
  g2063
  (
    n1835,
    n467,
    n423,
    n234,
    n595
  );


  or
  g2064
  (
    KeyWire_0_39,
    n165,
    n465,
    n461,
    n215
  );


  xnor
  g2065
  (
    n1345,
    n350,
    n468,
    n251,
    n374
  );


  xor
  g2066
  (
    n731,
    n355,
    n354,
    n400,
    n654
  );


  nor
  g2067
  (
    n1776,
    n625,
    n435,
    n597,
    n420
  );


  and
  g2068
  (
    n1422,
    n272,
    n632,
    n335,
    n433
  );


  or
  g2069
  (
    n780,
    n555,
    n507,
    n337,
    n524
  );


  nand
  g2070
  (
    n1858,
    n322,
    n637,
    n399,
    n245
  );


  nor
  g2071
  (
    n793,
    n255,
    n314,
    n258,
    n544
  );


  nand
  g2072
  (
    n1690,
    n259,
    n203,
    n388,
    n292
  );


  xor
  g2073
  (
    n1226,
    n438,
    n331,
    n357,
    n650
  );


  xnor
  g2074
  (
    n943,
    n490,
    n311,
    n180,
    n207
  );


  or
  g2075
  (
    n2051,
    n334,
    n303,
    n496,
    n553
  );


  xor
  g2076
  (
    n1141,
    n532,
    n398,
    n253,
    n406
  );


  xor
  g2077
  (
    n1168,
    n209,
    n551,
    n553,
    n472
  );


  nor
  g2078
  (
    n923,
    n523,
    n389,
    n586,
    n342
  );


  or
  g2079
  (
    n1850,
    n179,
    n279,
    n185,
    n224
  );


  xor
  g2080
  (
    KeyWire_0_58,
    n459,
    n627,
    n260,
    n265
  );


  or
  g2081
  (
    n1561,
    n458,
    n443,
    n374,
    n344
  );


  or
  g2082
  (
    n930,
    n293,
    n648,
    n192,
    n451
  );


  nand
  g2083
  (
    n1423,
    n451,
    n193,
    n338,
    n182
  );


  nor
  g2084
  (
    n697,
    n564,
    n492,
    n591,
    n314
  );


  or
  g2085
  (
    n1900,
    n492,
    n517,
    n552,
    n445
  );


  nand
  g2086
  (
    n1985,
    n538,
    n500,
    n346,
    n414
  );


  xnor
  g2087
  (
    n1866,
    n670,
    n202,
    n628,
    n438
  );


  nor
  g2088
  (
    n1531,
    n342,
    n498,
    n641,
    n537
  );


  and
  g2089
  (
    n1924,
    n640,
    n532,
    n301,
    n543
  );


  xor
  g2090
  (
    n1060,
    n579,
    n557,
    n474,
    n267
  );


  nor
  g2091
  (
    n1045,
    n408,
    n579,
    n271,
    n552
  );


  nand
  g2092
  (
    n2119,
    n578,
    n205,
    n464,
    n599
  );


  xnor
  g2093
  (
    n1128,
    n420,
    n273,
    n514,
    n666
  );


  xnor
  g2094
  (
    n672,
    n521,
    n517,
    n379,
    n381
  );


  nor
  g2095
  (
    n932,
    n328,
    n548,
    n404,
    n386
  );


  xor
  g2096
  (
    n1813,
    n447,
    n349,
    n183,
    n533
  );


  nor
  g2097
  (
    n1003,
    n499,
    n247,
    n176,
    n489
  );


  xor
  g2098
  (
    n1949,
    n321,
    n290,
    n450,
    n257
  );


  and
  g2099
  (
    n1894,
    n656,
    n351,
    n470,
    n645
  );


  nand
  g2100
  (
    n1920,
    n577,
    n571,
    n473,
    n444
  );


  and
  g2101
  (
    n1030,
    n332,
    n170,
    n244,
    n187
  );


  and
  g2102
  (
    n1773,
    n415,
    n239,
    n650,
    n180
  );


  nor
  g2103
  (
    n831,
    n339,
    n653,
    n604,
    n666
  );


  or
  g2104
  (
    n1570,
    n545,
    n268,
    n358,
    n597
  );


  xor
  g2105
  (
    n1272,
    n244,
    n474,
    n486,
    n600
  );


  xnor
  g2106
  (
    n1114,
    n223,
    n359,
    n295,
    n361
  );


  and
  g2107
  (
    n891,
    n309,
    n417,
    n376,
    n184
  );


  or
  g2108
  (
    n1863,
    n226,
    n194,
    n654,
    n628
  );


  xor
  g2109
  (
    n1067,
    n526,
    n417,
    n201,
    n239
  );


  xor
  g2110
  (
    n1648,
    n615,
    n392,
    n177,
    n512
  );


  nor
  g2111
  (
    n1968,
    n314,
    n344,
    n659,
    n669
  );


  xnor
  g2112
  (
    n698,
    n531,
    n210,
    n214,
    n525
  );


  xor
  g2113
  (
    n1407,
    n502,
    n362,
    n302,
    n404
  );


  nor
  g2114
  (
    n2057,
    n605,
    n327,
    n523,
    n291
  );


  xor
  g2115
  (
    n719,
    n212,
    n211,
    n506,
    n462
  );


  or
  g2116
  (
    n2097,
    n210,
    n476,
    n589,
    n573
  );


  xor
  g2117
  (
    n1660,
    n616,
    n610,
    n270,
    n636
  );


  nand
  g2118
  (
    n2126,
    n458,
    n222,
    n165,
    n280
  );


  and
  g2119
  (
    n2029,
    n189,
    n264,
    n249,
    n636
  );


  or
  g2120
  (
    n777,
    n431,
    n371,
    n280,
    n658
  );


  or
  g2121
  (
    n690,
    n569,
    n464,
    n268,
    n606
  );


  xnor
  g2122
  (
    KeyWire_0_50,
    n580,
    n390,
    n345,
    n366
  );


  nor
  g2123
  (
    n1500,
    n629,
    n572,
    n551,
    n658
  );


  or
  g2124
  (
    n689,
    n529,
    n433,
    n300,
    n548
  );


  nand
  g2125
  (
    n2099,
    n588,
    n217,
    n404,
    n272
  );


  nor
  g2126
  (
    n972,
    n612,
    n602,
    n451,
    n494
  );


  xnor
  g2127
  (
    n1954,
    n305,
    n328,
    n253,
    n546
  );


  nor
  g2128
  (
    n1493,
    n427,
    n600,
    n590,
    n281
  );


  xnor
  g2129
  (
    n732,
    n609,
    n485,
    n460,
    n299
  );


  nand
  g2130
  (
    n786,
    n529,
    n449,
    n446,
    n306
  );


  nor
  g2131
  (
    n1351,
    n267,
    n258,
    n535,
    n433
  );


  nor
  g2132
  (
    n778,
    n545,
    n447,
    n500,
    n207
  );


  and
  g2133
  (
    n1510,
    n555,
    n333,
    n170,
    n341
  );


  nor
  g2134
  (
    n1770,
    n637,
    n385,
    n671,
    n210
  );


  xnor
  g2135
  (
    n2207,
    n1220,
    n1190,
    n1441,
    n911
  );


  and
  g2136
  (
    n2503,
    n1067,
    n1447,
    n1461,
    n1473
  );


  nand
  g2137
  (
    n2468,
    n1640,
    n1587,
    n989,
    n1716
  );


  and
  g2138
  (
    n2628,
    n1490,
    n1242,
    n1559,
    n1356
  );


  nor
  g2139
  (
    n2703,
    n1350,
    n1456,
    n1207,
    n1827
  );


  xor
  g2140
  (
    n2345,
    n1338,
    n1878,
    n1420,
    n895
  );


  nor
  g2141
  (
    n2293,
    n1691,
    n1074,
    n1507,
    n1516
  );


  nand
  g2142
  (
    n2266,
    n1033,
    n1739,
    n1868,
    n729
  );


  xor
  g2143
  (
    n2457,
    n1779,
    n1221,
    n1421,
    n1753
  );


  xnor
  g2144
  (
    n2182,
    n1510,
    n1622,
    n1334,
    n724
  );


  nand
  g2145
  (
    n2411,
    n1636,
    n1800,
    n1507,
    n1395
  );


  xnor
  g2146
  (
    n2520,
    n1085,
    n1256,
    n1643,
    n1846
  );


  nand
  g2147
  (
    n2607,
    n1049,
    n1093,
    n1326,
    n1685
  );


  nor
  g2148
  (
    n2561,
    n1050,
    n780,
    n1651,
    n1061
  );


  and
  g2149
  (
    n2343,
    n1291,
    n1655,
    n1643,
    n1179
  );


  nor
  g2150
  (
    n2716,
    n1392,
    n1695,
    n1732,
    n1842
  );


  or
  g2151
  (
    n2603,
    n1758,
    n1883,
    n1605,
    n994
  );


  nor
  g2152
  (
    n2178,
    n1876,
    n1029,
    n1606,
    n1865
  );


  nor
  g2153
  (
    n2385,
    n784,
    n1870,
    n1518,
    n1301
  );


  or
  g2154
  (
    n2682,
    n1321,
    n1861,
    n1705,
    n1844
  );


  or
  g2155
  (
    n2202,
    n1849,
    n1497,
    n1311,
    n1418
  );


  nand
  g2156
  (
    n2240,
    n733,
    n984,
    n830,
    n876
  );


  nor
  g2157
  (
    n2514,
    n1233,
    n1607,
    n1650,
    n1388
  );


  nor
  g2158
  (
    n2461,
    n1553,
    n858,
    n970,
    n1929
  );


  nand
  g2159
  (
    n2495,
    n856,
    n1874,
    n1833,
    n1097
  );


  nand
  g2160
  (
    n2516,
    n1239,
    n1565,
    n1887,
    n1456
  );


  nor
  g2161
  (
    n2253,
    n1342,
    n1381,
    n1028,
    n1555
  );


  and
  g2162
  (
    n2233,
    n725,
    n1740,
    n1661,
    n1254
  );


  nand
  g2163
  (
    n2595,
    n1585,
    n1913,
    n1096,
    n1856
  );


  or
  g2164
  (
    n2307,
    n1766,
    n1147,
    n1729,
    n813
  );


  nor
  g2165
  (
    n2579,
    n1664,
    n1056,
    n1257,
    n719
  );


  nand
  g2166
  (
    n2494,
    n1901,
    n1112,
    n1888,
    n700
  );


  xnor
  g2167
  (
    n2277,
    n772,
    n689,
    n1168,
    n1072
  );


  or
  g2168
  (
    n2365,
    n1827,
    n1455,
    n1040,
    n898
  );


  xor
  g2169
  (
    n2690,
    n1441,
    n743,
    n1836,
    n839
  );


  and
  g2170
  (
    n2535,
    n1750,
    n1744,
    n756,
    n1761
  );


  or
  g2171
  (
    n2545,
    n1267,
    n889,
    n1646,
    n1124
  );


  xnor
  g2172
  (
    n2416,
    n1926,
    n703,
    n1307,
    n1272
  );


  or
  g2173
  (
    n2509,
    n1675,
    n770,
    n964,
    n1197
  );


  or
  g2174
  (
    n2356,
    n1708,
    n1584,
    n1647,
    n1414
  );


  nor
  g2175
  (
    n2212,
    n753,
    n1812,
    n991,
    n1901
  );


  nand
  g2176
  (
    n2215,
    n1206,
    n1723,
    n1757,
    n1873
  );


  nand
  g2177
  (
    n2281,
    n1026,
    n1563,
    n1076,
    n1271
  );


  or
  g2178
  (
    n2189,
    n1180,
    n861,
    n1368,
    n853
  );


  and
  g2179
  (
    n2219,
    n696,
    n1482,
    n1048,
    n1871
  );


  xor
  g2180
  (
    n2467,
    n737,
    n680,
    n1698,
    n1599
  );


  or
  g2181
  (
    n2476,
    n964,
    n1063,
    n920,
    n1357
  );


  nor
  g2182
  (
    n2501,
    n882,
    n1494,
    n1138,
    n898
  );


  or
  g2183
  (
    n2239,
    n1128,
    n1776,
    n1527,
    n1305
  );


  or
  g2184
  (
    n2632,
    n915,
    n1583,
    n1431,
    n1010
  );


  xnor
  g2185
  (
    n2705,
    n1017,
    n1155,
    n1368,
    n1748
  );


  xnor
  g2186
  (
    KeyWire_0_6,
    n1281,
    n1073,
    n939,
    n1751
  );


  xnor
  g2187
  (
    n2335,
    n1354,
    n1721,
    n1100,
    n1808
  );


  xor
  g2188
  (
    n2496,
    n1866,
    n1694,
    n1194,
    n1003
  );


  and
  g2189
  (
    n2491,
    n1439,
    n1390,
    n1183,
    n1656
  );


  and
  g2190
  (
    n2643,
    n1681,
    n1227,
    n1748,
    n1082
  );


  and
  g2191
  (
    n2729,
    n1771,
    n1225,
    n1452,
    n1726
  );


  and
  g2192
  (
    n2247,
    n1250,
    n1863,
    n1818,
    n996
  );


  and
  g2193
  (
    n2386,
    n1678,
    n1544,
    n1580,
    n1875
  );


  or
  g2194
  (
    n2500,
    n938,
    n823,
    n1370,
    n849
  );


  or
  g2195
  (
    n2342,
    n693,
    n891,
    n1911,
    n1501
  );


  and
  g2196
  (
    n2663,
    n1212,
    n1447,
    n1143,
    n1927
  );


  or
  g2197
  (
    n2480,
    n1335,
    n801,
    n1769,
    n1032
  );


  xnor
  g2198
  (
    n2572,
    n1300,
    n1334,
    n675,
    n914
  );


  nor
  g2199
  (
    n2388,
    n1749,
    n1642,
    n1156,
    n1803
  );


  and
  g2200
  (
    n2581,
    n899,
    n688,
    n1022,
    n1154
  );


  and
  g2201
  (
    n2554,
    n1062,
    n1135,
    n909,
    n1498
  );


  xnor
  g2202
  (
    n2217,
    n1360,
    n881,
    n1769,
    n1755
  );


  and
  g2203
  (
    n2534,
    n1536,
    n1919,
    n1810,
    n1309
  );


  and
  g2204
  (
    n2488,
    n1927,
    n1658,
    n1211,
    n1524
  );


  and
  g2205
  (
    n2324,
    n1073,
    n1600,
    n1094,
    n1214
  );


  and
  g2206
  (
    n2466,
    n1213,
    n759,
    n1517,
    n1036
  );


  and
  g2207
  (
    n2601,
    n1290,
    n1467,
    n1068,
    n1046
  );


  xnor
  g2208
  (
    n2400,
    n1069,
    n1332,
    n715,
    n1245
  );


  and
  g2209
  (
    n2513,
    n1538,
    n1255,
    n758,
    n1776
  );


  nand
  g2210
  (
    n2733,
    n1201,
    n933,
    n1162,
    n1616
  );


  nor
  g2211
  (
    n2325,
    n1611,
    n692,
    n1688,
    n971
  );


  or
  g2212
  (
    n2357,
    n720,
    n1796,
    n1757,
    n1400
  );


  nor
  g2213
  (
    n2506,
    n1157,
    n1072,
    n1336,
    n1194
  );


  nand
  g2214
  (
    n2186,
    n1416,
    n1787,
    n1315,
    n1716
  );


  and
  g2215
  (
    n2599,
    n1589,
    n1686,
    n1107,
    n1061
  );


  and
  g2216
  (
    n2348,
    n1581,
    n791,
    n1833,
    n1293
  );


  xnor
  g2217
  (
    n2731,
    n1427,
    n1620,
    n1184,
    n1032
  );


  and
  g2218
  (
    n2726,
    n775,
    n1105,
    n1730,
    n1262
  );


  xnor
  g2219
  (
    n2521,
    n1270,
    n1876,
    n904,
    n1785
  );


  or
  g2220
  (
    n2519,
    n1824,
    n1180,
    n1613,
    n1831
  );


  nor
  g2221
  (
    n2364,
    n1391,
    n1812,
    n1556,
    n1223
  );


  xnor
  g2222
  (
    n2683,
    n1305,
    n1390,
    n1383,
    n1163
  );


  and
  g2223
  (
    n2543,
    n1858,
    n1546,
    n829,
    n928
  );


  or
  g2224
  (
    n2449,
    n1014,
    n1567,
    n943,
    n1488
  );


  xnor
  g2225
  (
    n2575,
    n1582,
    n1303,
    n1512,
    n1735
  );


  nand
  g2226
  (
    n2228,
    n1289,
    n1098,
    n1001,
    n906
  );


  nor
  g2227
  (
    n2619,
    n1839,
    n1470,
    n799,
    n1261
  );


  xnor
  g2228
  (
    n2313,
    n1515,
    n1013,
    n986,
    n1711
  );


  nor
  g2229
  (
    n2674,
    n1464,
    n1079,
    n1299,
    n1663
  );


  nand
  g2230
  (
    n2713,
    n1896,
    n1574,
    n956,
    n1628
  );


  and
  g2231
  (
    n2314,
    n1403,
    n957,
    n1352,
    n900
  );


  or
  g2232
  (
    n2662,
    n919,
    n678,
    n1540,
    n1151
  );


  and
  g2233
  (
    KeyWire_0_23,
    n1668,
    n1840,
    n796,
    n1193
  );


  or
  g2234
  (
    n2490,
    n1551,
    n1641,
    n934,
    n1000
  );


  nor
  g2235
  (
    n2409,
    n1712,
    n894,
    n953,
    n1131
  );


  or
  g2236
  (
    n2743,
    n1905,
    n1176,
    n819,
    n815
  );


  nor
  g2237
  (
    n2340,
    n1634,
    n748,
    n1471,
    n685
  );


  xnor
  g2238
  (
    n2223,
    n1577,
    n1554,
    n1572,
    n1220
  );


  nor
  g2239
  (
    n2332,
    n1008,
    n1603,
    n1798,
    n1081
  );


  and
  g2240
  (
    n2242,
    n1468,
    n1113,
    n1754,
    n1701
  );


  and
  g2241
  (
    n2642,
    n1174,
    n942,
    n871,
    n873
  );


  and
  g2242
  (
    n2620,
    n790,
    n935,
    n1721,
    n1428
  );


  or
  g2243
  (
    n2611,
    n1672,
    n1600,
    n1185,
    n1236
  );


  xor
  g2244
  (
    n2232,
    n1837,
    n1397,
    n1138,
    n1164
  );


  or
  g2245
  (
    n2434,
    n1343,
    n1241,
    n1638,
    n903
  );


  and
  g2246
  (
    n2708,
    n1202,
    n1615,
    n892,
    n1843
  );


  nand
  g2247
  (
    n2511,
    n1171,
    n1638,
    n1133,
    n884
  );


  nor
  g2248
  (
    n2608,
    n1885,
    n927,
    n1337,
    n1434
  );


  or
  g2249
  (
    KeyWire_0_3,
    n1500,
    n765,
    n1276,
    n1230
  );


  nand
  g2250
  (
    n2594,
    n1449,
    n766,
    n1267,
    n988
  );


  or
  g2251
  (
    n2195,
    n1074,
    n1756,
    n1400,
    n807
  );


  xor
  g2252
  (
    n2523,
    n1653,
    n1905,
    n1367,
    n1075
  );


  nor
  g2253
  (
    n2586,
    n1534,
    n1450,
    n1497,
    n1426
  );


  and
  g2254
  (
    n2531,
    n1777,
    n1202,
    n1783,
    n1668
  );


  xor
  g2255
  (
    n2290,
    n691,
    n1584,
    n1188,
    n1532
  );


  or
  g2256
  (
    n2359,
    n1604,
    n1118,
    n1692,
    n1304
  );


  or
  g2257
  (
    n2471,
    n1792,
    n1453,
    n1801,
    n998
  );


  nor
  g2258
  (
    n2261,
    n1624,
    n1183,
    n1353,
    n902
  );


  nor
  g2259
  (
    n2241,
    n1055,
    n1790,
    n1496,
    n1459
  );


  xor
  g2260
  (
    n2697,
    n1199,
    n1070,
    n1345,
    n1897
  );


  nand
  g2261
  (
    n2634,
    n1788,
    n1579,
    n750,
    n1389
  );


  nand
  g2262
  (
    n2486,
    n926,
    n1355,
    n1733,
    n954
  );


  or
  g2263
  (
    n2688,
    n1190,
    n912,
    n901,
    n1423
  );


  nor
  g2264
  (
    n2270,
    n1834,
    n1119,
    n1256,
    n916
  );


  nand
  g2265
  (
    n2463,
    n1696,
    n1411,
    n1004,
    n930
  );


  or
  g2266
  (
    n2537,
    n1091,
    n1454,
    n751,
    n951
  );


  xnor
  g2267
  (
    n2473,
    n1719,
    n1528,
    n1777,
    n1333
  );


  nand
  g2268
  (
    n2533,
    n1434,
    n1921,
    n1793,
    n1140
  );


  nor
  g2269
  (
    n2738,
    n1234,
    n1505,
    n1406,
    n1438
  );


  nand
  g2270
  (
    n2483,
    n1903,
    n1107,
    n1730,
    n1666
  );


  and
  g2271
  (
    n2251,
    n1853,
    n1181,
    n1173,
    n930
  );


  xnor
  g2272
  (
    n2263,
    n1868,
    n1802,
    n1872,
    n1101
  );


  nand
  g2273
  (
    n2742,
    n1187,
    n1113,
    n903,
    n1636
  );


  or
  g2274
  (
    n2374,
    n937,
    n1744,
    n1075,
    n1698
  );


  xor
  g2275
  (
    n2191,
    n929,
    n1650,
    n959,
    n883
  );


  and
  g2276
  (
    n2464,
    n1182,
    n1060,
    n944,
    n1265
  );


  and
  g2277
  (
    n2724,
    n1756,
    n1741,
    n1502,
    n1595
  );


  nor
  g2278
  (
    n2727,
    n1570,
    n1153,
    n1049,
    n1859
  );


  nor
  g2279
  (
    n2320,
    n975,
    n1701,
    n1347,
    n1817
  );


  nand
  g2280
  (
    n2423,
    n1114,
    n1619,
    n1141,
    n1023
  );


  nand
  g2281
  (
    n2508,
    n1687,
    n1213,
    n1566,
    n1217
  );


  xnor
  g2282
  (
    n2719,
    n911,
    n1626,
    n1348,
    n687
  );


  or
  g2283
  (
    KeyWire_0_35,
    n1376,
    n1723,
    n1175,
    n1520
  );


  or
  g2284
  (
    n2275,
    n710,
    n1619,
    n924,
    n1116
  );


  nand
  g2285
  (
    n2709,
    n1492,
    n1851,
    n913,
    n1919
  );


  and
  g2286
  (
    n2585,
    n962,
    n1709,
    n1578,
    n1416
  );


  nor
  g2287
  (
    n2677,
    n1768,
    n1200,
    n1102,
    n1084
  );


  and
  g2288
  (
    n2437,
    n1057,
    n1093,
    n1811,
    n1733
  );


  nor
  g2289
  (
    n2640,
    n1676,
    n1795,
    n1423,
    n1747
  );


  and
  g2290
  (
    n2369,
    n1381,
    n1487,
    n1593,
    n1151
  );


  and
  g2291
  (
    n2265,
    n1759,
    n1419,
    n1504,
    n673
  );


  xnor
  g2292
  (
    n2484,
    n1737,
    n1725,
    n1665,
    n1850
  );


  and
  g2293
  (
    n2334,
    n810,
    n922,
    n1294,
    n1667
  );


  nor
  g2294
  (
    n2499,
    n1345,
    n1399,
    n968,
    n1264
  );


  xnor
  g2295
  (
    n2502,
    n763,
    n1637,
    n1519,
    n682
  );


  xnor
  g2296
  (
    n2451,
    n1370,
    n1286,
    n1011,
    n1278
  );


  and
  g2297
  (
    n2197,
    n1627,
    n771,
    n1099,
    n1064
  );


  nor
  g2298
  (
    n2273,
    n1435,
    n1389,
    n1019,
    n1258
  );


  nand
  g2299
  (
    n2378,
    n1654,
    n1013,
    n1911,
    n1854
  );


  and
  g2300
  (
    KeyWire_0_12,
    n1511,
    n1550,
    n1244,
    n960
  );


  nand
  g2301
  (
    n2406,
    n1822,
    n1644,
    n1797,
    n1912
  );


  xnor
  g2302
  (
    n2200,
    n1564,
    n1710,
    n1621,
    n1065
  );


  or
  g2303
  (
    n2542,
    n1677,
    n1167,
    n1541,
    n1881
  );


  nor
  g2304
  (
    n2412,
    n1552,
    n948,
    n811,
    n1458
  );


  or
  g2305
  (
    n2422,
    n958,
    n1020,
    n1204,
    n716
  );


  and
  g2306
  (
    n2597,
    n1306,
    n1465,
    n1117,
    n1128
  );


  nor
  g2307
  (
    n2699,
    n940,
    n1035,
    n795,
    n1293
  );


  nand
  g2308
  (
    n2629,
    n1781,
    n1575,
    n1618,
    n789
  );


  nand
  g2309
  (
    n2210,
    n1899,
    n1214,
    n874,
    n1720
  );


  and
  g2310
  (
    n2322,
    n1473,
    n679,
    n757,
    n1165
  );


  or
  g2311
  (
    n2211,
    n1526,
    n1566,
    n1172,
    n1727
  );


  and
  g2312
  (
    n2188,
    n1465,
    n1050,
    n929,
    n1627
  );


  xor
  g2313
  (
    n2551,
    n1608,
    n1126,
    n1308,
    n1734
  );


  xnor
  g2314
  (
    n2321,
    n865,
    n972,
    n1163,
    n1118
  );


  or
  g2315
  (
    n2673,
    n1612,
    n1532,
    n981,
    n1022
  );


  or
  g2316
  (
    n2655,
    n993,
    n1359,
    n1143,
    n992
  );


  xor
  g2317
  (
    n2527,
    n1880,
    n998,
    n1656,
    n1660
  );


  and
  g2318
  (
    n2390,
    n912,
    n747,
    n1778,
    n886
  );


  xnor
  g2319
  (
    n2518,
    n1678,
    n974,
    n1906,
    n1296
  );


  xnor
  g2320
  (
    n2544,
    n1123,
    n1610,
    n1796,
    n1405
  );


  xor
  g2321
  (
    n2671,
    n1167,
    n1377,
    n1920,
    n1845
  );


  nand
  g2322
  (
    n2613,
    n1711,
    n1433,
    n1051,
    n727
  );


  nand
  g2323
  (
    n2363,
    n1316,
    n1144,
    n1235,
    n1692
  );


  xnor
  g2324
  (
    n2237,
    n1274,
    n1646,
    n1752,
    n1444
  );


  or
  g2325
  (
    n2735,
    n1524,
    n1499,
    n1485,
    n1282
  );


  or
  g2326
  (
    n2375,
    n816,
    n740,
    n1828,
    n1739
  );


  and
  g2327
  (
    n2646,
    n1886,
    n1307,
    n1686,
    n1522
  );


  xnor
  g2328
  (
    n2627,
    n1523,
    n1031,
    n932,
    n1543
  );


  or
  g2329
  (
    n2548,
    n1374,
    n1795,
    n1396,
    n1645
  );


  nor
  g2330
  (
    n2458,
    n1448,
    n1915,
    n1044,
    n1040
  );


  xnor
  g2331
  (
    n2658,
    n1700,
    n1039,
    n1890,
    n1047
  );


  nor
  g2332
  (
    n2339,
    n1883,
    n1550,
    n1426,
    n1830
  );


  xor
  g2333
  (
    n2558,
    n1684,
    n1358,
    n1153,
    n1140
  );


  nand
  g2334
  (
    n2685,
    n1502,
    n1341,
    n1648,
    n1673
  );


  or
  g2335
  (
    n2360,
    n1682,
    n1904,
    n1683,
    n1161
  );


  nand
  g2336
  (
    n2669,
    n1586,
    n1216,
    n1884,
    n1042
  );


  xnor
  g2337
  (
    n2722,
    n1106,
    n1240,
    n1742,
    n1298
  );


  or
  g2338
  (
    n2672,
    n1697,
    n1740,
    n1110,
    n847
  );


  xor
  g2339
  (
    n2338,
    n1057,
    n1436,
    n1325,
    n1514
  );


  xor
  g2340
  (
    n2612,
    n709,
    n1258,
    n1098,
    n883
  );


  or
  g2341
  (
    n2303,
    n681,
    n1268,
    n1283,
    n1640
  );


  nor
  g2342
  (
    n2425,
    n1707,
    n1384,
    n1145,
    n1523
  );


  xnor
  g2343
  (
    n2510,
    n1869,
    n1533,
    n888,
    n1719
  );


  xor
  g2344
  (
    n2169,
    n988,
    n1366,
    n1495,
    n1404
  );


  nor
  g2345
  (
    n2700,
    n1152,
    n1763,
    n1923,
    n918
  );


  nand
  g2346
  (
    n2712,
    n966,
    n1092,
    n1297,
    n1573
  );


  and
  g2347
  (
    n2584,
    n712,
    n1443,
    n1359,
    n969
  );


  nor
  g2348
  (
    n2598,
    n1521,
    n1017,
    n1809,
    n695
  );


  and
  g2349
  (
    n2234,
    n1565,
    n1171,
    n1743,
    n1331
  );


  xor
  g2350
  (
    n2497,
    n1782,
    n1340,
    n958,
    n1204
  );


  and
  g2351
  (
    n2282,
    n1383,
    n1841,
    n1925,
    n1736
  );


  and
  g2352
  (
    n2556,
    n1178,
    n1251,
    n1462,
    n1682
  );


  nand
  g2353
  (
    n2730,
    n1148,
    n1433,
    n1580,
    n1902
  );


  or
  g2354
  (
    n2564,
    n1314,
    n1463,
    n1225,
    n1001
  );


  xor
  g2355
  (
    n2446,
    n1015,
    n1666,
    n1382,
    n1509
  );


  nand
  g2356
  (
    n2291,
    n1271,
    n936,
    n1534,
    n1326
  );


  and
  g2357
  (
    n2465,
    n923,
    n1884,
    n1703,
    n1208
  );


  xor
  g2358
  (
    n2689,
    n1048,
    n1380,
    n1484,
    n741
  );


  xnor
  g2359
  (
    n2659,
    n1688,
    n674,
    n940,
    n981
  );


  xnor
  g2360
  (
    n2350,
    n802,
    n1690,
    n1870,
    n982
  );


  nor
  g2361
  (
    n2260,
    n1229,
    n985,
    n1800,
    n1615
  );


  and
  g2362
  (
    n2589,
    n843,
    n1864,
    n1891,
    n1437
  );


  xnor
  g2363
  (
    n2373,
    n945,
    n1860,
    n1839,
    n1546
  );


  nor
  g2364
  (
    n2331,
    n1218,
    n1525,
    n960,
    n1555
  );


  xor
  g2365
  (
    n2230,
    n1705,
    n1517,
    n1481,
    n735
  );


  nand
  g2366
  (
    n2653,
    n1596,
    n1309,
    n1819,
    n1018
  );


  nand
  g2367
  (
    n2580,
    n781,
    n938,
    n1483,
    n1614
  );


  nand
  g2368
  (
    n2204,
    n868,
    n1878,
    n1734,
    n1823
  );


  xor
  g2369
  (
    n2487,
    n1585,
    n1298,
    n711,
    n826
  );


  and
  g2370
  (
    n2590,
    n1247,
    n1422,
    n1336,
    n1133
  );


  nor
  g2371
  (
    n2298,
    n906,
    n852,
    n774,
    n1758
  );


  xnor
  g2372
  (
    n2278,
    n1055,
    n1590,
    n1877,
    n1425
  );


  xor
  g2373
  (
    n2701,
    n1228,
    n1012,
    n1867,
    n1280
  );


  xor
  g2374
  (
    n2257,
    n1205,
    n965,
    n910,
    n1691
  );


  xnor
  g2375
  (
    n2238,
    n1710,
    n1439,
    n1385,
    n1454
  );


  xor
  g2376
  (
    n2454,
    n1243,
    n1821,
    n1924,
    n1142
  );


  or
  g2377
  (
    n2617,
    n1409,
    n1030,
    n803,
    n1475
  );


  and
  g2378
  (
    n2341,
    n1630,
    n1125,
    n1086,
    n1363
  );


  and
  g2379
  (
    n2557,
    n1568,
    n900,
    n1895,
    n1713
  );


  and
  g2380
  (
    n2408,
    n1743,
    n1054,
    n1671,
    n1622
  );


  nand
  g2381
  (
    n2546,
    n1722,
    n1918,
    n1284,
    n901
  );


  nand
  g2382
  (
    n2456,
    n1303,
    n1898,
    n1016,
    n1030
  );


  nand
  g2383
  (
    n2517,
    n1373,
    n1571,
    n1629,
    n1377
  );


  or
  g2384
  (
    n2582,
    n1853,
    n1038,
    n746,
    n728
  );


  nor
  g2385
  (
    n2433,
    n1505,
    n1900,
    n1160,
    n1846
  );


  xnor
  g2386
  (
    n2498,
    n738,
    n1158,
    n970,
    n1684
  );


  xor
  g2387
  (
    n2698,
    n844,
    n825,
    n1058,
    n1568
  );


  and
  g2388
  (
    n2286,
    n1602,
    n1396,
    n1770,
    n1431
  );


  nor
  g2389
  (
    n2553,
    n1879,
    n1365,
    n1854,
    n1221
  );


  and
  g2390
  (
    n2246,
    n1764,
    n997,
    n1091,
    n996
  );


  nor
  g2391
  (
    n2184,
    n1814,
    n1011,
    n1417,
    n1144
  );


  nand
  g2392
  (
    n2256,
    n884,
    n1602,
    n723,
    n1357
  );


  and
  g2393
  (
    n2306,
    n1921,
    n1811,
    n1071,
    n1451
  );


  nand
  g2394
  (
    n2489,
    n1391,
    n1794,
    n1287,
    n1569
  );


  nand
  g2395
  (
    n2475,
    n1087,
    n1561,
    n1609,
    n1717
  );


  xnor
  g2396
  (
    n2272,
    n1674,
    n1618,
    n887,
    n1209
  );


  and
  g2397
  (
    n2606,
    n885,
    n1347,
    n925,
    n1493
  );


  nor
  g2398
  (
    n2714,
    n1549,
    n1766,
    n1026,
    n1387
  );


  and
  g2399
  (
    n2668,
    n1841,
    n965,
    n1489,
    n794
  );


  nor
  g2400
  (
    n2288,
    n1358,
    n817,
    n1567,
    n1288
  );


  or
  g2401
  (
    n2255,
    n1727,
    n1302,
    n1226,
    n890
  );


  or
  g2402
  (
    n2630,
    n1486,
    n1378,
    n1880,
    n1587
  );


  xor
  g2403
  (
    n2172,
    n1457,
    n1799,
    n1651,
    n1411
  );


  nand
  g2404
  (
    n2192,
    n1909,
    n1210,
    n1525,
    n1159
  );


  or
  g2405
  (
    n2720,
    n1393,
    n980,
    n832,
    n821
  );


  and
  g2406
  (
    n2292,
    n1560,
    n1635,
    n1102,
    n1855
  );


  or
  g2407
  (
    n2440,
    n1110,
    n1322,
    n1852,
    n818
  );


  nor
  g2408
  (
    n2644,
    n1556,
    n1319,
    n704,
    n1012
  );


  xor
  g2409
  (
    n2573,
    n833,
    n1428,
    n1860,
    n862
  );


  nand
  g2410
  (
    n2391,
    n1683,
    n1637,
    n1770,
    n1625
  );


  xnor
  g2411
  (
    n2269,
    n1005,
    n1908,
    n1675,
    n1773
  );


  xor
  g2412
  (
    n2185,
    n995,
    n1351,
    n1895,
    n1544
  );


  nand
  g2413
  (
    n2295,
    n1315,
    n1286,
    n1007,
    n979
  );


  nand
  g2414
  (
    n2604,
    n1815,
    n973,
    n1548,
    n1025
  );


  xnor
  g2415
  (
    KeyWire_0_24,
    n1531,
    n1372,
    n1674,
    n925
  );


  or
  g2416
  (
    n2648,
    n792,
    n908,
    n1669,
    n1184
  );


  and
  g2417
  (
    n2221,
    n1816,
    n1467,
    n989,
    n1591
  );


  xor
  g2418
  (
    n2702,
    n1045,
    n1625,
    n1393,
    n1761
  );


  or
  g2419
  (
    n2337,
    n1867,
    n1177,
    n1672,
    n1406
  );


  xnor
  g2420
  (
    n2300,
    n1559,
    n1623,
    n1632,
    n1247
  );


  xor
  g2421
  (
    n2168,
    n957,
    n1344,
    n677,
    n927
  );


  xnor
  g2422
  (
    n2578,
    n1408,
    n1362,
    n1327,
    n1765
  );


  and
  g2423
  (
    n2326,
    n1610,
    n1122,
    n1332,
    n736
  );


  xor
  g2424
  (
    n2530,
    n967,
    n926,
    n936,
    n1707
  );


  nor
  g2425
  (
    n2526,
    n1277,
    n1412,
    n1851,
    n1457
  );


  xnor
  g2426
  (
    n2444,
    n1275,
    n1313,
    n1297,
    n1395
  );


  and
  g2427
  (
    n2460,
    n1120,
    n1240,
    n1914,
    n1139
  );


  or
  g2428
  (
    n2279,
    n1449,
    n690,
    n977,
    n694
  );


  nand
  g2429
  (
    n2289,
    n977,
    n954,
    n1135,
    n1244
  );


  or
  g2430
  (
    n2216,
    n714,
    n944,
    n1891,
    n1440
  );


  xor
  g2431
  (
    n2243,
    n1229,
    n1892,
    n1052,
    n1269
  );


  xnor
  g2432
  (
    n2686,
    n1246,
    n1825,
    n1388,
    n1237
  );


  and
  g2433
  (
    n2213,
    n842,
    n1781,
    n885,
    n782
  );


  nand
  g2434
  (
    n2308,
    n1401,
    n1174,
    n1409,
    n1485
  );


  and
  g2435
  (
    n2354,
    n730,
    n1659,
    n1284,
    n1127
  );


  and
  g2436
  (
    n2283,
    n893,
    n1189,
    n1599,
    n1245
  );


  and
  g2437
  (
    KeyWire_0_1,
    n1767,
    n1725,
    n1592,
    n1676
  );


  nor
  g2438
  (
    n2419,
    n1222,
    n1810,
    n872,
    n992
  );


  xor
  g2439
  (
    n2417,
    n1318,
    n1915,
    n1382,
    n840
  );


  nand
  g2440
  (
    n2355,
    n1205,
    n1784,
    n722,
    n961
  );


  nor
  g2441
  (
    n2442,
    n1530,
    n971,
    n1224,
    n1772
  );


  and
  g2442
  (
    n2244,
    n896,
    n1324,
    n1312,
    n1834
  );


  xor
  g2443
  (
    n2512,
    n1474,
    n1037,
    n1459,
    n932
  );


  nor
  g2444
  (
    n2652,
    n1461,
    n972,
    n1775,
    n1019
  );


  and
  g2445
  (
    n2621,
    n1134,
    n1772,
    n1132,
    n1364
  );


  xor
  g2446
  (
    n2665,
    n1826,
    n1436,
    n1161,
    n1193
  );


  and
  g2447
  (
    n2428,
    n1603,
    n1097,
    n1096,
    n1166
  );


  or
  g2448
  (
    n2687,
    n1907,
    n1547,
    n1037,
    n914
  );


  nor
  g2449
  (
    n2194,
    n1442,
    n1488,
    n1617,
    n1006
  );


  nor
  g2450
  (
    n2171,
    n1823,
    n1480,
    n986,
    n1402
  );


  or
  g2451
  (
    n2377,
    n1552,
    n1607,
    n718,
    n1134
  );


  nor
  g2452
  (
    n2249,
    n1689,
    n951,
    n1693,
    n1299
  );


  or
  g2453
  (
    n2301,
    n1300,
    n1340,
    n1589,
    n1386
  );


  xor
  g2454
  (
    n2576,
    n1317,
    n1889,
    n1660,
    n788
  );


  xnor
  g2455
  (
    n2368,
    n1415,
    n1100,
    n1492,
    n1070
  );


  xnor
  g2456
  (
    n2276,
    n1557,
    n918,
    n760,
    n1859
  );


  and
  g2457
  (
    n2505,
    n1139,
    n1376,
    n1071,
    n1529
  );


  nor
  g2458
  (
    n2208,
    n1662,
    n1386,
    n1594,
    n1430
  );


  and
  g2459
  (
    n2274,
    n1477,
    n1338,
    n1145,
    n749
  );


  and
  g2460
  (
    n2448,
    n1664,
    n1504,
    n1196,
    n1088
  );


  and
  g2461
  (
    n2399,
    n1545,
    n945,
    n1330,
    n1415
  );


  nand
  g2462
  (
    n2236,
    n767,
    n793,
    n1541,
    n1200
  );


  nand
  g2463
  (
    n2482,
    n1747,
    n1703,
    n1192,
    n1653
  );


  nor
  g2464
  (
    n2566,
    n1264,
    n1629,
    n1168,
    n787
  );


  xnor
  g2465
  (
    n2218,
    n1548,
    n806,
    n1422,
    n1387
  );


  nand
  g2466
  (
    n2622,
    n1437,
    n1665,
    n1407,
    n1857
  );


  nor
  g2467
  (
    n2224,
    n1750,
    n1410,
    n1058,
    n1731
  );


  nor
  g2468
  (
    n2593,
    n1899,
    n917,
    n1385,
    n1738
  );


  xor
  g2469
  (
    n2173,
    n1542,
    n1106,
    n1474,
    n991
  );


  or
  g2470
  (
    n2389,
    n1080,
    n1355,
    n1706,
    n1361
  );


  xor
  g2471
  (
    n2667,
    n1900,
    n1241,
    n1188,
    n1379
  );


  nand
  g2472
  (
    n2614,
    n1374,
    n1004,
    n1369,
    n1402
  );


  and
  g2473
  (
    n2414,
    n983,
    n1179,
    n1598,
    n1087
  );


  xor
  g2474
  (
    n2392,
    n1348,
    n894,
    n1874,
    n1445
  );


  xnor
  g2475
  (
    n2455,
    n798,
    n1611,
    n961,
    n1519
  );


  xnor
  g2476
  (
    n2344,
    n785,
    n1728,
    n1122,
    n1253
  );


  and
  g2477
  (
    n2430,
    n1237,
    n1528,
    n1789,
    n1760
  );


  or
  g2478
  (
    n2431,
    n888,
    n1125,
    n1223,
    n1704
  );


  or
  g2479
  (
    n2179,
    n1913,
    n1136,
    n1199,
    n1255
  );


  or
  g2480
  (
    n2397,
    n1558,
    n1639,
    n1596,
    n1506
  );


  nand
  g2481
  (
    n2717,
    n1273,
    n1077,
    n1630,
    n1835
  );


  xor
  g2482
  (
    n2199,
    n1281,
    n1060,
    n1902,
    n1279
  );


  nand
  g2483
  (
    n2524,
    n1918,
    n1130,
    n1331,
    n1371
  );


  nand
  g2484
  (
    n2174,
    n1312,
    n1169,
    n1804,
    n1432
  );


  nand
  g2485
  (
    n2504,
    n1801,
    n1896,
    n1226,
    n838
  );


  nand
  g2486
  (
    n2311,
    n1574,
    n947,
    n812,
    n1321
  );


  or
  g2487
  (
    n2447,
    n1538,
    n1259,
    n1228,
    n1910
  );


  xor
  g2488
  (
    n2367,
    n1155,
    n1443,
    n1418,
    n1715
  );


  nor
  g2489
  (
    n2470,
    n1304,
    n1661,
    n1024,
    n1002
  );


  xor
  g2490
  (
    n2296,
    n1557,
    n1086,
    n1509,
    n1774
  );


  nand
  g2491
  (
    n2439,
    n1249,
    n985,
    n1537,
    n1814
  );


  nor
  g2492
  (
    n2227,
    n731,
    n1786,
    n1469,
    n1150
  );


  or
  g2493
  (
    n2715,
    n1018,
    n1176,
    n1708,
    n973
  );


  nor
  g2494
  (
    n2262,
    n1285,
    n1438,
    n1510,
    n1890
  );


  nand
  g2495
  (
    n2631,
    n1121,
    n1494,
    n1791,
    n1039
  );


  nor
  g2496
  (
    n2571,
    n1469,
    n1251,
    n822,
    n1886
  );


  xor
  g2497
  (
    n2459,
    n1067,
    n805,
    n1917,
    n836
  );


  or
  g2498
  (
    n2231,
    n1794,
    n1832,
    n699,
    n726
  );


  xnor
  g2499
  (
    n2387,
    n1114,
    n950,
    n1000,
    n1815
  );


  and
  g2500
  (
    n2577,
    n1289,
    n1130,
    n1657,
    n1206
  );


  xnor
  g2501
  (
    n2493,
    n1268,
    n1481,
    n1483,
    n1718
  );


  and
  g2502
  (
    n2588,
    n978,
    n1083,
    n1460,
    n1009
  );


  nor
  g2503
  (
    n2623,
    n937,
    n907,
    n1413,
    n1522
  );


  xnor
  g2504
  (
    n2383,
    n1709,
    n935,
    n1677,
    n869
  );


  nor
  g2505
  (
    n2404,
    n952,
    n1126,
    n946,
    n877
  );


  or
  g2506
  (
    n2248,
    n1824,
    n1906,
    n1838,
    n854
  );


  xor
  g2507
  (
    n2319,
    n828,
    n1080,
    n978,
    n776
  );


  and
  g2508
  (
    n2175,
    n1501,
    n1893,
    n997,
    n1864
  );


  xnor
  g2509
  (
    n2694,
    n1076,
    n1908,
    n1361,
    n1121
  );


  xnor
  g2510
  (
    n2381,
    n1690,
    n980,
    n1771,
    n1224
  );


  and
  g2511
  (
    n2707,
    n1432,
    n713,
    n892,
    n1275
  );


  nor
  g2512
  (
    n2327,
    n1215,
    n1274,
    n1111,
    n1597
  );


  nor
  g2513
  (
    n2615,
    n1349,
    n850,
    n1346,
    n1606
  );


  or
  g2514
  (
    n2299,
    n1282,
    n1455,
    n1327,
    n1263
  );


  and
  g2515
  (
    n2316,
    n1084,
    n808,
    n739,
    n1366
  );


  nor
  g2516
  (
    n2267,
    n1732,
    n1569,
    n1545,
    n1464
  );


  xor
  g2517
  (
    n2268,
    n950,
    n1380,
    n1375,
    n1591
  );


  nand
  g2518
  (
    n2725,
    n1211,
    n1490,
    n1498,
    n1046
  );


  and
  g2519
  (
    n2616,
    n983,
    n1530,
    n1453,
    n1542
  );


  xnor
  g2520
  (
    n2453,
    n1806,
    n1105,
    n1687,
    n1132
  );


  nand
  g2521
  (
    n2271,
    n1549,
    n968,
    n984,
    n1169
  );


  and
  g2522
  (
    n2462,
    n1177,
    n933,
    n1261,
    n1570
  );


  and
  g2523
  (
    n2395,
    n982,
    n993,
    n1320,
    n1503
  );


  xnor
  g2524
  (
    n2170,
    n754,
    n1576,
    n1583,
    n1478
  );


  xnor
  g2525
  (
    n2692,
    n947,
    n1590,
    n1626,
    n1573
  );


  and
  g2526
  (
    n2424,
    n1717,
    n1156,
    n1543,
    n1216
  );


  and
  g2527
  (
    n2734,
    n1273,
    n1146,
    n745,
    n1581
  );


  nor
  g2528
  (
    n2552,
    n1466,
    n1924,
    n797,
    n1446
  );


  or
  g2529
  (
    n2284,
    n1446,
    n1922,
    n1792,
    n1746
  );


  or
  g2530
  (
    n2176,
    n1742,
    n1413,
    n924,
    n1754
  );


  and
  g2531
  (
    n2402,
    n1762,
    n1533,
    n1025,
    n1137
  );


  and
  g2532
  (
    n2264,
    n1724,
    n921,
    n1344,
    n1117
  );


  or
  g2533
  (
    n2441,
    n1265,
    n1187,
    n1916,
    n1773
  );


  nand
  g2534
  (
    n2651,
    n1410,
    n1628,
    n1137,
    n1036
  );


  and
  g2535
  (
    n2618,
    n1196,
    n1028,
    n1082,
    n1491
  );


  or
  g2536
  (
    n2294,
    n890,
    n1328,
    n1601,
    n1421
  );


  xor
  g2537
  (
    n2741,
    n1015,
    n846,
    n1310,
    n824
  );


  or
  g2538
  (
    n2225,
    n1476,
    n1790,
    n1910,
    n1068
  );


  or
  g2539
  (
    n2181,
    n1219,
    n1364,
    n1238,
    n1034
  );


  xor
  g2540
  (
    n2401,
    n1535,
    n1612,
    n1077,
    n1749
  );


  or
  g2541
  (
    n2183,
    n1460,
    n1115,
    n1313,
    n1920
  );


  and
  g2542
  (
    n2650,
    n886,
    n1010,
    n1825,
    n1604
  );


  or
  g2543
  (
    n2675,
    n1805,
    n1624,
    n1427,
    n1123
  );


  nor
  g2544
  (
    KeyWire_0_48,
    n1266,
    n994,
    n1430,
    n1914
  );


  xor
  g2545
  (
    n2203,
    n1472,
    n1782,
    n1616,
    n1065
  );


  or
  g2546
  (
    n2229,
    n1041,
    n1478,
    n1806,
    n1207
  );


  xnor
  g2547
  (
    n2472,
    n1363,
    n1620,
    n1090,
    n834
  );


  nand
  g2548
  (
    n2568,
    n916,
    n1515,
    n1405,
    n1002
  );


  or
  g2549
  (
    n2600,
    n1768,
    n1407,
    n1480,
    n1679
  );


  and
  g2550
  (
    n2190,
    n1232,
    n1718,
    n899,
    n786
  );


  xor
  g2551
  (
    n2609,
    n1835,
    n708,
    n1605,
    n1903
  );


  or
  g2552
  (
    n2384,
    n1149,
    n1697,
    n1063,
    n919
  );


  nand
  g2553
  (
    n2681,
    n827,
    n1575,
    n1513,
    n1785
  );


  nand
  g2554
  (
    n2647,
    n1894,
    n1553,
    n922,
    n897
  );


  or
  g2555
  (
    n2550,
    n1491,
    n1027,
    n1866,
    n962
  );


  and
  g2556
  (
    n2235,
    n1186,
    n684,
    n1609,
    n1003
  );


  and
  g2557
  (
    n2435,
    n987,
    n923,
    n1445,
    n1172
  );


  or
  g2558
  (
    n2538,
    n1352,
    n1598,
    n864,
    n1146
  );


  xor
  g2559
  (
    n2522,
    n1203,
    n895,
    n1649,
    n1746
  );


  xor
  g2560
  (
    n2180,
    n1694,
    n1079,
    n896,
    n1219
  );


  xor
  g2561
  (
    n2222,
    n974,
    n1798,
    n1760,
    n702
  );


  xnor
  g2562
  (
    n2515,
    n762,
    n1269,
    n1311,
    n1889
  );


  xor
  g2563
  (
    n2610,
    n764,
    n1248,
    n1008,
    n1681
  );


  nand
  g2564
  (
    n2696,
    n1857,
    n1828,
    n893,
    n1633
  );


  nand
  g2565
  (
    n2684,
    n1809,
    n1817,
    n1813,
    n1078
  );


  nand
  g2566
  (
    n2418,
    n941,
    n1712,
    n1365,
    n1745
  );


  and
  g2567
  (
    n2507,
    n1043,
    n1539,
    n732,
    n1350
  );


  nand
  g2568
  (
    n2670,
    n1832,
    n1536,
    n1512,
    n1016
  );


  xor
  g2569
  (
    n2721,
    n1005,
    n1477,
    n1558,
    n1775
  );


  xor
  g2570
  (
    n2254,
    n999,
    n1527,
    n1294,
    n1847
  );


  xnor
  g2571
  (
    n2318,
    n880,
    n1862,
    n897,
    n1208
  );


  and
  g2572
  (
    n2280,
    n1826,
    n1339,
    n1252,
    n1158
  );


  and
  g2573
  (
    n2587,
    n1192,
    n1246,
    n857,
    n676
  );


  xor
  g2574
  (
    n2361,
    n1562,
    n1472,
    n1540,
    n1316
  );


  nor
  g2575
  (
    n2656,
    n1572,
    n1829,
    n1041,
    n948
  );


  nand
  g2576
  (
    n2201,
    n835,
    n683,
    n1577,
    n1341
  );


  and
  g2577
  (
    n2209,
    n1227,
    n1753,
    n1066,
    n1330
  );


  nor
  g2578
  (
    n2567,
    n1412,
    n1173,
    n1713,
    n1784
  );


  and
  g2579
  (
    n2426,
    n1054,
    n701,
    n1819,
    n1129
  );


  xnor
  g2580
  (
    n2372,
    n1818,
    n1152,
    n1329,
    n1807
  );


  nor
  g2581
  (
    n2347,
    n1793,
    n1053,
    n1526,
    n1639
  );


  nor
  g2582
  (
    n2711,
    n1259,
    n1185,
    n1652,
    n1090
  );


  xor
  g2583
  (
    n2336,
    n1218,
    n1898,
    n976,
    n1367
  );


  nor
  g2584
  (
    n2333,
    n1621,
    n1807,
    n1845,
    n1343
  );


  nor
  g2585
  (
    n2549,
    n1820,
    n1328,
    n1855,
    n1295
  );


  nor
  g2586
  (
    n2198,
    n1210,
    n1252,
    n963,
    n1877
  );


  xnor
  g2587
  (
    n2596,
    n809,
    n1803,
    n1821,
    n1059
  );


  nand
  g2588
  (
    n2639,
    n867,
    n1378,
    n1287,
    n939
  );


  xor
  g2589
  (
    n2680,
    n1508,
    n1513,
    n1243,
    n820
  );


  nor
  g2590
  (
    n2250,
    n1322,
    n1181,
    n1634,
    n1066
  );


  nor
  g2591
  (
    n2625,
    n1408,
    n1263,
    n1837,
    n1601
  );


  xor
  g2592
  (
    n2432,
    n1006,
    n1318,
    n1500,
    n1787
  );


  and
  g2593
  (
    n2706,
    n949,
    n1657,
    n1511,
    n1508
  );


  nor
  g2594
  (
    n2664,
    n1319,
    n1435,
    n1371,
    n1493
  );


  and
  g2595
  (
    n2358,
    n1928,
    n1147,
    n1759,
    n1822
  );


  nor
  g2596
  (
    n2310,
    n955,
    n1317,
    n1780,
    n1053
  );


  and
  g2597
  (
    n2559,
    n1608,
    n831,
    n1335,
    n1325
  );


  nand
  g2598
  (
    n2485,
    n1056,
    n1645,
    n1182,
    n1641
  );


  xnor
  g2599
  (
    n2704,
    n1907,
    n941,
    n1232,
    n1162
  );


  and
  g2600
  (
    n2536,
    n1131,
    n1195,
    n1238,
    n1353
  );


  xnor
  g2601
  (
    n2695,
    n1260,
    n1198,
    n1588,
    n1023
  );


  nand
  g2602
  (
    n2737,
    n934,
    n1462,
    n1875,
    n1044
  );


  xor
  g2603
  (
    n2732,
    n1021,
    n1486,
    n1253,
    n1849
  );


  nand
  g2604
  (
    n2304,
    n1164,
    n1203,
    n1197,
    n1191
  );


  nor
  g2605
  (
    n2626,
    n1279,
    n1178,
    n1394,
    n889
  );


  nor
  g2606
  (
    n2583,
    n1879,
    n969,
    n1170,
    n1654
  );


  xor
  g2607
  (
    n2477,
    n841,
    n1882,
    n1021,
    n1116
  );


  nor
  g2608
  (
    n2591,
    n1699,
    n990,
    n1671,
    n946
  );


  or
  g2609
  (
    n2259,
    n721,
    n1658,
    n1922,
    n1670
  );


  xnor
  g2610
  (
    n2693,
    n1495,
    n1052,
    n1731,
    n755
  );


  or
  g2611
  (
    n2403,
    n851,
    n1551,
    n1452,
    n1081
  );


  xnor
  g2612
  (
    n2560,
    n1916,
    n1379,
    n913,
    n1780
  );


  nor
  g2613
  (
    n2649,
    n1693,
    n1414,
    n1337,
    n1231
  );


  nor
  g2614
  (
    n2452,
    n917,
    n1593,
    n1403,
    n837
  );


  and
  g2615
  (
    n2718,
    n1642,
    n1362,
    n1234,
    n1695
  );


  and
  g2616
  (
    n2450,
    n1563,
    n717,
    n1360,
    n1516
  );


  nor
  g2617
  (
    n2479,
    n1444,
    n1115,
    n1863,
    n1149
  );


  and
  g2618
  (
    n2379,
    n975,
    n1865,
    n1451,
    n866
  );


  and
  g2619
  (
    n2723,
    n1484,
    n1617,
    n1235,
    n1425
  );


  nor
  g2620
  (
    n2206,
    n1649,
    n1829,
    n1285,
    n1373
  );


  or
  g2621
  (
    n2370,
    n1791,
    n1112,
    n769,
    n1613
  );


  and
  g2622
  (
    n2205,
    n1813,
    n1323,
    n1108,
    n1597
  );


  or
  g2623
  (
    n2226,
    n859,
    n1735,
    n1850,
    n1154
  );


  or
  g2624
  (
    n2654,
    n955,
    n1136,
    n1881,
    n1129
  );


  and
  g2625
  (
    n2362,
    n1805,
    n1339,
    n1764,
    n1064
  );


  xnor
  g2626
  (
    n2220,
    n953,
    n1333,
    n1356,
    n1272
  );


  xor
  g2627
  (
    n2635,
    n1260,
    n1292,
    n1894,
    n1848
  );


  or
  g2628
  (
    n2736,
    n773,
    n976,
    n1231,
    n1254
  );


  and
  g2629
  (
    n2532,
    n1189,
    n1506,
    n1736,
    n1767
  );


  xor
  g2630
  (
    n2258,
    n1262,
    n1236,
    n1869,
    n1397
  );


  nand
  g2631
  (
    n2371,
    n1195,
    n987,
    n1398,
    n1104
  );


  nor
  g2632
  (
    n2592,
    n1239,
    n1419,
    n1062,
    n1160
  );


  xnor
  g2633
  (
    n2315,
    n1887,
    n1230,
    n1429,
    n1514
  );


  xnor
  g2634
  (
    n2547,
    n1476,
    n1662,
    n1324,
    n1458
  );


  nand
  g2635
  (
    n2678,
    n1926,
    n1520,
    n1089,
    n1644
  );


  xor
  g2636
  (
    n2330,
    n1463,
    n1007,
    n1020,
    n1804
  );


  nand
  g2637
  (
    n2380,
    n1862,
    n1816,
    n1560,
    n879
  );


  xor
  g2638
  (
    n2445,
    n1783,
    n1450,
    n1669,
    n1897
  );


  and
  g2639
  (
    n2562,
    n1215,
    n956,
    n1280,
    n1586
  );


  and
  g2640
  (
    n2287,
    n1861,
    n1840,
    n1831,
    n952
  );


  or
  g2641
  (
    n2474,
    n1024,
    n1420,
    n1537,
    n1799
  );


  nor
  g2642
  (
    n2676,
    n1375,
    n1045,
    n1470,
    n1033
  );


  xor
  g2643
  (
    n2196,
    n1404,
    n1296,
    n686,
    n1696
  );


  xor
  g2644
  (
    n2478,
    n1475,
    n1892,
    n779,
    n1529
  );


  or
  g2645
  (
    n2602,
    n1124,
    n1872,
    n1858,
    n1094
  );


  or
  g2646
  (
    n2396,
    n1424,
    n1372,
    n1741,
    n1035
  );


  xor
  g2647
  (
    n2187,
    n777,
    n1078,
    n1346,
    n1043
  );


  nand
  g2648
  (
    n2528,
    n1165,
    n959,
    n1085,
    n1290
  );


  nand
  g2649
  (
    n2541,
    n707,
    n1830,
    n1471,
    n1401
  );


  or
  g2650
  (
    n2302,
    n1250,
    n1487,
    n1201,
    n1852
  );


  and
  g2651
  (
    n2177,
    n1270,
    n1917,
    n1083,
    n1301
  );


  xnor
  g2652
  (
    n2353,
    n1521,
    n1349,
    n1448,
    n1212
  );


  xor
  g2653
  (
    n2443,
    n1842,
    n1009,
    n1351,
    n1198
  );


  xor
  g2654
  (
    n2376,
    n1276,
    n1329,
    n1489,
    n1680
  );


  and
  g2655
  (
    n2633,
    n1925,
    n1248,
    n706,
    n902
  );


  or
  g2656
  (
    n2438,
    n1702,
    n1673,
    n1394,
    n1763
  );


  xnor
  g2657
  (
    n2405,
    n1689,
    n1175,
    n1871,
    n1706
  );


  xnor
  g2658
  (
    n2421,
    n1893,
    n949,
    n1820,
    n1802
  );


  and
  g2659
  (
    n2570,
    n1667,
    n1479,
    n1166,
    n908
  );


  nor
  g2660
  (
    n2563,
    n878,
    n1635,
    n1751,
    n1789
  );


  nand
  g2661
  (
    n2346,
    n1217,
    n1142,
    n1923,
    n1314
  );


  nor
  g2662
  (
    n2252,
    n1778,
    n1222,
    n963,
    n1479
  );


  nand
  g2663
  (
    n2193,
    n966,
    n1856,
    n1554,
    n942
  );


  xor
  g2664
  (
    n2393,
    n1844,
    n905,
    n1847,
    n742
  );


  or
  g2665
  (
    n2555,
    n1729,
    n860,
    n1614,
    n1429
  );


  nand
  g2666
  (
    n2398,
    n1728,
    n1588,
    n1249,
    n1468
  );


  xnor
  g2667
  (
    n2407,
    n1089,
    n1127,
    n1466,
    n1499
  );


  or
  g2668
  (
    n2624,
    n1059,
    n1714,
    n1027,
    n1141
  );


  xnor
  g2669
  (
    n2679,
    n1582,
    n1595,
    n1369,
    n1631
  );


  or
  g2670
  (
    n2349,
    n1663,
    n1904,
    n1042,
    n870
  );


  or
  g2671
  (
    n2312,
    n1571,
    n1157,
    n1700,
    n967
  );


  xnor
  g2672
  (
    n2525,
    n995,
    n1539,
    n875,
    n1774
  );


  xnor
  g2673
  (
    n2637,
    n848,
    n1051,
    n1120,
    n1384
  );


  or
  g2674
  (
    n2469,
    n1888,
    n1101,
    n1150,
    n1424
  );


  or
  g2675
  (
    n2660,
    n1745,
    n1442,
    n1797,
    n1034
  );


  and
  g2676
  (
    n2436,
    n1295,
    n1392,
    n931,
    n1417
  );


  nor
  g2677
  (
    n2317,
    n1278,
    n1659,
    n979,
    n990
  );


  xnor
  g2678
  (
    n2481,
    n1108,
    n1014,
    n1788,
    n1702
  );


  nor
  g2679
  (
    n2540,
    n1564,
    n1283,
    n845,
    n1578
  );


  or
  g2680
  (
    n2394,
    n920,
    n1031,
    n1576,
    n1738
  );


  and
  g2681
  (
    n2728,
    n855,
    n1069,
    n905,
    n1302
  );


  nor
  g2682
  (
    n2413,
    n1779,
    n1836,
    n1720,
    n1579
  );


  xnor
  g2683
  (
    n2382,
    n1095,
    n768,
    n1323,
    n1148
  );


  or
  g2684
  (
    n2329,
    n672,
    n800,
    n1496,
    n1762
  );


  xnor
  g2685
  (
    n2420,
    n1562,
    n734,
    n907,
    n1535
  );


  xnor
  g2686
  (
    n2636,
    n1755,
    n1715,
    n863,
    n1170
  );


  or
  g2687
  (
    n2638,
    n1092,
    n1266,
    n804,
    n752
  );


  nand
  g2688
  (
    n2410,
    n1561,
    n1699,
    n1632,
    n761
  );


  nor
  g2689
  (
    n2529,
    n1726,
    n1594,
    n1647,
    n1685
  );


  nor
  g2690
  (
    n2214,
    n1885,
    n1320,
    n1843,
    n921
  );


  nor
  g2691
  (
    n2352,
    n1503,
    n1109,
    n1398,
    n783
  );


  nand
  g2692
  (
    n2641,
    n1714,
    n1873,
    n1342,
    n1038
  );


  xor
  g2693
  (
    n2605,
    n698,
    n1722,
    n1119,
    n910
  );


  xnor
  g2694
  (
    n2245,
    n1633,
    n1088,
    n1095,
    n744
  );


  nor
  g2695
  (
    n2645,
    n928,
    n1399,
    n1288,
    n1724
  );


  or
  g2696
  (
    n2309,
    n1848,
    n1233,
    n1209,
    n1440
  );


  or
  g2697
  (
    n2565,
    n891,
    n697,
    n1029,
    n1306
  );


  nand
  g2698
  (
    n2492,
    n1655,
    n1752,
    n1648,
    n1518
  );


  nor
  g2699
  (
    n2691,
    n1191,
    n1737,
    n1242,
    n1277
  );


  xnor
  g2700
  (
    n2323,
    n814,
    n1099,
    n909,
    n904
  );


  xor
  g2701
  (
    n2661,
    n1652,
    n1838,
    n1704,
    n1291
  );


  and
  g2702
  (
    n2666,
    n1482,
    n943,
    n1592,
    n1104
  );


  nor
  g2703
  (
    n2415,
    n1310,
    n1909,
    n1103,
    n1186
  );


  nor
  g2704
  (
    n2328,
    n915,
    n1808,
    n887,
    n1308
  );


  nor
  g2705
  (
    n2427,
    n1103,
    n1786,
    n1679,
    n1928
  );


  xor
  g2706
  (
    n2740,
    n1912,
    n1047,
    n999,
    n1680
  );


  nor
  g2707
  (
    n2305,
    n1623,
    n1547,
    n1765,
    n705
  );


  xor
  g2708
  (
    n2539,
    n1111,
    n1292,
    n778,
    n931
  );


  or
  g2709
  (
    n2351,
    n1354,
    n1631,
    n1109,
    n1531
  );


  or
  g2710
  (
    n2366,
    n1882,
    n1257,
    n1670,
    n1159
  );


  buf
  g2711
  (
    n2824,
    n2272
  );


  buf
  g2712
  (
    n2780,
    n2252
  );


  not
  g2713
  (
    n2787,
    n2176
  );


  buf
  g2714
  (
    n2775,
    n2289
  );


  buf
  g2715
  (
    n2786,
    n2196
  );


  buf
  g2716
  (
    n2794,
    n2188
  );


  buf
  g2717
  (
    n2801,
    n2230
  );


  buf
  g2718
  (
    n2798,
    n2215
  );


  not
  g2719
  (
    n2744,
    n2301
  );


  buf
  g2720
  (
    n2747,
    n2298
  );


  not
  g2721
  (
    n2746,
    n2197
  );


  buf
  g2722
  (
    n2750,
    n2293
  );


  buf
  g2723
  (
    n2777,
    n2204
  );


  buf
  g2724
  (
    n2779,
    n2285
  );


  buf
  g2725
  (
    n2754,
    n2304
  );


  not
  g2726
  (
    n2772,
    n2286
  );


  buf
  g2727
  (
    n2764,
    n2294
  );


  buf
  g2728
  (
    n2808,
    n2295
  );


  buf
  g2729
  (
    n2763,
    n2271
  );


  buf
  g2730
  (
    n2773,
    n2193
  );


  not
  g2731
  (
    n2792,
    n2280
  );


  not
  g2732
  (
    n2759,
    n2290
  );


  not
  g2733
  (
    n2778,
    n2273
  );


  not
  g2734
  (
    n2819,
    n2263
  );


  not
  g2735
  (
    n2805,
    n2278
  );


  buf
  g2736
  (
    n2811,
    n2190
  );


  buf
  g2737
  (
    n2823,
    n2282
  );


  not
  g2738
  (
    n2762,
    n2232
  );


  not
  g2739
  (
    n2753,
    n2276
  );


  not
  g2740
  (
    n2766,
    n2266
  );


  buf
  g2741
  (
    n2781,
    n2241
  );


  not
  g2742
  (
    n2771,
    n2251
  );


  buf
  g2743
  (
    n2761,
    n2271
  );


  not
  g2744
  (
    n2800,
    n2283
  );


  buf
  g2745
  (
    n2758,
    n2179
  );


  buf
  g2746
  (
    n2812,
    n2249
  );


  buf
  g2747
  (
    KeyWire_0_9,
    n2297
  );


  buf
  g2748
  (
    n2769,
    n2284
  );


  buf
  g2749
  (
    n2799,
    n2213
  );


  buf
  g2750
  (
    n2807,
    n2223
  );


  buf
  g2751
  (
    n2803,
    n2282
  );


  buf
  g2752
  (
    n2751,
    n2226
  );


  buf
  g2753
  (
    n2748,
    n2289
  );


  not
  g2754
  (
    n2796,
    n2205
  );


  not
  g2755
  (
    n2788,
    n2211
  );


  buf
  g2756
  (
    n2765,
    n2180
  );


  not
  g2757
  (
    n2815,
    n2260
  );


  buf
  g2758
  (
    n2817,
    n2247
  );


  buf
  g2759
  (
    n2770,
    n2288
  );


  buf
  g2760
  (
    n2768,
    n2183
  );


  buf
  g2761
  (
    n2784,
    n2206
  );


  buf
  g2762
  (
    n2814,
    n2261
  );


  buf
  g2763
  (
    n2816,
    n2255
  );


  not
  g2764
  (
    n2804,
    n2250
  );


  xnor
  g2765
  (
    n2752,
    n2234,
    n2295,
    n2184,
    n2279
  );


  nand
  g2766
  (
    n2810,
    n2292,
    n2207,
    n2224,
    n2283
  );


  xor
  g2767
  (
    n2809,
    n2292,
    n2228,
    n2177,
    n2202
  );


  nor
  g2768
  (
    n2820,
    n2240,
    n2178,
    n2181,
    n2264
  );


  nor
  g2769
  (
    n2749,
    n2278,
    n2218,
    n2274,
    n2237
  );


  and
  g2770
  (
    n2827,
    n2209,
    n2245,
    n2287,
    n2254
  );


  xor
  g2771
  (
    n2793,
    n2298,
    n2303,
    n2187,
    n2273
  );


  nand
  g2772
  (
    n2789,
    n2199,
    n2189,
    n2299,
    n2301
  );


  or
  g2773
  (
    n2782,
    n2216,
    n2229,
    n2267,
    n2274
  );


  nor
  g2774
  (
    n2756,
    n2210,
    n2279,
    n2222,
    n2217
  );


  xnor
  g2775
  (
    n2745,
    n2239,
    n2175,
    n2269,
    n2265
  );


  nand
  g2776
  (
    n2757,
    n2277,
    n2172,
    n2168,
    n2191
  );


  nor
  g2777
  (
    n2755,
    n2300,
    n2238,
    n2195,
    n2275
  );


  xnor
  g2778
  (
    n2774,
    n2280,
    n2235,
    n2296,
    n2198
  );


  nand
  g2779
  (
    n2783,
    n2272,
    n2227,
    n2256,
    n2233
  );


  nor
  g2780
  (
    n2813,
    n2171,
    n2299,
    n2225,
    n2244
  );


  nand
  g2781
  (
    n2790,
    n2262,
    n2302,
    n2291,
    n2288
  );


  nand
  g2782
  (
    n2826,
    n2246,
    n2220,
    n2169,
    n2200
  );


  nand
  g2783
  (
    n2802,
    n2276,
    n2275,
    n2192,
    n2194
  );


  or
  g2784
  (
    n2825,
    n2248,
    n2300,
    n2243,
    n2293
  );


  and
  g2785
  (
    n2818,
    n2173,
    n2270,
    n2291,
    n2170
  );


  and
  g2786
  (
    n2760,
    n2212,
    n2242,
    n2236,
    n2296
  );


  xor
  g2787
  (
    n2767,
    n2174,
    n2290,
    n2186,
    n2267
  );


  nor
  g2788
  (
    n2791,
    n2285,
    n2268,
    n2214,
    n2286
  );


  nand
  g2789
  (
    n2821,
    n2258,
    n2201,
    n2268,
    n2284
  );


  xnor
  g2790
  (
    n2785,
    n2270,
    n2259,
    n2302,
    n2257
  );


  nand
  g2791
  (
    n2806,
    n2221,
    n2294,
    n2287,
    n2281
  );


  nor
  g2792
  (
    n2822,
    n2281,
    n2277,
    n2231,
    n2185
  );


  xnor
  g2793
  (
    n2797,
    n2219,
    n2269,
    n2303,
    n2253
  );


  or
  g2794
  (
    n2776,
    n2203,
    n2208,
    n2297,
    n2182
  );


  not
  g2795
  (
    n2831,
    n2745
  );


  buf
  g2796
  (
    n2836,
    n2747
  );


  not
  g2797
  (
    n2835,
    n2744
  );


  buf
  g2798
  (
    n2832,
    n1931
  );


  xor
  g2799
  (
    n2838,
    n2744,
    n1932,
    n2745,
    n2747
  );


  and
  g2800
  (
    n2837,
    n2748,
    n1935,
    n1934,
    n2746
  );


  xnor
  g2801
  (
    n2829,
    n1932,
    n1933,
    n2748,
    n1930
  );


  and
  g2802
  (
    n2830,
    n2747,
    n1930,
    n1933,
    n2744
  );


  or
  g2803
  (
    n2834,
    n2748,
    n2747,
    n2745,
    n2746
  );


  nand
  g2804
  (
    n2833,
    n1934,
    n2746,
    n1935
  );


  or
  g2805
  (
    n2828,
    n2745,
    n1929,
    n2744,
    n1931
  );


  or
  g2806
  (
    n2855,
    n1966,
    n1951,
    n1941,
    n1936
  );


  nand
  g2807
  (
    n2846,
    n2830,
    n1969,
    n2832,
    n1939
  );


  and
  g2808
  (
    n2852,
    n2833,
    n1945,
    n1952,
    n1940
  );


  and
  g2809
  (
    n2848,
    n1942,
    n1943,
    n2836,
    n1949
  );


  xor
  g2810
  (
    n2859,
    n1964,
    n2832,
    n1960,
    n1947
  );


  xnor
  g2811
  (
    n2842,
    n2831,
    n1959,
    n2837
  );


  and
  g2812
  (
    n2858,
    n1975,
    n2836,
    n1954,
    n1972
  );


  xnor
  g2813
  (
    n2841,
    n2831,
    n1962,
    n1963,
    n1969
  );


  xor
  g2814
  (
    n2857,
    n2834,
    n1964,
    n2831,
    n1938
  );


  xnor
  g2815
  (
    n2844,
    n1965,
    n1968,
    n2828,
    n1946
  );


  and
  g2816
  (
    n2863,
    n2833,
    n1974,
    n1939,
    n1953
  );


  or
  g2817
  (
    n2860,
    n1960,
    n2829,
    n1950,
    n1948
  );


  or
  g2818
  (
    n2845,
    n1954,
    n1951,
    n1973,
    n2829
  );


  nor
  g2819
  (
    n2854,
    n1963,
    n1952,
    n1970,
    n1965
  );


  nand
  g2820
  (
    n2865,
    n1938,
    n1967,
    n1943,
    n1956
  );


  nor
  g2821
  (
    n2849,
    n1949,
    n1957,
    n2830,
    n1948
  );


  or
  g2822
  (
    n2843,
    n1955,
    n1961,
    n1958,
    n1976
  );


  or
  g2823
  (
    n2856,
    n1957,
    n2832,
    n2833,
    n1936
  );


  nand
  g2824
  (
    n2861,
    n2835,
    n1961,
    n1953,
    n1975
  );


  nand
  g2825
  (
    n2839,
    n1937,
    n1971,
    n1968,
    n1941
  );


  nand
  g2826
  (
    n2853,
    n2835,
    n2837,
    n1962,
    n1944
  );


  xnor
  g2827
  (
    n2850,
    n1959,
    n2836,
    n1944,
    n1955
  );


  nand
  g2828
  (
    n2847,
    n1974,
    n1966,
    n1972,
    n1946
  );


  xnor
  g2829
  (
    n2851,
    n2835,
    n1970,
    n1950,
    n1973
  );


  xnor
  g2830
  (
    n2864,
    n2834,
    n1937,
    n1947,
    n1967
  );


  or
  g2831
  (
    n2862,
    n1956,
    n1940,
    n2834,
    n1945
  );


  xor
  g2832
  (
    n2840,
    n1971,
    n1942,
    n2836,
    n1958
  );


  and
  g2833
  (
    n2883,
    n2345,
    n2362,
    n2351,
    n2310
  );


  nor
  g2834
  (
    n2905,
    n2845,
    n2846,
    n2345,
    n2307
  );


  and
  g2835
  (
    n2870,
    n2338,
    n2850,
    n2351,
    n2340
  );


  nor
  g2836
  (
    n2880,
    n2841,
    n2353,
    n2848,
    n2324
  );


  nand
  g2837
  (
    n2876,
    n2352,
    n2357,
    n2319,
    n2314
  );


  xnor
  g2838
  (
    n2887,
    n2332,
    n2316,
    n2846,
    n2327
  );


  nor
  g2839
  (
    n2877,
    n2850,
    n2319,
    n2330,
    n2341
  );


  and
  g2840
  (
    n2884,
    n2343,
    n2350,
    n2316,
    n2845
  );


  nand
  g2841
  (
    n2889,
    n2306,
    n2317,
    n2330,
    n2346
  );


  or
  g2842
  (
    n2866,
    n2314,
    n2325,
    n2344,
    n2847
  );


  or
  g2843
  (
    n2894,
    n2323,
    n2355,
    n2356,
    n2841
  );


  nor
  g2844
  (
    n2892,
    n2359,
    n2849,
    n2842,
    n2355
  );


  or
  g2845
  (
    n2897,
    n2328,
    n2361,
    n2317,
    n2352
  );


  and
  g2846
  (
    n2868,
    n2304,
    n2360,
    n2329,
    n2363
  );


  and
  g2847
  (
    n2895,
    n2840,
    n2327,
    n2318,
    n2848
  );


  nor
  g2848
  (
    n2878,
    n2308,
    n2849,
    n2329,
    n2346
  );


  nand
  g2849
  (
    n2881,
    n2348,
    n2847,
    n2305,
    n2320
  );


  nand
  g2850
  (
    n2896,
    n2305,
    n2846,
    n2326,
    n2322
  );


  nand
  g2851
  (
    n2900,
    n2318,
    n2349,
    n2315
  );


  and
  g2852
  (
    n2902,
    n2332,
    n2336,
    n2334,
    n2342
  );


  or
  g2853
  (
    n2890,
    n2851,
    n2360,
    n2337,
    n2846
  );


  xor
  g2854
  (
    n2867,
    n2354,
    n2348,
    n2335,
    n2358
  );


  nor
  g2855
  (
    n2904,
    n2839,
    n2333,
    n2354,
    n2331
  );


  nand
  g2856
  (
    n2899,
    n2307,
    n2322,
    n2311,
    n2358
  );


  and
  g2857
  (
    n2869,
    n2339,
    n2315,
    n2321,
    n2848
  );


  nand
  g2858
  (
    n2891,
    n2844,
    n2331,
    n2309,
    n2353
  );


  xor
  g2859
  (
    n2871,
    n2338,
    n2321,
    n2333,
    n2344
  );


  nand
  g2860
  (
    n2882,
    n2842,
    n2356,
    n2357,
    n2325
  );


  nand
  g2861
  (
    n2885,
    n2308,
    n2335,
    n2343,
    n2313
  );


  nand
  g2862
  (
    n2873,
    n2840,
    n2845,
    n2312
  );


  xnor
  g2863
  (
    n2875,
    n2362,
    n2361,
    n2334,
    n2336
  );


  or
  g2864
  (
    n2898,
    n2849,
    n2847,
    n2848,
    n2341
  );


  xor
  g2865
  (
    n2886,
    n2313,
    n2849,
    n2320,
    n2347
  );


  or
  g2866
  (
    n2893,
    n2843,
    n2844
  );


  xor
  g2867
  (
    n2901,
    n2347,
    n2851,
    n2350,
    n2306
  );


  and
  g2868
  (
    n2874,
    n2839,
    n2843,
    n2359,
    n1976
  );


  or
  g2869
  (
    n2872,
    n2328,
    n2850,
    n2340,
    n2845
  );


  nor
  g2870
  (
    n2903,
    n2342,
    n2326,
    n2363,
    n2337
  );


  and
  g2871
  (
    n2879,
    n2310,
    n2324,
    n2309,
    n2311
  );


  xnor
  g2872
  (
    n2888,
    n2850,
    n2847,
    n2339,
    n2323
  );


  not
  g2873
  (
    n2947,
    n2889
  );


  buf
  g2874
  (
    n2951,
    n1989
  );


  not
  g2875
  (
    n2938,
    n1998
  );


  buf
  g2876
  (
    n2935,
    n2874
  );


  not
  g2877
  (
    n2942,
    n2020
  );


  buf
  g2878
  (
    n2939,
    n1999
  );


  not
  g2879
  (
    n2911,
    n2016
  );


  not
  g2880
  (
    n2927,
    n2019
  );


  not
  g2881
  (
    n2906,
    n2887
  );


  not
  g2882
  (
    n2910,
    n2005
  );


  buf
  g2883
  (
    n2921,
    n1994
  );


  not
  g2884
  (
    n2909,
    n1999
  );


  buf
  g2885
  (
    n2922,
    n2883
  );


  buf
  g2886
  (
    n2928,
    n2008
  );


  not
  g2887
  (
    n2913,
    n2867
  );


  not
  g2888
  (
    n2932,
    n2014
  );


  buf
  g2889
  (
    n2936,
    n1983
  );


  buf
  g2890
  (
    n2916,
    n2875
  );


  buf
  g2891
  (
    n2920,
    n2872
  );


  buf
  g2892
  (
    n2941,
    n1993
  );


  buf
  g2893
  (
    n2944,
    n2884
  );


  buf
  g2894
  (
    n2923,
    n1980
  );


  nand
  g2895
  (
    n2954,
    n1983,
    n2876,
    n1980,
    n2006
  );


  and
  g2896
  (
    n2914,
    n1982,
    n2881,
    n1994,
    n2873
  );


  and
  g2897
  (
    n2956,
    n2008,
    n1996,
    n1979,
    n2887
  );


  xor
  g2898
  (
    n2943,
    n1988,
    n1984,
    n2888,
    n2000
  );


  nor
  g2899
  (
    n2926,
    n2887,
    n1981,
    n2001,
    n2871
  );


  nand
  g2900
  (
    n2933,
    n2874,
    n1993,
    n2882,
    n2009
  );


  and
  g2901
  (
    n2958,
    n1989,
    n2869,
    n1997,
    n1987
  );


  or
  g2902
  (
    n2937,
    n2888,
    n2010,
    n2877,
    n1982
  );


  xnor
  g2903
  (
    n2917,
    n1988,
    n1995,
    n2015,
    n1984
  );


  xnor
  g2904
  (
    n2907,
    n2886,
    n1978,
    n2876,
    n2880
  );


  nand
  g2905
  (
    n2945,
    n2000,
    n2017,
    n2013,
    n2870
  );


  xor
  g2906
  (
    n2915,
    n2885,
    n1998,
    n1977,
    n2003
  );


  or
  g2907
  (
    n2931,
    n2877,
    n2004,
    n2017,
    n1990
  );


  nor
  g2908
  (
    n2949,
    n2888,
    n2888,
    n2023,
    n1992
  );


  and
  g2909
  (
    n2940,
    n2889,
    n2007,
    n2004,
    n2011
  );


  xnor
  g2910
  (
    n2934,
    n1997,
    n2889,
    n2870,
    n2013
  );


  or
  g2911
  (
    n2948,
    n2001,
    n2007,
    n2878,
    n2018
  );


  nor
  g2912
  (
    n2930,
    n2011,
    n2016,
    n2873,
    n2009
  );


  nand
  g2913
  (
    n2950,
    n2021,
    n2002,
    n2875,
    n1986
  );


  nor
  g2914
  (
    n2955,
    n1979,
    n1985,
    n2021,
    n2006
  );


  nor
  g2915
  (
    n2925,
    n2019,
    n2885,
    n2882,
    n1987
  );


  or
  g2916
  (
    n2953,
    n2872,
    n1986,
    n2883,
    n2002
  );


  xnor
  g2917
  (
    n2918,
    n1991,
    n2005,
    n1977,
    n1996
  );


  nand
  g2918
  (
    n2912,
    n2018,
    n2871,
    n2012,
    n2879
  );


  xor
  g2919
  (
    n2908,
    n2012,
    n2022,
    n2867,
    n1985
  );


  xor
  g2920
  (
    n2924,
    n1991,
    n2003,
    n2880,
    n2869
  );


  or
  g2921
  (
    n2929,
    n2884,
    n2022,
    n2020,
    n2881
  );


  and
  g2922
  (
    n2946,
    n2878,
    n2866,
    n1990,
    n2010
  );


  nor
  g2923
  (
    n2952,
    n1981,
    n2866,
    n2014,
    n2868
  );


  nand
  g2924
  (
    n2957,
    n2879,
    n2868,
    n2015,
    n2889
  );


  and
  g2925
  (
    n2919,
    n2886,
    n1995,
    n1978,
    n1992
  );


  nand
  g2926
  (
    n3164,
    n2495,
    n2942,
    n2385,
    n2925
  );


  and
  g2927
  (
    n3018,
    n2587,
    n2438,
    n2929,
    n2443
  );


  and
  g2928
  (
    n3135,
    n2937,
    n2917,
    n2426,
    n2912
  );


  xnor
  g2929
  (
    n2964,
    n2468,
    n2506,
    n2672,
    n2406
  );


  nor
  g2930
  (
    n3149,
    n2502,
    n2442,
    n2639,
    n2447
  );


  nor
  g2931
  (
    n3145,
    n2372,
    n2507,
    n2466,
    n2405
  );


  nand
  g2932
  (
    n3054,
    n2487,
    n2573,
    n2641,
    n2624
  );


  and
  g2933
  (
    n3074,
    n2486,
    n2651,
    n2944,
    n2918
  );


  and
  g2934
  (
    n3006,
    n2675,
    n2942,
    n2374,
    n2514
  );


  nor
  g2935
  (
    n3142,
    n2456,
    n2481,
    n2666,
    n2469
  );


  xor
  g2936
  (
    n3098,
    n2638,
    n2471,
    n2630,
    n2947
  );


  or
  g2937
  (
    n2969,
    n2928,
    n2378,
    n2956,
    n2550
  );


  nand
  g2938
  (
    n3073,
    n2399,
    n2931,
    n2448,
    n2911
  );


  nand
  g2939
  (
    n3124,
    n2457,
    n2583,
    n2498,
    n2909
  );


  or
  g2940
  (
    n3119,
    n2390,
    n2944,
    n2954,
    n2488
  );


  or
  g2941
  (
    n3058,
    n2608,
    n2654,
    n2502,
    n2462
  );


  nor
  g2942
  (
    n3050,
    n2934,
    n2513,
    n2933,
    n2376
  );


  nand
  g2943
  (
    n3117,
    n2385,
    n2583,
    n2529,
    n2941
  );


  xnor
  g2944
  (
    n3072,
    n2521,
    n2490,
    n2416,
    n2436
  );


  or
  g2945
  (
    n3107,
    n2926,
    n2586,
    n2928,
    n2521
  );


  nor
  g2946
  (
    n3140,
    n2674,
    n2918,
    n2659,
    n2490
  );


  xor
  g2947
  (
    n3043,
    n2413,
    n2955,
    n2598,
    n2667
  );


  and
  g2948
  (
    n2960,
    n2430,
    n2571,
    n2919,
    n2922
  );


  xnor
  g2949
  (
    n3045,
    n2564,
    n2486,
    n2948,
    n2366
  );


  nor
  g2950
  (
    n3166,
    n2915,
    n2457,
    n2621,
    n2454
  );


  and
  g2951
  (
    n3115,
    n2491,
    n2560,
    n2632,
    n2956
  );


  or
  g2952
  (
    n3026,
    n2927,
    n2933,
    n2439,
    n2665
  );


  nand
  g2953
  (
    n3136,
    n2569,
    n2451,
    n2943,
    n2669
  );


  or
  g2954
  (
    n3034,
    n2428,
    n2474,
    n2914,
    n2946
  );


  xnor
  g2955
  (
    n3063,
    n2941,
    n2365,
    n2562
  );


  and
  g2956
  (
    n3023,
    n2403,
    n2617,
    n2652,
    n2561
  );


  or
  g2957
  (
    n3061,
    n2601,
    n2545,
    n2574,
    n2438
  );


  and
  g2958
  (
    n2984,
    n2506,
    n2378,
    n2665,
    n2594
  );


  nand
  g2959
  (
    n3070,
    n2595,
    n2650,
    n2955,
    n2503
  );


  xor
  g2960
  (
    n3082,
    n2676,
    n2570,
    n2633,
    n2946
  );


  and
  g2961
  (
    n3031,
    n2910,
    n2462,
    n2550,
    n2541
  );


  nand
  g2962
  (
    n3127,
    n2383,
    n2620,
    n2402,
    n2482
  );


  and
  g2963
  (
    n3170,
    n2549,
    n2935,
    n2645,
    n2954
  );


  xor
  g2964
  (
    n3116,
    n2446,
    n2924,
    n2459,
    n2400
  );


  xor
  g2965
  (
    n3081,
    n2417,
    n2436,
    n2592,
    n2610
  );


  nor
  g2966
  (
    n3032,
    n2367,
    n2451,
    n2948,
    n2516
  );


  xor
  g2967
  (
    n3134,
    n2626,
    n2911,
    n2919,
    n2414
  );


  nor
  g2968
  (
    n2985,
    n2916,
    n2464,
    n2910,
    n2608
  );


  and
  g2969
  (
    n3151,
    n2540,
    n2393,
    n2444,
    n2950
  );


  nor
  g2970
  (
    n3088,
    n2388,
    n2954,
    n2463,
    n2370
  );


  xor
  g2971
  (
    n2970,
    n2475,
    n2371,
    n2952,
    n2403
  );


  and
  g2972
  (
    n3017,
    n2542,
    n2413,
    n2400,
    n2441
  );


  nand
  g2973
  (
    n3113,
    n2477,
    n2924,
    n2588,
    n2489
  );


  xnor
  g2974
  (
    n2965,
    n2909,
    n2398,
    n2519,
    n2558
  );


  nor
  g2975
  (
    n3048,
    n2620,
    n2377,
    n2406,
    n2650
  );


  xnor
  g2976
  (
    n3019,
    n2437,
    n2531,
    n2933,
    n2643
  );


  nand
  g2977
  (
    KeyWire_0_60,
    n2596,
    n2372,
    n2460,
    n2510
  );


  and
  g2978
  (
    n3097,
    n2472,
    n2373,
    n2409,
    n2386
  );


  nand
  g2979
  (
    n3051,
    n2929,
    n2611,
    n2596,
    n2652
  );


  or
  g2980
  (
    n3010,
    n2926,
    n2671,
    n2528,
    n2572
  );


  xnor
  g2981
  (
    n2999,
    n2487,
    n2567,
    n2584,
    n2638
  );


  or
  g2982
  (
    n3131,
    n2483,
    n2401,
    n2635,
    n2643
  );


  and
  g2983
  (
    n3004,
    n2524,
    n2419,
    n2609,
    n2379
  );


  nor
  g2984
  (
    n3085,
    n2375,
    n2401,
    n2609,
    n2919
  );


  or
  g2985
  (
    n3062,
    n2408,
    n2649,
    n2568,
    n2517
  );


  and
  g2986
  (
    KeyWire_0_37,
    n2480,
    n2613,
    n2576,
    n2590
  );


  nand
  g2987
  (
    n3167,
    n2622,
    n2442,
    n2938,
    n2470
  );


  nand
  g2988
  (
    n3020,
    n2472,
    n2454,
    n2674,
    n2582
  );


  nand
  g2989
  (
    n2975,
    n2931,
    n2933,
    n2481,
    n2422
  );


  nor
  g2990
  (
    n2993,
    n2614,
    n2936,
    n2368,
    n2443
  );


  nand
  g2991
  (
    n3021,
    n2952,
    n2402,
    n2464,
    n2404
  );


  and
  g2992
  (
    n3013,
    n2493,
    n2425,
    n2597,
    n2412
  );


  nor
  g2993
  (
    n3089,
    n2526,
    n2927,
    n2950
  );


  or
  g2994
  (
    KeyWire_0_5,
    n2509,
    n2544,
    n2559,
    n2910
  );


  or
  g2995
  (
    n3122,
    n2629,
    n2635,
    n2364,
    n2661
  );


  xnor
  g2996
  (
    n3037,
    n2662,
    n2477,
    n2908,
    n2536
  );


  nand
  g2997
  (
    n3016,
    n2618,
    n2921,
    n2418,
    n2947
  );


  xnor
  g2998
  (
    n3039,
    n2585,
    n2591,
    n2581,
    n2613
  );


  xnor
  g2999
  (
    n3160,
    n2610,
    n2432,
    n2604,
    n2578
  );


  and
  g3000
  (
    n3156,
    n2578,
    n2605,
    n2935,
    n2922
  );


  nor
  g3001
  (
    n3087,
    n2367,
    n2389,
    n2515,
    n2936
  );


  and
  g3002
  (
    KeyWire_0_49,
    n2430,
    n2409,
    n2653
  );


  nand
  g3003
  (
    n2998,
    n2431,
    n2673,
    n2628,
    n2458
  );


  xor
  g3004
  (
    n3007,
    n2658,
    n2949,
    n2636,
    n2412
  );


  or
  g3005
  (
    n3041,
    n2657,
    n2541,
    n2917,
    n2507
  );


  xnor
  g3006
  (
    n2968,
    n2600,
    n2957,
    n2394,
    n2946
  );


  xnor
  g3007
  (
    n3143,
    n2476,
    n2552,
    n2673,
    n2917
  );


  or
  g3008
  (
    n3025,
    n2557,
    n2912,
    n2906,
    n2953
  );


  xnor
  g3009
  (
    n2980,
    n2384,
    n2951,
    n2424,
    n2644
  );


  xor
  g3010
  (
    n2982,
    n2572,
    n2423,
    n2602,
    n2912
  );


  nand
  g3011
  (
    n3102,
    n2410,
    n2924,
    n2554,
    n2548
  );


  xor
  g3012
  (
    n3093,
    n2664,
    n2423,
    n2508,
    n2425
  );


  xnor
  g3013
  (
    n3157,
    n2953,
    n2592,
    n2938,
    n2543
  );


  xor
  g3014
  (
    n3014,
    n2663,
    n2545,
    n2571,
    n2679
  );


  xor
  g3015
  (
    n3159,
    n2469,
    n2957,
    n2510,
    n2634
  );


  xnor
  g3016
  (
    n3064,
    n2911,
    n2931,
    n2937,
    n2636
  );


  xor
  g3017
  (
    n3078,
    n2551,
    n2681,
    n2935,
    n2916
  );


  nand
  g3018
  (
    n3155,
    n2478,
    n2623,
    n2399,
    n2928
  );


  or
  g3019
  (
    n3012,
    n2920,
    n2532,
    n2463,
    n2516
  );


  nor
  g3020
  (
    n2961,
    n2582,
    n2433,
    n2680,
    n2570
  );


  or
  g3021
  (
    n3150,
    n2476,
    n2503,
    n2420,
    n2515
  );


  xnor
  g3022
  (
    n2966,
    n2384,
    n2598,
    n2639,
    n2566
  );


  or
  g3023
  (
    n3101,
    n2930,
    n2606,
    n2577,
    n2544
  );


  nand
  g3024
  (
    n3146,
    n2595,
    n2611,
    n2629,
    n2957
  );


  and
  g3025
  (
    n3108,
    n2561,
    n2419,
    n2913,
    n2539
  );


  xor
  g3026
  (
    n2962,
    n2658,
    n2663,
    n2422,
    n2642
  );


  xor
  g3027
  (
    n3125,
    n2573,
    n2612,
    n2479,
    n2369
  );


  nor
  g3028
  (
    n3152,
    n2953,
    n2392,
    n2921,
    n2522
  );


  and
  g3029
  (
    n3110,
    n2536,
    n2539,
    n2915,
    n2526
  );


  xnor
  g3030
  (
    n3106,
    n2630,
    n2459,
    n2415,
    n2654
  );


  nand
  g3031
  (
    n3065,
    n2505,
    n2512,
    n2932,
    n2614
  );


  and
  g3032
  (
    n3153,
    n2942,
    n2511,
    n2500,
    n2518
  );


  xor
  g3033
  (
    n3096,
    n2915,
    n2567,
    n2563,
    n2648
  );


  xnor
  g3034
  (
    n3079,
    n2656,
    n2645,
    n2483,
    n2435
  );


  xnor
  g3035
  (
    n3118,
    n2634,
    n2492,
    n2940,
    n2525
  );


  nor
  g3036
  (
    n3092,
    n2666,
    n2920,
    n2655,
    n2593
  );


  or
  g3037
  (
    n3137,
    n2559,
    n2947,
    n2948,
    n2927
  );


  xnor
  g3038
  (
    n3128,
    n2475,
    n2605,
    n2915,
    n2599
  );


  xor
  g3039
  (
    n2986,
    n2589,
    n2466,
    n2568,
    n2379
  );


  nor
  g3040
  (
    n3022,
    n2919,
    n2922,
    n2640,
    n2644
  );


  xor
  g3041
  (
    n3120,
    n2628,
    n2624,
    n2404,
    n2371
  );


  or
  g3042
  (
    n3047,
    n2599,
    n2952,
    n2907,
    n2505
  );


  and
  g3043
  (
    n2983,
    n2530,
    n2924,
    n2556,
    n2955
  );


  xnor
  g3044
  (
    n3008,
    n2945,
    n2411,
    n2648,
    n2681
  );


  nand
  g3045
  (
    n3060,
    n2579,
    n2649,
    n2512,
    n2427
  );


  nor
  g3046
  (
    n2997,
    n2575,
    n2918,
    n2433,
    n2377
  );


  and
  g3047
  (
    n3042,
    n2388,
    n2956,
    n2484,
    n2547
  );


  nor
  g3048
  (
    n2963,
    n2563,
    n2467,
    n2434,
    n2580
  );


  or
  g3049
  (
    n3040,
    n2514,
    n2940,
    n2944,
    n2518
  );


  nor
  g3050
  (
    n2959,
    n2677,
    n2485,
    n2391,
    n2951
  );


  xnor
  g3051
  (
    n3133,
    n2930,
    n2591,
    n2553,
    n2560
  );


  xnor
  g3052
  (
    n3138,
    n2479,
    n2524,
    n2489,
    n2942
  );


  nand
  g3053
  (
    n3030,
    n2918,
    n2627,
    n2934,
    n2533
  );


  nand
  g3054
  (
    n3036,
    n2523,
    n2432,
    n2375,
    n2549
  );


  or
  g3055
  (
    n2995,
    n2491,
    n2945,
    n2911,
    n2452
  );


  or
  g3056
  (
    n3028,
    n2498,
    n2411,
    n2656,
    n2492
  );


  xnor
  g3057
  (
    n3105,
    n2621,
    n2397,
    n2954,
    n2467
  );


  or
  g3058
  (
    n3100,
    n2647,
    n2937,
    n2943,
    n2659
  );


  or
  g3059
  (
    n3162,
    n2452,
    n2923,
    n2525,
    n2535
  );


  nand
  g3060
  (
    n3056,
    n2947,
    n2435,
    n2380,
    n2537
  );


  nor
  g3061
  (
    n3038,
    n2538,
    n2387,
    n2470,
    n2532
  );


  or
  g3062
  (
    n3027,
    n2450,
    n2939,
    n2641,
    n2424
  );


  xnor
  g3063
  (
    n3068,
    n2677,
    n2374,
    n2923,
    n2940
  );


  xnor
  g3064
  (
    n3147,
    n2917,
    n2499,
    n2407,
    n2569
  );


  nor
  g3065
  (
    n3114,
    n2581,
    n2382,
    n2908,
    n2936
  );


  nand
  g3066
  (
    n3009,
    n2660,
    n2678,
    n2943,
    n2957
  );


  nor
  g3067
  (
    n3069,
    n2906,
    n2932,
    n2495,
    n2937
  );


  xor
  g3068
  (
    n3161,
    n2543,
    n2535,
    n2458,
    n2394
  );


  nand
  g3069
  (
    n3130,
    n2523,
    n2511,
    n2445,
    n2939
  );


  and
  g3070
  (
    n3126,
    n2908,
    n2364,
    n2565,
    n2907
  );


  and
  g3071
  (
    n3154,
    n2589,
    n2393,
    n2386,
    n2540
  );


  xor
  g3072
  (
    n3066,
    n2449,
    n2626,
    n2465,
    n2916
  );


  nor
  g3073
  (
    n3129,
    n2392,
    n2678,
    n2434,
    n2615
  );


  and
  g3074
  (
    n2977,
    n2934,
    n2390,
    n2485,
    n2657
  );


  nand
  g3075
  (
    n3083,
    n2580,
    n2429,
    n2431,
    n2615
  );


  and
  g3076
  (
    n2992,
    n2439,
    n2565,
    n2497,
    n2418
  );


  nand
  g3077
  (
    n3111,
    n2395,
    n2574,
    n2637,
    n2934
  );


  and
  g3078
  (
    n3033,
    n2948,
    n2389,
    n2909,
    n2445
  );


  nand
  g3079
  (
    n3059,
    n2922,
    n2950,
    n2496,
    n2923
  );


  nor
  g3080
  (
    n3044,
    n2670,
    n2529,
    n2932,
    n2675
  );


  xor
  g3081
  (
    n3141,
    n2522,
    n2437,
    n2428,
    n2504
  );


  or
  g3082
  (
    n3003,
    n2955,
    n2662,
    n2943,
    n2622
  );


  xnor
  g3083
  (
    n2987,
    n2546,
    n2421,
    n2557,
    n2642
  );


  and
  g3084
  (
    n2974,
    n2368,
    n2493,
    n2936,
    n2956
  );


  xor
  g3085
  (
    n3103,
    n2909,
    n2935,
    n2387,
    n2547
  );


  nor
  g3086
  (
    n3091,
    n2920,
    n2555,
    n2494,
    n2930
  );


  nand
  g3087
  (
    n3158,
    n2554,
    n2921,
    n2585,
    n2456
  );


  xnor
  g3088
  (
    n3099,
    n2551,
    n2958,
    n2509,
    n2553
  );


  xor
  g3089
  (
    n2967,
    n2461,
    n2449,
    n2912,
    n2427
  );


  xnor
  g3090
  (
    n3168,
    n2417,
    n2606,
    n2941,
    n2637
  );


  xor
  g3091
  (
    n3090,
    n2906,
    n2501,
    n2474,
    n2414
  );


  xnor
  g3092
  (
    n3080,
    n2929,
    n2415,
    n2546,
    n2616
  );


  or
  g3093
  (
    n3139,
    n2651,
    n2625,
    n2416,
    n2670
  );


  or
  g3094
  (
    n2994,
    n2627,
    n2527,
    n2945,
    n2944
  );


  and
  g3095
  (
    n3086,
    n2939,
    n2504,
    n2468,
    n2920
  );


  xor
  g3096
  (
    n3169,
    n2564,
    n2533,
    n2914,
    n2473
  );


  xor
  g3097
  (
    n3112,
    n2517,
    n2548,
    n2566,
    n2926
  );


  xor
  g3098
  (
    n3015,
    n2906,
    n2369,
    n2382,
    n2447
  );


  xor
  g3099
  (
    n3011,
    n2680,
    n2616,
    n2930,
    n2631
  );


  and
  g3100
  (
    n2972,
    n2440,
    n2664,
    n2603,
    n2932
  );


  and
  g3101
  (
    n3123,
    n2531,
    n2952,
    n2604,
    n2669
  );


  xnor
  g3102
  (
    n3094,
    n2646,
    n2625,
    n2672,
    n2576
  );


  and
  g3103
  (
    n2976,
    n2667,
    n2380,
    n2397,
    n2913
  );


  nor
  g3104
  (
    n2978,
    n2938,
    n2601,
    n2668,
    n2453
  );


  xor
  g3105
  (
    n3071,
    n2908,
    n2671,
    n2446,
    n2448
  );


  nor
  g3106
  (
    n3144,
    n2958,
    n2593,
    n2480,
    n2588
  );


  xor
  g3107
  (
    n3049,
    n2668,
    n2429,
    n2958,
    n2907
  );


  nor
  g3108
  (
    n3076,
    n2632,
    n2366,
    n2676,
    n2381
  );


  xnor
  g3109
  (
    n3046,
    n2494,
    n2617,
    n2552,
    n2914
  );


  nor
  g3110
  (
    n2990,
    n2453,
    n2619,
    n2602,
    n2497
  );


  xor
  g3111
  (
    n3035,
    n2577,
    n2949,
    n2365,
    n2450
  );


  nand
  g3112
  (
    n3121,
    n2496,
    n2420,
    n2538,
    n2558
  );


  nand
  g3113
  (
    n3067,
    n2927,
    n2513,
    n2555,
    n2542
  );


  or
  g3114
  (
    n2991,
    n2612,
    n2410,
    n2391,
    n2440
  );


  xor
  g3115
  (
    n3055,
    n2618,
    n2929,
    n2590,
    n2951
  );


  and
  g3116
  (
    n3077,
    n2603,
    n2679,
    n2925,
    n2484
  );


  nand
  g3117
  (
    n2971,
    n2594,
    n2655,
    n2623,
    n2534
  );


  nand
  g3118
  (
    n3084,
    n2407,
    n2949,
    n2619,
    n2421
  );


  or
  g3119
  (
    n3052,
    n2426,
    n2923,
    n2519,
    n2660
  );


  xor
  g3120
  (
    n3148,
    n2508,
    n2925,
    n2376,
    n2600
  );


  xor
  g3121
  (
    n3002,
    n2478,
    n2482,
    n2913,
    n2534
  );


  and
  g3122
  (
    n2988,
    n2500,
    n2455,
    n2938,
    n2395
  );


  xnor
  g3123
  (
    n3165,
    n2461,
    n2527,
    n2607,
    n2953
  );


  and
  g3124
  (
    n3057,
    n2441,
    n2640,
    n2383,
    n2373
  );


  and
  g3125
  (
    n2996,
    n2597,
    n2584,
    n2926,
    n2579
  );


  nor
  g3126
  (
    n3095,
    n2455,
    n2646,
    n2931,
    n2586
  );


  xor
  g3127
  (
    n3005,
    n2499,
    n2488,
    n2465,
    n2913
  );


  nor
  g3128
  (
    n3000,
    n2914,
    n2528,
    n2530,
    n2396
  );


  and
  g3129
  (
    n3053,
    n2370,
    n2575,
    n2928,
    n2939
  );


  and
  g3130
  (
    n3104,
    n2520,
    n2587,
    n2949,
    n2556
  );


  xnor
  g3131
  (
    n2973,
    n2940,
    n2381,
    n2473,
    n2396
  );


  and
  g3132
  (
    n2981,
    n2958,
    n2925,
    n2460,
    n2537
  );


  xnor
  g3133
  (
    n3075,
    n2921,
    n2444,
    n2945,
    n2607
  );


  xor
  g3134
  (
    n3001,
    n2633,
    n2910,
    n2907,
    n2631
  );


  nand
  g3135
  (
    n3109,
    n2398,
    n2501,
    n2916,
    n2408
  );


  xor
  g3136
  (
    n2989,
    n2951,
    n2946,
    n2941,
    n2520
  );


  and
  g3137
  (
    n3163,
    n2405,
    n2647,
    n2471,
    n2661
  );


  buf
  g3138
  (
    n3322,
    n2778
  );


  buf
  g3139
  (
    n3314,
    n2753
  );


  not
  g3140
  (
    n3256,
    n3086
  );


  buf
  g3141
  (
    n3286,
    n2762
  );


  buf
  g3142
  (
    KeyWire_0_42,
    n2989
  );


  xnor
  g3143
  (
    n3363,
    n2775,
    n3075
  );


  xnor
  g3144
  (
    n3390,
    n2805,
    n2976
  );


  xor
  g3145
  (
    n3270,
    n2767,
    n2979
  );


  nand
  g3146
  (
    n3232,
    n3013,
    n3024
  );


  nand
  g3147
  (
    n3196,
    n3011,
    n3026,
    n3102,
    n2825
  );


  and
  g3148
  (
    n3371,
    n3071,
    n2780,
    n3006,
    n3022
  );


  xnor
  g3149
  (
    n3295,
    n2752,
    n2811,
    n2965,
    n3008
  );


  xnor
  g3150
  (
    n3220,
    n3019,
    n2794,
    n3066,
    n2815
  );


  or
  g3151
  (
    n3377,
    n2798,
    n2975,
    n3007,
    n3091
  );


  and
  g3152
  (
    n3187,
    n2782,
    n2770,
    n2825,
    n2974
  );


  nand
  g3153
  (
    n3215,
    n2758,
    n2838,
    n3093,
    n2990
  );


  nor
  g3154
  (
    n3317,
    n2802,
    n3070,
    n3021,
    n3047
  );


  nor
  g3155
  (
    n3367,
    n3019,
    n3015,
    n3049,
    n3032
  );


  xnor
  g3156
  (
    n3223,
    n2968,
    n3001,
    n2987,
    n2964
  );


  and
  g3157
  (
    n3321,
    n2771,
    n2990,
    n3052,
    n3041
  );


  nor
  g3158
  (
    n3344,
    n2796,
    n3023,
    n3080,
    n3076
  );


  or
  g3159
  (
    n3179,
    n2764,
    n3064,
    n2992,
    n2816
  );


  xnor
  g3160
  (
    n3374,
    n2991,
    n2761,
    n3094,
    n2993
  );


  and
  g3161
  (
    n3289,
    n3067,
    n2755,
    n2989,
    n3042
  );


  nor
  g3162
  (
    n3181,
    n3042,
    n3078,
    n2821,
    n2978
  );


  nor
  g3163
  (
    n3231,
    n2971,
    n2817,
    n2789,
    n3009
  );


  nor
  g3164
  (
    n3199,
    n3068,
    n3041,
    n3033,
    n2857
  );


  or
  g3165
  (
    n3233,
    n2750,
    n3051,
    n2959,
    n2024
  );


  xnor
  g3166
  (
    n3209,
    n2799,
    n2979,
    n3008,
    n2824
  );


  nor
  g3167
  (
    n3357,
    n2765,
    n2976,
    n3091,
    n2855
  );


  and
  g3168
  (
    KeyWire_0_36,
    n2959,
    n2813,
    n2996,
    n2769
  );


  and
  g3169
  (
    n3361,
    n2823,
    n2817,
    n2779,
    n2784
  );


  xnor
  g3170
  (
    n3251,
    n2812,
    n2777,
    n3088,
    n2991
  );


  and
  g3171
  (
    n3408,
    n2816,
    n3013,
    n3081,
    n2819
  );


  or
  g3172
  (
    n3253,
    n2749,
    n2803,
    n3086,
    n3044
  );


  nand
  g3173
  (
    n3405,
    n2821,
    n2851,
    n3053,
    n3034
  );


  xnor
  g3174
  (
    n3189,
    n3004,
    n2981,
    n2762,
    n2785
  );


  or
  g3175
  (
    n3393,
    n3000,
    n3103,
    n3043,
    n3029
  );


  nand
  g3176
  (
    n3207,
    n3011,
    n2974,
    n3003,
    n2758
  );


  nand
  g3177
  (
    n3358,
    n3075,
    n2822,
    n3063,
    n2794
  );


  nor
  g3178
  (
    n3210,
    n3013,
    n3052,
    n3078,
    n2985
  );


  xor
  g3179
  (
    n3254,
    n2853,
    n2984,
    n2790,
    n2822
  );


  or
  g3180
  (
    n3269,
    n2977,
    n3005,
    n2758,
    n3078
  );


  and
  g3181
  (
    n3288,
    n3085,
    n3050,
    n2855,
    n3017
  );


  nor
  g3182
  (
    n3388,
    n3061,
    n3035,
    n2026,
    n3029
  );


  nand
  g3183
  (
    n3303,
    n2792,
    n3010,
    n2821,
    n3027
  );


  nor
  g3184
  (
    n3175,
    n3073,
    n2994,
    n2806,
    n2985
  );


  and
  g3185
  (
    n3287,
    n2962,
    n2994,
    n3066,
    n2854
  );


  or
  g3186
  (
    n3171,
    n3074,
    n3054,
    n2786,
    n3024
  );


  xnor
  g3187
  (
    n3261,
    n2782,
    n2989,
    n2980,
    n3033
  );


  nor
  g3188
  (
    n3308,
    n2026,
    n3076,
    n2857,
    n2858
  );


  nand
  g3189
  (
    n3197,
    n2827,
    n3060,
    n2687,
    n3067
  );


  and
  g3190
  (
    n3258,
    n3009,
    n3025,
    n2752,
    n2820
  );


  xor
  g3191
  (
    n3283,
    n2759,
    n2967,
    n2811,
    n3074
  );


  or
  g3192
  (
    n3176,
    n2977,
    n2978,
    n2804,
    n3091
  );


  xor
  g3193
  (
    n3402,
    n3024,
    n3083,
    n2752,
    n3040
  );


  xor
  g3194
  (
    n3264,
    n2769,
    n2970,
    n2858,
    n2791
  );


  or
  g3195
  (
    n3279,
    n3077,
    n2856,
    n3039,
    n3021
  );


  and
  g3196
  (
    n3315,
    n3012,
    n2755,
    n2966,
    n2857
  );


  xnor
  g3197
  (
    n3304,
    n3093,
    n3079,
    n3088,
    n2970
  );


  nor
  g3198
  (
    n3359,
    n3037,
    n3026,
    n3097,
    n3038
  );


  and
  g3199
  (
    n3312,
    n3003,
    n3063,
    n3035,
    n2024
  );


  nand
  g3200
  (
    n3240,
    n3014,
    n2789,
    n2992,
    n2800
  );


  or
  g3201
  (
    n3205,
    n3027,
    n2981,
    n3015,
    n3044
  );


  nor
  g3202
  (
    n3190,
    n2814,
    n3085,
    n3073,
    n3099
  );


  and
  g3203
  (
    n3297,
    n2971,
    n3043,
    n2980,
    n2961
  );


  nand
  g3204
  (
    n3296,
    n2995,
    n2997,
    n3047
  );


  xnor
  g3205
  (
    n3360,
    n3038,
    n3008,
    n2764,
    n2795
  );


  and
  g3206
  (
    n3330,
    n2813,
    n2854,
    n3017,
    n2802
  );


  xor
  g3207
  (
    n3395,
    n2814,
    n2804,
    n3060,
    n3095
  );


  xor
  g3208
  (
    n3242,
    n3045,
    n3097,
    n3002,
    n2983
  );


  and
  g3209
  (
    n3234,
    n2777,
    n2993,
    n2774,
    n2023
  );


  and
  g3210
  (
    n3352,
    n3061,
    n2807,
    n3031,
    n2987
  );


  or
  g3211
  (
    n3403,
    n3004,
    n3032,
    n2795,
    n2784
  );


  xor
  g3212
  (
    n3218,
    n3016,
    n3090,
    n2996,
    n2982
  );


  nand
  g3213
  (
    n3338,
    n2754,
    n3011,
    n3070,
    n3075
  );


  xor
  g3214
  (
    n3309,
    n2782,
    n3083,
    n3047,
    n3069
  );


  nand
  g3215
  (
    n3318,
    n3079,
    n3101,
    n3010,
    n2760
  );


  xor
  g3216
  (
    n3356,
    n3099,
    n2814,
    n3102,
    n2974
  );


  or
  g3217
  (
    n3227,
    n2783,
    n2975,
    n3012
  );


  nor
  g3218
  (
    n3277,
    n2852,
    n2979,
    n2989,
    n3017
  );


  nand
  g3219
  (
    n3248,
    n3067,
    n3044,
    n2757,
    n2780
  );


  or
  g3220
  (
    n3406,
    n2852,
    n3065,
    n3039,
    n3040
  );


  xor
  g3221
  (
    n3307,
    n3077,
    n2996,
    n2791,
    n2990
  );


  xnor
  g3222
  (
    n3306,
    n2803,
    n2797,
    n2994,
    n3079
  );


  xor
  g3223
  (
    n3213,
    n2767,
    n2770,
    n3072,
    n3023
  );


  xor
  g3224
  (
    n3226,
    n3011,
    n2977,
    n2755,
    n3073
  );


  and
  g3225
  (
    n3222,
    n2685,
    n3084,
    n2793,
    n3098
  );


  and
  g3226
  (
    n3183,
    n3099,
    n3012,
    n2853,
    n2969
  );


  nand
  g3227
  (
    n3345,
    n3001,
    n2827,
    n2791,
    n2859
  );


  or
  g3228
  (
    n3397,
    n3030,
    n2964,
    n2801,
    n3048
  );


  or
  g3229
  (
    n3362,
    n2987,
    n3053,
    n2803,
    n2752
  );


  or
  g3230
  (
    n3347,
    n2753,
    n3089,
    n2790,
    n3070
  );


  and
  g3231
  (
    n3219,
    n3021,
    n2797,
    n3015,
    n2751
  );


  and
  g3232
  (
    n3381,
    n2795,
    n2819,
    n3049,
    n2972
  );


  and
  g3233
  (
    n3228,
    n2988,
    n3099,
    n3055,
    n3007
  );


  xnor
  g3234
  (
    n3243,
    n2753,
    n3065,
    n2787,
    n3040
  );


  or
  g3235
  (
    n3300,
    n2808,
    n2858,
    n2823,
    n2817
  );


  xnor
  g3236
  (
    n3409,
    n3016,
    n3036,
    n2807,
    n3078
  );


  xnor
  g3237
  (
    n3259,
    n3076,
    n2855,
    n3052,
    n3023
  );


  xnor
  g3238
  (
    n3186,
    n2756,
    n3021,
    n3057,
    n2972
  );


  nor
  g3239
  (
    n3255,
    n3079,
    n2826,
    n3081
  );


  nand
  g3240
  (
    n3244,
    n3056,
    n3012,
    n3089,
    n2999
  );


  and
  g3241
  (
    n3291,
    n3082,
    n2826,
    n2766,
    n2856
  );


  xnor
  g3242
  (
    n3400,
    n2781,
    n2755,
    n2778,
    n3054
  );


  xor
  g3243
  (
    n3342,
    n2798,
    n2969,
    n2985,
    n3034
  );


  nor
  g3244
  (
    n3336,
    n2751,
    n3069,
    n3059,
    n3006
  );


  and
  g3245
  (
    n3208,
    n2979,
    n2815,
    n3014,
    n3029
  );


  xor
  g3246
  (
    n3364,
    n2764,
    n3072,
    n2798,
    n2799
  );


  xor
  g3247
  (
    n3247,
    n3037,
    n2800,
    n3048,
    n2820
  );


  xor
  g3248
  (
    n3294,
    n3056,
    n3089,
    n2781,
    n3018
  );


  or
  g3249
  (
    n3346,
    n3041,
    n3030,
    n2999,
    n2808
  );


  and
  g3250
  (
    n3194,
    n2851,
    n2968,
    n3050,
    n3062
  );


  xnor
  g3251
  (
    n3236,
    n3045,
    n3096,
    n2757,
    n2800
  );


  xor
  g3252
  (
    n3333,
    n2815,
    n3073,
    n2795,
    n2773
  );


  or
  g3253
  (
    n3173,
    n3005,
    n3056,
    n3024,
    n3027
  );


  nand
  g3254
  (
    n3373,
    n3084,
    n3077,
    n3005,
    n2972
  );


  xnor
  g3255
  (
    n3365,
    n3018,
    n3071,
    n2814,
    n2998
  );


  xnor
  g3256
  (
    n3262,
    n2775,
    n2991,
    n2768,
    n3016
  );


  or
  g3257
  (
    n3177,
    n3095,
    n3074,
    n3001,
    n2789
  );


  nand
  g3258
  (
    n3326,
    n3008,
    n2775,
    n2999,
    n2754
  );


  or
  g3259
  (
    n3246,
    n2806,
    n2992,
    n2750,
    n3084
  );


  xor
  g3260
  (
    n3266,
    n2983,
    n2810,
    n3083,
    n3003
  );


  nand
  g3261
  (
    n3201,
    n3071,
    n3000,
    n2766,
    n2796
  );


  and
  g3262
  (
    n3221,
    n2765,
    n2980,
    n3056,
    n3053
  );


  nand
  g3263
  (
    n3298,
    n3049,
    n2788,
    n2824,
    n2749
  );


  and
  g3264
  (
    n3305,
    n2800,
    n3098,
    n3002,
    n2994
  );


  xor
  g3265
  (
    n3339,
    n3102,
    n2962,
    n3086,
    n2760
  );


  xor
  g3266
  (
    n3274,
    n2792,
    n3015,
    n2978,
    n2775
  );


  xor
  g3267
  (
    n3252,
    n3006,
    n2785,
    n2992,
    n2682
  );


  nand
  g3268
  (
    n3313,
    n2779,
    n2768,
    n3018,
    n2776
  );


  or
  g3269
  (
    n3214,
    n2816,
    n2804,
    n2806,
    n3014
  );


  or
  g3270
  (
    n3216,
    n2966,
    n3062,
    n2688,
    n3093
  );


  nand
  g3271
  (
    n3276,
    n3063,
    n2761,
    n2973,
    n3066
  );


  nor
  g3272
  (
    n3260,
    n3043,
    n3040,
    n3041,
    n3081
  );


  nand
  g3273
  (
    n3250,
    n2855,
    n2852,
    n3082,
    n3086
  );


  nand
  g3274
  (
    n3372,
    n3088,
    n2822,
    n2799,
    n3084
  );


  or
  g3275
  (
    n3401,
    n3075,
    n2827,
    n3019,
    n2751
  );


  xnor
  g3276
  (
    n3350,
    n2817,
    n2788,
    n2790,
    n3037
  );


  nor
  g3277
  (
    n3206,
    n2987,
    n3101,
    n3061,
    n2983
  );


  xor
  g3278
  (
    n3384,
    n3030,
    n3087,
    n3058,
    n3050
  );


  nand
  g3279
  (
    n3378,
    n2812,
    n2769,
    n2773,
    n2770
  );


  nand
  g3280
  (
    n3178,
    n2791,
    n3039,
    n2772,
    n3091
  );


  and
  g3281
  (
    n3323,
    n3035,
    n3004,
    n2683,
    n2978
  );


  or
  g3282
  (
    n3238,
    n3047,
    n3005,
    n2995,
    n3097
  );


  nor
  g3283
  (
    n3324,
    n3089,
    n2801,
    n2756,
    n3096
  );


  xnor
  g3284
  (
    n3267,
    n3034,
    n3069,
    n2785,
    n2794
  );


  or
  g3285
  (
    n3217,
    n2769,
    n3097,
    n2856,
    n2767
  );


  nor
  g3286
  (
    n3376,
    n2765,
    n2826,
    n2753,
    n3003
  );


  nand
  g3287
  (
    n3235,
    n3072,
    n2790,
    n3036,
    n2984
  );


  or
  g3288
  (
    n3265,
    n2805,
    n3085,
    n3080,
    n2776
  );


  nor
  g3289
  (
    n3281,
    n3006,
    n3083,
    n3101,
    n3031
  );


  nand
  g3290
  (
    n3380,
    n2818,
    n3098,
    n3100,
    n2810
  );


  or
  g3291
  (
    n3182,
    n3032,
    n2961,
    n2786,
    n3022
  );


  nand
  g3292
  (
    n3188,
    n2760,
    n2788,
    n3030,
    n3009
  );


  nand
  g3293
  (
    n3319,
    n3025,
    n3020,
    n2824,
    n2857
  );


  xnor
  g3294
  (
    n3349,
    n2750,
    n2768,
    n3031,
    n3059
  );


  nand
  g3295
  (
    n3387,
    n2778,
    n3032,
    n3022,
    n3087
  );


  xnor
  g3296
  (
    n3392,
    n3043,
    n3068,
    n2985,
    n2818
  );


  xnor
  g3297
  (
    n3328,
    n2774,
    n3053,
    n2998,
    n2787
  );


  and
  g3298
  (
    n3399,
    n2793,
    n3090,
    n2854,
    n3067
  );


  and
  g3299
  (
    n3211,
    n2998,
    n2824,
    n2756,
    n2770
  );


  and
  g3300
  (
    n3192,
    n2986,
    n2805,
    n2779,
    n2815
  );


  nand
  g3301
  (
    n3172,
    n2960,
    n3077,
    n2805,
    n2982
  );


  xor
  g3302
  (
    n3334,
    n3103,
    n2821,
    n3020,
    n2984
  );


  xnor
  g3303
  (
    n3329,
    n3058,
    n2777,
    n2768,
    n3029
  );


  nand
  g3304
  (
    n3348,
    n2786,
    n2963,
    n3002,
    n2999
  );


  and
  g3305
  (
    n3293,
    n2990,
    n2802,
    n3058,
    n3028
  );


  nor
  g3306
  (
    n3337,
    n2682,
    n2784,
    n2804,
    n3065
  );


  xnor
  g3307
  (
    n3272,
    n3080,
    n3090,
    n3094,
    n2763
  );


  xnor
  g3308
  (
    n3263,
    n2754,
    n3038,
    n2852,
    n2859
  );


  nand
  g3309
  (
    n3379,
    n3101,
    n3037,
    n3026,
    n3059
  );


  nor
  g3310
  (
    n3355,
    n3071,
    n3013,
    n2858,
    n3085
  );


  nand
  g3311
  (
    n3239,
    n2759,
    n2776,
    n2802
  );


  xnor
  g3312
  (
    n3299,
    n2764,
    n3014,
    n2787,
    n2784
  );


  nor
  g3313
  (
    n3282,
    n3025,
    n2771,
    n2758,
    n2827
  );


  or
  g3314
  (
    n3354,
    n2982,
    n3087,
    n3022,
    n2789
  );


  nor
  g3315
  (
    n3341,
    n2970,
    n3087,
    n3048,
    n2748
  );


  or
  g3316
  (
    n3353,
    n2792,
    n2688,
    n2809,
    n3057
  );


  nand
  g3317
  (
    n3273,
    n3055,
    n2797,
    n3100,
    n2799
  );


  and
  g3318
  (
    n3268,
    n2766,
    n2854,
    n2762,
    n2809
  );


  xor
  g3319
  (
    n3174,
    n3045,
    n2967,
    n2813,
    n2984
  );


  and
  g3320
  (
    n3335,
    n2756,
    n2749,
    n2765,
    n3052
  );


  nor
  g3321
  (
    n3369,
    n3088,
    n3054,
    n3046,
    n2773
  );


  nor
  g3322
  (
    n3284,
    n3028,
    n2812,
    n2785,
    n2997
  );


  nor
  g3323
  (
    n3331,
    n3048,
    n3055,
    n2820,
    n2986
  );


  nor
  g3324
  (
    n3404,
    n2997,
    n2771,
    n2971,
    n3050
  );


  nand
  g3325
  (
    n3391,
    n2977,
    n3092,
    n2684,
    n2793
  );


  and
  g3326
  (
    n3325,
    n3068,
    n2968,
    n2778,
    n2797
  );


  xnor
  g3327
  (
    n3271,
    n2808,
    n2986,
    n3038,
    n2818
  );


  and
  g3328
  (
    n3275,
    n2980,
    n2983,
    n2803,
    n2683
  );


  or
  g3329
  (
    n3386,
    n2853,
    n2796,
    n2859,
    n3082
  );


  xnor
  g3330
  (
    n3310,
    n2998,
    n2969,
    n2793,
    n3019
  );


  xor
  g3331
  (
    n3204,
    n3068,
    n2809,
    n2819,
    n2780
  );


  xor
  g3332
  (
    n3280,
    n3020,
    n2767,
    n3001,
    n2761
  );


  xnor
  g3333
  (
    n3202,
    n3082,
    n3044,
    n3016,
    n3098
  );


  or
  g3334
  (
    n3366,
    n2801,
    n3100,
    n3033
  );


  xnor
  g3335
  (
    n3193,
    n2783,
    n3065,
    n2749,
    n2808
  );


  xor
  g3336
  (
    n3292,
    n2757,
    n2801,
    n2771,
    n3000
  );


  xnor
  g3337
  (
    n3198,
    n2787,
    n2751,
    n3034,
    n2968
  );


  nand
  g3338
  (
    n3382,
    n3092,
    n3093,
    n2991,
    n2973
  );


  nor
  g3339
  (
    n3249,
    n2988,
    n2750,
    n2782,
    n2686
  );


  nor
  g3340
  (
    n3301,
    n2772,
    n2825,
    n3020,
    n3072
  );


  xor
  g3341
  (
    KeyWire_0_27,
    n3051,
    n3092,
    n2993
  );


  xor
  g3342
  (
    n3195,
    n3055,
    n2969,
    n2981,
    n2780
  );


  or
  g3343
  (
    n3278,
    n3042,
    n3095,
    n2995,
    n3064
  );


  nor
  g3344
  (
    n3398,
    n2816,
    n3076,
    n3000,
    n3063
  );


  xnor
  g3345
  (
    n3290,
    n2763,
    n3036,
    n2820,
    n3027
  );


  and
  g3346
  (
    n3332,
    n2810,
    n2783,
    n2686,
    n2974
  );


  xnor
  g3347
  (
    n3375,
    n2976,
    n3062,
    n3064,
    n3033
  );


  xor
  g3348
  (
    n3316,
    n2759,
    n2773,
    n2779,
    n3090
  );


  and
  g3349
  (
    n3389,
    n2988,
    n2988,
    n2856,
    n2993
  );


  nor
  g3350
  (
    n3185,
    n3039,
    n3080,
    n2783,
    n3066
  );


  and
  g3351
  (
    n3285,
    n2819,
    n2786,
    n2812,
    n2685
  );


  xnor
  g3352
  (
    n3407,
    n2794,
    n3017,
    n3094,
    n3051
  );


  or
  g3353
  (
    n3180,
    n3051,
    n3081,
    n2772,
    n3046
  );


  xnor
  g3354
  (
    n3257,
    n2798,
    n3096,
    n2754
  );


  or
  g3355
  (
    n3212,
    n2759,
    n2766,
    n2760,
    n3028
  );


  nand
  g3356
  (
    n3241,
    n2792,
    n3045,
    n3060,
    n3007
  );


  xnor
  g3357
  (
    n3224,
    n3009,
    n3046,
    n3058,
    n2970
  );


  nand
  g3358
  (
    n3396,
    n2986,
    n2973,
    n2971,
    n3059
  );


  xor
  g3359
  (
    n3327,
    n2976,
    n3002,
    n3057,
    n2853
  );


  nor
  g3360
  (
    n3311,
    n3094,
    n2687,
    n2761,
    n3028
  );


  xor
  g3361
  (
    n3351,
    n3062,
    n2837,
    n2763,
    n3057
  );


  xor
  g3362
  (
    n3230,
    n2825,
    n3018,
    n2982,
    n3060
  );


  or
  g3363
  (
    n3383,
    n3061,
    n3069,
    n2781,
    n3036
  );


  xor
  g3364
  (
    n3394,
    n2996,
    n2807,
    n2995,
    n2762
  );


  and
  g3365
  (
    n3203,
    n2818,
    n2975,
    n3074,
    n2025
  );


  xnor
  g3366
  (
    n3229,
    n3102,
    n2774,
    n3095,
    n3049
  );


  xnor
  g3367
  (
    n3385,
    n3031,
    n2823,
    n2777
  );


  or
  g3368
  (
    n3370,
    n3042,
    n3064,
    n2963,
    n2772
  );


  nor
  g3369
  (
    n3237,
    n2981,
    n2796,
    n3026,
    n3046
  );


  xnor
  g3370
  (
    n3225,
    n2811,
    n3035,
    n2972,
    n3010
  );


  nand
  g3371
  (
    n3245,
    n3004,
    n3054,
    n3070,
    n2774
  );


  nand
  g3372
  (
    n3340,
    n2781,
    n2025,
    n2813,
    n2807
  );


  xor
  g3373
  (
    n3343,
    n2822,
    n3007,
    n2763,
    n2684
  );


  nand
  g3374
  (
    n3184,
    n3023,
    n2806,
    n3025,
    n2965
  );


  or
  g3375
  (
    n3302,
    n2810,
    n2757,
    n2809,
    n2960
  );


  nor
  g3376
  (
    n3320,
    n3010,
    n2973,
    n2788,
    n2811
  );


  and
  g3377
  (
    n3416,
    n3180,
    n3197,
    n3193,
    n3183
  );


  nor
  g3378
  (
    n3411,
    n3189,
    n3182,
    n3191,
    n3200
  );


  xnor
  g3379
  (
    n3412,
    n3185,
    n3186,
    n3201,
    n3188
  );


  nor
  g3380
  (
    n3414,
    n3173,
    n3172,
    n3174,
    n3199
  );


  or
  g3381
  (
    n3417,
    n3196,
    n3194,
    n3195,
    n3198
  );


  xor
  g3382
  (
    n3415,
    n3176,
    n3184,
    n3192,
    n3177
  );


  xor
  g3383
  (
    n3413,
    n3187,
    n3178,
    n3190,
    n3181
  );


  xnor
  g3384
  (
    n3410,
    n3171,
    n3202,
    n3175,
    n3179
  );


  nand
  g3385
  (
    n3433,
    n3414,
    n2692
  );


  nor
  g3386
  (
    n3426,
    n2861,
    n3417
  );


  nand
  g3387
  (
    n3438,
    n3415,
    n2691
  );


  xor
  g3388
  (
    n3435,
    n2863,
    n3417
  );


  buf
  g3389
  (
    n3428,
    n2690
  );


  xor
  g3390
  (
    n3420,
    n3204,
    n3412
  );


  xnor
  g3391
  (
    n3431,
    n3416,
    n3203
  );


  xnor
  g3392
  (
    n3425,
    n2694,
    n2696
  );


  xor
  g3393
  (
    n3440,
    n2865,
    n3211
  );


  xnor
  g3394
  (
    n3442,
    n3206,
    n2695,
    n2862,
    n2027
  );


  and
  g3395
  (
    n3437,
    n3213,
    n3416,
    n3411,
    n3414
  );


  xor
  g3396
  (
    n3423,
    n3414,
    n2697,
    n3417,
    n3415
  );


  or
  g3397
  (
    n3443,
    n2865,
    n2689,
    n3205,
    n3413
  );


  or
  g3398
  (
    n3436,
    n2694,
    n3214,
    n3209,
    n2865
  );


  and
  g3399
  (
    n3418,
    n2698,
    n3212,
    n2691,
    n2860
  );


  xor
  g3400
  (
    n3427,
    n3416,
    n2695,
    n2862,
    n2860
  );


  xnor
  g3401
  (
    n3429,
    n3413,
    n2861,
    n3415
  );


  nand
  g3402
  (
    n3432,
    n3411,
    n2698,
    n3412,
    n2028
  );


  nand
  g3403
  (
    n3444,
    n2860,
    n2027,
    n2863,
    n3410
  );


  and
  g3404
  (
    n3430,
    n2693,
    n2863,
    n3417,
    n3415
  );


  or
  g3405
  (
    n3424,
    n3414,
    n3413,
    n2693,
    n2862
  );


  xnor
  g3406
  (
    n3421,
    n3216,
    n2864,
    n3416,
    n3412
  );


  xnor
  g3407
  (
    n3422,
    n3412,
    n3413,
    n2862,
    n2865
  );


  nand
  g3408
  (
    n3434,
    n3208,
    n2861,
    n2864,
    n3217
  );


  nor
  g3409
  (
    n3439,
    n2863,
    n3210,
    n2860,
    n2689
  );


  xor
  g3410
  (
    n3441,
    n2864,
    n3215,
    n2859,
    n2696
  );


  nand
  g3411
  (
    n3419,
    n3207,
    n2697,
    n2692,
    n2864
  );


  xnor
  g3412
  (
    n3464,
    n2895,
    n3140,
    n3139,
    n3116
  );


  or
  g3413
  (
    n3455,
    n3425,
    n3151,
    n2902,
    n3142
  );


  xor
  g3414
  (
    n3462,
    n2905,
    n3107,
    n2030,
    n3130
  );


  xnor
  g3415
  (
    n3456,
    n2029,
    n3127,
    n3428,
    n3161
  );


  xor
  g3416
  (
    KeyWire_0_51,
    n3429,
    n3147,
    n3143,
    n3432
  );


  xor
  g3417
  (
    n3543,
    n3138,
    n2031,
    n3419,
    n3136
  );


  xnor
  g3418
  (
    n3493,
    n3442,
    n3432,
    n3431,
    n3437
  );


  and
  g3419
  (
    n3496,
    n3103,
    n3131,
    n3148,
    n3162
  );


  and
  g3420
  (
    n3482,
    n3125,
    n3157,
    n3160,
    n3444
  );


  xnor
  g3421
  (
    n3519,
    n2028,
    n3440,
    n3429,
    n3110
  );


  xnor
  g3422
  (
    n3507,
    n3436,
    n3158,
    n3154,
    n3428
  );


  or
  g3423
  (
    n3520,
    n3154,
    n3140,
    n3118,
    n2897
  );


  nor
  g3424
  (
    n3514,
    n2031,
    n3119,
    n3159,
    n3109
  );


  or
  g3425
  (
    n3501,
    n3122,
    n3142,
    n3432,
    n3111
  );


  xnor
  g3426
  (
    n3466,
    n3155,
    n3123,
    n3427
  );


  xor
  g3427
  (
    n3459,
    n3424,
    n3114,
    n3141,
    n3419
  );


  or
  g3428
  (
    n3517,
    n3104,
    n3129,
    n2902,
    n3117
  );


  xor
  g3429
  (
    n3502,
    n3113,
    n3109,
    n3420,
    n2900
  );


  or
  g3430
  (
    n3535,
    n3436,
    n3130,
    n3157,
    n3144
  );


  and
  g3431
  (
    n3508,
    n3433,
    n3124,
    n3161,
    n3117
  );


  and
  g3432
  (
    n3481,
    n3107,
    n3442,
    n3424,
    n3440
  );


  nor
  g3433
  (
    n3523,
    n3442,
    n3149,
    n3422,
    n3122
  );


  xnor
  g3434
  (
    n3542,
    n2896,
    n2897,
    n3432,
    n3418
  );


  nand
  g3435
  (
    n3448,
    n3159,
    n2039,
    n3117,
    n3104
  );


  nand
  g3436
  (
    n3536,
    n3106,
    n3132,
    n2892,
    n2903
  );


  xnor
  g3437
  (
    n3479,
    n3425,
    n3132,
    n3143,
    n2898
  );


  xor
  g3438
  (
    n3494,
    n3127,
    n3428,
    n2040,
    n3140
  );


  or
  g3439
  (
    n3503,
    n3114,
    n2898,
    n2900,
    n3423
  );


  or
  g3440
  (
    n3518,
    n2894,
    n2035,
    n3444,
    n3437
  );


  xor
  g3441
  (
    n3546,
    n3131,
    n3430,
    n2901,
    n3128
  );


  nand
  g3442
  (
    n3510,
    n2900,
    n2899,
    n3106,
    n3119
  );


  nor
  g3443
  (
    n3537,
    n3421,
    n3139,
    n3441
  );


  xnor
  g3444
  (
    KeyWire_0_55,
    n3422,
    n3127,
    n2903,
    n3154
  );


  xor
  g3445
  (
    n3526,
    n3121,
    n3126,
    n3438,
    n2893
  );


  xor
  g3446
  (
    n3528,
    n3421,
    n3109,
    n3120,
    n3150
  );


  and
  g3447
  (
    n3495,
    n2901,
    n2029,
    n3107,
    n3142
  );


  or
  g3448
  (
    n3498,
    n3443,
    n3126,
    n3160,
    n2895
  );


  and
  g3449
  (
    n3445,
    n3123,
    n3137,
    n2902,
    n3145
  );


  xor
  g3450
  (
    n3463,
    n3126,
    n3434,
    n3142,
    n3443
  );


  xnor
  g3451
  (
    n3506,
    n3122,
    n3158,
    n3146,
    n3126
  );


  nor
  g3452
  (
    n3516,
    n3149,
    n3431,
    n3108,
    n3133
  );


  xnor
  g3453
  (
    n3468,
    n3158,
    n3135,
    n3439,
    n3111
  );


  xor
  g3454
  (
    n3487,
    n3137,
    n3141,
    n3160,
    n3427
  );


  and
  g3455
  (
    n3476,
    n3149,
    n3438,
    n3139,
    n3158
  );


  nor
  g3456
  (
    n3451,
    n3151,
    n3156,
    n3145,
    n3112
  );


  or
  g3457
  (
    n3458,
    n3145,
    n3161,
    n3425,
    n2032
  );


  nand
  g3458
  (
    n3497,
    n3116,
    n3120,
    n3441,
    n3149
  );


  nor
  g3459
  (
    n3469,
    n2890,
    n3440,
    n3115,
    n3121
  );


  xor
  g3460
  (
    n3533,
    n3160,
    n3116,
    n3431,
    n2904
  );


  xnor
  g3461
  (
    n3488,
    n2902,
    n2037,
    n3433,
    n3144
  );


  nand
  g3462
  (
    n3515,
    n2903,
    n3108,
    n3104,
    n3419
  );


  xor
  g3463
  (
    n3484,
    n3138,
    n3105,
    n2893,
    n3418
  );


  xor
  g3464
  (
    n3473,
    n2035,
    n3443,
    n3155,
    n3138
  );


  nand
  g3465
  (
    n3499,
    n2901,
    n3136,
    n3121,
    n2033
  );


  xor
  g3466
  (
    n3477,
    n2899,
    n3103,
    n3118,
    n3128
  );


  xor
  g3467
  (
    n3449,
    n3106,
    n3424,
    n3146,
    n3150
  );


  or
  g3468
  (
    n3511,
    n3125,
    n3117,
    n3157,
    n2905
  );


  or
  g3469
  (
    n3551,
    n2894,
    n3155,
    n3436,
    n3146
  );


  xor
  g3470
  (
    n3478,
    n2040,
    n2904,
    n3424,
    n3148
  );


  or
  g3471
  (
    n3544,
    n3426,
    n3423,
    n3113,
    n2897
  );


  nand
  g3472
  (
    n3483,
    n3130,
    n3439,
    n3133,
    n3105
  );


  xor
  g3473
  (
    n3491,
    n3147,
    n3147,
    n2037,
    n3429
  );


  or
  g3474
  (
    n3525,
    n2036,
    n3423,
    n3129,
    n3444
  );


  nand
  g3475
  (
    n3490,
    n3440,
    n3121,
    n3157,
    n3134
  );


  nor
  g3476
  (
    n3540,
    n2895,
    n3422,
    n3443,
    n3420
  );


  xnor
  g3477
  (
    n3538,
    n2893,
    n2892,
    n3427,
    n3435
  );


  nand
  g3478
  (
    n3549,
    n3120,
    n3131,
    n3430,
    n3115
  );


  nor
  g3479
  (
    n3545,
    n3426,
    n3116,
    n3132,
    n3433
  );


  nor
  g3480
  (
    n3492,
    n3104,
    n2894,
    n3430,
    n3441
  );


  and
  g3481
  (
    n3457,
    n3111,
    n3110,
    n3127,
    n3135
  );


  nand
  g3482
  (
    n3539,
    n3437,
    n3133,
    n3153,
    n2036
  );


  nor
  g3483
  (
    n3552,
    n3156,
    n3435,
    n3430,
    n2901
  );


  xnor
  g3484
  (
    n3472,
    n3423,
    n3156,
    n3153,
    n3124
  );


  nor
  g3485
  (
    n3504,
    n3131,
    n3136,
    n3159,
    n3418
  );


  xor
  g3486
  (
    n3446,
    n2890,
    n3426,
    n3122,
    n3141
  );


  xor
  g3487
  (
    n3447,
    n3114,
    n3439,
    n2891,
    n3124
  );


  nor
  g3488
  (
    n3461,
    n3439,
    n3145,
    n3438,
    n2896
  );


  xnor
  g3489
  (
    n3470,
    n2895,
    n3146,
    n3108,
    n2898
  );


  and
  g3490
  (
    n3534,
    n3128,
    n3435,
    n2900,
    n3151
  );


  nor
  g3491
  (
    n3454,
    n3110,
    n3115,
    n3109,
    n3130
  );


  xnor
  g3492
  (
    n3460,
    n3159,
    n2893,
    n3444,
    n3111
  );


  xor
  g3493
  (
    n3550,
    n2897,
    n3429,
    n2033,
    n3426
  );


  xor
  g3494
  (
    n3527,
    n3140,
    n3152,
    n3132,
    n3115
  );


  xor
  g3495
  (
    n3541,
    n3148,
    n3112,
    n2896,
    n3161
  );


  xnor
  g3496
  (
    n3521,
    n3144,
    n3125,
    n2894,
    n2030
  );


  xnor
  g3497
  (
    n3547,
    n2038,
    n2891,
    n2898,
    n2904
  );


  xor
  g3498
  (
    n3512,
    n2892,
    n3139,
    n3418,
    n2891
  );


  or
  g3499
  (
    n3509,
    n3138,
    n3136,
    n3420,
    n3118
  );


  xor
  g3500
  (
    n3452,
    n3133,
    n3129,
    n3421,
    n2905
  );


  nand
  g3501
  (
    n3450,
    n3107,
    n3434,
    n3105,
    n3151
  );


  and
  g3502
  (
    n3548,
    n3425,
    n3436,
    n3144,
    n2038
  );


  nor
  g3503
  (
    n3453,
    n3119,
    n3152,
    n3438,
    n3112
  );


  xnor
  g3504
  (
    n3500,
    n3152,
    n3125,
    n2899,
    n3427
  );


  xnor
  g3505
  (
    n3489,
    n3134,
    n3421,
    n2039,
    n3150
  );


  and
  g3506
  (
    n3474,
    n3123,
    n3143,
    n3113,
    n2034
  );


  xor
  g3507
  (
    n3486,
    n3431,
    n3141,
    n3134,
    n2903
  );


  or
  g3508
  (
    n3532,
    n3108,
    n2892,
    n3154,
    n3135
  );


  nor
  g3509
  (
    n3505,
    n3106,
    n3153,
    n3437,
    n3112
  );


  nand
  g3510
  (
    n3485,
    n3143,
    n3152,
    n3434,
    n3433
  );


  or
  g3511
  (
    n3531,
    n2891,
    n3124,
    n2905,
    n3442
  );


  xor
  g3512
  (
    n3513,
    n2899,
    n3148,
    n3128,
    n3137
  );


  nor
  g3513
  (
    n3467,
    n3134,
    n3155,
    n3150,
    n2032
  );


  nand
  g3514
  (
    n3480,
    n3120,
    n3110,
    n3428,
    n3420
  );


  nor
  g3515
  (
    n3530,
    n3114,
    n2904,
    n3422,
    n3434
  );


  xnor
  g3516
  (
    n3522,
    n3419,
    n2890,
    n3119
  );


  nand
  g3517
  (
    n3529,
    n3147,
    n2034,
    n3137,
    n3156
  );


  xor
  g3518
  (
    n3471,
    n2896,
    n3105,
    n3129,
    n3435
  );


  or
  g3519
  (
    n3475,
    n3153,
    n3135,
    n3113,
    n3118
  );


  xor
  g3520
  (
    n3571,
    n3243,
    n3266,
    n3288,
    n3225
  );


  nand
  g3521
  (
    n3561,
    n3261,
    n3295,
    n3287,
    n3257
  );


  nor
  g3522
  (
    n3553,
    n3256,
    n3464,
    n3234,
    n3300
  );


  xnor
  g3523
  (
    n3564,
    n3451,
    n3228,
    n3246,
    n3263
  );


  xnor
  g3524
  (
    n3569,
    n3283,
    n3239,
    n3463,
    n3231
  );


  nand
  g3525
  (
    n3573,
    n3455,
    n3218,
    n3469,
    n3279
  );


  nand
  g3526
  (
    n3580,
    n3230,
    n3268,
    n3277,
    n3249
  );


  xnor
  g3527
  (
    n3566,
    n3294,
    n3456,
    n3301,
    n3220
  );


  xor
  g3528
  (
    n3563,
    n3445,
    n3298,
    n3252,
    n3258
  );


  xor
  g3529
  (
    n3554,
    n3461,
    n3465,
    n3267,
    n3269
  );


  nand
  g3530
  (
    n3576,
    n3253,
    n3285,
    n3470,
    n3289
  );


  or
  g3531
  (
    n3578,
    n3227,
    n3238,
    n3233,
    n3471
  );


  or
  g3532
  (
    n3556,
    n3254,
    n3453,
    n3275,
    n3292
  );


  xnor
  g3533
  (
    KeyWire_0_57,
    n3222,
    n3458,
    n3280,
    n3446
  );


  nand
  g3534
  (
    n3562,
    n3235,
    n3457,
    n3251,
    n3255
  );


  and
  g3535
  (
    n3570,
    n3448,
    n3274,
    n3223,
    n3472
  );


  nor
  g3536
  (
    n3567,
    n3242,
    n3449,
    n3260,
    n3270
  );


  nand
  g3537
  (
    n3558,
    n3454,
    n3286,
    n3293,
    n3241
  );


  or
  g3538
  (
    n3579,
    n3265,
    n3447,
    n3467,
    n3229
  );


  and
  g3539
  (
    n3557,
    n3276,
    n3297,
    n3272,
    n3262
  );


  xor
  g3540
  (
    n3565,
    n3466,
    n3245,
    n3450,
    n3460
  );


  and
  g3541
  (
    n3572,
    n3278,
    n3299,
    n3248,
    n3271
  );


  nand
  g3542
  (
    n3575,
    n3459,
    n3250,
    n3226,
    n3462
  );


  or
  g3543
  (
    n3568,
    n3264,
    n3247,
    n3290,
    n3244
  );


  xnor
  g3544
  (
    n3555,
    n3273,
    n3284,
    n3468,
    n3221
  );


  xor
  g3545
  (
    n3574,
    n3224,
    n3240,
    n3291,
    n3282
  );


  nand
  g3546
  (
    n3577,
    n3232,
    n3237,
    n3296,
    n3219
  );


  xor
  g3547
  (
    n3560,
    n3281,
    n3259,
    n3236,
    n3452
  );


  or
  g3548
  (
    n3591,
    n3328,
    n3341,
    n3168,
    n3558
  );


  xor
  g3549
  (
    n3583,
    n3553,
    n3165,
    n3166,
    n3557
  );


  nor
  g3550
  (
    n3615,
    n3342,
    n3163,
    n3333,
    n3560
  );


  nand
  g3551
  (
    n3587,
    n3556,
    n3312,
    n3554,
    n3162
  );


  xnor
  g3552
  (
    n3593,
    n3553,
    n3332,
    n3559,
    n3162
  );


  nor
  g3553
  (
    n3588,
    n3555,
    n3307,
    n3319,
    n2046
  );


  nor
  g3554
  (
    n3611,
    n2045,
    n3559,
    n3308,
    n3553
  );


  xnor
  g3555
  (
    n3605,
    n3344,
    n3169,
    n3555
  );


  xnor
  g3556
  (
    n3601,
    n3346,
    n2048,
    n3560,
    n3164
  );


  or
  g3557
  (
    n3612,
    n3315,
    n3556,
    n3320,
    n3561
  );


  xnor
  g3558
  (
    n3594,
    n3349,
    n3554,
    n3316,
    n2044
  );


  or
  g3559
  (
    n3604,
    n2044,
    n3559,
    n3167,
    n3168
  );


  nor
  g3560
  (
    n3586,
    n3339,
    n3350,
    n3164,
    n3170
  );


  xnor
  g3561
  (
    n3597,
    n3555,
    n3167,
    n3325,
    n3304
  );


  xor
  g3562
  (
    n3596,
    n2045,
    n3166,
    n3354,
    n3330
  );


  nor
  g3563
  (
    n3606,
    n3168,
    n3554,
    n2041,
    n2043
  );


  nand
  g3564
  (
    n3610,
    n3170,
    n2049,
    n2047,
    n3322
  );


  xnor
  g3565
  (
    n3599,
    n2041,
    n3311,
    n3556,
    n3318
  );


  or
  g3566
  (
    n3598,
    n3557,
    n3351,
    n3561,
    n3163
  );


  nor
  g3567
  (
    n3600,
    n3347,
    n3164,
    n3167,
    n3336
  );


  xnor
  g3568
  (
    n3585,
    n3560,
    n3303,
    n3165,
    n3553
  );


  xor
  g3569
  (
    n3581,
    n3313,
    n3166,
    n3340,
    n3326
  );


  nand
  g3570
  (
    n3608,
    n3164,
    n3337,
    n3556,
    n3331
  );


  and
  g3571
  (
    n3603,
    n2043,
    n3317,
    n3558,
    n3321
  );


  nor
  g3572
  (
    n3609,
    n3163,
    n3348,
    n3558,
    n3306
  );


  xnor
  g3573
  (
    n3602,
    n3302,
    n3168,
    n3352,
    n3335
  );


  or
  g3574
  (
    n3607,
    n3560,
    n3305,
    n3167,
    n3169
  );


  or
  g3575
  (
    n3614,
    n3323,
    n2047,
    n3165,
    n3345
  );


  and
  g3576
  (
    n3584,
    n2042,
    n3163,
    n2048,
    n3559
  );


  nand
  g3577
  (
    n3613,
    n3329,
    n3314,
    n2042,
    n3169
  );


  or
  g3578
  (
    n3592,
    n3561,
    n3310,
    n3309,
    n3324
  );


  nand
  g3579
  (
    n3595,
    n3170,
    n3353,
    n3338,
    n3557
  );


  nand
  g3580
  (
    n3582,
    n2046,
    n3166,
    n3169,
    n3327
  );


  and
  g3581
  (
    n3589,
    n3558,
    n3343,
    n3162,
    n3334
  );


  xor
  g3582
  (
    n3590,
    n3170,
    n3554,
    n3165,
    n3557
  );


  and
  g3583
  (
    n3624,
    n3586,
    n3367,
    n3371,
    n3361
  );


  nand
  g3584
  (
    n3628,
    n3586,
    n3378,
    n3581,
    n3377
  );


  or
  g3585
  (
    n3621,
    n3357,
    n3583,
    n3355,
    n3371
  );


  nand
  g3586
  (
    n3629,
    n3368,
    n3374,
    n3369,
    n3375
  );


  or
  g3587
  (
    n3625,
    n3361,
    n3582,
    n3360
  );


  xnor
  g3588
  (
    n3626,
    n3369,
    n3588,
    n3364,
    n3376
  );


  nor
  g3589
  (
    n3630,
    n3583,
    n3368,
    n3582,
    n3359
  );


  and
  g3590
  (
    n3617,
    n3584,
    n3373,
    n3367,
    n3376
  );


  and
  g3591
  (
    n3616,
    n3374,
    n3363,
    n3378,
    n3366
  );


  xnor
  g3592
  (
    n3623,
    n3365,
    n3363,
    n3581,
    n3375
  );


  xor
  g3593
  (
    n3622,
    n3587,
    n3372,
    n3365,
    n3585
  );


  or
  g3594
  (
    n3618,
    n3370,
    n3366,
    n3377,
    n3373
  );


  xor
  g3595
  (
    n3627,
    n3370,
    n3364,
    n3372,
    n3587
  );


  xor
  g3596
  (
    n3620,
    n3585,
    n3356,
    n3358
  );


  and
  g3597
  (
    n3619,
    n3362,
    n3362,
    n3584,
    n3359
  );


  and
  g3598
  (
    n3641,
    n3630,
    n3482,
    n2052,
    n3487
  );


  xor
  g3599
  (
    n3631,
    n3476,
    n3626,
    n3499,
    n2699
  );


  xnor
  g3600
  (
    n3637,
    n3620,
    n3491,
    n3477,
    n3501
  );


  xor
  g3601
  (
    n3642,
    n3497,
    n2055,
    n3624,
    n3621
  );


  nand
  g3602
  (
    n3640,
    n3622,
    n3625,
    n2054,
    n3478
  );


  and
  g3603
  (
    n3636,
    n2051,
    n3492,
    n3488,
    n3474
  );


  nor
  g3604
  (
    n3635,
    n3623,
    n3481,
    n3480,
    n3617
  );


  nor
  g3605
  (
    n3634,
    n3628,
    n3485,
    n3479,
    n3494
  );


  and
  g3606
  (
    n3646,
    n2701,
    n3616,
    n3619,
    n3629
  );


  xor
  g3607
  (
    n3633,
    n2055,
    n2053,
    n2056,
    n3484
  );


  xnor
  g3608
  (
    n3632,
    n2050,
    n3486,
    n2700,
    n3618
  );


  and
  g3609
  (
    n3638,
    n2050,
    n3496,
    n3627,
    n2052
  );


  xor
  g3610
  (
    n3643,
    n2049,
    n3489,
    n3498,
    n3493
  );


  xor
  g3611
  (
    n3639,
    n2700,
    n2056,
    n3500,
    n3502
  );


  xnor
  g3612
  (
    n3645,
    n3495,
    n2701,
    n3483,
    n2054
  );


  or
  g3613
  (
    n3647,
    n3630,
    n2053,
    n3490,
    n2699
  );


  nor
  g3614
  (
    n3644,
    n2051,
    n3475,
    n3630,
    n3473
  );


  nand
  g3615
  (
    n3658,
    n3637,
    n2059,
    n3644,
    n2078
  );


  and
  g3616
  (
    n3661,
    n3638,
    n2060,
    n2069,
    n3633
  );


  and
  g3617
  (
    n3650,
    n2069,
    n3642,
    n2072,
    n2066
  );


  nand
  g3618
  (
    n3654,
    n2072,
    n2078,
    n3632,
    n2057
  );


  nor
  g3619
  (
    n3657,
    n3645,
    n2079,
    n3639,
    n2076
  );


  nand
  g3620
  (
    n3653,
    n2057,
    n2071,
    n2063
  );


  nor
  g3621
  (
    KeyWire_0_53,
    n2063,
    n2075,
    n2058,
    n2068
  );


  and
  g3622
  (
    n3659,
    n3643,
    n2061,
    n2073,
    n3634
  );


  xnor
  g3623
  (
    n3660,
    n2070,
    n2068,
    n2064,
    n3635
  );


  nand
  g3624
  (
    n3662,
    n2073,
    n2061,
    n2065,
    n2066
  );


  xor
  g3625
  (
    n3655,
    n2058,
    n2064,
    n2062,
    n3631
  );


  nor
  g3626
  (
    n3648,
    n2077,
    n2074,
    n3641,
    n2059
  );


  and
  g3627
  (
    n3649,
    n2070,
    n2067,
    n2077
  );


  nor
  g3628
  (
    n3651,
    n2075,
    n2074,
    n3636,
    n2060
  );


  or
  g3629
  (
    n3656,
    n2065,
    n2076,
    n3640,
    n2062
  );


  xor
  g3630
  (
    n3676,
    n3655,
    n3660,
    n3593,
    n2706
  );


  nand
  g3631
  (
    n3675,
    n3661,
    n3662,
    n3594,
    n3589
  );


  and
  g3632
  (
    n3672,
    n3591,
    n3594,
    n2708,
    n3658
  );


  nor
  g3633
  (
    n3677,
    n2708,
    n3592,
    n3653,
    n3648
  );


  nor
  g3634
  (
    n3664,
    n3600,
    n2704,
    n3651,
    n3597
  );


  xor
  g3635
  (
    n3668,
    n3593,
    n3592,
    n3590,
    n2709
  );


  nor
  g3636
  (
    n3669,
    n2702,
    n2707,
    n2709,
    n3591
  );


  xnor
  g3637
  (
    n3674,
    n2705,
    n3588,
    n2706,
    n3601
  );


  xor
  g3638
  (
    n3667,
    n3600,
    n3657,
    n3589,
    n3596
  );


  or
  g3639
  (
    n3671,
    n3598,
    n3595,
    n3590,
    n3654
  );


  xor
  g3640
  (
    n3673,
    n2707,
    n2702,
    n3598,
    n3652
  );


  nand
  g3641
  (
    n3670,
    n3596,
    n3659,
    n3595,
    n3656
  );


  or
  g3642
  (
    n3663,
    n3650,
    n2703,
    n3597,
    n3649
  );


  nor
  g3643
  (
    n3665,
    n2703,
    n3599,
    n2704,
    n2711
  );


  or
  g3644
  (
    n3666,
    n3599,
    n2705,
    n2710
  );


  not
  g3645
  (
    n3734,
    n3677
  );


  not
  g3646
  (
    n3726,
    n3575
  );


  not
  g3647
  (
    n3721,
    n3676
  );


  not
  g3648
  (
    n3717,
    n3615
  );


  buf
  g3649
  (
    n3678,
    n2080
  );


  not
  g3650
  (
    n3687,
    n2717
  );


  not
  g3651
  (
    n3684,
    n3666
  );


  not
  g3652
  (
    n3703,
    n3606
  );


  not
  g3653
  (
    n3730,
    n3568
  );


  nand
  g3654
  (
    n3695,
    n3579,
    n3670,
    n3610,
    n3561
  );


  or
  g3655
  (
    n3714,
    n3665,
    n3565,
    n3675,
    n2718
  );


  nor
  g3656
  (
    n3682,
    n3673,
    n3674,
    n3580,
    n3614
  );


  nor
  g3657
  (
    n3693,
    n3675,
    n3570,
    n2083,
    n2724
  );


  xnor
  g3658
  (
    n3735,
    n3665,
    n3563,
    n3663,
    n3664
  );


  xor
  g3659
  (
    n3696,
    n3564,
    n3601,
    n3607,
    n3565
  );


  xnor
  g3660
  (
    n3722,
    n2718,
    n3580,
    n3677,
    n2716
  );


  xor
  g3661
  (
    n3718,
    n3664,
    n3672,
    n2079,
    n3669
  );


  nor
  g3662
  (
    n3725,
    n2712,
    n3669,
    n3665,
    n3668
  );


  nor
  g3663
  (
    n3731,
    n3674,
    n3576,
    n3577,
    n3663
  );


  nor
  g3664
  (
    n3698,
    n3577,
    n3562,
    n3612,
    n2084
  );


  nor
  g3665
  (
    n3681,
    n3672,
    n3673,
    n3578,
    n2713
  );


  xnor
  g3666
  (
    n3729,
    n3675,
    n2086,
    n3562,
    n2081
  );


  xnor
  g3667
  (
    n3700,
    n3673,
    n3568,
    n3603,
    n3612
  );


  xnor
  g3668
  (
    n3716,
    n3574,
    n2086,
    n3673,
    n3668
  );


  xnor
  g3669
  (
    n3715,
    n2724,
    n3669,
    n3572,
    n3609
  );


  nor
  g3670
  (
    n3683,
    n3563,
    n3602,
    n3575,
    n3670
  );


  nor
  g3671
  (
    n3724,
    n3667,
    n2719,
    n3569,
    n3611
  );


  nor
  g3672
  (
    n3733,
    n3603,
    n3604,
    n3569,
    n3564
  );


  or
  g3673
  (
    n3719,
    n3571,
    n2725,
    n2719,
    n3573
  );


  or
  g3674
  (
    n3697,
    n3573,
    n3609,
    n3666,
    n3571
  );


  xnor
  g3675
  (
    n3723,
    n2713,
    n3663,
    n3615,
    n3607
  );


  xnor
  g3676
  (
    n3680,
    n3665,
    n3577,
    n3674,
    n3576
  );


  and
  g3677
  (
    n3701,
    n3567,
    n2715,
    n3572,
    n3671
  );


  or
  g3678
  (
    n3685,
    n2726,
    n2726,
    n3663,
    n3578
  );


  xor
  g3679
  (
    n3707,
    n3572,
    n3675,
    n3613,
    n3564
  );


  nor
  g3680
  (
    n3705,
    n3578,
    n2722,
    n3566,
    n3574
  );


  xnor
  g3681
  (
    n3709,
    n3569,
    n3564,
    n3608,
    n3570
  );


  nor
  g3682
  (
    n3712,
    n3677,
    n3566,
    n2081,
    n3576
  );


  nand
  g3683
  (
    n3688,
    n3575,
    n3608,
    n3677,
    n3570
  );


  nor
  g3684
  (
    n3720,
    n3574,
    n2722,
    n3606,
    n3666
  );


  and
  g3685
  (
    n3692,
    n2714,
    n3670,
    n3580,
    n3566
  );


  and
  g3686
  (
    n3708,
    n2720,
    n3574,
    n3563,
    n3613
  );


  xor
  g3687
  (
    n3689,
    n2085,
    n3567,
    n2723,
    n3569
  );


  xor
  g3688
  (
    n3737,
    n3670,
    n3571,
    n3580,
    n2083
  );


  and
  g3689
  (
    n3728,
    n3563,
    n3667,
    n3614,
    n3570
  );


  nand
  g3690
  (
    n3686,
    n3562,
    n3579,
    n3566,
    n2723
  );


  or
  g3691
  (
    n3710,
    n3578,
    n2727,
    n2082,
    n3664
  );


  or
  g3692
  (
    n3713,
    n3669,
    n3571,
    n3602,
    n3667
  );


  xnor
  g3693
  (
    n3727,
    n2717,
    n2714,
    n3573,
    n3562
  );


  xor
  g3694
  (
    n3679,
    n2720,
    n2082,
    n3676,
    n3573
  );


  nand
  g3695
  (
    n3690,
    n2711,
    n3610,
    n2725,
    n3674
  );


  or
  g3696
  (
    n3736,
    n3671,
    n3671,
    n3576,
    n3572
  );


  nor
  g3697
  (
    n3691,
    n2716,
    n3567,
    n3568,
    n2721
  );


  or
  g3698
  (
    n3699,
    n3671,
    n3568,
    n2721,
    n3565
  );


  xor
  g3699
  (
    n3702,
    n3672,
    n3605,
    n3575,
    n3668
  );


  xnor
  g3700
  (
    n3706,
    n3579,
    n3604,
    n3664,
    n2712
  );


  or
  g3701
  (
    n3704,
    n2715,
    n3567,
    n3577,
    n3565
  );


  xor
  g3702
  (
    n3711,
    n3672,
    n3668,
    n3676,
    n3667
  );


  xor
  g3703
  (
    n3694,
    n2085,
    n3579,
    n2084,
    n3676
  );


  nand
  g3704
  (
    n3732,
    n3666,
    n3611,
    n2080,
    n3605
  );


  nand
  g3705
  (
    n3757,
    n3723,
    n3727
  );


  or
  g3706
  (
    n3759,
    n3717,
    n3726
  );


  or
  g3707
  (
    n3738,
    n3679,
    n3694
  );


  nor
  g3708
  (
    KeyWire_0_45,
    n3682,
    n3727
  );


  xor
  g3709
  (
    n3760,
    n3708,
    n3701
  );


  nand
  g3710
  (
    n3762,
    n3716,
    n3725
  );


  or
  g3711
  (
    n3766,
    n3692,
    n3721
  );


  xor
  g3712
  (
    n3741,
    n3695,
    n3726
  );


  xor
  g3713
  (
    n3742,
    n3728,
    n3687
  );


  or
  g3714
  (
    n3761,
    n3711,
    n3683
  );


  xnor
  g3715
  (
    n3749,
    n3693,
    n3691
  );


  nor
  g3716
  (
    n3746,
    n3718,
    n3714
  );


  and
  g3717
  (
    n3740,
    n3696,
    n3724
  );


  xnor
  g3718
  (
    n3752,
    n3715,
    n3689
  );


  or
  g3719
  (
    n3755,
    n3713,
    n3710
  );


  nand
  g3720
  (
    n3739,
    n3702,
    n3681
  );


  and
  g3721
  (
    n3753,
    n3697,
    n3690
  );


  xnor
  g3722
  (
    n3751,
    n3685,
    n3727
  );


  nand
  g3723
  (
    n3764,
    n3709,
    n3719
  );


  nand
  g3724
  (
    n3747,
    n3678,
    n3712
  );


  xor
  g3725
  (
    n3748,
    n3686,
    n3722
  );


  xor
  g3726
  (
    n3758,
    n3728,
    n3684
  );


  and
  g3727
  (
    n3763,
    n3726,
    n3688
  );


  and
  g3728
  (
    n3745,
    n3707,
    n3720
  );


  xor
  g3729
  (
    KeyWire_0_25,
    n3698,
    n3680
  );


  or
  g3730
  (
    n3765,
    n3705,
    n3727
  );


  xor
  g3731
  (
    n3754,
    n3706,
    n3699
  );


  nand
  g3732
  (
    n3744,
    n3726,
    n3704
  );


  and
  g3733
  (
    n3743,
    n3703,
    n3700
  );


  and
  g3734
  (
    n3776,
    n3738,
    n2733,
    n3753,
    n3755
  );


  and
  g3735
  (
    n3773,
    n2727,
    n3761,
    n2732,
    n2728
  );


  xor
  g3736
  (
    n3771,
    n3744,
    n3759,
    n3745,
    n2730
  );


  xor
  g3737
  (
    n3770,
    n2729,
    n3749,
    n3742,
    n3746
  );


  nand
  g3738
  (
    n3772,
    n2731,
    n3756,
    n2732,
    n3760
  );


  or
  g3739
  (
    n3774,
    n3751,
    n2731,
    n3757,
    n3747
  );


  nand
  g3740
  (
    n3767,
    n3748,
    n3740,
    n2734
  );


  or
  g3741
  (
    n3769,
    n3750,
    n3739,
    n2735,
    n2733
  );


  and
  g3742
  (
    n3768,
    n3754,
    n2728,
    n3752,
    n3758
  );


  or
  g3743
  (
    n3775,
    n3743,
    n2729,
    n2730,
    n3741
  );


  buf
  g3744
  (
    n3781,
    n3772
  );


  buf
  g3745
  (
    n3778,
    n3646
  );


  buf
  g3746
  (
    n3777,
    n3647
  );


  buf
  g3747
  (
    n3782,
    n3773
  );


  xnor
  g3748
  (
    n3779,
    n2088,
    n2087,
    n3769,
    n3774
  );


  xnor
  g3749
  (
    n3780,
    n2088,
    n2087,
    n3770,
    n3771
  );


  or
  g3750
  (
    n3793,
    n3778,
    n3733,
    n3730,
    n3777
  );


  and
  g3751
  (
    n3788,
    n3737,
    n3729,
    n3734,
    n3732
  );


  and
  g3752
  (
    n3786,
    n3733,
    n3782,
    n3729,
    n3732
  );


  or
  g3753
  (
    n3784,
    n3735,
    n3778,
    n3730,
    n3728
  );


  or
  g3754
  (
    n3785,
    n3731,
    n3732,
    n3736,
    n3733
  );


  and
  g3755
  (
    n3790,
    n3781,
    n3781,
    n3736,
    n3780
  );


  or
  g3756
  (
    n3794,
    n3779,
    n3731,
    n3735
  );


  xnor
  g3757
  (
    n3789,
    n3728,
    n3736,
    n3780,
    n3731
  );


  xor
  g3758
  (
    n3792,
    n3735,
    n3730,
    n3733,
    n3779
  );


  xnor
  g3759
  (
    n3783,
    n3734,
    n3777,
    n3730,
    n3729
  );


  or
  g3760
  (
    n3791,
    n3734,
    n3737,
    n3736,
    n3732
  );


  or
  g3761
  (
    n3787,
    n3735,
    n3729,
    n3782,
    n3734
  );


  buf
  g3762
  (
    n3797,
    n3793
  );


  not
  g3763
  (
    n3798,
    n3790
  );


  not
  g3764
  (
    n3796,
    n3792
  );


  or
  g3765
  (
    n3795,
    n3791,
    n2089
  );


  and
  g3766
  (
    n3807,
    n2096,
    n3387,
    n3798,
    n3385
  );


  xnor
  g3767
  (
    n3802,
    n3797,
    n3795,
    n3384,
    n2095
  );


  xnor
  g3768
  (
    n3805,
    n3392,
    n2094,
    n3388
  );


  or
  g3769
  (
    n3801,
    n3390,
    n2090,
    n3386,
    n3392
  );


  nand
  g3770
  (
    KeyWire_0_15,
    n3380,
    n3379,
    n3383,
    n3387
  );


  xor
  g3771
  (
    n3799,
    n3389,
    n3389,
    n3380,
    n2735
  );


  or
  g3772
  (
    n3809,
    n3798,
    n3797,
    n3382
  );


  xnor
  g3773
  (
    n3810,
    n3391,
    n3383,
    n2090,
    n3795
  );


  nand
  g3774
  (
    n3813,
    n3796,
    n3382,
    n3798,
    n3795
  );


  xor
  g3775
  (
    n3806,
    n2091,
    n3385,
    n3390,
    n2096
  );


  or
  g3776
  (
    n3811,
    n3388,
    n2093,
    n3379,
    n3796
  );


  or
  g3777
  (
    n3803,
    n3384,
    n2092,
    n2089,
    n3386
  );


  xnor
  g3778
  (
    n3800,
    n3381,
    n3391,
    n3798,
    n3796
  );


  and
  g3779
  (
    n3808,
    n2091,
    n3381,
    n3797,
    n2097
  );


  and
  g3780
  (
    n3804,
    n2093,
    n2095,
    n3796,
    n2092
  );


  not
  g3781
  (
    n3821,
    n3799
  );


  buf
  g3782
  (
    n3828,
    n3800
  );


  buf
  g3783
  (
    n3826,
    n2103
  );


  buf
  g3784
  (
    n3823,
    n3802
  );


  and
  g3785
  (
    n3820,
    n3804,
    n3800
  );


  and
  g3786
  (
    n3816,
    n3799,
    n3762
  );


  xor
  g3787
  (
    n3825,
    n2098,
    n3801
  );


  nand
  g3788
  (
    n3814,
    n3801,
    n3802
  );


  nand
  g3789
  (
    n3818,
    n3804,
    n3803
  );


  nand
  g3790
  (
    n3824,
    n2101,
    n2100
  );


  nor
  g3791
  (
    n3829,
    n3800,
    n2098
  );


  nand
  g3792
  (
    n3827,
    n3803,
    n2100
  );


  xnor
  g3793
  (
    n3822,
    n3801,
    n3802
  );


  nand
  g3794
  (
    n3830,
    n3799,
    n2102
  );


  nand
  g3795
  (
    n3817,
    n3804,
    n2099
  );


  xnor
  g3796
  (
    n3815,
    n2101,
    n3803
  );


  and
  g3797
  (
    n3831,
    n3804,
    n2102
  );


  nor
  g3798
  (
    n3819,
    n2099,
    n2097
  );


  not
  g3799
  (
    n3841,
    n3831
  );


  buf
  g3800
  (
    n3840,
    n3830
  );


  not
  g3801
  (
    n3851,
    n2838
  );


  not
  g3802
  (
    KeyWire_0_31,
    n3819
  );


  not
  g3803
  (
    n3846,
    n3818
  );


  not
  g3804
  (
    n3842,
    n3823
  );


  not
  g3805
  (
    n3858,
    n3830
  );


  buf
  g3806
  (
    n3874,
    n2838
  );


  buf
  g3807
  (
    n3854,
    n3831
  );


  buf
  g3808
  (
    n3857,
    n3828
  );


  not
  g3809
  (
    n3868,
    n3824
  );


  not
  g3810
  (
    n3875,
    n3829
  );


  buf
  g3811
  (
    n3869,
    n3817
  );


  not
  g3812
  (
    n3876,
    n3820
  );


  not
  g3813
  (
    n3862,
    n3826
  );


  not
  g3814
  (
    n3852,
    n3825
  );


  not
  g3815
  (
    n3845,
    n3829
  );


  not
  g3816
  (
    n3871,
    n3817
  );


  not
  g3817
  (
    n3878,
    n3824
  );


  not
  g3818
  (
    n3835,
    n3776
  );


  buf
  g3819
  (
    n3832,
    n3825
  );


  not
  g3820
  (
    n3850,
    n3814
  );


  not
  g3821
  (
    n3870,
    n3815
  );


  buf
  g3822
  (
    n3859,
    n3822
  );


  buf
  g3823
  (
    n3863,
    n3826
  );


  buf
  g3824
  (
    n3847,
    n3822
  );


  buf
  g3825
  (
    n3856,
    n3827
  );


  not
  g3826
  (
    n3864,
    n3821
  );


  not
  g3827
  (
    n3837,
    n3828
  );


  buf
  g3828
  (
    n3839,
    n3794
  );


  buf
  g3829
  (
    n3836,
    n3827
  );


  not
  g3830
  (
    n3867,
    n3829
  );


  not
  g3831
  (
    n3877,
    n3819
  );


  buf
  g3832
  (
    n3843,
    n3823
  );


  buf
  g3833
  (
    n3838,
    n3826
  );


  buf
  g3834
  (
    n3873,
    n3827
  );


  not
  g3835
  (
    n3860,
    n3826
  );


  buf
  g3836
  (
    n3855,
    n3828
  );


  not
  g3837
  (
    n3861,
    n3822
  );


  not
  g3838
  (
    n3866,
    n3775
  );


  buf
  g3839
  (
    n3833,
    n3829
  );


  not
  g3840
  (
    n3853,
    n3831
  );


  xnor
  g3841
  (
    n3844,
    n3820,
    n3816,
    n3823,
    n3825
  );


  nand
  g3842
  (
    n3834,
    n3830,
    n3824,
    n3818,
    n3821
  );


  and
  g3843
  (
    n3848,
    n3831,
    n3823,
    n3824,
    n3828
  );


  xor
  g3844
  (
    n3849,
    n2838,
    n3815,
    n2103,
    n3827
  );


  nand
  g3845
  (
    KeyWire_0_2,
    n3822,
    n3830,
    n3816,
    n3825
  );


  xnor
  g3846
  (
    n3922,
    n3851,
    n3835,
    n3507,
    n3540
  );


  xnor
  g3847
  (
    n3890,
    n3548,
    n3841,
    n3534,
    n3539
  );


  xor
  g3848
  (
    n3886,
    n3547,
    n3506,
    n3533,
    n3513
  );


  or
  g3849
  (
    n3894,
    n3550,
    n3515,
    n3837,
    n3542
  );


  nor
  g3850
  (
    n3918,
    n3525,
    n3870,
    n2104,
    n3542
  );


  or
  g3851
  (
    n3888,
    n3836,
    n3527,
    n3505,
    n3541
  );


  nor
  g3852
  (
    n3900,
    n3536,
    n3876,
    n3856,
    n3535
  );


  xor
  g3853
  (
    n3889,
    n3529,
    n3543,
    n3538,
    n3874
  );


  or
  g3854
  (
    n3911,
    n3548,
    n3540,
    n3397,
    n3398
  );


  nor
  g3855
  (
    n3905,
    n3518,
    n3842,
    n3550,
    n3538
  );


  nor
  g3856
  (
    n3917,
    n3549,
    n3852,
    n3504,
    n3544
  );


  xor
  g3857
  (
    n3899,
    n3539,
    n3551,
    n3523,
    n3516
  );


  and
  g3858
  (
    n3893,
    n3843,
    n3858,
    n3867,
    n3549
  );


  xor
  g3859
  (
    n3892,
    n2104,
    n3537,
    n3551,
    n3538
  );


  nand
  g3860
  (
    n3903,
    n3869,
    n3546,
    n3541,
    n3547
  );


  xor
  g3861
  (
    n3923,
    n3530,
    n3526,
    n3514,
    n3517
  );


  nor
  g3862
  (
    n3914,
    n3548,
    n3832,
    n3530,
    n3552
  );


  nand
  g3863
  (
    n3884,
    n3549,
    n3850,
    n3552,
    n3547
  );


  or
  g3864
  (
    n3916,
    n3534,
    n3551,
    n3543,
    n3549
  );


  nor
  g3865
  (
    n3904,
    n3848,
    n3547,
    n3860,
    n3845
  );


  nand
  g3866
  (
    n3879,
    n3849,
    n3545,
    n3878,
    n3537
  );


  and
  g3867
  (
    n3901,
    n3846,
    n3520,
    n3518,
    n3543
  );


  or
  g3868
  (
    n3920,
    n3782,
    n3527,
    n3528,
    n3855
  );


  nand
  g3869
  (
    n3919,
    n3522,
    n3526,
    n3545,
    n3541
  );


  xnor
  g3870
  (
    n3883,
    n3550,
    n3847,
    n3539,
    n3551
  );


  nor
  g3871
  (
    n3882,
    n3840,
    n3521,
    n3546,
    n3519
  );


  nand
  g3872
  (
    n3913,
    n3873,
    n3394,
    n3393,
    n3521
  );


  xor
  g3873
  (
    n3915,
    n3397,
    n3865,
    n3511,
    n3857
  );


  and
  g3874
  (
    n3924,
    n3540,
    n3523,
    n3395
  );


  xor
  g3875
  (
    n3880,
    n3838,
    n3508,
    n3541,
    n3394
  );


  or
  g3876
  (
    n3912,
    n3531,
    n3550,
    n3866,
    n3509
  );


  xnor
  g3877
  (
    n3881,
    n3546,
    n3545,
    n3839,
    n3853
  );


  xor
  g3878
  (
    n3902,
    n3871,
    n3544,
    n3878,
    n3517
  );


  nand
  g3879
  (
    n3909,
    n3533,
    n3400,
    n3396,
    n3877
  );


  xor
  g3880
  (
    n3895,
    n3512,
    n3520,
    n3519,
    n3535
  );


  xnor
  g3881
  (
    n3897,
    n3834,
    n3398,
    n3515,
    n3542
  );


  xnor
  g3882
  (
    n3898,
    n3514,
    n3393,
    n3531,
    n3516
  );


  and
  g3883
  (
    n3921,
    n3844,
    n3522,
    n3833,
    n3861
  );


  and
  g3884
  (
    n3885,
    n3544,
    n3532,
    n3546,
    n3524
  );


  and
  g3885
  (
    n3896,
    n3864,
    n3862,
    n3863,
    n3525
  );


  nand
  g3886
  (
    n3910,
    n3399,
    n3552,
    n3539,
    n3859
  );


  and
  g3887
  (
    n3887,
    n3399,
    n3528,
    n3503,
    n3872
  );


  xor
  g3888
  (
    n3906,
    n3543,
    n3538,
    n3396,
    n3544
  );


  nand
  g3889
  (
    n3908,
    n3524,
    n3868,
    n3548,
    n3540
  );


  or
  g3890
  (
    n3891,
    n3510,
    n3875,
    n3545,
    n3532
  );


  nor
  g3891
  (
    n3907,
    n3854,
    n3542,
    n3529,
    n3536
  );


  xnor
  g3892
  (
    n3932,
    n2160,
    n2107,
    n3808,
    n3894
  );


  and
  g3893
  (
    n3959,
    n2137,
    n2140,
    n3883,
    n3906
  );


  xor
  g3894
  (
    n3969,
    n2105,
    n2130,
    n2145,
    n3903
  );


  nor
  g3895
  (
    n3930,
    n2147,
    n3884,
    n3905,
    n2131
  );


  or
  g3896
  (
    n3956,
    n2109,
    n2149,
    n2148,
    n3912
  );


  or
  g3897
  (
    n3950,
    n3809,
    n3924,
    n2151,
    n2156
  );


  nand
  g3898
  (
    n3970,
    n3810,
    n3806,
    n3909,
    n2159
  );


  xor
  g3899
  (
    n3940,
    n3805,
    n2140,
    n2106
  );


  or
  g3900
  (
    n3943,
    n2115,
    n3809,
    n3916,
    n3908
  );


  xor
  g3901
  (
    n3962,
    n2138,
    n2127,
    n2134,
    n2150
  );


  nand
  g3902
  (
    n3971,
    n3902,
    n2113,
    n2122,
    n3806
  );


  or
  g3903
  (
    n3925,
    n3896,
    n2152,
    n2112,
    n3808
  );


  nor
  g3904
  (
    n3935,
    n2111,
    n2111,
    n2123,
    n3805
  );


  nor
  g3905
  (
    n3951,
    n2156,
    n2132,
    n2116,
    n3913
  );


  nor
  g3906
  (
    n3961,
    n3890,
    n3892,
    n3907,
    n2151
  );


  nor
  g3907
  (
    n3963,
    n2148,
    n3810,
    n3880,
    n3807
  );


  and
  g3908
  (
    KeyWire_0_54,
    n2158,
    n3811,
    n2132,
    n2149
  );


  and
  g3909
  (
    n3946,
    n3895,
    n3921,
    n2128,
    n2124
  );


  and
  g3910
  (
    n3937,
    n3810,
    n2141,
    n3806,
    n2108
  );


  nand
  g3911
  (
    n3945,
    n2109,
    n2128,
    n2144,
    n3899
  );


  xor
  g3912
  (
    n3954,
    n3901,
    n2121,
    n2114,
    n2155
  );


  and
  g3913
  (
    n3948,
    n2137,
    n3924,
    n2117
  );


  xor
  g3914
  (
    n3939,
    n2157,
    n2144,
    n3922,
    n2122
  );


  xnor
  g3915
  (
    n3933,
    n2158,
    n2142,
    n3893,
    n3911
  );


  nor
  g3916
  (
    n3944,
    n2126,
    n3809,
    n3888,
    n3808
  );


  xor
  g3917
  (
    KeyWire_0_16,
    n2157,
    n2154,
    n2110,
    n2139
  );


  and
  g3918
  (
    n3942,
    n2133,
    n2130,
    n3805,
    n2153
  );


  nor
  g3919
  (
    n3938,
    n2119,
    n2136,
    n3889,
    n2114
  );


  nor
  g3920
  (
    n3928,
    n2135,
    n2121,
    n3891,
    n2120
  );


  and
  g3921
  (
    n3934,
    n2150,
    n2124,
    n3881,
    n2127
  );


  xnor
  g3922
  (
    n3927,
    n2107,
    n3810,
    n2123,
    n3898
  );


  nor
  g3923
  (
    n3936,
    n2146,
    n3886,
    n2112,
    n2105
  );


  xor
  g3924
  (
    n3960,
    n3914,
    n3897,
    n3915,
    n2129
  );


  nand
  g3925
  (
    n3958,
    n2113,
    n3885,
    n2160,
    n3811
  );


  nor
  g3926
  (
    n3929,
    n3811,
    n3879,
    n2134,
    n2133
  );


  xnor
  g3927
  (
    n3955,
    n3900,
    n2153,
    n2139,
    n2152
  );


  xnor
  g3928
  (
    n3957,
    n2135,
    n3910,
    n2115,
    n2155
  );


  xnor
  g3929
  (
    n3952,
    n2143,
    n2154,
    n2141,
    n2147
  );


  xnor
  g3930
  (
    n3965,
    n3923,
    n2161,
    n2146,
    n3806
  );


  nand
  g3931
  (
    n3931,
    n3918,
    n2143,
    n2145,
    n2120
  );


  or
  g3932
  (
    n3968,
    n2110,
    n3887,
    n2118,
    n2142
  );


  nand
  g3933
  (
    n3947,
    n2126,
    n3807,
    n2159,
    n3904
  );


  or
  g3934
  (
    n3941,
    n2118,
    n3808,
    n3807,
    n3917
  );


  or
  g3935
  (
    n3966,
    n3805,
    n2136,
    n2119,
    n3920
  );


  nand
  g3936
  (
    n3953,
    n2125,
    n2125,
    n3807,
    n2129
  );


  xnor
  g3937
  (
    n3926,
    n2116,
    n3811,
    n3882,
    n2108
  );


  nand
  g3938
  (
    n3949,
    n2138,
    n2131,
    n3919,
    n3809
  );


  buf
  g3939
  (
    n3979,
    n3931
  );


  not
  g3940
  (
    n3976,
    n3933
  );


  not
  g3941
  (
    n3982,
    n3930
  );


  buf
  g3942
  (
    n3974,
    n3932
  );


  not
  g3943
  (
    n3983,
    n3937
  );


  not
  g3944
  (
    n3977,
    n3936
  );


  buf
  g3945
  (
    n3981,
    n3925
  );


  buf
  g3946
  (
    n3984,
    n3934
  );


  buf
  g3947
  (
    n3978,
    n3927
  );


  buf
  g3948
  (
    n3975,
    n3926
  );


  not
  g3949
  (
    n3972,
    n3929
  );


  not
  g3950
  (
    n3980,
    n3928
  );


  not
  g3951
  (
    n3973,
    n3935
  );


  xor
  g3952
  (
    n3986,
    n3972,
    n3977,
    n3813,
    n3982
  );


  xor
  g3953
  (
    n3987,
    n3981,
    n3976,
    n3405,
    n3400
  );


  and
  g3954
  (
    n3990,
    n2738,
    n3976,
    n3975,
    n3980
  );


  or
  g3955
  (
    n3988,
    n3976,
    n3979,
    n3401,
    n3403
  );


  xor
  g3956
  (
    n3995,
    n2739,
    n3401,
    n3980,
    n3977
  );


  xnor
  g3957
  (
    n3994,
    n2740,
    n3978,
    n3812
  );


  and
  g3958
  (
    n4000,
    n3972,
    n3404,
    n3813,
    n3979
  );


  and
  g3959
  (
    n3989,
    n3976,
    n3981,
    n3980
  );


  xor
  g3960
  (
    n3985,
    n3974,
    n2737,
    n3402,
    n3975
  );


  nand
  g3961
  (
    n3999,
    n2742,
    n3978,
    n2739,
    n2736
  );


  nor
  g3962
  (
    n3998,
    n3978,
    n3973,
    n3975,
    n2741
  );


  nor
  g3963
  (
    n3992,
    n3975,
    n3402,
    n2737,
    n3982
  );


  xnor
  g3964
  (
    n3996,
    n3979,
    n3812
  );


  or
  g3965
  (
    n3991,
    n3980,
    n3978,
    n2738,
    n3405
  );


  or
  g3966
  (
    n3993,
    n2736,
    n3403,
    n2741,
    n3404
  );


  nand
  g3967
  (
    n3997,
    n3977,
    n2741,
    n3981,
    n3813
  );


  or
  g3968
  (
    n4002,
    n3974,
    n3982,
    n2740,
    n3977
  );


  xnor
  g3969
  (
    n4001,
    n3813,
    n2740,
    n3737,
    n3973
  );


  xnor
  g3970
  (
    n4005,
    n4001,
    n2162,
    n3406
  );


  or
  g3971
  (
    n4003,
    n2163,
    n2163,
    n2161,
    n3407
  );


  or
  g3972
  (
    n4004,
    n3407,
    n4000,
    n3406,
    n4002
  );


  or
  g3973
  (
    n4009,
    n3941,
    n3951,
    n3946,
    n4004
  );


  nor
  g3974
  (
    n4012,
    n3958,
    n3968,
    n3942,
    n3944
  );


  nand
  g3975
  (
    n4008,
    n3965,
    n4003,
    n3953
  );


  nor
  g3976
  (
    n4017,
    n4005,
    n3948,
    n4004,
    n3962
  );


  xor
  g3977
  (
    n4016,
    n3939,
    n4005,
    n4004
  );


  or
  g3978
  (
    n4006,
    n3964,
    n4004,
    n3954,
    n3966
  );


  xnor
  g3979
  (
    n4015,
    n3959,
    n3947,
    n3961,
    n3963
  );


  nand
  g3980
  (
    n4007,
    n4003,
    n4003,
    n4005,
    n3969
  );


  or
  g3981
  (
    n4014,
    n3969,
    n2164,
    n3970,
    n3952
  );


  xor
  g3982
  (
    n4011,
    n3950,
    n3940,
    n3967,
    n3945
  );


  xnor
  g3983
  (
    n4013,
    n3957,
    n3949,
    n3955,
    n3943
  );


  xor
  g3984
  (
    n4010,
    n3956,
    n3968,
    n3960,
    n3938
  );


  xor
  g3985
  (
    n4024,
    n4011,
    n4015,
    n3984,
    n4017
  );


  xnor
  g3986
  (
    n4019,
    n4009,
    n4017,
    n4008
  );


  nor
  g3987
  (
    n4022,
    n4016,
    n4010,
    n4006,
    n3982
  );


  xnor
  g3988
  (
    n4023,
    n3983,
    n3984,
    n2743,
    n4007
  );


  nand
  g3989
  (
    n4018,
    n3983,
    n4014,
    n3409,
    n2742
  );


  nand
  g3990
  (
    n4025,
    n3984,
    n3408
  );


  nor
  g3991
  (
    n4020,
    n4012,
    n3409,
    n2743,
    n3983
  );


  or
  g3992
  (
    n4021,
    n4013,
    n3983,
    n2743,
    n2742
  );


  xnor
  g3993
  (
    n4026,
    n4025,
    n3970,
    n3971
  );


  xor
  g3994
  (
    n4029,
    n3552,
    n4026,
    n3766,
    n671
  );


  nor
  g3995
  (
    n4028,
    n671,
    n4026,
    n3765,
    n2164
  );


  xnor
  g3996
  (
    n4027,
    n4026,
    n2165,
    n3764,
    n3763
  );


  and
  g3997
  (
    n4030,
    n2165,
    n2167,
    n2166
  );


  nand
  g3998
  (
    n4031,
    n4027,
    n4029,
    n4028,
    n2166
  );


  nand
  g3999
  (
    n4032,
    n3737,
    n160,
    n4031,
    n4030
  );


  xnor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n1462,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n2285,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n3865,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n2739,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n655,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n2979,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n2574,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n1372,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n35,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n2795,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n2047,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n133,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n2569,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n595,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n421,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n3812,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n3964,
    KeyNOTWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1658,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n634,
    KeyNOTWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n469,
    keyIn_0_19,
    KeyWire_0_19
  );


  xor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n1348,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n452,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n461,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n2657,
    KeyNOTWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n2297,
    KeyNOTWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n3756,
    KeyNOTWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n2072,
    keyIn_0_26,
    KeyWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n3191,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n1343,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n888,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n789,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n3872,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n1425,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n1244,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n1710,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    KeyNOTWire_0_35,
    keyIn_0_35,
    KeyWire_0_35
  );


  not
  KeyNOTGate_0_35
  (
    n2710,
    KeyNOTWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n3368,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n3024,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n1608,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n1519,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n1997,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n964,
    keyIn_0_41,
    KeyWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    n3200,
    keyIn_0_42,
    KeyWire_0_42
  );


  xor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n1887,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n1752,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n3750,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n2061,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n1167,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n2429,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n3029,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n1580,
    KeyNOTWire_0_50
  );


  xor
  KeyGate_0_51
  (
    n3524,
    keyIn_0_51,
    KeyWire_0_51
  );


  xor
  KeyGate_0_52
  (
    n1802,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n3652,
    KeyNOTWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n3967,
    keyIn_0_54,
    KeyWire_0_54
  );


  xor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n3465,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n76,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n3559,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n726,
    keyIn_0_58,
    KeyWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n924,
    KeyNOTWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n3132,
    keyIn_0_60,
    KeyWire_0_60
  );


  xnor
  KeyGate_0_61
  (
    n1397,
    keyIn_0_61,
    KeyWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n1783,
    KeyNOTWire_0_62
  );


  xor
  KeyGate_0_63
  (
    KeyNOTWire_0_63,
    keyIn_0_63,
    KeyWire_0_63
  );


  not
  KeyNOTGate_0_63
  (
    n1373,
    KeyNOTWire_0_63
  );


endmodule

