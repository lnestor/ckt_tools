

module Stat_804_2825
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n398,
  n413,
  n409,
  n419,
  n415,
  n417,
  n421,
  n410,
  n420,
  n422,
  n412,
  n418,
  n414,
  n832,
  n829,
  n828,
  n827,
  n834,
  n836,
  n835,
  n831,
  n830,
  n833,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n398;
  output n413;
  output n409;
  output n419;
  output n415;
  output n417;
  output n421;
  output n410;
  output n420;
  output n422;
  output n412;
  output n418;
  output n414;
  output n832;
  output n829;
  output n828;
  output n827;
  output n834;
  output n836;
  output n835;
  output n831;
  output n830;
  output n833;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n411;
  wire n416;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n129,
    n14
  );


  not
  g1
  (
    n87,
    n9
  );


  buf
  g2
  (
    n100,
    n1
  );


  not
  g3
  (
    n50,
    n11
  );


  buf
  g4
  (
    n36,
    n4
  );


  not
  g5
  (
    n82,
    n5
  );


  buf
  g6
  (
    n139,
    n15
  );


  buf
  g7
  (
    n120,
    n15
  );


  not
  g8
  (
    n138,
    n9
  );


  not
  g9
  (
    n89,
    n26
  );


  buf
  g10
  (
    n47,
    n25
  );


  not
  g11
  (
    n140,
    n19
  );


  buf
  g12
  (
    n155,
    n13
  );


  buf
  g13
  (
    n40,
    n23
  );


  buf
  g14
  (
    n119,
    n11
  );


  not
  g15
  (
    n33,
    n2
  );


  not
  g16
  (
    n148,
    n32
  );


  not
  g17
  (
    n66,
    n24
  );


  not
  g18
  (
    n114,
    n2
  );


  buf
  g19
  (
    n68,
    n4
  );


  buf
  g20
  (
    n77,
    n19
  );


  buf
  g21
  (
    n81,
    n17
  );


  not
  g22
  (
    n54,
    n12
  );


  not
  g23
  (
    n154,
    n6
  );


  buf
  g24
  (
    n37,
    n16
  );


  buf
  g25
  (
    n64,
    n17
  );


  not
  g26
  (
    n57,
    n5
  );


  not
  g27
  (
    n159,
    n29
  );


  buf
  g28
  (
    n75,
    n26
  );


  not
  g29
  (
    n109,
    n22
  );


  not
  g30
  (
    n101,
    n25
  );


  not
  g31
  (
    n98,
    n28
  );


  buf
  g32
  (
    n111,
    n8
  );


  buf
  g33
  (
    n147,
    n19
  );


  buf
  g34
  (
    n115,
    n18
  );


  not
  g35
  (
    n110,
    n3
  );


  buf
  g36
  (
    KeyWire_0_6,
    n16
  );


  buf
  g37
  (
    n42,
    n20
  );


  buf
  g38
  (
    n92,
    n23
  );


  buf
  g39
  (
    n151,
    n7
  );


  buf
  g40
  (
    n104,
    n7
  );


  not
  g41
  (
    n45,
    n4
  );


  not
  g42
  (
    KeyWire_0_0,
    n5
  );


  buf
  g43
  (
    n38,
    n8
  );


  not
  g44
  (
    n62,
    n20
  );


  not
  g45
  (
    n131,
    n18
  );


  not
  g46
  (
    n46,
    n31
  );


  not
  g47
  (
    n53,
    n6
  );


  not
  g48
  (
    n145,
    n2
  );


  buf
  g49
  (
    n39,
    n17
  );


  not
  g50
  (
    n127,
    n11
  );


  not
  g51
  (
    n152,
    n32
  );


  buf
  g52
  (
    n43,
    n26
  );


  buf
  g53
  (
    n126,
    n19
  );


  buf
  g54
  (
    n103,
    n27
  );


  buf
  g55
  (
    n149,
    n28
  );


  not
  g56
  (
    n143,
    n15
  );


  not
  g57
  (
    n107,
    n11
  );


  buf
  g58
  (
    n63,
    n21
  );


  buf
  g59
  (
    n74,
    n27
  );


  not
  g60
  (
    n146,
    n27
  );


  not
  g61
  (
    n123,
    n16
  );


  buf
  g62
  (
    n52,
    n9
  );


  not
  g63
  (
    n142,
    n25
  );


  not
  g64
  (
    n76,
    n10
  );


  buf
  g65
  (
    n49,
    n15
  );


  buf
  g66
  (
    n130,
    n29
  );


  buf
  g67
  (
    n91,
    n29
  );


  buf
  g68
  (
    n84,
    n32
  );


  not
  g69
  (
    n34,
    n31
  );


  buf
  g70
  (
    n113,
    n22
  );


  not
  g71
  (
    n83,
    n14
  );


  not
  g72
  (
    n133,
    n13
  );


  buf
  g73
  (
    n78,
    n6
  );


  not
  g74
  (
    n144,
    n30
  );


  not
  g75
  (
    n60,
    n24
  );


  buf
  g76
  (
    n71,
    n6
  );


  buf
  g77
  (
    n150,
    n31
  );


  buf
  g78
  (
    n69,
    n12
  );


  not
  g79
  (
    n135,
    n29
  );


  buf
  g80
  (
    n128,
    n10
  );


  not
  g81
  (
    n116,
    n30
  );


  buf
  g82
  (
    n108,
    n18
  );


  not
  g83
  (
    n93,
    n25
  );


  buf
  g84
  (
    n160,
    n3
  );


  buf
  g85
  (
    n85,
    n1
  );


  not
  g86
  (
    n118,
    n32
  );


  not
  g87
  (
    n136,
    n17
  );


  buf
  g88
  (
    n102,
    n14
  );


  not
  g89
  (
    n157,
    n21
  );


  buf
  g90
  (
    n134,
    n27
  );


  not
  g91
  (
    n61,
    n8
  );


  buf
  g92
  (
    n79,
    n5
  );


  not
  g93
  (
    n105,
    n10
  );


  not
  g94
  (
    n153,
    n12
  );


  not
  g95
  (
    n65,
    n13
  );


  buf
  g96
  (
    n132,
    n28
  );


  buf
  g97
  (
    n156,
    n13
  );


  buf
  g98
  (
    n141,
    n1
  );


  buf
  g99
  (
    n51,
    n4
  );


  not
  g100
  (
    n106,
    n21
  );


  buf
  g101
  (
    n122,
    n10
  );


  buf
  g102
  (
    n58,
    n8
  );


  not
  g103
  (
    n44,
    n20
  );


  buf
  g104
  (
    n137,
    n20
  );


  not
  g105
  (
    n117,
    n18
  );


  buf
  g106
  (
    n67,
    n1
  );


  not
  g107
  (
    n124,
    n12
  );


  not
  g108
  (
    n86,
    n30
  );


  not
  g109
  (
    n56,
    n31
  );


  not
  g110
  (
    n90,
    n16
  );


  not
  g111
  (
    n80,
    n3
  );


  buf
  g112
  (
    n72,
    n3
  );


  buf
  g113
  (
    n158,
    n7
  );


  buf
  g114
  (
    n73,
    n30
  );


  not
  g115
  (
    n59,
    n14
  );


  not
  g116
  (
    n99,
    n9
  );


  buf
  g117
  (
    n55,
    n22
  );


  buf
  g118
  (
    n88,
    n21
  );


  buf
  g119
  (
    n121,
    n2
  );


  not
  g120
  (
    n41,
    n28
  );


  not
  g121
  (
    n97,
    n22
  );


  not
  g122
  (
    n95,
    n24
  );


  not
  g123
  (
    n112,
    n23
  );


  not
  g124
  (
    n70,
    n24
  );


  not
  g125
  (
    n125,
    n26
  );


  buf
  g126
  (
    n35,
    n7
  );


  not
  g127
  (
    n96,
    n23
  );


  not
  g128
  (
    n259,
    n34
  );


  not
  g129
  (
    n264,
    n81
  );


  not
  g130
  (
    n302,
    n82
  );


  not
  g131
  (
    n177,
    n72
  );


  not
  g132
  (
    n164,
    n110
  );


  buf
  g133
  (
    n229,
    n136
  );


  buf
  g134
  (
    n263,
    n91
  );


  buf
  g135
  (
    n306,
    n129
  );


  not
  g136
  (
    n294,
    n151
  );


  buf
  g137
  (
    n269,
    n102
  );


  not
  g138
  (
    n167,
    n142
  );


  not
  g139
  (
    n312,
    n58
  );


  not
  g140
  (
    n296,
    n67
  );


  buf
  g141
  (
    n198,
    n160
  );


  not
  g142
  (
    n199,
    n73
  );


  buf
  g143
  (
    n318,
    n144
  );


  not
  g144
  (
    n328,
    n47
  );


  buf
  g145
  (
    n174,
    n135
  );


  not
  g146
  (
    n211,
    n49
  );


  not
  g147
  (
    n256,
    n89
  );


  buf
  g148
  (
    n289,
    n126
  );


  not
  g149
  (
    n310,
    n130
  );


  not
  g150
  (
    n253,
    n147
  );


  not
  g151
  (
    n245,
    n41
  );


  not
  g152
  (
    n243,
    n76
  );


  not
  g153
  (
    n257,
    n80
  );


  buf
  g154
  (
    n309,
    n125
  );


  not
  g155
  (
    n239,
    n137
  );


  buf
  g156
  (
    n179,
    n138
  );


  not
  g157
  (
    n237,
    n125
  );


  buf
  g158
  (
    n324,
    n81
  );


  not
  g159
  (
    n226,
    n44
  );


  not
  g160
  (
    n180,
    n107
  );


  not
  g161
  (
    n248,
    n118
  );


  buf
  g162
  (
    n295,
    n128
  );


  not
  g163
  (
    n304,
    n97
  );


  buf
  g164
  (
    n218,
    n68
  );


  buf
  g165
  (
    n250,
    n94
  );


  not
  g166
  (
    n166,
    n117
  );


  not
  g167
  (
    n191,
    n107
  );


  buf
  g168
  (
    n298,
    n133
  );


  buf
  g169
  (
    n238,
    n145
  );


  not
  g170
  (
    n216,
    n100
  );


  not
  g171
  (
    n215,
    n127
  );


  not
  g172
  (
    n262,
    n124
  );


  not
  g173
  (
    n225,
    n88
  );


  not
  g174
  (
    n284,
    n67
  );


  buf
  g175
  (
    n285,
    n49
  );


  buf
  g176
  (
    n279,
    n54
  );


  buf
  g177
  (
    n183,
    n107
  );


  buf
  g178
  (
    n273,
    n117
  );


  not
  g179
  (
    n249,
    n94
  );


  not
  g180
  (
    n173,
    n83
  );


  not
  g181
  (
    n247,
    n143
  );


  not
  g182
  (
    n317,
    n132
  );


  not
  g183
  (
    n277,
    n103
  );


  xnor
  g184
  (
    n197,
    n122,
    n126,
    n103,
    n160
  );


  xnor
  g185
  (
    n202,
    n58,
    n49,
    n97,
    n121
  );


  or
  g186
  (
    n299,
    n107,
    n94,
    n90,
    n65
  );


  and
  g187
  (
    KeyWire_0_10,
    n54,
    n157,
    n117,
    n127
  );


  and
  g188
  (
    n188,
    n36,
    n108,
    n90,
    n45
  );


  and
  g189
  (
    n233,
    n141,
    n139,
    n144,
    n89
  );


  or
  g190
  (
    KeyWire_0_13,
    n156,
    n54,
    n82,
    n44
  );


  xor
  g191
  (
    n176,
    n154,
    n134,
    n146,
    n132
  );


  nor
  g192
  (
    n236,
    n43,
    n113,
    n35,
    n62
  );


  or
  g193
  (
    n293,
    n92,
    n95,
    n88,
    n44
  );


  or
  g194
  (
    n187,
    n159,
    n55,
    n96,
    n70
  );


  nand
  g195
  (
    n290,
    n141,
    n73,
    n71,
    n66
  );


  nor
  g196
  (
    n330,
    n149,
    n155,
    n93,
    n134
  );


  or
  g197
  (
    n244,
    n74,
    n35,
    n153,
    n42
  );


  nor
  g198
  (
    n246,
    n124,
    n57,
    n105,
    n104
  );


  and
  g199
  (
    n320,
    n131,
    n123,
    n88,
    n111
  );


  xnor
  g200
  (
    n292,
    n100,
    n111,
    n80,
    n85
  );


  nor
  g201
  (
    n186,
    n119,
    n145,
    n77,
    n144
  );


  nand
  g202
  (
    n181,
    n116,
    n39,
    n60,
    n87
  );


  or
  g203
  (
    n276,
    n137,
    n98,
    n116,
    n87
  );


  or
  g204
  (
    n316,
    n119,
    n136,
    n135,
    n130
  );


  xor
  g205
  (
    n267,
    n144,
    n146,
    n101,
    n158
  );


  xnor
  g206
  (
    n240,
    n69,
    n81,
    n153,
    n87
  );


  or
  g207
  (
    n195,
    n155,
    n91,
    n140,
    n120
  );


  nor
  g208
  (
    n228,
    n157,
    n104,
    n74,
    n82
  );


  nand
  g209
  (
    n169,
    n154,
    n160,
    n112,
    n35
  );


  or
  g210
  (
    n297,
    n124,
    n74,
    n158,
    n121
  );


  or
  g211
  (
    n221,
    n108,
    n115,
    n46,
    n33
  );


  nand
  g212
  (
    n190,
    n142,
    n103,
    n56,
    n92
  );


  xor
  g213
  (
    n252,
    n76,
    n148,
    n121,
    n33
  );


  xor
  g214
  (
    n274,
    n45,
    n108,
    n104,
    n64
  );


  xnor
  g215
  (
    n268,
    n57,
    n87,
    n62,
    n151
  );


  xor
  g216
  (
    n205,
    n75,
    n34,
    n61,
    n49
  );


  and
  g217
  (
    n283,
    n56,
    n149,
    n60,
    n70
  );


  nand
  g218
  (
    n213,
    n89,
    n151,
    n40,
    n111
  );


  xor
  g219
  (
    n311,
    n105,
    n109,
    n59,
    n53
  );


  xor
  g220
  (
    n203,
    n142,
    n39,
    n84,
    n56
  );


  nor
  g221
  (
    n321,
    n61,
    n100,
    n148,
    n159
  );


  and
  g222
  (
    n162,
    n86,
    n71,
    n122,
    n160
  );


  nand
  g223
  (
    n163,
    n128,
    n73,
    n101,
    n110
  );


  nor
  g224
  (
    n255,
    n106,
    n79,
    n110
  );


  or
  g225
  (
    n326,
    n105,
    n63,
    n108,
    n151
  );


  xnor
  g226
  (
    n242,
    n65,
    n51,
    n63,
    n66
  );


  nand
  g227
  (
    n288,
    n44,
    n125,
    n153,
    n114
  );


  xor
  g228
  (
    n275,
    n99,
    n42,
    n37,
    n33
  );


  nor
  g229
  (
    n185,
    n46,
    n92,
    n40,
    n127
  );


  xnor
  g230
  (
    n270,
    n66,
    n152,
    n136,
    n55
  );


  and
  g231
  (
    n300,
    n115,
    n36,
    n145,
    n96
  );


  xor
  g232
  (
    n278,
    n146,
    n47,
    n147,
    n102
  );


  and
  g233
  (
    n214,
    n124,
    n98,
    n155,
    n64
  );


  nand
  g234
  (
    n307,
    n42,
    n56,
    n154,
    n140
  );


  xor
  g235
  (
    n266,
    n88,
    n72,
    n58,
    n80
  );


  nand
  g236
  (
    n325,
    n47,
    n46,
    n130,
    n155
  );


  or
  g237
  (
    n281,
    n76,
    n55,
    n138,
    n96
  );


  xor
  g238
  (
    n303,
    n77,
    n94,
    n149,
    n65
  );


  nand
  g239
  (
    n308,
    n156,
    n156,
    n93,
    n100
  );


  or
  g240
  (
    n189,
    n106,
    n156,
    n38,
    n53
  );


  and
  g241
  (
    n261,
    n45,
    n93,
    n97,
    n42
  );


  or
  g242
  (
    n265,
    n121,
    n115,
    n84,
    n118
  );


  xor
  g243
  (
    n313,
    n39,
    n157,
    n129,
    n112
  );


  xnor
  g244
  (
    n329,
    n51,
    n132,
    n103,
    n101
  );


  xor
  g245
  (
    n171,
    n71,
    n123,
    n41,
    n113
  );


  and
  g246
  (
    n206,
    n95,
    n118,
    n54,
    n68
  );


  or
  g247
  (
    n232,
    n99,
    n59,
    n63,
    n35
  );


  or
  g248
  (
    n193,
    n130,
    n114,
    n37,
    n83
  );


  xnor
  g249
  (
    n231,
    n128,
    n152,
    n133,
    n60
  );


  nand
  g250
  (
    n217,
    n142,
    n146,
    n75,
    n59
  );


  nor
  g251
  (
    n208,
    n143,
    n43,
    n150
  );


  xnor
  g252
  (
    n305,
    n57,
    n48,
    n79,
    n92
  );


  nor
  g253
  (
    n301,
    n95,
    n143,
    n120,
    n152
  );


  xor
  g254
  (
    n260,
    n101,
    n159,
    n74,
    n41
  );


  xnor
  g255
  (
    n258,
    n47,
    n67,
    n134,
    n120
  );


  or
  g256
  (
    n220,
    n122,
    n86,
    n78,
    n82
  );


  xor
  g257
  (
    n314,
    n91,
    n110,
    n38,
    n137
  );


  or
  g258
  (
    n223,
    n48,
    n158,
    n93,
    n90
  );


  nor
  g259
  (
    n182,
    n137,
    n99,
    n65,
    n150
  );


  xnor
  g260
  (
    n323,
    n158,
    n119,
    n38,
    n150
  );


  or
  g261
  (
    n230,
    n43,
    n37,
    n58
  );


  xor
  g262
  (
    n172,
    n38,
    n39,
    n154,
    n78
  );


  or
  g263
  (
    n224,
    n105,
    n85,
    n73,
    n118
  );


  or
  g264
  (
    n192,
    n70,
    n126,
    n50,
    n78
  );


  xor
  g265
  (
    n271,
    n117,
    n106,
    n62,
    n75
  );


  xnor
  g266
  (
    n235,
    n36,
    n52,
    n126
  );


  xnor
  g267
  (
    n194,
    n123,
    n63,
    n50,
    n127
  );


  nor
  g268
  (
    n286,
    n72,
    n115,
    n116,
    n45
  );


  xor
  g269
  (
    n175,
    n85,
    n131,
    n125,
    n68
  );


  or
  g270
  (
    n315,
    n148,
    n52,
    n98,
    n84
  );


  nand
  g271
  (
    n319,
    n75,
    n86,
    n157,
    n69
  );


  or
  g272
  (
    n272,
    n139,
    n61,
    n129,
    n132
  );


  xor
  g273
  (
    n251,
    n145,
    n55,
    n78,
    n50
  );


  nand
  g274
  (
    n204,
    n138,
    n61,
    n81,
    n84
  );


  xor
  g275
  (
    n254,
    n128,
    n79,
    n57,
    n33
  );


  nand
  g276
  (
    n212,
    n68,
    n104,
    n135,
    n34
  );


  or
  g277
  (
    n165,
    n109,
    n52,
    n72,
    n114
  );


  nor
  g278
  (
    n170,
    n85,
    n77,
    n53,
    n153
  );


  xor
  g279
  (
    n219,
    n143,
    n112,
    n139,
    n89
  );


  and
  g280
  (
    n322,
    n97,
    n131,
    n40,
    n66
  );


  xor
  g281
  (
    n196,
    n51,
    n95,
    n86,
    n77
  );


  xnor
  g282
  (
    n234,
    n69,
    n116,
    n112,
    n41
  );


  xnor
  g283
  (
    n184,
    n152,
    n64,
    n50,
    n80
  );


  nand
  g284
  (
    n168,
    n98,
    n149,
    n60,
    n109
  );


  xor
  g285
  (
    n207,
    n83,
    n148,
    n139,
    n71
  );


  and
  g286
  (
    n161,
    n51,
    n48,
    n90,
    n46
  );


  and
  g287
  (
    n282,
    n64,
    n147,
    n83,
    n122
  );


  and
  g288
  (
    n210,
    n59,
    n106,
    n133,
    n48
  );


  or
  g289
  (
    n287,
    n134,
    n40,
    n147,
    n133
  );


  xnor
  g290
  (
    n241,
    n34,
    n113,
    n119,
    n114
  );


  and
  g291
  (
    n209,
    n140,
    n102,
    n69,
    n53
  );


  nand
  g292
  (
    n280,
    n131,
    n91,
    n99,
    n62
  );


  xor
  g293
  (
    n178,
    n159,
    n102,
    n123,
    n135
  );


  xor
  g294
  (
    n327,
    n36,
    n96,
    n111,
    n138
  );


  nand
  g295
  (
    n291,
    n150,
    n140,
    n120,
    n129
  );


  xnor
  g296
  (
    n222,
    n67,
    n109,
    n76,
    n141
  );


  xnor
  g297
  (
    KeyWire_0_14,
    n136,
    n113,
    n141,
    n70
  );


  nor
  g298
  (
    n372,
    n219,
    n275,
    n181,
    n175
  );


  xor
  g299
  (
    n381,
    n233,
    n165,
    n245,
    n271
  );


  or
  g300
  (
    n358,
    n258,
    n179,
    n251,
    n173
  );


  or
  g301
  (
    n365,
    n255,
    n256,
    n264,
    n213
  );


  and
  g302
  (
    n333,
    n283,
    n300,
    n296,
    n284
  );


  nor
  g303
  (
    n331,
    n166,
    n288,
    n204,
    n197
  );


  and
  g304
  (
    KeyWire_0_5,
    n187,
    n281,
    n294,
    n238
  );


  nand
  g305
  (
    n374,
    n226,
    n243,
    n201,
    n206
  );


  xor
  g306
  (
    n345,
    n225,
    n266,
    n278,
    n170
  );


  or
  g307
  (
    n377,
    n259,
    n280,
    n253,
    n203
  );


  or
  g308
  (
    n346,
    n164,
    n281,
    n282,
    n210
  );


  xor
  g309
  (
    n362,
    n241,
    n192,
    n178,
    n265
  );


  or
  g310
  (
    n371,
    n286,
    n276,
    n176,
    n272
  );


  nor
  g311
  (
    n332,
    n168,
    n260,
    n237,
    n214
  );


  xor
  g312
  (
    n338,
    n230,
    n291,
    n261,
    n227
  );


  nor
  g313
  (
    n347,
    n234,
    n266,
    n247,
    n225
  );


  or
  g314
  (
    n355,
    n167,
    n242,
    n185,
    n263
  );


  nand
  g315
  (
    n334,
    n247,
    n268,
    n299,
    n258
  );


  nand
  g316
  (
    n343,
    n248,
    n235,
    n264,
    n282
  );


  nor
  g317
  (
    n339,
    n193,
    n298,
    n291,
    n262
  );


  xnor
  g318
  (
    n349,
    n286,
    n243,
    n200,
    n207
  );


  and
  g319
  (
    n336,
    n232,
    n259,
    n244,
    n228
  );


  nand
  g320
  (
    n335,
    n194,
    n161,
    n287,
    n240
  );


  xor
  g321
  (
    n342,
    n249,
    n285,
    n251,
    n274
  );


  nor
  g322
  (
    n373,
    n232,
    n299,
    n231,
    n300
  );


  and
  g323
  (
    n348,
    n287,
    n276,
    n278,
    n221
  );


  or
  g324
  (
    n384,
    n267,
    n217,
    n231,
    n216
  );


  or
  g325
  (
    n356,
    n229,
    n196,
    n257,
    n227
  );


  or
  g326
  (
    n386,
    n297,
    n235,
    n239,
    n244
  );


  nand
  g327
  (
    n352,
    n162,
    n289,
    n228,
    n284
  );


  and
  g328
  (
    n364,
    n279,
    n224,
    n295,
    n180
  );


  nor
  g329
  (
    n379,
    n238,
    n279,
    n220,
    n270
  );


  and
  g330
  (
    n383,
    n252,
    n236,
    n223
  );


  xor
  g331
  (
    n369,
    n202,
    n205,
    n239,
    n269
  );


  xor
  g332
  (
    n353,
    n293,
    n292,
    n199,
    n222
  );


  nor
  g333
  (
    n370,
    n280,
    n191,
    n241,
    n250
  );


  xnor
  g334
  (
    n366,
    n198,
    n186,
    n294,
    n290
  );


  nor
  g335
  (
    n378,
    n174,
    n217,
    n172,
    n269
  );


  xor
  g336
  (
    n376,
    n246,
    n261,
    n283,
    n219
  );


  xor
  g337
  (
    n337,
    n274,
    n289,
    n262,
    n298
  );


  or
  g338
  (
    n380,
    n211,
    n226,
    n250,
    n222
  );


  xnor
  g339
  (
    n385,
    n218,
    n208,
    n265,
    n268
  );


  or
  g340
  (
    n357,
    n183,
    n218,
    n301,
    n236
  );


  xor
  g341
  (
    n359,
    n288,
    n242,
    n229,
    n254
  );


  and
  g342
  (
    n344,
    n255,
    n190,
    n263,
    n245
  );


  and
  g343
  (
    n382,
    n270,
    n293,
    n214,
    n240
  );


  xnor
  g344
  (
    n361,
    n277,
    n252,
    n234,
    n253
  );


  xnor
  g345
  (
    n354,
    n169,
    n285,
    n248,
    n184
  );


  xnor
  g346
  (
    n363,
    n177,
    n233,
    n220,
    n275
  );


  or
  g347
  (
    n341,
    n221,
    n254,
    n212,
    n224
  );


  nor
  g348
  (
    n387,
    n171,
    n272,
    n297,
    n209
  );


  and
  g349
  (
    n350,
    n257,
    n249,
    n273,
    n182
  );


  nor
  g350
  (
    n375,
    n195,
    n267,
    n215,
    n230
  );


  or
  g351
  (
    n351,
    n215,
    n273,
    n188,
    n237
  );


  xnor
  g352
  (
    n367,
    n216,
    n292,
    n296,
    n163
  );


  xnor
  g353
  (
    n340,
    n271,
    n246,
    n295,
    n256
  );


  nand
  g354
  (
    n360,
    n189,
    n277,
    n290,
    n260
  );


  buf
  g355
  (
    n400,
    n331
  );


  buf
  g356
  (
    n404,
    n345
  );


  not
  g357
  (
    n395,
    n336
  );


  not
  g358
  (
    n396,
    n333
  );


  buf
  g359
  (
    n394,
    n334
  );


  not
  g360
  (
    n397,
    n348
  );


  buf
  g361
  (
    n392,
    n337
  );


  not
  g362
  (
    n405,
    n340
  );


  buf
  g363
  (
    n402,
    n341
  );


  not
  g364
  (
    n399,
    n343
  );


  not
  g365
  (
    n390,
    n344
  );


  buf
  g366
  (
    n389,
    n346
  );


  not
  g367
  (
    n401,
    n347
  );


  not
  g368
  (
    n393,
    n332
  );


  buf
  g369
  (
    n388,
    n339
  );


  not
  g370
  (
    n403,
    n338
  );


  not
  g371
  (
    n398,
    n342
  );


  not
  g372
  (
    n391,
    n335
  );


  buf
  g373
  (
    n407,
    n398
  );


  buf
  g374
  (
    n406,
    n397
  );


  buf
  g375
  (
    n415,
    n403
  );


  not
  g376
  (
    n420,
    n400
  );


  buf
  g377
  (
    n412,
    n394
  );


  buf
  g378
  (
    n418,
    n402
  );


  buf
  g379
  (
    n408,
    n396
  );


  buf
  g380
  (
    n416,
    n404
  );


  buf
  g381
  (
    n422,
    n401
  );


  buf
  g382
  (
    n417,
    n393
  );


  not
  g383
  (
    n414,
    n399
  );


  not
  g384
  (
    n419,
    n392
  );


  not
  g385
  (
    n421,
    n391
  );


  not
  g386
  (
    n410,
    n390
  );


  not
  g387
  (
    n413,
    n395
  );


  buf
  g388
  (
    n409,
    n389
  );


  buf
  g389
  (
    n411,
    n405
  );


  buf
  g390
  (
    n424,
    n411
  );


  buf
  g391
  (
    n426,
    n422
  );


  buf
  g392
  (
    n433,
    n414
  );


  not
  g393
  (
    n423,
    n412
  );


  not
  g394
  (
    n437,
    n416
  );


  not
  g395
  (
    n432,
    n422
  );


  not
  g396
  (
    n438,
    n419
  );


  not
  g397
  (
    n425,
    n421
  );


  not
  g398
  (
    n436,
    n421
  );


  buf
  g399
  (
    n428,
    n417
  );


  buf
  g400
  (
    n430,
    n418
  );


  not
  g401
  (
    n434,
    n410
  );


  buf
  g402
  (
    n431,
    n420
  );


  not
  g403
  (
    n429,
    n420
  );


  not
  g404
  (
    n427,
    n415
  );


  not
  g405
  (
    n435,
    n413
  );


  not
  g406
  (
    n443,
    n427
  );


  not
  g407
  (
    n439,
    n429
  );


  not
  g408
  (
    n440,
    n431
  );


  not
  g409
  (
    n444,
    n425
  );


  not
  g410
  (
    n446,
    n432
  );


  nor
  g411
  (
    n445,
    n424,
    n430,
    n432,
    n423
  );


  xnor
  g412
  (
    n442,
    n431,
    n424,
    n429,
    n432
  );


  or
  g413
  (
    n441,
    n423,
    n428,
    n426
  );


  and
  g414
  (
    n447,
    n430,
    n427,
    n425,
    n428
  );


  not
  g415
  (
    n449,
    n442
  );


  not
  g416
  (
    n453,
    n443
  );


  buf
  g417
  (
    n454,
    n441
  );


  not
  g418
  (
    n448,
    n442
  );


  buf
  g419
  (
    n450,
    n443
  );


  not
  g420
  (
    n455,
    n440
  );


  buf
  g421
  (
    n451,
    n441
  );


  not
  g422
  (
    n452,
    n440
  );


  not
  g423
  (
    n465,
    n451
  );


  buf
  g424
  (
    n458,
    n357
  );


  buf
  g425
  (
    n467,
    n450
  );


  buf
  g426
  (
    n468,
    n349
  );


  buf
  g427
  (
    n456,
    n350
  );


  not
  g428
  (
    n460,
    n448
  );


  buf
  g429
  (
    n462,
    n455
  );


  buf
  g430
  (
    n471,
    n449
  );


  buf
  g431
  (
    n463,
    n455
  );


  buf
  g432
  (
    n470,
    n448
  );


  buf
  g433
  (
    n461,
    n453
  );


  not
  g434
  (
    n469,
    n356
  );


  not
  g435
  (
    n464,
    n353
  );


  nand
  g436
  (
    n459,
    n450,
    n452,
    n351,
    n352
  );


  nor
  g437
  (
    n457,
    n451,
    n452,
    n449,
    n454
  );


  xor
  g438
  (
    n466,
    n453,
    n355,
    n354,
    n454
  );


  buf
  g439
  (
    n473,
    n456
  );


  not
  g440
  (
    n472,
    n456
  );


  and
  g441
  (
    n474,
    n473,
    n472
  );


  not
  g442
  (
    n478,
    n474
  );


  not
  g443
  (
    n477,
    n474
  );


  not
  g444
  (
    n475,
    n474
  );


  not
  g445
  (
    n476,
    n474
  );


  buf
  g446
  (
    n480,
    n475
  );


  not
  g447
  (
    n479,
    n475
  );


  not
  g448
  (
    n482,
    n479
  );


  not
  g449
  (
    n483,
    n480
  );


  xor
  g450
  (
    n481,
    n480,
    n444
  );


  xnor
  g451
  (
    n484,
    n479,
    n445,
    n444
  );


  nand
  g452
  (
    n485,
    n456,
    n481
  );


  nor
  g453
  (
    n486,
    n482,
    n481
  );


  buf
  g454
  (
    n487,
    n485
  );


  buf
  g455
  (
    n489,
    n487
  );


  not
  g456
  (
    n488,
    n487
  );


  buf
  g457
  (
    n490,
    n488
  );


  buf
  g458
  (
    n492,
    n490
  );


  buf
  g459
  (
    n491,
    n490
  );


  not
  g460
  (
    n494,
    n482
  );


  not
  g461
  (
    n496,
    n358
  );


  buf
  g462
  (
    n498,
    n483
  );


  not
  g463
  (
    n493,
    n363
  );


  nand
  g464
  (
    n495,
    n483,
    n361,
    n491,
    n360
  );


  xnor
  g465
  (
    n500,
    n432,
    n491,
    n362
  );


  not
  g466
  (
    n497,
    n492
  );


  or
  g467
  (
    n499,
    n359,
    n491,
    n484
  );


  and
  g468
  (
    n507,
    n437,
    n433,
    n497
  );


  xnor
  g469
  (
    n508,
    n500,
    n434,
    n499
  );


  and
  g470
  (
    n516,
    n496,
    n494,
    n436,
    n446
  );


  xor
  g471
  (
    n515,
    n500,
    n434,
    n495,
    n496
  );


  xnor
  g472
  (
    n501,
    n447,
    n493,
    n435
  );


  nor
  g473
  (
    n503,
    n494,
    n498,
    n434,
    n500
  );


  xor
  g474
  (
    n514,
    n493,
    n498,
    n433,
    n434
  );


  xnor
  g475
  (
    n505,
    n498,
    n500,
    n438,
    n497
  );


  or
  g476
  (
    n506,
    n498,
    n494,
    n433,
    n496
  );


  xnor
  g477
  (
    n502,
    n497,
    n495
  );


  nand
  g478
  (
    n511,
    n493,
    n436,
    n437,
    n446
  );


  xor
  g479
  (
    n510,
    n499,
    n438,
    n433,
    n437
  );


  and
  g480
  (
    n509,
    n497,
    n493,
    n499,
    n494
  );


  or
  g481
  (
    n512,
    n486,
    n436,
    n447
  );


  xnor
  g482
  (
    n513,
    n301,
    n438,
    n435,
    n437
  );


  and
  g483
  (
    n504,
    n499,
    n435,
    n496,
    n438
  );


  not
  g484
  (
    n517,
    n503
  );


  not
  g485
  (
    n518,
    n503
  );


  not
  g486
  (
    n525,
    n517
  );


  buf
  g487
  (
    n523,
    n517
  );


  not
  g488
  (
    n520,
    n518
  );


  not
  g489
  (
    n524,
    n517
  );


  not
  g490
  (
    n522,
    n518
  );


  buf
  g491
  (
    n521,
    n518
  );


  not
  g492
  (
    n526,
    n517
  );


  not
  g493
  (
    n519,
    n518
  );


  not
  g494
  (
    n541,
    n506
  );


  buf
  g495
  (
    n545,
    n506
  );


  not
  g496
  (
    n528,
    n526
  );


  not
  g497
  (
    n540,
    n507
  );


  buf
  g498
  (
    n544,
    n524
  );


  buf
  g499
  (
    n543,
    n513
  );


  buf
  g500
  (
    n534,
    n508
  );


  not
  g501
  (
    n539,
    n519
  );


  buf
  g502
  (
    n537,
    n523
  );


  buf
  g503
  (
    n532,
    n512
  );


  and
  g504
  (
    n538,
    n505,
    n511
  );


  buf
  g505
  (
    n536,
    n522
  );


  xnor
  g506
  (
    n542,
    n524,
    n512,
    n510,
    n507
  );


  or
  g507
  (
    n535,
    n526,
    n526,
    n525,
    n514
  );


  nor
  g508
  (
    n530,
    n525,
    n519,
    n505,
    n515
  );


  xnor
  g509
  (
    n546,
    n516,
    n504,
    n514,
    n511
  );


  xnor
  g510
  (
    n533,
    n525,
    n525,
    n520,
    n513
  );


  or
  g511
  (
    KeyWire_0_2,
    n526,
    n504,
    n520,
    n523
  );


  nand
  g512
  (
    n531,
    n521,
    n509,
    n516
  );


  or
  g513
  (
    n527,
    n515,
    n521,
    n510,
    n508
  );


  not
  g514
  (
    n614,
    n527
  );


  buf
  g515
  (
    KeyWire_0_12,
    n303
  );


  not
  g516
  (
    n574,
    n546
  );


  not
  g517
  (
    n619,
    n312
  );


  buf
  g518
  (
    n605,
    n304
  );


  buf
  g519
  (
    n616,
    n537
  );


  not
  g520
  (
    n568,
    n329
  );


  buf
  g521
  (
    n577,
    n540
  );


  not
  g522
  (
    n587,
    n545
  );


  buf
  g523
  (
    n626,
    n530
  );


  buf
  g524
  (
    n558,
    n314
  );


  not
  g525
  (
    n552,
    n539
  );


  buf
  g526
  (
    n553,
    n316
  );


  buf
  g527
  (
    n590,
    n305
  );


  buf
  g528
  (
    n576,
    n324
  );


  buf
  g529
  (
    n565,
    n543
  );


  buf
  g530
  (
    n550,
    n538
  );


  not
  g531
  (
    n600,
    n537
  );


  buf
  g532
  (
    n588,
    n327
  );


  buf
  g533
  (
    n602,
    n545
  );


  not
  g534
  (
    n604,
    n539
  );


  not
  g535
  (
    n548,
    n546
  );


  not
  g536
  (
    n585,
    n527
  );


  not
  g537
  (
    n607,
    n540
  );


  not
  g538
  (
    n589,
    n313
  );


  not
  g539
  (
    n555,
    n531
  );


  buf
  g540
  (
    n615,
    n529
  );


  not
  g541
  (
    n613,
    n324
  );


  not
  g542
  (
    n595,
    n302
  );


  buf
  g543
  (
    n579,
    n316
  );


  not
  g544
  (
    n559,
    n545
  );


  not
  g545
  (
    n625,
    n328
  );


  not
  g546
  (
    n556,
    n326
  );


  not
  g547
  (
    n572,
    n308
  );


  not
  g548
  (
    n591,
    n532
  );


  not
  g549
  (
    n561,
    n536
  );


  not
  g550
  (
    n586,
    n528
  );


  not
  g551
  (
    n564,
    n329
  );


  buf
  g552
  (
    n617,
    n541
  );


  not
  g553
  (
    n563,
    n533
  );


  buf
  g554
  (
    n599,
    n304
  );


  not
  g555
  (
    n584,
    n529
  );


  not
  g556
  (
    n623,
    n540
  );


  buf
  g557
  (
    n583,
    n541
  );


  buf
  g558
  (
    n573,
    n325
  );


  buf
  g559
  (
    n609,
    n323
  );


  not
  g560
  (
    n569,
    n534
  );


  not
  g561
  (
    KeyWire_0_3,
    n322
  );


  not
  g562
  (
    n557,
    n327
  );


  not
  g563
  (
    n549,
    n307
  );


  not
  g564
  (
    n608,
    n527
  );


  buf
  g565
  (
    n594,
    n310
  );


  buf
  g566
  (
    n598,
    n330
  );


  buf
  g567
  (
    n618,
    n531
  );


  not
  g568
  (
    n580,
    n319
  );


  not
  g569
  (
    n611,
    n533
  );


  not
  g570
  (
    n603,
    n538
  );


  buf
  g571
  (
    n606,
    n311
  );


  buf
  g572
  (
    n592,
    n531
  );


  buf
  g573
  (
    n601,
    n530
  );


  xor
  g574
  (
    n610,
    n306,
    n321,
    n538
  );


  and
  g575
  (
    n566,
    n532,
    n544,
    n320,
    n315
  );


  xor
  g576
  (
    n624,
    n330,
    n532,
    n544,
    n540
  );


  xnor
  g577
  (
    n597,
    n541,
    n535,
    n317,
    n536
  );


  or
  g578
  (
    n578,
    n528,
    n305,
    n535,
    n530
  );


  xnor
  g579
  (
    n593,
    n535,
    n529,
    n318,
    n323
  );


  nor
  g580
  (
    n554,
    n314,
    n309,
    n534,
    n487
  );


  xnor
  g581
  (
    n575,
    n532,
    n326,
    n542,
    n303
  );


  nor
  g582
  (
    n620,
    n537,
    n536,
    n539
  );


  xnor
  g583
  (
    n570,
    n543,
    n537,
    n534
  );


  and
  g584
  (
    n560,
    n543,
    n328,
    n322,
    n528
  );


  or
  g585
  (
    n612,
    n318,
    n308,
    n320,
    n542
  );


  nor
  g586
  (
    n596,
    n541,
    n313,
    n312,
    n546
  );


  and
  g587
  (
    n567,
    n544,
    n545,
    n528,
    n487
  );


  xnor
  g588
  (
    n562,
    n531,
    n539,
    n302,
    n530
  );


  nand
  g589
  (
    n571,
    n533,
    n533,
    n529,
    n306
  );


  xnor
  g590
  (
    n622,
    n546,
    n317,
    n527,
    n309
  );


  or
  g591
  (
    n621,
    n535,
    n319,
    n538,
    n325
  );


  xor
  g592
  (
    n582,
    n311,
    n542,
    n315,
    n307
  );


  or
  g593
  (
    n551,
    n543,
    n310,
    n542,
    n544
  );


  not
  g594
  (
    n776,
    n587
  );


  not
  g595
  (
    n674,
    n624
  );


  buf
  g596
  (
    n685,
    n488
  );


  not
  g597
  (
    n682,
    n467
  );


  buf
  g598
  (
    n767,
    n553
  );


  buf
  g599
  (
    n735,
    n577
  );


  not
  g600
  (
    n733,
    n383
  );


  buf
  g601
  (
    n680,
    n561
  );


  not
  g602
  (
    n744,
    n567
  );


  not
  g603
  (
    n724,
    n565
  );


  not
  g604
  (
    n713,
    n365
  );


  not
  g605
  (
    n719,
    n561
  );


  not
  g606
  (
    n649,
    n606
  );


  not
  g607
  (
    n645,
    n568
  );


  buf
  g608
  (
    n750,
    n373
  );


  not
  g609
  (
    n730,
    n624
  );


  buf
  g610
  (
    n656,
    n580
  );


  buf
  g611
  (
    n707,
    n554
  );


  buf
  g612
  (
    n742,
    n478
  );


  buf
  g613
  (
    n691,
    n588
  );


  not
  g614
  (
    n630,
    n548
  );


  not
  g615
  (
    n749,
    n601
  );


  buf
  g616
  (
    n640,
    n458
  );


  not
  g617
  (
    n709,
    n588
  );


  not
  g618
  (
    n696,
    n458
  );


  buf
  g619
  (
    n648,
    n465
  );


  buf
  g620
  (
    n771,
    n571
  );


  not
  g621
  (
    n720,
    n551
  );


  not
  g622
  (
    n659,
    n596
  );


  not
  g623
  (
    n756,
    n571
  );


  not
  g624
  (
    n688,
    n605
  );


  buf
  g625
  (
    n670,
    n556
  );


  not
  g626
  (
    n689,
    n573
  );


  buf
  g627
  (
    n651,
    n547
  );


  buf
  g628
  (
    n716,
    n614
  );


  buf
  g629
  (
    n676,
    n457
  );


  buf
  g630
  (
    n705,
    n619
  );


  not
  g631
  (
    n740,
    n564
  );


  not
  g632
  (
    n710,
    n551
  );


  buf
  g633
  (
    n660,
    n606
  );


  buf
  g634
  (
    n667,
    n573
  );


  not
  g635
  (
    n732,
    n488
  );


  not
  g636
  (
    n769,
    n379
  );


  not
  g637
  (
    n647,
    n573
  );


  not
  g638
  (
    n754,
    n581
  );


  buf
  g639
  (
    n761,
    n624
  );


  buf
  g640
  (
    n700,
    n575
  );


  buf
  g641
  (
    n655,
    n606
  );


  not
  g642
  (
    n706,
    n603
  );


  buf
  g643
  (
    n755,
    n466
  );


  buf
  g644
  (
    n753,
    n560
  );


  not
  g645
  (
    n748,
    n470
  );


  buf
  g646
  (
    n775,
    n599
  );


  buf
  g647
  (
    n784,
    n466
  );


  buf
  g648
  (
    n665,
    n555
  );


  not
  g649
  (
    n677,
    n586
  );


  buf
  g650
  (
    n736,
    n587
  );


  not
  g651
  (
    n638,
    n567
  );


  buf
  g652
  (
    n652,
    n591
  );


  buf
  g653
  (
    n758,
    n607
  );


  not
  g654
  (
    n639,
    n571
  );


  not
  g655
  (
    n686,
    n615
  );


  buf
  g656
  (
    n702,
    n557
  );


  buf
  g657
  (
    n701,
    n489
  );


  buf
  g658
  (
    n773,
    n600
  );


  not
  g659
  (
    n778,
    n557
  );


  buf
  g660
  (
    n687,
    n590
  );


  not
  g661
  (
    n658,
    n367
  );


  buf
  g662
  (
    n781,
    n580
  );


  not
  g663
  (
    n727,
    n620
  );


  buf
  g664
  (
    KeyWire_0_1,
    n622
  );


  not
  g665
  (
    n650,
    n457
  );


  not
  g666
  (
    n734,
    n600
  );


  not
  g667
  (
    n721,
    n460
  );


  or
  g668
  (
    n698,
    n586,
    n385,
    n610,
    n598
  );


  nor
  g669
  (
    n671,
    n468,
    n614,
    n615,
    n622
  );


  or
  g670
  (
    n783,
    n597,
    n591,
    n462,
    n607
  );


  xnor
  g671
  (
    n693,
    n470,
    n590,
    n460,
    n551
  );


  nand
  g672
  (
    n695,
    n581,
    n567,
    n376,
    n571
  );


  or
  g673
  (
    n627,
    n619,
    n582,
    n565,
    n461
  );


  and
  g674
  (
    n729,
    n570,
    n581,
    n584,
    n489
  );


  nand
  g675
  (
    n643,
    n595,
    n575,
    n626,
    n558
  );


  nor
  g676
  (
    n715,
    n583,
    n620,
    n464,
    n567
  );


  xor
  g677
  (
    n703,
    n489,
    n613,
    n611,
    n596
  );


  xnor
  g678
  (
    n739,
    n613,
    n607,
    n461,
    n366
  );


  xnor
  g679
  (
    n664,
    n464,
    n622,
    n370,
    n469
  );


  xnor
  g680
  (
    n722,
    n466,
    n574,
    n595,
    n550
  );


  nor
  g681
  (
    n768,
    n621,
    n461,
    n564,
    n593
  );


  xor
  g682
  (
    n766,
    n574,
    n597,
    n570,
    n623
  );


  xnor
  g683
  (
    n780,
    n547,
    n465,
    n590,
    n626
  );


  xor
  g684
  (
    n637,
    n604,
    n575,
    n611,
    n580
  );


  nand
  g685
  (
    n673,
    n586,
    n601,
    n550,
    n559
  );


  nand
  g686
  (
    n708,
    n549,
    n609,
    n604,
    n566
  );


  or
  g687
  (
    n681,
    n592,
    n471,
    n589,
    n603
  );


  xor
  g688
  (
    n770,
    n625,
    n462,
    n378,
    n548
  );


  and
  g689
  (
    KeyWire_0_9,
    n471,
    n562,
    n578,
    n458
  );


  or
  g690
  (
    n697,
    n583,
    n563,
    n605,
    n553
  );


  nor
  g691
  (
    n772,
    n589,
    n603,
    n608,
    n621
  );


  and
  g692
  (
    n636,
    n596,
    n467,
    n561,
    n562
  );


  nand
  g693
  (
    n728,
    n618,
    n616,
    n467,
    n476
  );


  nand
  g694
  (
    n712,
    n586,
    n555,
    n585,
    n556
  );


  or
  g695
  (
    n762,
    n558,
    n566,
    n565,
    n605
  );


  and
  g696
  (
    n774,
    n620,
    n461,
    n602
  );


  or
  g697
  (
    n631,
    n562,
    n614,
    n578,
    n457
  );


  nand
  g698
  (
    n760,
    n613,
    n551,
    n575,
    n563
  );


  and
  g699
  (
    n642,
    n587,
    n549,
    n372,
    n550
  );


  xnor
  g700
  (
    n690,
    n599,
    n572,
    n384,
    n489
  );


  and
  g701
  (
    n741,
    n612,
    n465,
    n471,
    n469
  );


  and
  g702
  (
    n725,
    n466,
    n377,
    n615,
    n374
  );


  or
  g703
  (
    n747,
    n604,
    n610,
    n569,
    n548
  );


  and
  g704
  (
    n633,
    n622,
    n582,
    n585,
    n547
  );


  xor
  g705
  (
    n711,
    n605,
    n582,
    n554,
    n588
  );


  and
  g706
  (
    n678,
    n460,
    n617,
    n588,
    n610
  );


  xnor
  g707
  (
    n629,
    n555,
    n598,
    n553,
    n602
  );


  nand
  g708
  (
    n692,
    n566,
    n566,
    n460,
    n477
  );


  xor
  g709
  (
    n752,
    n596,
    n387,
    n623,
    n589
  );


  or
  g710
  (
    n779,
    n612,
    n560,
    n579,
    n584
  );


  or
  g711
  (
    n666,
    n577,
    n618,
    n591,
    n601
  );


  nand
  g712
  (
    n763,
    n582,
    n463,
    n459,
    n469
  );


  xor
  g713
  (
    n737,
    n469,
    n600,
    n458,
    n568
  );


  xnor
  g714
  (
    n731,
    n616,
    n611,
    n464,
    n547
  );


  nand
  g715
  (
    n699,
    n459,
    n570,
    n478,
    n624
  );


  nand
  g716
  (
    n717,
    n457,
    n578,
    n548,
    n615
  );


  nor
  g717
  (
    n684,
    n557,
    n568,
    n572,
    n625
  );


  or
  g718
  (
    n746,
    n580,
    n462,
    n554,
    n626
  );


  xnor
  g719
  (
    n661,
    n561,
    n467,
    n564,
    n593
  );


  and
  g720
  (
    n757,
    n599,
    n623,
    n597,
    n618
  );


  nor
  g721
  (
    n679,
    n609,
    n562,
    n563,
    n612
  );


  nor
  g722
  (
    n714,
    n570,
    n604,
    n368,
    n463
  );


  or
  g723
  (
    n765,
    n364,
    n581,
    n552,
    n602
  );


  and
  g724
  (
    n718,
    n618,
    n584,
    n555,
    n620
  );


  and
  g725
  (
    n704,
    n565,
    n559,
    n556,
    n619
  );


  xnor
  g726
  (
    n785,
    n594,
    n463,
    n574,
    n576
  );


  nor
  g727
  (
    n653,
    n568,
    n599,
    n608,
    n593
  );


  or
  g728
  (
    n777,
    n577,
    n552,
    n549,
    n550
  );


  xor
  g729
  (
    n759,
    n584,
    n606,
    n557,
    n585
  );


  and
  g730
  (
    n669,
    n592,
    n552,
    n470,
    n625
  );


  and
  g731
  (
    n675,
    n583,
    n381,
    n616,
    n577
  );


  nand
  g732
  (
    n632,
    n614,
    n576,
    n558,
    n598
  );


  xor
  g733
  (
    n634,
    n592,
    n600,
    n576,
    n569
  );


  and
  g734
  (
    n743,
    n558,
    n371,
    n598,
    n590
  );


  nand
  g735
  (
    n662,
    n476,
    n463,
    n613,
    n459
  );


  nand
  g736
  (
    n672,
    n623,
    n608,
    n369,
    n552
  );


  nor
  g737
  (
    n764,
    n585,
    n559,
    n462,
    n587
  );


  nand
  g738
  (
    n635,
    n564,
    n609,
    n569,
    n553
  );


  nand
  g739
  (
    n694,
    n456,
    n612,
    n601,
    n576
  );


  and
  g740
  (
    n663,
    n616,
    n617,
    n574,
    n468
  );


  or
  g741
  (
    n786,
    n560,
    n603,
    n465,
    n594
  );


  and
  g742
  (
    n628,
    n607,
    n464,
    n593,
    n621
  );


  and
  g743
  (
    KeyWire_0_8,
    n611,
    n556,
    n595,
    n594
  );


  and
  g744
  (
    n668,
    n563,
    n572,
    n470,
    n573
  );


  xnor
  g745
  (
    KeyWire_0_15,
    n589,
    n609,
    n583,
    n387
  );


  xor
  g746
  (
    n654,
    n560,
    n578,
    n375,
    n382
  );


  and
  g747
  (
    n738,
    n468,
    n569,
    n554,
    n386
  );


  and
  g748
  (
    n723,
    n591,
    n617,
    n621,
    n595
  );


  and
  g749
  (
    n644,
    n579,
    n617,
    n471,
    n619
  );


  xor
  g750
  (
    n646,
    n579,
    n594,
    n549,
    n625
  );


  and
  g751
  (
    n641,
    n579,
    n559,
    n459,
    n610
  );


  xor
  g752
  (
    n726,
    n572,
    n592,
    n468,
    n626
  );


  nand
  g753
  (
    n782,
    n608,
    n477,
    n380,
    n597
  );


  and
  g754
  (
    n814,
    n752,
    n629,
    n663,
    n755
  );


  or
  g755
  (
    n790,
    n747,
    n742,
    n709,
    n776
  );


  nor
  g756
  (
    n808,
    n711,
    n702,
    n745,
    n638
  );


  or
  g757
  (
    n822,
    n763,
    n769,
    n675,
    n647
  );


  nand
  g758
  (
    n810,
    n665,
    n631,
    n715,
    n782
  );


  nor
  g759
  (
    n793,
    n785,
    n771,
    n720,
    n768
  );


  xor
  g760
  (
    n817,
    n764,
    n698,
    n700,
    n693
  );


  or
  g761
  (
    KeyWire_0_7,
    n646,
    n632,
    n744,
    n657
  );


  nor
  g762
  (
    n823,
    n682,
    n681,
    n740,
    n724
  );


  or
  g763
  (
    n792,
    n659,
    n666,
    n680,
    n777
  );


  and
  g764
  (
    KeyWire_0_4,
    n718,
    n651,
    n635,
    n759
  );


  or
  g765
  (
    n815,
    n705,
    n754,
    n684,
    n630
  );


  nor
  g766
  (
    n819,
    n670,
    n689,
    n644,
    n673
  );


  or
  g767
  (
    KeyWire_0_11,
    n712,
    n733,
    n726,
    n750
  );


  xnor
  g768
  (
    n807,
    n645,
    n784,
    n654,
    n757
  );


  and
  g769
  (
    n821,
    n737,
    n761,
    n655,
    n643
  );


  or
  g770
  (
    n799,
    n692,
    n708,
    n767,
    n739
  );


  xnor
  g771
  (
    n803,
    n628,
    n751,
    n649,
    n719
  );


  nor
  g772
  (
    n811,
    n773,
    n694,
    n753,
    n701
  );


  nor
  g773
  (
    n816,
    n674,
    n721,
    n710,
    n687
  );


  and
  g774
  (
    n802,
    n770,
    n738,
    n662,
    n717
  );


  xor
  g775
  (
    n806,
    n671,
    n778,
    n648,
    n633
  );


  nor
  g776
  (
    n787,
    n716,
    n758,
    n762,
    n735
  );


  and
  g777
  (
    n798,
    n697,
    n756,
    n690,
    n704
  );


  nor
  g778
  (
    n794,
    n730,
    n783,
    n713,
    n660
  );


  xnor
  g779
  (
    n824,
    n736,
    n696,
    n652,
    n766
  );


  nand
  g780
  (
    n813,
    n781,
    n748,
    n683,
    n707
  );


  xor
  g781
  (
    n818,
    n685,
    n637,
    n634,
    n760
  );


  xnor
  g782
  (
    n797,
    n786,
    n722,
    n775,
    n765
  );


  and
  g783
  (
    n805,
    n678,
    n639,
    n734,
    n691
  );


  or
  g784
  (
    n820,
    n636,
    n714,
    n743,
    n725
  );


  xnor
  g785
  (
    n795,
    n706,
    n668,
    n642,
    n664
  );


  xor
  g786
  (
    n809,
    n741,
    n661,
    n779,
    n627
  );


  xnor
  g787
  (
    n812,
    n729,
    n732,
    n772,
    n780
  );


  and
  g788
  (
    n804,
    n676,
    n723,
    n728,
    n650
  );


  nor
  g789
  (
    n826,
    n656,
    n672,
    n688,
    n667
  );


  nor
  g790
  (
    n788,
    n703,
    n727,
    n641,
    n658
  );


  xnor
  g791
  (
    n789,
    n746,
    n774,
    n686,
    n749
  );


  nor
  g792
  (
    n800,
    n699,
    n653,
    n640,
    n669
  );


  and
  g793
  (
    n801,
    n695,
    n679,
    n731,
    n677
  );


  nor
  g794
  (
    n833,
    n821,
    n805,
    n813,
    n815
  );


  xnor
  g795
  (
    n834,
    n807,
    n809,
    n803,
    n823
  );


  or
  g796
  (
    n831,
    n814,
    n822,
    n792,
    n812
  );


  xnor
  g797
  (
    n829,
    n818,
    n801,
    n798,
    n791
  );


  nor
  g798
  (
    n828,
    n816,
    n788,
    n806,
    n825
  );


  or
  g799
  (
    n832,
    n819,
    n789,
    n810,
    n790
  );


  or
  g800
  (
    n830,
    n811,
    n808,
    n794,
    n795
  );


  nand
  g801
  (
    n835,
    n802,
    n804,
    n796,
    n787
  );


  xnor
  g802
  (
    n836,
    n824,
    n793,
    n817,
    n826
  );


  nand
  g803
  (
    n827,
    n799,
    n820,
    n797,
    n800
  );


  xnor
  KeyGate_0_0
  (
    n94,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n657,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n529,
    KeyNOTWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n581,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n825,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n368,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n48,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n791,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n745,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n683,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n201,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n796,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n547,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n200,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n227,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n751,
    KeyNOTWire_0_15
  );


endmodule

