// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1436_31_3 written by SynthGen on 2021/05/24 19:45:40
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1436_31_3 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26,
 n1241, n1303, n1310, n1313, n1305, n1306, n1309, n1311,
 n1301, n1367, n1357, n1355, n1363, n1353, n1358, n1366,
 n1370, n1368, n1359, n1462);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26;

output n1241, n1303, n1310, n1313, n1305, n1306, n1309, n1311,
 n1301, n1367, n1357, n1355, n1363, n1353, n1358, n1366,
 n1370, n1368, n1359, n1462;

wire n27, n28, n29, n30, n31, n32, n33, n34,
 n35, n36, n37, n38, n39, n40, n41, n42,
 n43, n44, n45, n46, n47, n48, n49, n50,
 n51, n52, n53, n54, n55, n56, n57, n58,
 n59, n60, n61, n62, n63, n64, n65, n66,
 n67, n68, n69, n70, n71, n72, n73, n74,
 n75, n76, n77, n78, n79, n80, n81, n82,
 n83, n84, n85, n86, n87, n88, n89, n90,
 n91, n92, n93, n94, n95, n96, n97, n98,
 n99, n100, n101, n102, n103, n104, n105, n106,
 n107, n108, n109, n110, n111, n112, n113, n114,
 n115, n116, n117, n118, n119, n120, n121, n122,
 n123, n124, n125, n126, n127, n128, n129, n130,
 n131, n132, n133, n134, n135, n136, n137, n138,
 n139, n140, n141, n142, n143, n144, n145, n146,
 n147, n148, n149, n150, n151, n152, n153, n154,
 n155, n156, n157, n158, n159, n160, n161, n162,
 n163, n164, n165, n166, n167, n168, n169, n170,
 n171, n172, n173, n174, n175, n176, n177, n178,
 n179, n180, n181, n182, n183, n184, n185, n186,
 n187, n188, n189, n190, n191, n192, n193, n194,
 n195, n196, n197, n198, n199, n200, n201, n202,
 n203, n204, n205, n206, n207, n208, n209, n210,
 n211, n212, n213, n214, n215, n216, n217, n218,
 n219, n220, n221, n222, n223, n224, n225, n226,
 n227, n228, n229, n230, n231, n232, n233, n234,
 n235, n236, n237, n238, n239, n240, n241, n242,
 n243, n244, n245, n246, n247, n248, n249, n250,
 n251, n252, n253, n254, n255, n256, n257, n258,
 n259, n260, n261, n262, n263, n264, n265, n266,
 n267, n268, n269, n270, n271, n272, n273, n274,
 n275, n276, n277, n278, n279, n280, n281, n282,
 n283, n284, n285, n286, n287, n288, n289, n290,
 n291, n292, n293, n294, n295, n296, n297, n298,
 n299, n300, n301, n302, n303, n304, n305, n306,
 n307, n308, n309, n310, n311, n312, n313, n314,
 n315, n316, n317, n318, n319, n320, n321, n322,
 n323, n324, n325, n326, n327, n328, n329, n330,
 n331, n332, n333, n334, n335, n336, n337, n338,
 n339, n340, n341, n342, n343, n344, n345, n346,
 n347, n348, n349, n350, n351, n352, n353, n354,
 n355, n356, n357, n358, n359, n360, n361, n362,
 n363, n364, n365, n366, n367, n368, n369, n370,
 n371, n372, n373, n374, n375, n376, n377, n378,
 n379, n380, n381, n382, n383, n384, n385, n386,
 n387, n388, n389, n390, n391, n392, n393, n394,
 n395, n396, n397, n398, n399, n400, n401, n402,
 n403, n404, n405, n406, n407, n408, n409, n410,
 n411, n412, n413, n414, n415, n416, n417, n418,
 n419, n420, n421, n422, n423, n424, n425, n426,
 n427, n428, n429, n430, n431, n432, n433, n434,
 n435, n436, n437, n438, n439, n440, n441, n442,
 n443, n444, n445, n446, n447, n448, n449, n450,
 n451, n452, n453, n454, n455, n456, n457, n458,
 n459, n460, n461, n462, n463, n464, n465, n466,
 n467, n468, n469, n470, n471, n472, n473, n474,
 n475, n476, n477, n478, n479, n480, n481, n482,
 n483, n484, n485, n486, n487, n488, n489, n490,
 n491, n492, n493, n494, n495, n496, n497, n498,
 n499, n500, n501, n502, n503, n504, n505, n506,
 n507, n508, n509, n510, n511, n512, n513, n514,
 n515, n516, n517, n518, n519, n520, n521, n522,
 n523, n524, n525, n526, n527, n528, n529, n530,
 n531, n532, n533, n534, n535, n536, n537, n538,
 n539, n540, n541, n542, n543, n544, n545, n546,
 n547, n548, n549, n550, n551, n552, n553, n554,
 n555, n556, n557, n558, n559, n560, n561, n562,
 n563, n564, n565, n566, n567, n568, n569, n570,
 n571, n572, n573, n574, n575, n576, n577, n578,
 n579, n580, n581, n582, n583, n584, n585, n586,
 n587, n588, n589, n590, n591, n592, n593, n594,
 n595, n596, n597, n598, n599, n600, n601, n602,
 n603, n604, n605, n606, n607, n608, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n660, n661, n662, n663, n664, n665, n666,
 n667, n668, n669, n670, n671, n672, n673, n674,
 n675, n676, n677, n678, n679, n680, n681, n682,
 n683, n684, n685, n686, n687, n688, n689, n690,
 n691, n692, n693, n694, n695, n696, n697, n698,
 n699, n700, n701, n702, n703, n704, n705, n706,
 n707, n708, n709, n710, n711, n712, n713, n714,
 n715, n716, n717, n718, n719, n720, n721, n722,
 n723, n724, n725, n726, n727, n728, n729, n730,
 n731, n732, n733, n734, n735, n736, n737, n738,
 n739, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1242, n1243,
 n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
 n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
 n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
 n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
 n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
 n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
 n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
 n1300, n1302, n1304, n1307, n1308, n1312, n1314, n1315,
 n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
 n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
 n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
 n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
 n1348, n1349, n1350, n1351, n1352, n1354, n1356, n1360,
 n1361, n1362, n1364, n1365, n1369, n1371, n1372, n1373,
 n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
 n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
 n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
 n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
 n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
 n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
 n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
 n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
 n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
 n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
 n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461;

not  g0 (n96, n4);
buf  g1 (n35, n26);
not  g2 (n126, n2);
not  g3 (n38, n10);
not  g4 (n49, n5);
buf  g5 (n108, n24);
not  g6 (n82, n4);
not  g7 (n98, n19);
buf  g8 (n83, n26);
not  g9 (n41, n23);
not  g10 (n92, n11);
buf  g11 (n52, n12);
not  g12 (n53, n7);
buf  g13 (n84, n4);
buf  g14 (n47, n15);
buf  g15 (n91, n5);
buf  g16 (n94, n18);
buf  g17 (n33, n14);
not  g18 (n62, n17);
not  g19 (n70, n24);
buf  g20 (n37, n24);
not  g21 (n107, n2);
buf  g22 (n34, n21);
buf  g23 (n89, n16);
buf  g24 (n60, n19);
not  g25 (n28, n1);
buf  g26 (n43, n25);
buf  g27 (n90, n23);
not  g28 (n128, n11);
buf  g29 (n57, n9);
not  g30 (n30, n24);
not  g31 (n44, n18);
not  g32 (n120, n7);
buf  g33 (n95, n16);
buf  g34 (n106, n9);
not  g35 (n63, n19);
buf  g36 (n127, n15);
buf  g37 (n117, n10);
buf  g38 (n122, n3);
not  g39 (n125, n15);
not  g40 (n99, n25);
not  g41 (n58, n23);
not  g42 (n66, n20);
not  g43 (n65, n21);
not  g44 (n112, n22);
buf  g45 (n102, n21);
buf  g46 (n29, n1);
not  g47 (n67, n14);
buf  g48 (n85, n15);
not  g49 (n76, n6);
not  g50 (n45, n12);
buf  g51 (n74, n8);
not  g52 (n32, n6);
buf  g53 (n72, n20);
buf  g54 (n64, n26);
buf  g55 (n71, n8);
not  g56 (n68, n22);
not  g57 (n61, n11);
not  g58 (n55, n3);
not  g59 (n113, n5);
buf  g60 (n111, n18);
not  g61 (n97, n23);
not  g62 (n88, n11);
buf  g63 (n40, n3);
not  g64 (n39, n10);
buf  g65 (n86, n14);
buf  g66 (n105, n14);
buf  g67 (n118, n5);
buf  g68 (n115, n6);
not  g69 (n42, n1);
buf  g70 (n50, n12);
buf  g71 (n101, n19);
not  g72 (n114, n22);
buf  g73 (n79, n16);
buf  g74 (n110, n17);
buf  g75 (n103, n8);
not  g76 (n109, n20);
buf  g77 (n36, n8);
not  g78 (n81, n10);
not  g79 (n104, n9);
buf  g80 (n93, n21);
buf  g81 (n69, n25);
buf  g82 (n124, n9);
buf  g83 (n121, n13);
not  g84 (n75, n17);
not  g85 (n77, n1);
buf  g86 (n59, n26);
not  g87 (n80, n13);
buf  g88 (n78, n18);
not  g89 (n51, n25);
buf  g90 (n116, n17);
not  g91 (n129, n2);
buf  g92 (n100, n6);
buf  g93 (n31, n3);
not  g94 (n87, n7);
not  g95 (n73, n13);
buf  g96 (n54, n20);
buf  g97 (n48, n12);
not  g98 (n27, n2);
buf  g99 (n119, n4);
buf  g100 (n123, n13);
buf  g101 (n56, n7);
not  g102 (n46, n22);
buf  g103 (n130, n16);
not  g104 (n394, n124);
buf  g105 (n255, n70);
buf  g106 (n515, n95);
not  g107 (n299, n127);
buf  g108 (n423, n69);
not  g109 (n189, n65);
buf  g110 (n228, n39);
buf  g111 (n187, n30);
not  g112 (n356, n114);
not  g113 (n155, n112);
buf  g114 (n240, n73);
buf  g115 (n320, n77);
buf  g116 (n408, n129);
buf  g117 (n263, n85);
not  g118 (n289, n101);
buf  g119 (n424, n85);
buf  g120 (n333, n48);
not  g121 (n532, n50);
buf  g122 (n524, n51);
not  g123 (n301, n44);
buf  g124 (n416, n43);
not  g125 (n495, n119);
buf  g126 (n164, n70);
not  g127 (n251, n103);
not  g128 (n428, n67);
buf  g129 (n481, n127);
not  g130 (n150, n87);
not  g131 (n345, n31);
buf  g132 (n530, n62);
buf  g133 (n201, n105);
not  g134 (n279, n82);
buf  g135 (n519, n97);
buf  g136 (n329, n43);
not  g137 (n304, n35);
buf  g138 (n466, n29);
buf  g139 (n435, n56);
buf  g140 (n160, n44);
buf  g141 (n477, n51);
buf  g142 (n199, n108);
buf  g143 (n148, n33);
buf  g144 (n206, n111);
not  g145 (n382, n66);
not  g146 (n285, n40);
buf  g147 (n151, n53);
buf  g148 (n411, n65);
not  g149 (n476, n101);
not  g150 (n318, n98);
buf  g151 (n173, n122);
buf  g152 (n244, n113);
buf  g153 (n236, n68);
not  g154 (n305, n128);
not  g155 (n259, n74);
buf  g156 (n241, n30);
not  g157 (n494, n110);
not  g158 (n331, n40);
not  g159 (n439, n82);
buf  g160 (n312, n95);
not  g161 (n385, n37);
not  g162 (n488, n118);
buf  g163 (n268, n86);
buf  g164 (n499, n130);
not  g165 (n485, n91);
buf  g166 (n195, n57);
not  g167 (n307, n42);
buf  g168 (n438, n87);
not  g169 (n309, n105);
not  g170 (n487, n50);
buf  g171 (n483, n28);
not  g172 (n252, n80);
not  g173 (n381, n59);
buf  g174 (n321, n100);
not  g175 (n174, n56);
not  g176 (n194, n49);
not  g177 (n256, n98);
buf  g178 (n291, n74);
not  g179 (n462, n64);
not  g180 (n340, n79);
buf  g181 (n429, n113);
buf  g182 (n232, n100);
not  g183 (n288, n55);
not  g184 (n149, n122);
not  g185 (n544, n61);
buf  g186 (n358, n36);
buf  g187 (n425, n47);
not  g188 (n245, n89);
buf  g189 (n175, n83);
buf  g190 (n469, n94);
buf  g191 (n342, n128);
not  g192 (n351, n58);
buf  g193 (n503, n72);
buf  g194 (n498, n130);
not  g195 (n354, n102);
not  g196 (n242, n79);
buf  g197 (n138, n67);
buf  g198 (n541, n45);
not  g199 (n396, n92);
buf  g200 (n357, n64);
not  g201 (n190, n49);
buf  g202 (n296, n27);
buf  g203 (n426, n62);
buf  g204 (n414, n64);
not  g205 (n472, n111);
not  g206 (n520, n35);
not  g207 (n522, n109);
buf  g208 (n336, n124);
not  g209 (n440, n120);
buf  g210 (n311, n61);
not  g211 (n379, n54);
buf  g212 (n167, n59);
not  g213 (n225, n41);
not  g214 (n389, n59);
not  g215 (n172, n72);
not  g216 (n535, n47);
not  g217 (n516, n105);
not  g218 (n538, n115);
not  g219 (n184, n76);
not  g220 (n243, n92);
not  g221 (n412, n45);
not  g222 (n274, n111);
not  g223 (n267, n129);
buf  g224 (n310, n129);
buf  g225 (n334, n120);
not  g226 (n161, n112);
buf  g227 (n246, n116);
not  g228 (n393, n117);
not  g229 (n493, n75);
not  g230 (n168, n115);
buf  g231 (n355, n113);
buf  g232 (n276, n28);
buf  g233 (n534, n106);
buf  g234 (n402, n125);
not  g235 (n446, n121);
not  g236 (n528, n39);
not  g237 (n217, n93);
buf  g238 (n445, n70);
buf  g239 (n509, n96);
not  g240 (n459, n86);
not  g241 (n457, n117);
buf  g242 (n395, n93);
not  g243 (n529, n34);
buf  g244 (n480, n49);
not  g245 (n448, n29);
buf  g246 (n237, n121);
not  g247 (n332, n100);
not  g248 (n370, n93);
not  g249 (n227, n40);
buf  g250 (n341, n126);
not  g251 (n271, n71);
not  g252 (n364, n107);
not  g253 (n328, n52);
buf  g254 (n543, n102);
not  g255 (n162, n60);
buf  g256 (n359, n27);
not  g257 (n501, n113);
buf  g258 (n292, n57);
not  g259 (n421, n37);
buf  g260 (n514, n118);
not  g261 (n221, n95);
not  g262 (n506, n36);
buf  g263 (n179, n119);
buf  g264 (n399, n53);
buf  g265 (n275, n66);
buf  g266 (n250, n35);
not  g267 (n171, n52);
buf  g268 (n436, n73);
buf  g269 (n343, n109);
buf  g270 (n369, n41);
buf  g271 (n204, n74);
not  g272 (n239, n99);
not  g273 (n454, n46);
not  g274 (n475, n85);
not  g275 (n400, n109);
not  g276 (n388, n29);
buf  g277 (n461, n29);
buf  g278 (n384, n50);
buf  g279 (n234, n119);
not  g280 (n387, n77);
not  g281 (n193, n108);
not  g282 (n365, n94);
not  g283 (n492, n71);
not  g284 (n235, n32);
not  g285 (n473, n116);
buf  g286 (n185, n119);
buf  g287 (n135, n54);
buf  g288 (n441, n27);
not  g289 (n474, n91);
buf  g290 (n390, n89);
buf  g291 (n181, n111);
buf  g292 (n373, n64);
buf  g293 (n542, n103);
buf  g294 (n319, n92);
buf  g295 (n407, n74);
not  g296 (n266, n48);
not  g297 (n368, n99);
buf  g298 (n478, n75);
buf  g299 (n419, n31);
not  g300 (n417, n38);
not  g301 (n497, n90);
not  g302 (n323, n68);
not  g303 (n418, n83);
not  g304 (n208, n61);
not  g305 (n460, n97);
buf  g306 (n145, n46);
not  g307 (n451, n89);
buf  g308 (n360, n105);
buf  g309 (n484, n81);
buf  g310 (n152, n88);
buf  g311 (n182, n95);
buf  g312 (n437, n55);
buf  g313 (n410, n122);
not  g314 (n537, n110);
not  g315 (n264, n36);
buf  g316 (n531, n103);
not  g317 (n447, n77);
buf  g318 (n527, n125);
not  g319 (n479, n45);
not  g320 (n432, n94);
buf  g321 (n482, n86);
not  g322 (n330, n127);
buf  g323 (n386, n75);
buf  g324 (n363, n115);
not  g325 (n265, n54);
not  g326 (n504, n63);
buf  g327 (n324, n116);
buf  g328 (n218, n114);
not  g329 (n283, n97);
not  g330 (n362, n78);
not  g331 (n133, n32);
buf  g332 (n261, n126);
not  g333 (n219, n51);
not  g334 (n147, n104);
not  g335 (n545, n128);
buf  g336 (n391, n84);
buf  g337 (n293, n51);
buf  g338 (n280, n104);
buf  g339 (n202, n98);
not  g340 (n380, n33);
not  g341 (n361, n88);
not  g342 (n348, n116);
not  g343 (n282, n40);
not  g344 (n143, n27);
not  g345 (n372, n87);
buf  g346 (n486, n96);
buf  g347 (n277, n129);
not  g348 (n403, n126);
buf  g349 (n508, n54);
not  g350 (n347, n48);
buf  g351 (n231, n104);
buf  g352 (n525, n81);
not  g353 (n518, n124);
not  g354 (n196, n78);
not  g355 (n298, n32);
not  g356 (n287, n57);
buf  g357 (n496, n127);
buf  g358 (n316, n85);
buf  g359 (n270, n102);
not  g360 (n349, n91);
buf  g361 (n197, n120);
buf  g362 (n207, n88);
not  g363 (n213, n106);
buf  g364 (n546, n109);
buf  g365 (n353, n28);
buf  g366 (n502, n106);
not  g367 (n450, n44);
buf  g368 (n224, n82);
not  g369 (n470, n38);
buf  g370 (n272, n34);
buf  g371 (n339, n128);
not  g372 (n281, n117);
not  g373 (n183, n47);
buf  g374 (n452, n86);
not  g375 (n223, n94);
buf  g376 (n464, n34);
buf  g377 (n322, n50);
buf  g378 (n521, n48);
not  g379 (n453, n76);
not  g380 (n352, n110);
buf  g381 (n229, n58);
not  g382 (n415, n123);
not  g383 (n366, n39);
not  g384 (n286, n71);
not  g385 (n404, n102);
not  g386 (n378, n123);
not  g387 (n420, n120);
not  g388 (n203, n114);
buf  g389 (n533, n121);
buf  g390 (n490, n130);
buf  g391 (n491, n90);
not  g392 (n191, n38);
buf  g393 (n159, n130);
not  g394 (n401, n73);
not  g395 (n433, n83);
not  g396 (n313, n80);
buf  g397 (n434, n106);
not  g398 (n295, n108);
not  g399 (n297, n60);
not  g400 (n338, n55);
not  g401 (n214, n38);
buf  g402 (n269, n87);
buf  g403 (n489, n72);
buf  g404 (n383, n36);
not  g405 (n144, n117);
buf  g406 (n463, n30);
buf  g407 (n294, n96);
not  g408 (n146, n52);
not  g409 (n180, n69);
buf  g410 (n216, n41);
not  g411 (n539, n114);
buf  g412 (n156, n107);
buf  g413 (n377, n99);
buf  g414 (n376, n76);
not  g415 (n248, n98);
buf  g416 (n536, n62);
buf  g417 (n517, n83);
buf  g418 (n137, n80);
buf  g419 (n230, n67);
buf  g420 (n157, n122);
not  g421 (n317, n118);
not  g422 (n131, n79);
not  g423 (n211, n66);
not  g424 (n188, n53);
not  g425 (n176, n93);
buf  g426 (n284, n84);
buf  g427 (n468, n33);
buf  g428 (n247, n97);
buf  g429 (n507, n82);
not  g430 (n513, n79);
not  g431 (n153, n57);
not  g432 (n132, n110);
not  g433 (n178, n32);
not  g434 (n170, n72);
buf  g435 (n141, n60);
buf  g436 (n290, n43);
not  g437 (n413, n42);
buf  g438 (n215, n42);
buf  g439 (n158, n56);
not  g440 (n306, n107);
buf  g441 (n374, n69);
not  g442 (n371, n78);
not  g443 (n142, n77);
buf  g444 (n210, n104);
not  g445 (n262, n80);
buf  g446 (n200, n60);
buf  g447 (n136, n58);
buf  g448 (n273, n46);
not  g449 (n166, n90);
buf  g450 (n406, n53);
not  g451 (n505, n30);
not  g452 (n335, n35);
not  g453 (n222, n33);
buf  g454 (n163, n124);
not  g455 (n367, n121);
buf  g456 (n500, n107);
not  g457 (n212, n81);
buf  g458 (n327, n126);
not  g459 (n444, n49);
buf  g460 (n165, n84);
not  g461 (n465, n112);
buf  g462 (n430, n76);
not  g463 (n422, n123);
buf  g464 (n134, n63);
buf  g465 (n169, n75);
buf  g466 (n140, n103);
not  g467 (n409, n66);
buf  g468 (n375, n118);
buf  g469 (n467, n91);
not  g470 (n209, n34);
not  g471 (n392, n55);
not  g472 (n456, n52);
buf  g473 (n257, n28);
not  g474 (n337, n108);
buf  g475 (n192, n58);
buf  g476 (n302, n68);
not  g477 (n471, n39);
not  g478 (n238, n43);
buf  g479 (n512, n63);
not  g480 (n260, n96);
not  g481 (n249, n101);
buf  g482 (n300, n73);
buf  g483 (n540, n92);
not  g484 (n431, n41);
not  g485 (n398, n125);
buf  g486 (n346, n88);
buf  g487 (n177, n100);
buf  g488 (n186, n44);
not  g489 (n308, n84);
buf  g490 (n278, n61);
buf  g491 (n455, n37);
not  g492 (n427, n125);
buf  g493 (n314, n37);
buf  g494 (n258, n47);
not  g495 (n139, n31);
not  g496 (n233, n101);
not  g497 (n253, n46);
not  g498 (n458, n42);
buf  g499 (n325, n115);
buf  g500 (n326, n59);
buf  g501 (n198, n31);
not  g502 (n510, n68);
buf  g503 (n344, n112);
buf  g504 (n405, n99);
buf  g505 (n315, n70);
not  g506 (n205, n62);
not  g507 (n449, n45);
buf  g508 (n220, n69);
buf  g509 (n443, n78);
buf  g510 (n303, n90);
buf  g511 (n226, n71);
buf  g512 (n154, n65);
buf  g513 (n511, n65);
not  g514 (n523, n67);
not  g515 (n526, n81);
not  g516 (n254, n89);
buf  g517 (n397, n123);
not  g518 (n442, n63);
buf  g519 (n350, n56);
not  g520 (n547, n134);
buf  g521 (n550, n133);
buf  g522 (n549, n131);
buf  g523 (n548, n132);
nor  g524 (n553, n140, n168, n181, n550);
nand g525 (n560, n142, n138, n548, n148);
xor  g526 (n559, n139, n151, n150, n165);
nand g527 (n565, n170, n163, n167, n147);
xnor g528 (n556, n550, n145, n164, n547);
xor  g529 (n564, n160, n156, n161, n152);
xor  g530 (n561, n166, n171, n143, n182);
xnor g531 (n551, n175, n550, n548, n179);
xnor g532 (n554, n172, n153, n149, n169);
nor  g533 (n558, n155, n549, n141);
or   g534 (n563, n549, n548, n162, n146);
xnor g535 (n555, n144, n176, n549, n178);
nor  g536 (n562, n135, n137, n180, n548);
nand g537 (n557, n173, n174, n158, n547);
or   g538 (n566, n136, n547, n159);
and  g539 (n552, n154, n550, n177, n157);
buf  g540 (n587, n554);
not  g541 (n578, n561);
not  g542 (n576, n562);
buf  g543 (n608, n551);
not  g544 (n601, n557);
not  g545 (n589, n565);
buf  g546 (n583, n558);
buf  g547 (n597, n556);
not  g548 (n616, n560);
buf  g549 (n577, n556);
not  g550 (n595, n562);
buf  g551 (n584, n559);
not  g552 (n590, n563);
buf  g553 (n607, n562);
buf  g554 (n572, n565);
not  g555 (n586, n558);
not  g556 (n605, n555);
buf  g557 (n606, n558);
buf  g558 (n610, n555);
not  g559 (n594, n565);
buf  g560 (n588, n564);
not  g561 (n580, n552);
not  g562 (n573, n553);
not  g563 (n585, n557);
buf  g564 (n600, n566);
buf  g565 (n567, n183);
buf  g566 (n579, n564);
buf  g567 (n581, n557);
not  g568 (n603, n565);
buf  g569 (n582, n559);
not  g570 (n593, n564);
buf  g571 (n592, n563);
not  g572 (n599, n566);
buf  g573 (n571, n559);
buf  g574 (n609, n557);
buf  g575 (n602, n563);
not  g576 (n604, n564);
not  g577 (n598, n561);
not  g578 (n615, n560);
buf  g579 (n596, n563);
buf  g580 (n575, n560);
not  g581 (n611, n561);
not  g582 (n591, n561);
not  g583 (n569, n556);
not  g584 (n612, n562);
buf  g585 (n614, n559);
not  g586 (n570, n566);
buf  g587 (n568, n566);
buf  g588 (n574, n558);
xnor g589 (n613, n556, n560);
buf  g590 (n707, n611);
not  g591 (n728, n276);
buf  g592 (n665, n614);
buf  g593 (n810, n584);
buf  g594 (n736, n587);
buf  g595 (n759, n206);
buf  g596 (n708, n341);
not  g597 (n706, n603);
not  g598 (n625, n312);
buf  g599 (n714, n187);
buf  g600 (n619, n346);
not  g601 (n727, n259);
buf  g602 (n797, n610);
not  g603 (n656, n227);
not  g604 (n791, n243);
buf  g605 (n778, n280);
buf  g606 (n767, n256);
not  g607 (n667, n591);
buf  g608 (n768, n592);
buf  g609 (n765, n577);
buf  g610 (n723, n580);
not  g611 (n637, n609);
not  g612 (n772, n596);
buf  g613 (n648, n188);
buf  g614 (n636, n198);
not  g615 (n678, n260);
not  g616 (n710, n201);
not  g617 (n680, n594);
not  g618 (n682, n572);
not  g619 (n694, n569);
not  g620 (n660, n607);
not  g621 (n739, n615);
buf  g622 (n807, n599);
not  g623 (n734, n571);
buf  g624 (n691, n586);
not  g625 (n782, n599);
not  g626 (n779, n612);
buf  g627 (n679, n269);
buf  g628 (n742, n330);
buf  g629 (n649, n306);
buf  g630 (n731, n602);
not  g631 (n754, n342);
not  g632 (n787, n610);
not  g633 (n738, n345);
buf  g634 (n816, n594);
not  g635 (n662, n303);
buf  g636 (n716, n257);
buf  g637 (n666, n578);
buf  g638 (n645, n574);
buf  g639 (n766, n592);
not  g640 (n774, n592);
buf  g641 (n740, n604);
not  g642 (n663, n570);
buf  g643 (n659, n231);
not  g644 (n721, n321);
buf  g645 (n757, n229);
buf  g646 (n802, n262);
not  g647 (n642, n591);
not  g648 (n681, n576);
buf  g649 (n713, n598);
not  g650 (n805, n203);
buf  g651 (n755, n212);
not  g652 (n704, n241);
not  g653 (n777, n258);
buf  g654 (n758, n576);
buf  g655 (n812, n239);
not  g656 (n673, n595);
not  g657 (n633, n591);
buf  g658 (n654, n585);
buf  g659 (n630, n611);
not  g660 (n687, n593);
not  g661 (n719, n613);
buf  g662 (n617, n587);
buf  g663 (n690, n582);
not  g664 (n703, n214);
buf  g665 (n650, n605);
not  g666 (n792, n308);
not  g667 (n638, n592);
buf  g668 (n702, n249);
buf  g669 (n788, n575);
not  g670 (n697, n602);
not  g671 (n647, n573);
not  g672 (n726, n568);
not  g673 (n724, n254);
buf  g674 (n790, n590);
not  g675 (n733, n583);
not  g676 (n785, n575);
not  g677 (n641, n284);
buf  g678 (n770, n612);
not  g679 (n798, n593);
buf  g680 (n639, n317);
not  g681 (n669, n261);
not  g682 (n671, n577);
buf  g683 (n741, n604);
not  g684 (n756, n221);
not  g685 (n764, n586);
buf  g686 (n729, n574);
not  g687 (n701, n602);
not  g688 (n796, n235);
not  g689 (n622, n573);
buf  g690 (n709, n304);
not  g691 (n705, n607);
buf  g692 (n771, n596);
not  g693 (n711, n238);
buf  g694 (n811, n608);
not  g695 (n730, n323);
not  g696 (n813, n339);
not  g697 (n717, n216);
not  g698 (n676, n291);
not  g699 (n698, n237);
buf  g700 (n688, n287);
buf  g701 (n808, n614);
not  g702 (n794, n332);
buf  g703 (n735, n598);
not  g704 (n627, n596);
not  g705 (n699, n575);
buf  g706 (n786, n213);
or   g707 (n628, n606, n570);
nand g708 (n799, n574, n603, n569);
nor  g709 (n806, n185, n584, n211);
xnor g710 (n780, n275, n605, n616);
nand g711 (n763, n298, n589, n594);
or   g712 (n652, n606, n569, n571);
or   g713 (n775, n595, n322, n334);
xnor g714 (n675, n290, n593, n265);
nor  g715 (n651, n193, n587, n604);
or   g716 (n664, n293, n315, n569);
nor  g717 (n658, n347, n590, n319);
or   g718 (n684, n255, n210, n335);
nand g719 (n640, n578, n200, n307);
nor  g720 (n635, n197, n208, n190);
xnor g721 (n769, n314, n266, n595);
nand g722 (n624, n340, n209, n590);
or   g723 (n644, n612, n297, n609);
xor  g724 (n720, n585, n184, n601);
and  g725 (n693, n578, n600, n590);
and  g726 (n745, n609, n616, n604);
and  g727 (n631, n337, n348, n250);
nor  g728 (n781, n300, n274, n302);
nand g729 (n661, n199, n588, n584);
nand g730 (n689, n600, n579, n202);
and  g731 (n732, n615, n224, n582);
nand g732 (n696, n603, n244, n586);
nand g733 (n773, n613, n585, n606);
or   g734 (n683, n579, n233, n578);
and  g735 (n750, n579, n272, n207);
nand g736 (n695, n246, n600, n324);
nand g737 (n718, n597, n325, n277);
and  g738 (n621, n326, n616, n613);
xor  g739 (n747, n205, n567);
nor  g740 (n809, n316, n593, n226);
xor  g741 (n804, n572, n584, n601);
nand g742 (n795, n311, n583, n573);
nand g743 (n783, n613, n299, n248);
xor  g744 (n632, n601, n580, n264);
or   g745 (n634, n580, n286, n581);
xor  g746 (n801, n236, n570, n610);
nor  g747 (n712, n338, n279, n327);
xor  g748 (n629, n575, n587, n283);
or   g749 (n618, n245, n615, n567);
xnor g750 (n749, n242, n574, n252);
or   g751 (n653, n196, n582, n218);
nor  g752 (n762, n596, n570, n610);
xor  g753 (n753, n320, n605, n594);
xor  g754 (n743, n285, n597, n189);
or   g755 (n620, n599, n344, n568);
xor  g756 (n670, n586, n568, n605);
or   g757 (n751, n576, n278, n288);
and  g758 (n668, n294, n606, n585);
nand g759 (n672, n267, n607, n194);
and  g760 (n800, n295, n583, n331);
or   g761 (n776, n270, n230, n580);
nor  g762 (n815, n310, n318, n329);
xnor g763 (n643, n273, n577, n228);
and  g764 (n626, n232, n268, n296);
nor  g765 (n748, n333, n195, n271);
xor  g766 (n692, n215, n282, n225);
or   g767 (n646, n615, n598, n336);
and  g768 (n686, n616, n600, n191);
xnor g769 (n746, n234, n220, n263);
or   g770 (n715, n597, n222, n611);
xor  g771 (n744, n281, n614, n588);
or   g772 (n760, n253, n223, n599);
nand g773 (n700, n219, n589, n247);
xnor g774 (n674, n579, n589);
nand g775 (n737, n608, n595, n240);
nor  g776 (n752, n591, n289, n582);
xnor g777 (n623, n581, n301, n292);
or   g778 (n655, n609, n611, n572);
and  g779 (n803, n577, n572, n217);
and  g780 (n789, n305, n571, n614);
and  g781 (n814, n607, n309, n204);
xnor g782 (n677, n583, n588, n573);
and  g783 (n657, n608, n588, n612);
xor  g784 (n761, n598, n597, n576);
nand g785 (n725, n192, n567, n571);
xnor g786 (n793, n602, n603, n251);
nor  g787 (n784, n581, n186, n328);
nand g788 (n722, n581, n343, n313);
xor  g789 (n685, n568, n608, n601);
not  g790 (n935, n803);
buf  g791 (n884, n675);
buf  g792 (n998, n641);
not  g793 (n1134, n639);
buf  g794 (n1013, n791);
not  g795 (n1109, n808);
buf  g796 (n888, n759);
buf  g797 (n1062, n701);
not  g798 (n1161, n660);
not  g799 (n864, n624);
buf  g800 (n945, n807);
buf  g801 (n1046, n711);
buf  g802 (n1123, n623);
not  g803 (n1101, n702);
not  g804 (n970, n643);
buf  g805 (n1120, n721);
buf  g806 (n1107, n802);
buf  g807 (n876, n751);
not  g808 (n978, n763);
not  g809 (n1130, n634);
not  g810 (n880, n746);
not  g811 (n841, n727);
buf  g812 (n933, n638);
buf  g813 (n829, n693);
buf  g814 (n883, n729);
buf  g815 (n1063, n689);
buf  g816 (n999, n814);
buf  g817 (n1100, n790);
buf  g818 (n1069, n695);
buf  g819 (n895, n807);
not  g820 (n1086, n633);
buf  g821 (n1111, n631);
not  g822 (n832, n733);
buf  g823 (n1164, n699);
buf  g824 (n1000, n702);
not  g825 (n937, n741);
not  g826 (n866, n650);
not  g827 (n827, n645);
not  g828 (n911, n782);
not  g829 (n863, n658);
buf  g830 (n1048, n664);
buf  g831 (n965, n751);
buf  g832 (n1117, n739);
buf  g833 (n969, n640);
buf  g834 (n1124, n730);
buf  g835 (n861, n797);
not  g836 (n1168, n796);
buf  g837 (n878, n654);
buf  g838 (n862, n812);
not  g839 (n1078, n678);
buf  g840 (n957, n806);
buf  g841 (n1053, n808);
not  g842 (n1042, n730);
buf  g843 (n1068, n775);
not  g844 (n1080, n717);
buf  g845 (n1035, n685);
not  g846 (n1110, n683);
buf  g847 (n1025, n793);
not  g848 (n1137, n639);
not  g849 (n1064, n803);
not  g850 (n981, n788);
not  g851 (n1088, n689);
buf  g852 (n817, n735);
not  g853 (n870, n799);
not  g854 (n1039, n642);
buf  g855 (n995, n809);
not  g856 (n1106, n790);
buf  g857 (n865, n723);
buf  g858 (n1031, n793);
not  g859 (n843, n685);
not  g860 (n1082, n714);
buf  g861 (n906, n770);
not  g862 (n826, n729);
buf  g863 (n979, n816);
buf  g864 (n991, n794);
not  g865 (n1043, n790);
not  g866 (n1138, n686);
not  g867 (n1136, n719);
buf  g868 (n1028, n764);
buf  g869 (n836, n747);
buf  g870 (n925, n802);
not  g871 (n1151, n810);
buf  g872 (n1067, n724);
buf  g873 (n1006, n750);
buf  g874 (n856, n763);
not  g875 (n894, n649);
not  g876 (n1044, n745);
buf  g877 (n875, n694);
not  g878 (n907, n804);
not  g879 (n931, n751);
buf  g880 (n901, n681);
not  g881 (n873, n752);
buf  g882 (n1163, n719);
not  g883 (n958, n646);
not  g884 (n1089, n779);
not  g885 (n1122, n713);
not  g886 (n913, n770);
not  g887 (n909, n653);
buf  g888 (n1125, n656);
not  g889 (n1114, n765);
not  g890 (n908, n797);
buf  g891 (n960, n697);
not  g892 (n927, n666);
not  g893 (n919, n764);
buf  g894 (n1146, n815);
not  g895 (n1020, n655);
buf  g896 (n990, n666);
buf  g897 (n834, n630);
buf  g898 (n1143, n755);
buf  g899 (n917, n705);
buf  g900 (n892, n655);
buf  g901 (n975, n628);
not  g902 (n890, n681);
not  g903 (n986, n779);
buf  g904 (n1133, n718);
not  g905 (n1083, n688);
not  g906 (n1152, n804);
buf  g907 (n882, n792);
buf  g908 (n855, n816);
not  g909 (n842, n733);
not  g910 (n854, n637);
not  g911 (n859, n351);
buf  g912 (n889, n703);
not  g913 (n1169, n661);
not  g914 (n902, n736);
buf  g915 (n887, n793);
buf  g916 (n947, n671);
not  g917 (n845, n674);
not  g918 (n1144, n662);
buf  g919 (n1149, n722);
buf  g920 (n974, n692);
buf  g921 (n1096, n756);
buf  g922 (n1011, n691);
buf  g923 (n1085, n750);
not  g924 (n967, n731);
buf  g925 (n1166, n716);
not  g926 (n1059, n790);
buf  g927 (n938, n664);
not  g928 (n1016, n745);
not  g929 (n953, n680);
not  g930 (n1103, n715);
buf  g931 (n1115, n795);
buf  g932 (n932, n755);
buf  g933 (n983, n786);
buf  g934 (n1099, n767);
buf  g935 (n1056, n803);
not  g936 (n1104, n792);
buf  g937 (n1036, n774);
not  g938 (n837, n795);
not  g939 (n982, n703);
not  g940 (n1112, n754);
not  g941 (n1172, n811);
not  g942 (n1081, n630);
buf  g943 (n1127, n768);
not  g944 (n985, n733);
not  g945 (n853, n649);
buf  g946 (n1065, n648);
buf  g947 (n939, n684);
not  g948 (n1105, n713);
buf  g949 (n920, n798);
buf  g950 (n858, n768);
not  g951 (n1019, n668);
buf  g952 (n1148, n743);
not  g953 (n1090, n676);
buf  g954 (n914, n691);
not  g955 (n1029, n696);
buf  g956 (n1070, n814);
not  g957 (n1008, n737);
buf  g958 (n954, n777);
not  g959 (n1154, n763);
buf  g960 (n848, n617);
buf  g961 (n897, n671);
not  g962 (n1034, n736);
not  g963 (n891, n622);
not  g964 (n1093, n707);
buf  g965 (n893, n811);
buf  g966 (n984, n747);
buf  g967 (n1098, n647);
not  g968 (n1041, n744);
buf  g969 (n852, n651);
not  g970 (n903, n703);
not  g971 (n846, n797);
buf  g972 (n1061, n794);
not  g973 (n851, n694);
not  g974 (n963, n737);
not  g975 (n1030, n794);
buf  g976 (n879, n784);
not  g977 (n1057, n733);
buf  g978 (n819, n810);
not  g979 (n899, n699);
buf  g980 (n1076, n805);
not  g981 (n1171, n695);
not  g982 (n849, n788);
buf  g983 (n835, n644);
not  g984 (n962, n669);
not  g985 (n996, n657);
not  g986 (n867, n688);
not  g987 (n988, n649);
not  g988 (n1040, n748);
buf  g989 (n1139, n686);
not  g990 (n934, n754);
not  g991 (n1058, n670);
buf  g992 (n833, n783);
not  g993 (n1026, n714);
buf  g994 (n926, n663);
not  g995 (n910, n761);
not  g996 (n921, n656);
buf  g997 (n993, n682);
buf  g998 (n1170, n654);
buf  g999 (n900, n628);
not  g1000 (n940, n709);
buf  g1001 (n1047, n757);
nand g1002 (n1119, n633, n654, n787, n680);
xor  g1003 (n928, n696, n734, n760, n661);
xnor g1004 (n912, n801, n693, n762, n772);
or   g1005 (n821, n750, n669, n639, n770);
and  g1006 (n818, n781, n797, n774, n696);
xor  g1007 (n942, n789, n796, n731, n721);
nor  g1008 (n952, n692, n660, n364, n678);
nor  g1009 (n944, n637, n767, n811, n659);
nand g1010 (n924, n666, n787, n639, n775);
or   g1011 (n822, n670, n709, n722, n360);
xnor g1012 (n1045, n734, n656, n792, n354);
xor  g1013 (n1017, n696, n730, n644, n811);
and  g1014 (n1049, n647, n780, n721, n655);
xnor g1015 (n1001, n648, n798, n646, n704);
xor  g1016 (n997, n669, n682, n782, n748);
nor  g1017 (n923, n349, n715, n648, n804);
xor  g1018 (n966, n648, n668, n688, n722);
or   g1019 (n930, n697, n725, n719, n708);
nand g1020 (n1052, n805, n693, n712, n357);
and  g1021 (n1077, n717, n778, n692, n798);
nor  g1022 (n918, n766, n747, n728, n716);
and  g1023 (n1074, n728, n676, n699, n672);
and  g1024 (n1003, n749, n709, n725, n798);
nor  g1025 (n824, n706, n743, n739, n774);
nor  g1026 (n1128, n684, n752, n748, n712);
nor  g1027 (n1066, n629, n682, n670, n642);
nand g1028 (n1012, n796, n786, n631, n654);
or   g1029 (n1097, n675, n638, n781, n767);
nor  g1030 (n987, n695, n807, n638, n640);
and  g1031 (n1005, n814, n743, n638, n716);
or   g1032 (n968, n755, n641, n642, n715);
nor  g1033 (n886, n634, n749, n361, n713);
nand g1034 (n1027, n665, n750, n663, n766);
nand g1035 (n959, n674, n632, n743, n718);
and  g1036 (n830, n641, n757, n684, n628);
xnor g1037 (n964, n774, n753, n808, n684);
nor  g1038 (n955, n792, n812, n742, n771);
xnor g1039 (n828, n629, n725, n791, n783);
nand g1040 (n820, n751, n765, n675, n737);
xnor g1041 (n869, n745, n712, n627, n731);
and  g1042 (n850, n668, n796, n665, n746);
and  g1043 (n973, n704, n761, n779, n672);
or   g1044 (n1158, n703, n809, n739, n744);
xnor g1045 (n874, n715, n763, n662, n780);
nand g1046 (n1094, n643, n806, n780, n726);
nand g1047 (n972, n769, n711, n681, n666);
xor  g1048 (n971, n730, n636, n689, n738);
xor  g1049 (n1073, n707, n352, n717, n619);
or   g1050 (n1167, n801, n732, n710, n740);
nor  g1051 (n857, n700, n685, n778, n785);
nor  g1052 (n1132, n672, n711, n800, n657);
nand g1053 (n976, n636, n627, n753, n754);
or   g1054 (n1022, n679, n356, n769, n710);
and  g1055 (n1118, n783, n772, n778, n660);
nor  g1056 (n1162, n658, n816, n624, n664);
nand g1057 (n885, n765, n642, n769, n620);
and  g1058 (n847, n630, n688, n772, n653);
xor  g1059 (n1150, n626, n674, n732, n676);
and  g1060 (n1014, n754, n784, n651, n671);
nor  g1061 (n1092, n815, n744, n738, n745);
and  g1062 (n989, n362, n744, n717, n801);
and  g1063 (n1007, n789, n711, n746, n706);
and  g1064 (n1004, n700, n705, n782, n718);
and  g1065 (n1024, n752, n749, n651, n673);
xnor g1066 (n1009, n667, n775, n724, n762);
xnor g1067 (n877, n659, n640, n813, n637);
or   g1068 (n1155, n813, n698, n707, n786);
xor  g1069 (n868, n720, n624, n813, n697);
or   g1070 (n936, n660, n777, n806, n625);
or   g1071 (n994, n740, n629, n726, n793);
nor  g1072 (n977, n677, n810, n766, n679);
and  g1073 (n961, n726, n727, n771, n758);
nand g1074 (n980, n698, n634, n695, n770);
nor  g1075 (n1054, n803, n678, n732, n767);
xnor g1076 (n838, n640, n800, n700);
nor  g1077 (n949, n749, n759, n635);
and  g1078 (n1165, n674, n724, n657, n644);
xor  g1079 (n1126, n671, n759, n773, n736);
nor  g1080 (n916, n776, n633, n742, n701);
nor  g1081 (n1021, n773, n809, n687, n784);
or   g1082 (n1091, n635, n768, n658, n800);
xnor g1083 (n881, n704, n665, n788, n669);
nor  g1084 (n1051, n761, n804, n662, n659);
nor  g1085 (n1129, n718, n729, n690, n665);
xnor g1086 (n1050, n734, n704, n649, n791);
nand g1087 (n1159, n692, n701, n740, n813);
nand g1088 (n1157, n773, n721, n739, n787);
xnor g1089 (n839, n714, n728, n779, n756);
xor  g1090 (n1087, n650, n653, n771, n673);
nor  g1091 (n1147, n709, n723, n714, n753);
and  g1092 (n956, n651, n794, n636, n652);
or   g1093 (n1071, n689, n748, n355, n643);
nor  g1094 (n823, n756, n708, n764, n702);
xnor g1095 (n1135, n683, n780, n645, n686);
nor  g1096 (n860, n661, n816, n784, n752);
or   g1097 (n896, n728, n720, n687, n760);
or   g1098 (n1113, n809, n675, n656, n716);
nor  g1099 (n1102, n634, n777, n667, n753);
nand g1100 (n1037, n741, n762, n623, n740);
or   g1101 (n943, n782, n713, n802, n734);
xor  g1102 (n946, n727, n636, n707, n677);
nand g1103 (n840, n359, n678, n781, n812);
and  g1104 (n1131, n758, n668, n621, n736);
and  g1105 (n950, n677, n647, n758, n637);
nand g1106 (n1075, n732, n663, n775, n785);
nand g1107 (n1145, n679, n787, n738, n801);
or   g1108 (n1002, n737, n690, n757, n742);
xnor g1109 (n1095, n706, n653, n677, n663);
and  g1110 (n1140, n720, n723, n694, n699);
or   g1111 (n1023, n756, n785, n633, n710);
and  g1112 (n1141, n776, n667, n682, n686);
xnor g1113 (n1079, n363, n710, n766, n789);
xor  g1114 (n1018, n701, n776, n799, n781);
xor  g1115 (n1033, n746, n685, n741, n795);
and  g1116 (n1060, n708, n760, n627, n631);
xnor g1117 (n1116, n805, n643, n764, n652);
nand g1118 (n905, n723, n778, n658, n719);
xor  g1119 (n941, n690, n741, n765, n657);
or   g1120 (n1153, n762, n768, n673, n350);
xnor g1121 (n1121, n706, n805, n650, n799);
nor  g1122 (n1142, n814, n738, n755, n687);
xor  g1123 (n1015, n812, n769, n626, n786);
xor  g1124 (n844, n724, n772, n691, n698);
xor  g1125 (n825, n676, n680, n747, n806);
xor  g1126 (n831, n712, n662, n641, n694);
or   g1127 (n929, n726, n625, n785, n661);
nand g1128 (n871, n646, n720, n802, n679);
and  g1129 (n904, n771, n650, n697, n729);
nor  g1130 (n872, n683, n810, n632, n655);
nor  g1131 (n1010, n700, n731, n791, n758);
and  g1132 (n898, n789, n815, n795, n647);
nand g1133 (n992, n652, n708, n808, n644);
xnor g1134 (n915, n799, n646, n632, n777);
nor  g1135 (n1038, n760, n645, n358, n776);
nor  g1136 (n1160, n664, n698, n652, n687);
and  g1137 (n1156, n673, n702, n735);
nand g1138 (n922, n690, n815, n618, n788);
nor  g1139 (n1084, n807, n622, n705, n626);
xnor g1140 (n1055, n625, n645, n691, n759);
xnor g1141 (n1032, n672, n693, n722, n725);
xor  g1142 (n1072, n680, n635, n705, n761);
and  g1143 (n1108, n670, n683, n773, n742);
nor  g1144 (n948, n667, n783, n757, n735);
nand g1145 (n951, n727, n681, n659, n353);
not  g1146 (n1187, n817);
buf  g1147 (n1179, n828);
not  g1148 (n1176, n832);
not  g1149 (n1183, n829);
buf  g1150 (n1178, n826);
buf  g1151 (n1182, n830);
not  g1152 (n1177, n822);
not  g1153 (n1173, n831);
not  g1154 (n1185, n818);
not  g1155 (n1174, n823);
not  g1156 (n1186, n825);
not  g1157 (n1181, n819);
buf  g1158 (n1188, n820);
buf  g1159 (n1180, n827);
not  g1160 (n1184, n824);
not  g1161 (n1175, n821);
xnor g1162 (n1189, n1178, n1177, n1174, n1179);
xnor g1163 (n1190, n833, n1176, n1173, n1175);
buf  g1164 (n1191, n1190);
not  g1165 (n1192, n1180);
xor  g1166 (n1193, n1190, n1189);
not  g1167 (n1200, n846);
not  g1168 (n1195, n1191);
nor  g1169 (n1202, n371, n1193);
or   g1170 (n1201, n839, n367, n844, n847);
xnor g1171 (n1198, n838, n1192, n850);
nor  g1172 (n1197, n1191, n372, n1193, n840);
or   g1173 (n1199, n1181, n852, n843, n834);
or   g1174 (n1203, n1191, n368, n849, n365);
nor  g1175 (n1204, n845, n841, n837, n851);
xor  g1176 (n1196, n1191, n848, n836, n366);
xnor g1177 (n1194, n1192, n370, n842, n1193);
xnor g1178 (n1205, n835, n1192, n369, n1193);
nand g1179 (n1238, n413, n452, n436, n458);
or   g1180 (n1207, n394, n1199, n462, n473);
xnor g1181 (n1214, n423, n446, n1203, n380);
xnor g1182 (n1228, n442, n1205, n414, n392);
xor  g1183 (n1225, n1204, n476, n454, n417);
nand g1184 (n1222, n374, n467, n1195, n404);
xnor g1185 (n1218, n441, n477, n464, n1198);
and  g1186 (n1209, n449, n408, n470, n438);
xor  g1187 (n1206, n450, n475, n424, n466);
or   g1188 (n1239, n384, n402, n1202, n1204);
nand g1189 (n1236, n1201, n1200, n463, n397);
and  g1190 (n1230, n1197, n431, n382, n399);
xor  g1191 (n1220, n1199, n412, n383, n474);
xor  g1192 (n1229, n439, n444, n409, n1204);
and  g1193 (n1221, n451, n426, n447, n1203);
xnor g1194 (n1232, n387, n403, n1203, n448);
and  g1195 (n1235, n386, n1202, n1200, n440);
xor  g1196 (n1219, n1198, n427, n395, n1196);
nand g1197 (n1240, n381, n1197, n419, n1201);
xnor g1198 (n1210, n422, n469, n472, n391);
and  g1199 (n1226, n1194, n420, n407, n456);
or   g1200 (n1213, n421, n375, n400, n1205);
nand g1201 (n1223, n429, n418, n411, n459);
xor  g1202 (n1208, n455, n457, n432, n388);
nand g1203 (n1212, n435, n1205, n1201, n377);
and  g1204 (n1233, n1200, n1196, n471, n1204);
nor  g1205 (n1211, n390, n430, n1205, n406);
and  g1206 (n1231, n389, n1203, n443, n428);
or   g1207 (n1215, n385, n468, n1195, n410);
and  g1208 (n1224, n378, n437, n434, n396);
and  g1209 (n1227, n379, n433, n398, n465);
or   g1210 (n1216, n416, n1202, n376, n425);
nand g1211 (n1217, n393, n415, n1201, n461);
nor  g1212 (n1234, n373, n453, n1202, n1200);
xor  g1213 (n1237, n401, n460, n445, n405);
xnor g1214 (n1247, n1206, n1233, n1229, n1219);
nor  g1215 (n1241, n1218, n1212, n1234, n1223);
nand g1216 (n1242, n1234, n1210, n1232, n1228);
and  g1217 (n1245, n1214, n1230, n1225, n1227);
xor  g1218 (n1250, n1229, n1231, n1208);
nor  g1219 (n1246, n1220, n1232, n1221, n1217);
xnor g1220 (n1249, n1216, n1213, n1230, n1224);
xor  g1221 (n1243, n1235, n1211, n1215, n1228);
xor  g1222 (n1248, n1226, n1222, n1227, n1209);
xnor g1223 (n1244, n1226, n1233, n1235, n1207);
buf  g1224 (n1254, n854);
not  g1225 (n1253, n1244);
buf  g1226 (n1257, n1250);
buf  g1227 (n1255, n860);
not  g1228 (n1259, n1246);
buf  g1229 (n1256, n1243);
or   g1230 (n1251, n856, n1242, n1249, n1245);
or   g1231 (n1258, n853, n858, n859, n857);
xnor g1232 (n1252, n1248, n861, n855, n1247);
buf  g1233 (n1260, n1251);
buf  g1234 (n1261, n1251);
buf  g1235 (n1263, n1252);
buf  g1236 (n1262, n1251);
nand g1237 (n1270, n1252, n870, n1260, n865);
and  g1238 (n1265, n1253, n1253, n863, n1261);
xnor g1239 (n1268, n864, n478, n1254, n873);
xor  g1240 (n1266, n866, n868, n871, n1252);
nor  g1241 (n1264, n867, n1261, n1263, n1262);
nand g1242 (n1269, n1253, n1253, n1252, n869);
nor  g1243 (n1267, n1262, n872, n1263, n862);
buf  g1244 (n1274, n1265);
not  g1245 (n1273, n1264);
buf  g1246 (n1272, n1265);
buf  g1247 (n1271, n1264);
buf  g1248 (n1277, n880);
not  g1249 (n1276, n877);
buf  g1250 (n1278, n1273);
not  g1251 (n1282, n1272);
buf  g1252 (n1280, n1274);
or   g1253 (n1281, n879, n878, n1274);
xnor g1254 (n1275, n876, n874, n881, n1272);
xor  g1255 (n1279, n1273, n1271, n875);
nor  g1256 (n1296, n506, n487, n502, n481);
nand g1257 (n1283, n505, n1237, n508, n884);
xnor g1258 (n1289, n888, n1282, n482, n890);
or   g1259 (n1288, n490, n483, n1182, n495);
xnor g1260 (n1295, n503, n491, n498, n497);
nor  g1261 (n1300, n882, n1276, n1184, n1282);
and  g1262 (n1287, n1282, n496, n1281);
nand g1263 (n1285, n1188, n504, n886, n480);
xor  g1264 (n1292, n509, n510, n1278, n494);
or   g1265 (n1291, n885, n484, n1277, n501);
and  g1266 (n1293, n1279, n889, n1275, n1237);
nand g1267 (n1298, n887, n489, n1276, n492);
nand g1268 (n1284, n1183, n1275, n486, n500);
xor  g1269 (n1297, n485, n883, n479, n1278);
xor  g1270 (n1290, n1187, n1279, n507, n1277);
and  g1271 (n1299, n488, n1281, n499, n1186);
and  g1272 (n1286, n1280, n511, n493, n1236);
or   g1273 (n1294, n1280, n1280, n1185, n1236);
nand g1274 (n1310, n894, n534, n517, n515);
xor  g1275 (n1307, n1291, n1283, n1284, n891);
or   g1276 (n1308, n535, n536, n520, n530);
xnor g1277 (n1311, n519, n533, n526, n1256);
nand g1278 (n1306, n537, n1255, n516, n1292);
nand g1279 (n1316, n1296, n1255, n529, n1300);
and  g1280 (n1301, n538, n521, n892, n1299);
or   g1281 (n1305, n895, n522, n527, n1294);
and  g1282 (n1315, n1256, n1290, n1255, n1254);
xnor g1283 (n1304, n524, n525, n1254, n1298);
or   g1284 (n1303, n1286, n1287, n539, n528);
nand g1285 (n1309, n1256, n1285, n1288, n513);
nand g1286 (n1313, n1295, n531, n532, n523);
nor  g1287 (n1302, n1254, n897, n514, n1289);
xnor g1288 (n1314, n518, n896, n512, n898);
xnor g1289 (n1312, n1297, n893, n1293, n1255);
buf  g1290 (n1317, n1313);
not  g1291 (n1319, n900);
buf  g1292 (n1323, n903);
not  g1293 (n1320, n901);
not  g1294 (n1322, n1309);
xnor g1295 (n1324, n1310, n906, n905);
nand g1296 (n1318, n1316, n904, n1314, n899);
or   g1297 (n1321, n1311, n1312, n902, n1315);
not  g1298 (n1326, n1319);
buf  g1299 (n1327, n1318);
buf  g1300 (n1333, n1318);
buf  g1301 (n1329, n1320);
buf  g1302 (n1330, n1319);
buf  g1303 (n1335, n1317);
buf  g1304 (n1331, n1320);
not  g1305 (n1332, n1320);
not  g1306 (n1325, n1317);
xor  g1307 (n1328, n1320, n1318, n1319);
nor  g1308 (n1334, n1318, n1317, n1319);
xor  g1309 (n1344, n1332, n949, n944, n918);
or   g1310 (n1342, n917, n914, n921, n1327);
nor  g1311 (n1348, n1335, n1334, n951, n942);
nor  g1312 (n1338, n919, n1326, n911, n945);
xor  g1313 (n1351, n912, n952, n933, n943);
nand g1314 (n1350, n1331, n910, n927, n1334);
xor  g1315 (n1336, n950, n940, n928, n931);
xor  g1316 (n1340, n926, n1328, n908, n953);
and  g1317 (n1343, n924, n920, n938, n909);
nor  g1318 (n1349, n1325, n941, n1335, n937);
nor  g1319 (n1337, n916, n1335, n925, n1330);
xnor g1320 (n1339, n932, n934, n1329, n929);
xnor g1321 (n1346, n913, n939, n923, n1333);
or   g1322 (n1341, n947, n948, n954, n946);
xnor g1323 (n1347, n936, n915, n930, n1335);
xor  g1324 (n1345, n907, n1334, n935, n922);
or   g1325 (n1354, n970, n987, n964, n1348);
xor  g1326 (n1364, n1347, n1344, n961, n963);
nand g1327 (n1369, n991, n1347, n997, n990);
xnor g1328 (n1355, n1343, n1336, n1346, n979);
nor  g1329 (n1368, n992, n1345, n1337, n1341);
or   g1330 (n1366, n966, n975, n1344, n962);
xor  g1331 (n1353, n960, n984, n1346, n1343);
or   g1332 (n1367, n973, n1346, n1343, n996);
xnor g1333 (n1359, n980, n968, n1338, n981);
nand g1334 (n1363, n985, n994, n974, n965);
nand g1335 (n1362, n1342, n959, n1340, n1345);
xor  g1336 (n1361, n1344, n969, n978, n982);
nor  g1337 (n1360, n1341, n956, n998, n1342);
or   g1338 (n1358, n971, n989, n957, n1336);
and  g1339 (n1352, n993, n1345, n976, n986);
xor  g1340 (n1357, n972, n1348, n1337, n983);
xor  g1341 (n1370, n955, n1339, n1338, n988);
nand g1342 (n1365, n958, n1340, n995, n1342);
xor  g1343 (n1356, n1339, n967, n1347, n977);
or   g1344 (n1371, n1004, n1002, n1020, n1018);
xnor g1345 (n1374, n1013, n1367, n1000, n1369);
xor  g1346 (n1373, n1019, n1001, n1007, n1024);
nor  g1347 (n1376, n1022, n1005, n1009, n1015);
or   g1348 (n1375, n1014, n1366, n1370, n999);
and  g1349 (n1378, n1025, n1016, n1012, n1368);
nor  g1350 (n1372, n1362, n1023, n1011, n1003);
nor  g1351 (n1379, n1008, n1006, n1017, n1010);
and  g1352 (n1377, n1021, n1365, n1363, n1364);
xor  g1353 (n1396, n1053, n1068, n1103, n545);
or   g1354 (n1384, n1076, n1376, n1106, n1099);
nand g1355 (n1407, n1039, n1052, n1051, n1377);
xnor g1356 (n1403, n1082, n1038, n1373, n1379);
xor  g1357 (n1398, n1375, n1372, n1058, n1121);
xnor g1358 (n1409, n1120, n1060, n1266, n1037);
and  g1359 (n1386, n1054, n1044, n1375, n541);
xnor g1360 (n1395, n1100, n1371, n1108, n1116);
or   g1361 (n1402, n1034, n543, n1036, n1029);
nand g1362 (n1388, n1073, n1374, n1069);
nor  g1363 (n1408, n1096, n1372, n1041, n1378);
nand g1364 (n1412, n1375, n1055, n1118, n544);
nor  g1365 (n1414, n1374, n1373, n1045, n1091);
nand g1366 (n1411, n1088, n1090, n1085, n1061);
xnor g1367 (n1400, n1372, n546, n1105, n1028);
and  g1368 (n1410, n1084, n1075, n1070, n1378);
or   g1369 (n1392, n542, n1114, n1374, n1040);
nand g1370 (n1380, n1077, n1094, n1074, n1062);
xor  g1371 (n1391, n1050, n1373, n1372, n1072);
xnor g1372 (n1393, n1035, n1092, n1379, n1048);
or   g1373 (n1413, n1046, n1102, n1087, n1376);
or   g1374 (n1389, n1371, n540, n1111, n1375);
xnor g1375 (n1387, n1049, n1078, n1379, n1080);
or   g1376 (n1405, n1026, n1110, n1115, n1030);
nor  g1377 (n1397, n1378, n1047, n1064, n1377);
or   g1378 (n1394, n1081, n1376, n1043, n1104);
nor  g1379 (n1390, n1378, n1071, n1033, n1095);
nor  g1380 (n1401, n1379, n1032, n1119, n1059);
xor  g1381 (n1381, n1113, n1373, n1098, n1086);
xnor g1382 (n1406, n1027, n1097, n1067, n1109);
nand g1383 (n1399, n1063, n1089, n1056, n1065);
nand g1384 (n1383, n1101, n1107, n1079, n1117);
xor  g1385 (n1385, n1112, n1266, n1376, n1031);
nor  g1386 (n1382, n1093, n1377, n1042, n1066);
or   g1387 (n1404, n1377, n1057, n1371, n1083);
xor  g1388 (n1418, n1411, n1413, n1387, n1400);
or   g1389 (n1419, n1383, n1409, n1391, n1408);
nand g1390 (n1426, n1406, n1397, n1268, n1414);
and  g1391 (n1427, n1380, n1122, n1399, n1269);
or   g1392 (n1424, n1410, n1395, n1381, n1398);
and  g1393 (n1422, n1268, n1396, n1125, n1128);
nand g1394 (n1423, n1126, n1267, n1384);
nor  g1395 (n1417, n1393, n1270, n1124, n1403);
or   g1396 (n1420, n1412, n1269, n1385, n1386);
nor  g1397 (n1415, n1129, n1392, n1390, n1402);
nand g1398 (n1421, n1401, n1270, n1394, n1127);
nor  g1399 (n1416, n1270, n1407, n1388, n1382);
xor  g1400 (n1425, n1389, n1404, n1405, n1123);
nand g1401 (n1434, n1150, n1424, n1132, n1418);
nand g1402 (n1440, n1142, n1133, n1151, n1427);
nand g1403 (n1439, n1168, n1165, n1426, n1140);
nor  g1404 (n1436, n1167, n1131, n1154, n1415);
and  g1405 (n1435, n1157, n1161, n1158, n1425);
or   g1406 (n1441, n1416, n1171, n1419, n1135);
and  g1407 (n1437, n1170, n1417, n1420, n1166);
xor  g1408 (n1431, n1160, n1145, n1134, n1169);
xor  g1409 (n1432, n1423, n1144, n1427, n1159);
xnor g1410 (n1428, n1422, n1152, n1141, n1421);
xor  g1411 (n1433, n1137, n1162, n1163, n1139);
or   g1412 (n1429, n1136, n1138, n1147, n1146);
and  g1413 (n1430, n1156, n1155, n1164, n1148);
and  g1414 (n1438, n1153, n1149, n1130, n1143);
nand g1415 (n1449, n1239, n1257, n1322);
nand g1416 (n1454, n1350, n1323, n1349, n1429);
or   g1417 (n1446, n1438, n1322, n1351, n1324);
xnor g1418 (n1443, n1433, n1349, n1322, n1441);
nor  g1419 (n1445, n1257, n1240, n1258, n1440);
nor  g1420 (n1447, n1351, n1323, n1348, n1259);
nand g1421 (n1455, n1239, n1259, n1321, n1350);
and  g1422 (n1451, n1321, n1258, n1257);
xor  g1423 (n1456, n1350, n1435, n1259, n1172);
nand g1424 (n1448, n1436, n1434, n1321);
or   g1425 (n1457, n1238, n1324, n1240);
nand g1426 (n1442, n1259, n1323, n1258, n1441);
nand g1427 (n1444, n1431, n1437, n1351, n1349);
or   g1428 (n1452, n1256, n1432, n1240, n1323);
or   g1429 (n1450, n1430, n1238, n1428, n1324);
xnor g1430 (n1453, n1440, n1240, n1258, n1439);
nand g1431 (n1458, n1455, n1447, n1454, n1456);
and  g1432 (n1459, n1446, n1451, n1452, n1449);
or   g1433 (n1460, n1453, n1450, n1445, n1443);
xnor g1434 (n1461, n1442, n1448, n1457, n1444);
xor  g1435 (n1462, n1458, n1460, n1459, n1461);
endmodule
