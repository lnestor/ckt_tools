

module Stat_100_53
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n100,
  n93,
  n80,
  n114,
  n99,
  n110,
  n107,
  n92,
  n84,
  n86,
  n79,
  n115,
  n91,
  n95,
  n88,
  n112,
  n117,
  n89,
  n132,
  n129,
  n120,
  n124,
  n128,
  n127,
  n125,
  n123,
  n119,
  n126,
  n122,
  n121,
  n131,
  n130,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n100;
  output n93;
  output n80;
  output n114;
  output n99;
  output n110;
  output n107;
  output n92;
  output n84;
  output n86;
  output n79;
  output n115;
  output n91;
  output n95;
  output n88;
  output n112;
  output n117;
  output n89;
  output n132;
  output n129;
  output n120;
  output n124;
  output n128;
  output n127;
  output n125;
  output n123;
  output n119;
  output n126;
  output n122;
  output n121;
  output n131;
  output n130;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n81;
  wire n82;
  wire n83;
  wire n85;
  wire n87;
  wire n90;
  wire n94;
  wire n96;
  wire n97;
  wire n98;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n108;
  wire n109;
  wire n111;
  wire n113;
  wire n116;
  wire n118;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyNOTWire_0_4;
  wire KeyWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyNOTWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyWire_0_51;
  wire KeyNOTWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyNOTWire_0_54;
  wire KeyWire_0_55;
  wire KeyNOTWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n41,
    n2
  );


  buf
  g1
  (
    KeyWire_0_42,
    n2
  );


  not
  g2
  (
    KeyWire_0_36,
    n1
  );


  buf
  g3
  (
    KeyWire_0_15,
    n1
  );


  buf
  g4
  (
    KeyWire_0_47,
    n2
  );


  buf
  g5
  (
    KeyWire_0_26,
    n3
  );


  not
  g6
  (
    n42,
    n1
  );


  not
  g7
  (
    KeyWire_0_25,
    n2
  );


  buf
  g8
  (
    n40,
    n3
  );


  not
  g9
  (
    KeyWire_0_28,
    n1
  );


  not
  g10
  (
    KeyWire_0_60,
    n33
  );


  not
  g11
  (
    KeyWire_0_17,
    n34
  );


  buf
  g12
  (
    KeyWire_0_11,
    n34
  );


  buf
  g13
  (
    n46,
    n33
  );


  buf
  g14
  (
    KeyWire_0_23,
    n33
  );


  buf
  g15
  (
    KeyWire_0_56,
    n34
  );


  buf
  g16
  (
    n43,
    n34
  );


  buf
  g17
  (
    n44,
    n33
  );


  buf
  g18
  (
    KeyWire_0_5,
    n45
  );


  buf
  g19
  (
    KeyWire_0_18,
    n49
  );


  buf
  g20
  (
    KeyWire_0_3,
    n43
  );


  buf
  g21
  (
    n51,
    n44
  );


  buf
  g22
  (
    n52,
    n46
  );


  buf
  g23
  (
    KeyWire_0_19,
    n48
  );


  not
  g24
  (
    KeyWire_0_44,
    n44
  );


  buf
  g25
  (
    KeyWire_0_38,
    n35
  );


  not
  g26
  (
    KeyWire_0_43,
    n47
  );


  buf
  g27
  (
    KeyWire_0_7,
    n44
  );


  not
  g28
  (
    KeyWire_0_39,
    n45
  );


  buf
  g29
  (
    KeyWire_0_31,
    n47
  );


  xor
  g30
  (
    KeyWire_0_35,
    n44,
    n48
  );


  nor
  g31
  (
    KeyWire_0_2,
    n46,
    n47
  );


  or
  g32
  (
    KeyWire_0_13,
    n35,
    n35,
    n43,
    n48
  );


  nand
  g33
  (
    n62,
    n47,
    n45,
    n35,
    n46
  );


  nor
  g34
  (
    KeyWire_0_63,
    n43,
    n43,
    n48,
    n49
  );


  xor
  g35
  (
    n60,
    n46,
    n36,
    n45
  );


  xor
  g36
  (
    KeyWire_0_58,
    n62,
    n6
  );


  and
  g37
  (
    n94,
    n64,
    n29,
    n3,
    n32
  );


  nand
  g38
  (
    KeyWire_0_51,
    n20,
    n67,
    n12,
    n32
  );


  xnor
  g39
  (
    KeyWire_0_61,
    n67,
    n11,
    n30,
    n7
  );


  nor
  g40
  (
    n80,
    n15,
    n51,
    n29,
    n8
  );


  xnor
  g41
  (
    n91,
    n17,
    n61,
    n4
  );


  or
  g42
  (
    n72,
    n51,
    n49,
    n18,
    n50
  );


  xor
  g43
  (
    KeyWire_0_53,
    n56,
    n54,
    n27,
    n14
  );


  or
  g44
  (
    KeyWire_0_57,
    n16,
    n36,
    n60,
    n15
  );


  nor
  g45
  (
    KeyWire_0_27,
    n59,
    n10,
    n54,
    n12
  );


  nor
  g46
  (
    KeyWire_0_55,
    n67,
    n50,
    n15,
    n55
  );


  xnor
  g47
  (
    KeyWire_0_50,
    n26,
    n16,
    n27,
    n20
  );


  and
  g48
  (
    n107,
    n25,
    n64,
    n24,
    n58
  );


  or
  g49
  (
    n110,
    n63,
    n9,
    n22,
    n68
  );


  or
  g50
  (
    n99,
    n50,
    n6,
    n51,
    n8
  );


  xnor
  g51
  (
    n118,
    n68,
    n16,
    n14,
    n11
  );


  xor
  g52
  (
    KeyWire_0_40,
    n10,
    n5,
    n66,
    n28
  );


  xnor
  g53
  (
    KeyWire_0_8,
    n13,
    n57,
    n32,
    n7
  );


  nor
  g54
  (
    n84,
    n10,
    n23,
    n63,
    n58
  );


  and
  g55
  (
    n77,
    n13,
    n64,
    n14,
    n62
  );


  nor
  g56
  (
    KeyWire_0_24,
    n22,
    n24,
    n57,
    n66
  );


  or
  g57
  (
    KeyWire_0_1,
    n23,
    n8,
    n18,
    n59
  );


  xnor
  g58
  (
    KeyWire_0_21,
    n60,
    n64,
    n9,
    n4
  );


  nor
  g59
  (
    KeyWire_0_9,
    n65,
    n26,
    n66,
    n21
  );


  and
  g60
  (
    n112,
    n25,
    n55,
    n59,
    n23
  );


  xnor
  g61
  (
    KeyWire_0_37,
    n36,
    n49,
    n63,
    n8
  );


  xor
  g62
  (
    n88,
    n57,
    n12,
    n62,
    n18
  );


  and
  g63
  (
    n115,
    n52,
    n60,
    n25
  );


  xnor
  g64
  (
    n85,
    n18,
    n21,
    n50,
    n5
  );


  xnor
  g65
  (
    KeyWire_0_46,
    n25,
    n7,
    n13,
    n26
  );


  or
  g66
  (
    KeyWire_0_12,
    n61,
    n21,
    n27,
    n52
  );


  and
  g67
  (
    KeyWire_0_22,
    n61,
    n55,
    n4,
    n30
  );


  nor
  g68
  (
    KeyWire_0_14,
    n23,
    n59,
    n30
  );


  xor
  g69
  (
    KeyWire_0_52,
    n53,
    n62,
    n29,
    n10
  );


  and
  g70
  (
    KeyWire_0_54,
    n21,
    n4,
    n58,
    n13
  );


  xnor
  g71
  (
    KeyWire_0_62,
    n54,
    n56,
    n31,
    n65
  );


  or
  g72
  (
    n103,
    n52,
    n31,
    n54,
    n9
  );


  xor
  g73
  (
    KeyWire_0_0,
    n22,
    n6,
    n67,
    n17
  );


  and
  g74
  (
    n73,
    n20,
    n15,
    n11,
    n19
  );


  or
  g75
  (
    KeyWire_0_48,
    n65,
    n28,
    n5,
    n14
  );


  or
  g76
  (
    n114,
    n29,
    n31,
    n26,
    n68
  );


  and
  g77
  (
    KeyWire_0_49,
    n17,
    n19,
    n58
  );


  nand
  g78
  (
    KeyWire_0_30,
    n55,
    n5,
    n11,
    n53
  );


  or
  g79
  (
    KeyWire_0_32,
    n17,
    n63,
    n22,
    n9
  );


  xnor
  g80
  (
    KeyWire_0_20,
    n56,
    n27,
    n28,
    n66
  );


  or
  g81
  (
    n106,
    n56,
    n3,
    n53,
    n65
  );


  nor
  g82
  (
    n87,
    n32,
    n53,
    n68,
    n24
  );


  nor
  g83
  (
    KeyWire_0_10,
    n57,
    n24,
    n31,
    n52
  );


  or
  g84
  (
    KeyWire_0_29,
    n20,
    n7,
    n19,
    n6
  );


  nand
  g85
  (
    KeyWire_0_6,
    n16,
    n51,
    n12,
    n28
  );


  nor
  g86
  (
    KeyWire_0_41,
    n102,
    n41,
    n42
  );


  and
  g87
  (
    n127,
    n40,
    n106,
    n110,
    n88
  );


  nor
  g88
  (
    KeyWire_0_34,
    n91,
    n38,
    n101,
    n117
  );


  xor
  g89
  (
    KeyWire_0_16,
    n94,
    n90,
    n92,
    n111
  );


  nand
  g90
  (
    n132,
    n98,
    n118,
    n37,
    n113
  );


  xor
  g91
  (
    KeyWire_0_4,
    n95,
    n38,
    n87,
    n89
  );


  nor
  g92
  (
    KeyWire_0_45,
    n93,
    n41,
    n42
  );


  and
  g93
  (
    n126,
    n103,
    n97,
    n38,
    n37
  );


  and
  g94
  (
    n128,
    n40,
    n37,
    n38,
    n115
  );


  xor
  g95
  (
    n131,
    n40,
    n41,
    n104,
    n109
  );


  xor
  g96
  (
    KeyWire_0_59,
    n105,
    n41,
    n116,
    n114
  );


  and
  g97
  (
    n123,
    n39,
    n39,
    n107,
    n99
  );


  nor
  g98
  (
    KeyWire_0_33,
    n112,
    n37,
    n108,
    n39
  );


  and
  g99
  (
    n130,
    n40,
    n39,
    n96,
    n100
  );


  xor
  KeyGate_0_0
  (
    n76,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n71,
    KeyNOTWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n54,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n61,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n120,
    KeyNOTWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n57,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n81,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n58,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n82,
    keyIn_0_8,
    KeyWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n69,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n78,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n48,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n79,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n59,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n74,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n37,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n119,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n47,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n67,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n55,
    KeyNOTWire_0_19
  );


  xor
  KeyGate_0_20
  (
    n100,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n105,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n96,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n45,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    KeyNOTWire_0_24,
    keyIn_0_24,
    KeyWire_0_24
  );


  not
  KeyNOTGate_0_24
  (
    n93,
    KeyNOTWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n38,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n34,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    n113,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n33,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n90,
    KeyNOTWire_0_29
  );


  xor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n104,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n63,
    keyIn_0_31,
    KeyWire_0_31
  );


  xnor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n75,
    KeyNOTWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n122,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n124,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n66,
    keyIn_0_35,
    KeyWire_0_35
  );


  xnor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n35,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n98,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    n65,
    keyIn_0_38,
    KeyWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n56,
    keyIn_0_39,
    KeyWire_0_39
  );


  xor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n108,
    KeyNOTWire_0_40
  );


  xor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n129,
    KeyNOTWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n36,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n64,
    KeyNOTWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    n53,
    keyIn_0_44,
    KeyWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n125,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    n102,
    keyIn_0_46,
    KeyWire_0_46
  );


  xor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n39,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    n117,
    keyIn_0_48,
    KeyWire_0_48
  );


  xor
  KeyGate_0_49
  (
    n83,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    n95,
    keyIn_0_50,
    KeyWire_0_50
  );


  xor
  KeyGate_0_51
  (
    KeyNOTWire_0_51,
    keyIn_0_51,
    KeyWire_0_51
  );


  not
  KeyNOTGate_0_51
  (
    n70,
    KeyNOTWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n111,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n89,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    KeyNOTWire_0_54,
    keyIn_0_54,
    KeyWire_0_54
  );


  not
  KeyNOTGate_0_54
  (
    n101,
    KeyNOTWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    KeyNOTWire_0_55,
    keyIn_0_55,
    KeyWire_0_55
  );


  not
  KeyNOTGate_0_55
  (
    n116,
    KeyNOTWire_0_55
  );


  xor
  KeyGate_0_56
  (
    n49,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    n109,
    keyIn_0_57,
    KeyWire_0_57
  );


  xor
  KeyGate_0_58
  (
    n92,
    keyIn_0_58,
    KeyWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n121,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n50,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    n97,
    keyIn_0_61,
    KeyWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n86,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n68,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

