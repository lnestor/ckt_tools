

module Stat_377_1329
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n402,
  n405,
  n395,
  n392,
  n390,
  n397,
  n400,
  n393,
  n403,
  n399,
  n404,
  n401,
  n396,
  n391,
  n389,
  n398,
  n394
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n402;output n405;output n395;output n392;output n390;output n397;output n400;output n393;output n403;output n399;output n404;output n401;output n396;output n391;output n389;output n398;output n394;
  wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n102,
    n6
  );


  not
  g1
  (
    n88,
    n3
  );


  buf
  g2
  (
    n75,
    n12
  );


  not
  g3
  (
    n92,
    n15
  );


  buf
  g4
  (
    n85,
    n4
  );


  not
  g5
  (
    n47,
    n13
  );


  not
  g6
  (
    n90,
    n20
  );


  buf
  g7
  (
    n56,
    n9
  );


  buf
  g8
  (
    n77,
    n18
  );


  buf
  g9
  (
    n95,
    n8
  );


  buf
  g10
  (
    n65,
    n8
  );


  not
  g11
  (
    n29,
    n15
  );


  buf
  g12
  (
    n33,
    n3
  );


  not
  g13
  (
    n37,
    n12
  );


  buf
  g14
  (
    n101,
    n13
  );


  buf
  g15
  (
    n35,
    n2
  );


  buf
  g16
  (
    n32,
    n1
  );


  not
  g17
  (
    n70,
    n18
  );


  not
  g18
  (
    n103,
    n2
  );


  not
  g19
  (
    n96,
    n6
  );


  buf
  g20
  (
    n66,
    n7
  );


  not
  g21
  (
    n60,
    n17
  );


  buf
  g22
  (
    n43,
    n12
  );


  not
  g23
  (
    n64,
    n6
  );


  buf
  g24
  (
    n30,
    n17
  );


  not
  g25
  (
    n54,
    n2
  );


  not
  g26
  (
    n41,
    n13
  );


  buf
  g27
  (
    KeyWire_0_15,
    n8
  );


  not
  g28
  (
    n57,
    n17
  );


  not
  g29
  (
    KeyWire_0_2,
    n11
  );


  not
  g30
  (
    n80,
    n4
  );


  not
  g31
  (
    n104,
    n16
  );


  buf
  g32
  (
    n34,
    n7
  );


  not
  g33
  (
    n46,
    n9
  );


  buf
  g34
  (
    n51,
    n14
  );


  buf
  g35
  (
    n106,
    n10
  );


  not
  g36
  (
    n69,
    n11
  );


  buf
  g37
  (
    n44,
    n19
  );


  not
  g38
  (
    n84,
    n15
  );


  buf
  g39
  (
    n94,
    n19
  );


  buf
  g40
  (
    n72,
    n5
  );


  buf
  g41
  (
    n83,
    n15
  );


  not
  g42
  (
    n53,
    n9
  );


  not
  g43
  (
    n79,
    n17
  );


  buf
  g44
  (
    n38,
    n1
  );


  buf
  g45
  (
    n31,
    n5
  );


  buf
  g46
  (
    n55,
    n20
  );


  not
  g47
  (
    n93,
    n7
  );


  buf
  g48
  (
    n39,
    n11
  );


  buf
  g49
  (
    KeyWire_0_31,
    n5
  );


  not
  g50
  (
    n48,
    n4
  );


  buf
  g51
  (
    KeyWire_0_4,
    n8
  );


  not
  g52
  (
    n86,
    n12
  );


  not
  g53
  (
    n52,
    n10
  );


  not
  g54
  (
    n74,
    n13
  );


  not
  g55
  (
    n100,
    n11
  );


  not
  g56
  (
    n61,
    n14
  );


  not
  g57
  (
    n42,
    n18
  );


  not
  g58
  (
    n68,
    n10
  );


  not
  g59
  (
    n82,
    n6
  );


  not
  g60
  (
    n58,
    n14
  );


  not
  g61
  (
    n97,
    n1
  );


  not
  g62
  (
    n67,
    n18
  );


  buf
  g63
  (
    n49,
    n7
  );


  buf
  g64
  (
    n59,
    n16
  );


  not
  g65
  (
    n63,
    n9
  );


  buf
  g66
  (
    n40,
    n19
  );


  buf
  g67
  (
    KeyWire_0_26,
    n2
  );


  buf
  g68
  (
    n81,
    n14
  );


  not
  g69
  (
    n78,
    n10
  );


  buf
  g70
  (
    n87,
    n1
  );


  not
  g71
  (
    n76,
    n16
  );


  not
  g72
  (
    n71,
    n4
  );


  not
  g73
  (
    n36,
    n3
  );


  not
  g74
  (
    n73,
    n3
  );


  buf
  g75
  (
    n45,
    n5
  );


  not
  g76
  (
    n105,
    n19
  );


  buf
  g77
  (
    n98,
    n16
  );


  not
  g78
  (
    n113,
    n37
  );


  buf
  g79
  (
    n117,
    n39
  );


  buf
  g80
  (
    n118,
    n44
  );


  not
  g81
  (
    n110,
    n35
  );


  not
  g82
  (
    n114,
    n43
  );


  buf
  g83
  (
    n116,
    n32
  );


  buf
  g84
  (
    n120,
    n30
  );


  buf
  g85
  (
    KeyWire_0_12,
    n33
  );


  buf
  g86
  (
    n112,
    n36
  );


  buf
  g87
  (
    n121,
    n40
  );


  not
  g88
  (
    n119,
    n31
  );


  buf
  g89
  (
    n111,
    n38
  );


  not
  g90
  (
    KeyWire_0_9,
    n29
  );


  buf
  g91
  (
    n108,
    n45
  );


  not
  g92
  (
    n122,
    n41
  );


  buf
  g93
  (
    n107,
    n42
  );


  not
  g94
  (
    n109,
    n34
  );


  and
  g95
  (
    n124,
    n56,
    n63,
    n58,
    n48
  );


  or
  g96
  (
    n131,
    n112,
    n61,
    n47,
    n59
  );


  nand
  g97
  (
    n127,
    n51,
    n65,
    n62,
    n64
  );


  xnor
  g98
  (
    n130,
    n64,
    n108,
    n109,
    n50
  );


  xnor
  g99
  (
    n126,
    n54,
    n107,
    n49,
    n52
  );


  or
  g100
  (
    KeyWire_0_30,
    n66,
    n65,
    n55,
    n113
  );


  nor
  g101
  (
    KeyWire_0_20,
    n53,
    n46,
    n66,
    n57
  );


  or
  g102
  (
    n129,
    n114,
    n60,
    n110,
    n111
  );


  xnor
  g103
  (
    KeyWire_0_21,
    n68,
    n83,
    n128,
    n79
  );


  nand
  g104
  (
    n137,
    n75,
    n129,
    n81
  );


  xnor
  g105
  (
    n134,
    n90,
    n68,
    n127,
    n87
  );


  nor
  g106
  (
    n139,
    n89,
    n74,
    n82
  );


  and
  g107
  (
    n146,
    n78,
    n74,
    n131,
    n72
  );


  and
  g108
  (
    n135,
    n129,
    n76,
    n124,
    n72
  );


  nand
  g109
  (
    n140,
    n75,
    n87,
    n90,
    n67
  );


  nand
  g110
  (
    KeyWire_0_23,
    n85,
    n80,
    n88
  );


  and
  g111
  (
    n138,
    n76,
    n89,
    n73,
    n84
  );


  nand
  g112
  (
    n136,
    n125,
    n79,
    n78,
    n69
  );


  xor
  g113
  (
    n141,
    n73,
    n86,
    n127
  );


  xor
  g114
  (
    n143,
    n128,
    n70,
    n84
  );


  nand
  g115
  (
    n144,
    n71,
    n125,
    n77,
    n130
  );


  xnor
  g116
  (
    n145,
    n69,
    n124,
    n131,
    n85
  );


  nand
  g117
  (
    n132,
    n77,
    n67,
    n83,
    n126
  );


  and
  g118
  (
    n147,
    n130,
    n71,
    n126,
    n88
  );


  buf
  g119
  (
    n154,
    n20
  );


  buf
  g120
  (
    n150,
    n91
  );


  not
  g121
  (
    n157,
    n140
  );


  buf
  g122
  (
    n156,
    n20
  );


  buf
  g123
  (
    n149,
    n134
  );


  not
  g124
  (
    n153,
    n92
  );


  nor
  g125
  (
    n155,
    n135,
    n21,
    n94,
    n91
  );


  nor
  g126
  (
    n148,
    n93,
    n139,
    n92,
    n133
  );


  xnor
  g127
  (
    n152,
    n94,
    n132,
    n138,
    n93
  );


  nand
  g128
  (
    n151,
    n141,
    n137,
    n21,
    n136
  );


  buf
  g129
  (
    n167,
    n149
  );


  xnor
  g130
  (
    n170,
    n98,
    n99,
    n100,
    n96
  );


  or
  g131
  (
    n160,
    n97,
    n102,
    n98,
    n95
  );


  nand
  g132
  (
    KeyWire_0_16,
    n151,
    n103,
    n148
  );


  xor
  g133
  (
    n161,
    n149,
    n148,
    n97
  );


  nor
  g134
  (
    n159,
    n149,
    n97,
    n98,
    n150
  );


  nor
  g135
  (
    n164,
    n100,
    n150,
    n96,
    n103
  );


  and
  g136
  (
    n168,
    n99,
    n102,
    n151
  );


  nand
  g137
  (
    n169,
    n101,
    n151,
    n95,
    n99
  );


  nor
  g138
  (
    n166,
    n100,
    n149,
    n101,
    n96
  );


  xnor
  g139
  (
    n162,
    n95,
    n98,
    n150,
    n101
  );


  or
  g140
  (
    n163,
    n150,
    n100,
    n102,
    n96
  );


  xor
  g141
  (
    n158,
    n103,
    n101,
    n99,
    n95
  );


  not
  g142
  (
    n215,
    n170
  );


  not
  g143
  (
    n173,
    n156
  );


  buf
  g144
  (
    n174,
    n144
  );


  buf
  g145
  (
    n199,
    n146
  );


  not
  g146
  (
    n209,
    n163
  );


  buf
  g147
  (
    KeyWire_0_13,
    n155
  );


  not
  g148
  (
    n202,
    n162
  );


  not
  g149
  (
    n197,
    n166
  );


  not
  g150
  (
    n210,
    n159
  );


  not
  g151
  (
    n212,
    n119
  );


  buf
  g152
  (
    n213,
    n165
  );


  not
  g153
  (
    n205,
    n163
  );


  buf
  g154
  (
    n189,
    n160
  );


  buf
  g155
  (
    n187,
    n147
  );


  not
  g156
  (
    n176,
    n154
  );


  not
  g157
  (
    n185,
    n152
  );


  not
  g158
  (
    n192,
    n161
  );


  buf
  g159
  (
    n177,
    n163
  );


  not
  g160
  (
    n195,
    n167
  );


  not
  g161
  (
    KeyWire_0_29,
    n163
  );


  buf
  g162
  (
    n188,
    n151
  );


  not
  g163
  (
    n203,
    n161
  );


  buf
  g164
  (
    n219,
    n120
  );


  buf
  g165
  (
    n214,
    n152
  );


  buf
  g166
  (
    n186,
    n146
  );


  buf
  g167
  (
    n183,
    n156
  );


  not
  g168
  (
    n196,
    n160
  );


  not
  g169
  (
    n184,
    n145
  );


  buf
  g170
  (
    n182,
    n153
  );


  buf
  g171
  (
    KeyWire_0_8,
    n170
  );


  buf
  g172
  (
    n171,
    n169
  );


  not
  g173
  (
    KeyWire_0_6,
    n165
  );


  not
  g174
  (
    n216,
    n170
  );


  and
  g175
  (
    n200,
    n162,
    n166,
    n121
  );


  xnor
  g176
  (
    n208,
    n152,
    n162,
    n117,
    n146
  );


  xnor
  g177
  (
    n175,
    n147,
    n158,
    n152,
    n165
  );


  xor
  g178
  (
    n206,
    n155,
    n154,
    n167,
    n153
  );


  nor
  g179
  (
    n201,
    n155,
    n147,
    n168,
    n165
  );


  and
  g180
  (
    KeyWire_0_3,
    n166,
    n161,
    n146,
    n168
  );


  nor
  g181
  (
    n218,
    n116,
    n155,
    n153,
    n159
  );


  and
  g182
  (
    n191,
    n147,
    n157,
    n164,
    n166
  );


  or
  g183
  (
    n204,
    n167,
    n170,
    n161,
    n168
  );


  nor
  g184
  (
    n217,
    n157,
    n167,
    n115,
    n169
  );


  and
  g185
  (
    n207,
    n162,
    n169,
    n156,
    n131
  );


  nor
  g186
  (
    n194,
    n122,
    n157,
    n164,
    n154
  );


  or
  g187
  (
    n181,
    n142,
    n143,
    n154,
    n160
  );


  xor
  g188
  (
    n193,
    n157,
    n159,
    n164
  );


  and
  g189
  (
    KeyWire_0_22,
    n118,
    n159,
    n123,
    n169
  );


  xor
  g190
  (
    n180,
    n153,
    n160,
    n156,
    n168
  );


  not
  g191
  (
    n225,
    n175
  );


  buf
  g192
  (
    n228,
    n172
  );


  buf
  g193
  (
    KeyWire_0_0,
    n171
  );


  not
  g194
  (
    n230,
    n172
  );


  not
  g195
  (
    n227,
    n174
  );


  buf
  g196
  (
    n223,
    n174
  );


  buf
  g197
  (
    n235,
    n172
  );


  not
  g198
  (
    n221,
    n173
  );


  buf
  g199
  (
    n224,
    n173
  );


  not
  g200
  (
    n234,
    n171
  );


  buf
  g201
  (
    n232,
    n175
  );


  buf
  g202
  (
    n233,
    n174
  );


  buf
  g203
  (
    n222,
    n173
  );


  not
  g204
  (
    n231,
    n172
  );


  not
  g205
  (
    n237,
    n171
  );


  not
  g206
  (
    n220,
    n174
  );


  not
  g207
  (
    n226,
    n173
  );


  buf
  g208
  (
    n236,
    n171
  );


  xnor
  g209
  (
    n283,
    n206,
    n214,
    n226
  );


  xnor
  g210
  (
    KeyWire_0_19,
    n231,
    n196,
    n209
  );


  nor
  g211
  (
    n245,
    n25,
    n223,
    n234
  );


  or
  g212
  (
    n291,
    n212,
    n232,
    n236
  );


  and
  g213
  (
    n309,
    n235,
    n225,
    n183
  );


  nor
  g214
  (
    n242,
    n210,
    n28,
    n225
  );


  xnor
  g215
  (
    n300,
    n227,
    n191,
    n177
  );


  xor
  g216
  (
    n238,
    n223,
    n207,
    n200
  );


  and
  g217
  (
    KeyWire_0_7,
    n222,
    n176,
    n180
  );


  and
  g218
  (
    n290,
    n183,
    n201,
    n203
  );


  or
  g219
  (
    n241,
    n188,
    n190,
    n224
  );


  and
  g220
  (
    n307,
    n193,
    n188,
    n201
  );


  or
  g221
  (
    n284,
    n202,
    n177,
    n206
  );


  nand
  g222
  (
    n302,
    n224,
    n186,
    n237
  );


  nand
  g223
  (
    n270,
    n222,
    n184,
    n205,
    n194
  );


  or
  g224
  (
    n294,
    n229,
    n224,
    n220,
    n184
  );


  xor
  g225
  (
    n240,
    n184,
    n194,
    n197,
    n198
  );


  nor
  g226
  (
    n275,
    n231,
    n207,
    n183,
    n27
  );


  and
  g227
  (
    KeyWire_0_28,
    n184,
    n186,
    n196,
    n200
  );


  xnor
  g228
  (
    n239,
    n228,
    n225,
    n208,
    n209
  );


  nand
  g229
  (
    n263,
    n199,
    n221,
    n104,
    n209
  );


  nor
  g230
  (
    n258,
    n22,
    n21,
    n214,
    n199
  );


  xor
  g231
  (
    n260,
    n211,
    n178,
    n175,
    n234
  );


  or
  g232
  (
    n286,
    n188,
    n191,
    n204,
    n203
  );


  nor
  g233
  (
    n255,
    n203,
    n195,
    n193,
    n182
  );


  xor
  g234
  (
    n277,
    n181,
    n105,
    n234,
    n24
  );


  xor
  g235
  (
    n282,
    n105,
    n202,
    n180,
    n187
  );


  nand
  g236
  (
    n293,
    n211,
    n21,
    n192,
    n179
  );


  xor
  g237
  (
    n268,
    n213,
    n197,
    n235,
    n178
  );


  nor
  g238
  (
    n256,
    n209,
    n179,
    n195,
    n24
  );


  nand
  g239
  (
    n251,
    n198,
    n236,
    n212,
    n186
  );


  xor
  g240
  (
    n295,
    n207,
    n224,
    n23,
    n205
  );


  xor
  g241
  (
    n303,
    n28,
    n189,
    n232,
    n195
  );


  or
  g242
  (
    n274,
    n231,
    n208,
    n199,
    n28
  );


  xor
  g243
  (
    n244,
    n226,
    n208,
    n220,
    n178
  );


  nor
  g244
  (
    n281,
    n28,
    n179,
    n26,
    n197
  );


  xnor
  g245
  (
    n287,
    n213,
    n205,
    n189,
    n227
  );


  xor
  g246
  (
    n247,
    n223,
    n189,
    n205,
    n193
  );


  and
  g247
  (
    n269,
    n25,
    n24,
    n176,
    n180
  );


  nand
  g248
  (
    n253,
    n177,
    n22,
    n27,
    n181
  );


  nand
  g249
  (
    n248,
    n236,
    n104,
    n106,
    n176
  );


  nand
  g250
  (
    n257,
    n23,
    n215,
    n106,
    n229
  );


  nand
  g251
  (
    n265,
    n214,
    n237,
    n190,
    n26
  );


  and
  g252
  (
    n304,
    n233,
    n230,
    n194,
    n177
  );


  and
  g253
  (
    n261,
    n222,
    n202,
    n227,
    n231
  );


  and
  g254
  (
    n301,
    n180,
    n182,
    n196,
    n185
  );


  or
  g255
  (
    n264,
    n212,
    n178,
    n214,
    n22
  );


  nand
  g256
  (
    n250,
    n226,
    n233,
    n221
  );


  xnor
  g257
  (
    n273,
    n187,
    n228,
    n192,
    n229
  );


  xor
  g258
  (
    n298,
    n195,
    n189,
    n191,
    n235
  );


  nor
  g259
  (
    n267,
    n105,
    n228,
    n192,
    n210
  );


  nor
  g260
  (
    n297,
    n215,
    n24,
    n23,
    n106
  );


  and
  g261
  (
    n285,
    n194,
    n204,
    n232,
    n213
  );


  nand
  g262
  (
    n254,
    n192,
    n186,
    n206,
    n183
  );


  and
  g263
  (
    n246,
    n208,
    n181,
    n237,
    n221
  );


  and
  g264
  (
    KeyWire_0_14,
    n200,
    n237,
    n210,
    n220
  );


  nor
  g265
  (
    n279,
    n26,
    n210,
    n106,
    n212
  );


  xnor
  g266
  (
    n299,
    n200,
    n187,
    n26,
    n229
  );


  or
  g267
  (
    KeyWire_0_25,
    n23,
    n190,
    n207,
    n211
  );


  nor
  g268
  (
    n243,
    n193,
    n196,
    n211,
    n197
  );


  nand
  g269
  (
    n292,
    n228,
    n230,
    n181,
    n199
  );


  or
  g270
  (
    n276,
    n188,
    n27,
    n182
  );


  nor
  g271
  (
    n272,
    n203,
    n198,
    n226,
    n175
  );


  or
  g272
  (
    n288,
    n104,
    n201,
    n182,
    n206
  );


  xnor
  g273
  (
    n308,
    n191,
    n185,
    n221,
    n236
  );


  and
  g274
  (
    n262,
    n227,
    n105,
    n185,
    n190
  );


  xor
  g275
  (
    n259,
    n223,
    n230,
    n201,
    n233
  );


  nor
  g276
  (
    KeyWire_0_24,
    n25,
    n187,
    n222,
    n220
  );


  xnor
  g277
  (
    n296,
    n204,
    n176,
    n185,
    n179
  );


  nor
  g278
  (
    KeyWire_0_10,
    n225,
    n202,
    n230,
    n213
  );


  nand
  g279
  (
    n252,
    n198,
    n204,
    n25,
    n232
  );


  nor
  g280
  (
    n266,
    n235,
    n234,
    n22,
    n104
  );


  buf
  g281
  (
    n312,
    n239
  );


  not
  g282
  (
    n315,
    n238
  );


  buf
  g283
  (
    n313,
    n241
  );


  not
  g284
  (
    n311,
    n240
  );


  not
  g285
  (
    n314,
    n240
  );


  not
  g286
  (
    n310,
    n239
  );


  buf
  g287
  (
    n330,
    n248
  );


  buf
  g288
  (
    n331,
    n314
  );


  not
  g289
  (
    n325,
    n249
  );


  not
  g290
  (
    n321,
    n245
  );


  buf
  g291
  (
    n322,
    n243
  );


  buf
  g292
  (
    n316,
    n241
  );


  not
  g293
  (
    KeyWire_0_27,
    n247
  );


  buf
  g294
  (
    n328,
    n246
  );


  buf
  g295
  (
    n323,
    n244
  );


  xor
  g296
  (
    n326,
    n311,
    n250,
    n314
  );


  or
  g297
  (
    n329,
    n245,
    n251,
    n315,
    n312
  );


  nand
  g298
  (
    n327,
    n313,
    n242,
    n312
  );


  xor
  g299
  (
    n320,
    n247,
    n314,
    n315,
    n246
  );


  nand
  g300
  (
    n318,
    n244,
    n252,
    n313,
    n315
  );


  or
  g301
  (
    n332,
    n251,
    n250,
    n243,
    n242
  );


  or
  g302
  (
    n319,
    n314,
    n252,
    n313
  );


  xnor
  g303
  (
    n324,
    n312,
    n249,
    n248,
    n310
  );


  buf
  g304
  (
    n358,
    n282
  );


  not
  g305
  (
    n383,
    n293
  );


  not
  g306
  (
    n372,
    n289
  );


  nand
  g307
  (
    n385,
    n320,
    n259,
    n301,
    n292
  );


  xor
  g308
  (
    n360,
    n253,
    n284,
    n290,
    n282
  );


  or
  g309
  (
    n371,
    n257,
    n260,
    n295,
    n323
  );


  xnor
  g310
  (
    n357,
    n307,
    n299,
    n261,
    n303
  );


  xor
  g311
  (
    n381,
    n273,
    n257,
    n321,
    n265
  );


  nor
  g312
  (
    n380,
    n306,
    n295,
    n327,
    n309
  );


  nand
  g313
  (
    n343,
    n297,
    n280,
    n283
  );


  xnor
  g314
  (
    n349,
    n284,
    n308,
    n320,
    n303
  );


  nor
  g315
  (
    n373,
    n256,
    n272,
    n277,
    n309
  );


  and
  g316
  (
    n366,
    n266,
    n216,
    n323,
    n299
  );


  nor
  g317
  (
    n353,
    n300,
    n302,
    n217
  );


  nand
  g318
  (
    n375,
    n321,
    n306,
    n288,
    n305
  );


  xor
  g319
  (
    n374,
    n218,
    n318,
    n316,
    n300
  );


  xor
  g320
  (
    KeyWire_0_11,
    n218,
    n308,
    n219,
    n307
  );


  xnor
  g321
  (
    n370,
    n304,
    n269,
    n328,
    n216
  );


  or
  g322
  (
    n336,
    n323,
    n259,
    n262,
    n298
  );


  xor
  g323
  (
    n369,
    n305,
    n319,
    n329,
    n318
  );


  or
  g324
  (
    n362,
    n215,
    n319,
    n218,
    n287
  );


  xnor
  g325
  (
    n363,
    n291,
    n326,
    n278,
    n286
  );


  nand
  g326
  (
    n348,
    n306,
    n286,
    n267,
    n327
  );


  or
  g327
  (
    n342,
    n319,
    n325,
    n264
  );


  and
  g328
  (
    n350,
    n268,
    n318,
    n258,
    n299
  );


  and
  g329
  (
    n345,
    n279,
    n328,
    n219,
    n278
  );


  xnor
  g330
  (
    KeyWire_0_18,
    n276,
    n326,
    n325,
    n316
  );


  or
  g331
  (
    n347,
    n270,
    n300,
    n216,
    n298
  );


  nand
  g332
  (
    n387,
    n256,
    n215,
    n262,
    n289
  );


  xnor
  g333
  (
    n355,
    n261,
    n309,
    n303,
    n324
  );


  nand
  g334
  (
    n367,
    n321,
    n302,
    n254,
    n258
  );


  nor
  g335
  (
    n378,
    n301,
    n292,
    n304
  );


  or
  g336
  (
    n338,
    n273,
    n301,
    n328,
    n290
  );


  nand
  g337
  (
    n354,
    n307,
    n263,
    n293,
    n317
  );


  nand
  g338
  (
    n368,
    n327,
    n265,
    n302,
    n255
  );


  xor
  g339
  (
    n341,
    n219,
    n321,
    n324
  );


  and
  g340
  (
    n346,
    n285,
    n275,
    n320,
    n329
  );


  nand
  g341
  (
    n340,
    n322,
    n277,
    n316,
    n255
  );


  xor
  g342
  (
    n344,
    n325,
    n322,
    n253,
    n216
  );


  nor
  g343
  (
    n359,
    n298,
    n264,
    n274,
    n287
  );


  or
  g344
  (
    n333,
    n298,
    n303,
    n322,
    n327
  );


  and
  g345
  (
    n351,
    n296,
    n302,
    n299,
    n322
  );


  and
  g346
  (
    n379,
    n275,
    n276,
    n305,
    n324
  );


  xnor
  g347
  (
    n364,
    n297,
    n304,
    n294,
    n326
  );


  nand
  g348
  (
    n377,
    n300,
    n294,
    n320,
    n297
  );


  xor
  g349
  (
    n384,
    n308,
    n317,
    n296,
    n272
  );


  and
  g350
  (
    n388,
    n271,
    n266,
    n217,
    n269
  );


  nand
  g351
  (
    n386,
    n318,
    n297,
    n285,
    n319
  );


  xor
  g352
  (
    KeyWire_0_17,
    n328,
    n329,
    n288,
    n305
  );


  or
  g353
  (
    n365,
    n274,
    n268,
    n308,
    n317
  );


  and
  g354
  (
    KeyWire_0_5,
    n281,
    n279,
    n329,
    n263
  );


  xnor
  g355
  (
    n382,
    n326,
    n217,
    n218,
    n301
  );


  nand
  g356
  (
    n335,
    n307,
    n254,
    n323,
    n306
  );


  and
  g357
  (
    n356,
    n267,
    n260,
    n280,
    n291
  );


  xnor
  g358
  (
    n352,
    n281,
    n219,
    n315,
    n316
  );


  xnor
  g359
  (
    n376,
    n270,
    n309,
    n271,
    n317
  );


  nor
  g360
  (
    n393,
    n330,
    n346,
    n336,
    n376
  );


  or
  g361
  (
    n395,
    n373,
    n361,
    n332,
    n383
  );


  xor
  g362
  (
    n402,
    n368,
    n358,
    n348,
    n333
  );


  nor
  g363
  (
    KeyWire_0_1,
    n357,
    n371,
    n331,
    n365
  );


  xor
  g364
  (
    n405,
    n362,
    n387,
    n382,
    n388
  );


  nor
  g365
  (
    n391,
    n334,
    n332,
    n374
  );


  nand
  g366
  (
    n398,
    n330,
    n344,
    n375,
    n352
  );


  xnor
  g367
  (
    n389,
    n370,
    n341,
    n386,
    n343
  );


  or
  g368
  (
    n397,
    n332,
    n372,
    n331,
    n342
  );


  nor
  g369
  (
    n392,
    n359,
    n331,
    n355,
    n337
  );


  or
  g370
  (
    n400,
    n377,
    n384,
    n353,
    n380
  );


  nand
  g371
  (
    n396,
    n331,
    n350,
    n335,
    n345
  );


  nor
  g372
  (
    n390,
    n360,
    n356,
    n330,
    n369
  );


  nand
  g373
  (
    n399,
    n364,
    n379,
    n381,
    n347
  );


  nand
  g374
  (
    n403,
    n378,
    n363,
    n366,
    n351
  );


  xor
  g375
  (
    n394,
    n354,
    n385,
    n330,
    n367
  );


  or
  g376
  (
    n404,
    n339,
    n338,
    n349,
    n340
  );


  xnor
  KeyGate_0_0
  (
    n229,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n401,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n89,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n178,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n99,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n337,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n190,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n289,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    n198,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n123,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n249,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n361,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n115,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n211,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n271,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n62,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    n165,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n339,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n334,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n278,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n125,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n142,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n172,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    n133,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n306,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n305,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n91,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n317,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n280,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n179,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n128,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n50,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


