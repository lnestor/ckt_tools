

module Stat_221_421
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n231,
  n212,
  n208,
  n238,
  n207,
  n226,
  n218,
  n214,
  n220,
  n227,
  n234,
  n235,
  n228,
  n222,
  n223,
  n209,
  n230,
  n224,
  n221,
  n210,
  n233,
  n216,
  n219,
  n237,
  n236,
  n232,
  n217,
  n213,
  n229,
  n215,
  n211,
  n225,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n231;
  output n212;
  output n208;
  output n238;
  output n207;
  output n226;
  output n218;
  output n214;
  output n220;
  output n227;
  output n234;
  output n235;
  output n228;
  output n222;
  output n223;
  output n209;
  output n230;
  output n224;
  output n221;
  output n210;
  output n233;
  output n216;
  output n219;
  output n237;
  output n236;
  output n232;
  output n217;
  output n213;
  output n229;
  output n215;
  output n211;
  output n225;
  wire n18;
  wire n19;
  wire n20;
  wire n21;
  wire n22;
  wire n23;
  wire n24;
  wire n25;
  wire n26;
  wire n27;
  wire n28;
  wire n29;
  wire n30;
  wire n31;
  wire n32;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyWire_0_12;
  wire KeyWire_0_13;
  wire KeyNOTWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyNOTWire_0_16;
  wire KeyWire_0_17;
  wire KeyNOTWire_0_17;
  wire KeyWire_0_18;
  wire KeyWire_0_19;
  wire KeyNOTWire_0_19;
  wire KeyWire_0_20;
  wire KeyNOTWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyNOTWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyNOTWire_0_32;
  wire KeyWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyNOTWire_0_36;
  wire KeyWire_0_37;
  wire KeyNOTWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyNOTWire_0_39;
  wire KeyWire_0_40;
  wire KeyNOTWire_0_40;
  wire KeyWire_0_41;
  wire KeyNOTWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyNOTWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyNOTWire_0_45;
  wire KeyWire_0_46;
  wire KeyWire_0_47;
  wire KeyWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyWire_0_57;
  wire KeyNOTWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyNOTWire_0_62;
  wire KeyWire_0_63;

  not
  g0
  (
    n28,
    n2
  );


  buf
  g1
  (
    n18,
    n3
  );


  not
  g2
  (
    n26,
    n3
  );


  not
  g3
  (
    KeyWire_0_44,
    n1
  );


  buf
  g4
  (
    n22,
    n5
  );


  buf
  g5
  (
    n30,
    n1
  );


  buf
  g6
  (
    n23,
    n3
  );


  not
  g7
  (
    KeyWire_0_13,
    n5
  );


  buf
  g8
  (
    n19,
    n2
  );


  not
  g9
  (
    KeyWire_0_57,
    n5
  );


  not
  g10
  (
    n20,
    n1
  );


  buf
  g11
  (
    KeyWire_0_48,
    n4
  );


  buf
  g12
  (
    KeyWire_0_56,
    n2
  );


  buf
  g13
  (
    n27,
    n4
  );


  not
  g14
  (
    n24,
    n4
  );


  buf
  g15
  (
    n78,
    n23
  );


  not
  g16
  (
    n58,
    n21
  );


  not
  g17
  (
    KeyWire_0_54,
    n22
  );


  not
  g18
  (
    KeyWire_0_62,
    n32
  );


  not
  g19
  (
    KeyWire_0_41,
    n22
  );


  buf
  g20
  (
    KeyWire_0_21,
    n24
  );


  buf
  g21
  (
    n48,
    n21
  );


  buf
  g22
  (
    n61,
    n20
  );


  not
  g23
  (
    n67,
    n26
  );


  not
  g24
  (
    n65,
    n18
  );


  not
  g25
  (
    n52,
    n30
  );


  buf
  g26
  (
    KeyWire_0_61,
    n32
  );


  not
  g27
  (
    n73,
    n28
  );


  not
  g28
  (
    n40,
    n31
  );


  not
  g29
  (
    n50,
    n20
  );


  buf
  g30
  (
    n43,
    n23
  );


  not
  g31
  (
    n44,
    n19
  );


  not
  g32
  (
    n34,
    n18
  );


  buf
  g33
  (
    KeyWire_0_63,
    n29
  );


  buf
  g34
  (
    KeyWire_0_22,
    n25
  );


  not
  g35
  (
    n74,
    n28
  );


  not
  g36
  (
    KeyWire_0_49,
    n18
  );


  not
  g37
  (
    n41,
    n27
  );


  not
  g38
  (
    n47,
    n29
  );


  not
  g39
  (
    KeyWire_0_16,
    n24
  );


  buf
  g40
  (
    n55,
    n30
  );


  not
  g41
  (
    n68,
    n22
  );


  buf
  g42
  (
    n38,
    n20
  );


  buf
  g43
  (
    n64,
    n28
  );


  buf
  g44
  (
    n72,
    n24
  );


  not
  g45
  (
    KeyWire_0_8,
    n27
  );


  buf
  g46
  (
    n39,
    n26
  );


  buf
  g47
  (
    KeyWire_0_2,
    n19
  );


  buf
  g48
  (
    n54,
    n30
  );


  not
  g49
  (
    n63,
    n26
  );


  not
  g50
  (
    n45,
    n21
  );


  buf
  g51
  (
    n60,
    n27
  );


  buf
  g52
  (
    n75,
    n32
  );


  buf
  g53
  (
    n36,
    n19
  );


  buf
  g54
  (
    n71,
    n25
  );


  buf
  g55
  (
    n77,
    n31
  );


  buf
  g56
  (
    KeyWire_0_27,
    n23
  );


  not
  g57
  (
    n66,
    n32
  );


  not
  g58
  (
    n46,
    n29
  );


  not
  g59
  (
    n76,
    n31
  );


  buf
  g60
  (
    KeyWire_0_15,
    n25
  );


  buf
  g61
  (
    n174,
    n33
  );


  buf
  g62
  (
    KeyWire_0_59,
    n60
  );


  not
  g63
  (
    n94,
    n45
  );


  buf
  g64
  (
    n181,
    n77
  );


  buf
  g65
  (
    KeyWire_0_9,
    n48
  );


  not
  g66
  (
    KeyWire_0_53,
    n52
  );


  not
  g67
  (
    n201,
    n9
  );


  buf
  g68
  (
    n143,
    n76
  );


  not
  g69
  (
    n91,
    n71
  );


  buf
  g70
  (
    n165,
    n34
  );


  buf
  g71
  (
    n99,
    n35
  );


  not
  g72
  (
    KeyWire_0_50,
    n65
  );


  not
  g73
  (
    n106,
    n77
  );


  not
  g74
  (
    n98,
    n57
  );


  buf
  g75
  (
    KeyWire_0_39,
    n53
  );


  buf
  g76
  (
    n178,
    n75
  );


  not
  g77
  (
    n108,
    n17
  );


  not
  g78
  (
    n141,
    n59
  );


  buf
  g79
  (
    n150,
    n45
  );


  not
  g80
  (
    n124,
    n41
  );


  buf
  g81
  (
    KeyWire_0_46,
    n77
  );


  not
  g82
  (
    n128,
    n69
  );


  not
  g83
  (
    n196,
    n39
  );


  not
  g84
  (
    n102,
    n67
  );


  buf
  g85
  (
    n156,
    n46
  );


  buf
  g86
  (
    n139,
    n41
  );


  buf
  g87
  (
    KeyWire_0_37,
    n78
  );


  buf
  g88
  (
    n132,
    n47
  );


  not
  g89
  (
    n127,
    n50
  );


  not
  g90
  (
    KeyWire_0_31,
    n61
  );


  buf
  g91
  (
    n197,
    n60
  );


  buf
  g92
  (
    KeyWire_0_51,
    n69
  );


  not
  g93
  (
    KeyWire_0_10,
    n78
  );


  buf
  g94
  (
    n80,
    n65
  );


  buf
  g95
  (
    n125,
    n38
  );


  not
  g96
  (
    n182,
    n14
  );


  buf
  g97
  (
    n81,
    n41
  );


  buf
  g98
  (
    KeyWire_0_5,
    n7
  );


  buf
  g99
  (
    KeyWire_0_28,
    n66
  );


  not
  g100
  (
    n160,
    n14
  );


  buf
  g101
  (
    n87,
    n65
  );


  buf
  g102
  (
    n118,
    n55
  );


  buf
  g103
  (
    n138,
    n36
  );


  not
  g104
  (
    n170,
    n8
  );


  not
  g105
  (
    n154,
    n72
  );


  not
  g106
  (
    n188,
    n70
  );


  not
  g107
  (
    n145,
    n54
  );


  buf
  g108
  (
    KeyWire_0_23,
    n44
  );


  not
  g109
  (
    n130,
    n76
  );


  buf
  g110
  (
    n206,
    n73
  );


  buf
  g111
  (
    n149,
    n52
  );


  buf
  g112
  (
    n90,
    n35
  );


  not
  g113
  (
    n120,
    n42
  );


  not
  g114
  (
    n192,
    n8
  );


  not
  g115
  (
    n111,
    n74
  );


  buf
  g116
  (
    n117,
    n74
  );


  buf
  g117
  (
    KeyWire_0_30,
    n7
  );


  not
  g118
  (
    n202,
    n15
  );


  not
  g119
  (
    KeyWire_0_55,
    n49
  );


  buf
  g120
  (
    KeyWire_0_52,
    n6
  );


  buf
  g121
  (
    n126,
    n47
  );


  not
  g122
  (
    n142,
    n59
  );


  not
  g123
  (
    n96,
    n33
  );


  buf
  g124
  (
    n147,
    n15
  );


  buf
  g125
  (
    KeyWire_0_17,
    n53
  );


  not
  g126
  (
    KeyWire_0_32,
    n34
  );


  buf
  g127
  (
    KeyWire_0_34,
    n58
  );


  not
  g128
  (
    n183,
    n10
  );


  not
  g129
  (
    n185,
    n66
  );


  buf
  g130
  (
    n169,
    n64
  );


  buf
  g131
  (
    KeyWire_0_35,
    n45
  );


  not
  g132
  (
    KeyWire_0_26,
    n73
  );


  not
  g133
  (
    n109,
    n40
  );


  not
  g134
  (
    KeyWire_0_4,
    n59
  );


  buf
  g135
  (
    n85,
    n9
  );


  buf
  g136
  (
    n131,
    n74
  );


  not
  g137
  (
    KeyWire_0_0,
    n71
  );


  not
  g138
  (
    KeyWire_0_29,
    n51
  );


  buf
  g139
  (
    n88,
    n62
  );


  not
  g140
  (
    n82,
    n43
  );


  buf
  g141
  (
    KeyWire_0_36,
    n75
  );


  buf
  g142
  (
    n193,
    n40
  );


  buf
  g143
  (
    n158,
    n37
  );


  not
  g144
  (
    KeyWire_0_43,
    n50
  );


  buf
  g145
  (
    n100,
    n49
  );


  not
  g146
  (
    n140,
    n71
  );


  buf
  g147
  (
    n110,
    n49
  );


  buf
  g148
  (
    n186,
    n38
  );


  buf
  g149
  (
    n191,
    n57
  );


  not
  g150
  (
    n119,
    n43
  );


  not
  g151
  (
    KeyWire_0_11,
    n37
  );


  not
  g152
  (
    KeyWire_0_18,
    n37
  );


  not
  g153
  (
    KeyWire_0_45,
    n46
  );


  buf
  g154
  (
    n162,
    n48
  );


  buf
  g155
  (
    n83,
    n48
  );


  not
  g156
  (
    n148,
    n66
  );


  buf
  g157
  (
    n195,
    n13
  );


  not
  g158
  (
    n95,
    n54
  );


  not
  g159
  (
    n204,
    n10
  );


  buf
  g160
  (
    KeyWire_0_40,
    n14
  );


  buf
  g161
  (
    n189,
    n75
  );


  buf
  g162
  (
    KeyWire_0_12,
    n55
  );


  not
  g163
  (
    n187,
    n39
  );


  buf
  g164
  (
    n200,
    n35
  );


  buf
  g165
  (
    n168,
    n73
  );


  not
  g166
  (
    n172,
    n34
  );


  not
  g167
  (
    n190,
    n53
  );


  buf
  g168
  (
    KeyWire_0_60,
    n72
  );


  not
  g169
  (
    KeyWire_0_47,
    n68
  );


  not
  g170
  (
    KeyWire_0_42,
    n61
  );


  buf
  g171
  (
    n177,
    n15
  );


  not
  g172
  (
    n153,
    n33
  );


  nor
  g173
  (
    n144,
    n16,
    n17
  );


  xor
  g174
  (
    KeyWire_0_1,
    n57,
    n6,
    n38,
    n36
  );


  or
  g175
  (
    n164,
    n70,
    n56,
    n11,
    n50
  );


  xor
  g176
  (
    KeyWire_0_7,
    n70,
    n9,
    n12,
    n56
  );


  and
  g177
  (
    n103,
    n17,
    n55,
    n68,
    n46
  );


  nand
  g178
  (
    n179,
    n10,
    n78,
    n6,
    n16
  );


  nand
  g179
  (
    n116,
    n13,
    n44,
    n64,
    n42
  );


  and
  g180
  (
    n121,
    n7,
    n51,
    n64,
    n72
  );


  and
  g181
  (
    KeyWire_0_20,
    n39,
    n44,
    n8,
    n47
  );


  and
  g182
  (
    KeyWire_0_33,
    n68,
    n67,
    n54,
    n61
  );


  xor
  g183
  (
    n173,
    n60,
    n16,
    n58,
    n52
  );


  xor
  g184
  (
    n167,
    n76,
    n12,
    n63,
    n67
  );


  or
  g185
  (
    n134,
    n62,
    n63,
    n69
  );


  xor
  g186
  (
    n113,
    n56,
    n36,
    n12,
    n51
  );


  nor
  g187
  (
    n135,
    n43,
    n11,
    n62,
    n58
  );


  xnor
  g188
  (
    n89,
    n13,
    n40,
    n11,
    n42
  );


  xnor
  g189
  (
    n220,
    n121,
    n135,
    n101,
    n184
  );


  and
  g190
  (
    n222,
    n204,
    n199,
    n196,
    n119
  );


  nand
  g191
  (
    n213,
    n87,
    n126,
    n206,
    n194
  );


  or
  g192
  (
    n208,
    n139,
    n120,
    n92,
    n183
  );


  and
  g193
  (
    KeyWire_0_14,
    n154,
    n198,
    n202,
    n163
  );


  and
  g194
  (
    n232,
    n109,
    n107,
    n96,
    n146
  );


  and
  g195
  (
    n225,
    n178,
    n158,
    n160,
    n102
  );


  xnor
  g196
  (
    n227,
    n179,
    n157,
    n145,
    n192
  );


  nand
  g197
  (
    n210,
    n83,
    n85,
    n193,
    n190
  );


  and
  g198
  (
    n218,
    n86,
    n182,
    n156,
    n148
  );


  xnor
  g199
  (
    n231,
    n99,
    n162,
    n128,
    n147
  );


  xor
  g200
  (
    n214,
    n169,
    n116,
    n88,
    n165
  );


  and
  g201
  (
    n224,
    n98,
    n79,
    n123,
    n143
  );


  and
  g202
  (
    n238,
    n104,
    n134,
    n132,
    n108
  );


  nand
  g203
  (
    KeyWire_0_58,
    n136,
    n131,
    n176,
    n172
  );


  or
  g204
  (
    n223,
    n170,
    n175,
    n106,
    n140
  );


  or
  g205
  (
    KeyWire_0_38,
    n186,
    n166,
    n168,
    n82
  );


  and
  g206
  (
    KeyWire_0_3,
    n110,
    n94,
    n173,
    n124
  );


  and
  g207
  (
    n211,
    n115,
    n138,
    n153,
    n149
  );


  and
  g208
  (
    n215,
    n195,
    n111,
    n137,
    n100
  );


  nand
  g209
  (
    KeyWire_0_19,
    n129,
    n197,
    n114,
    n95
  );


  xnor
  g210
  (
    n234,
    n151,
    n122,
    n91,
    n81
  );


  nand
  g211
  (
    KeyWire_0_24,
    n167,
    n150,
    n185,
    n171
  );


  xnor
  g212
  (
    n217,
    n187,
    n103,
    n152,
    n203
  );


  and
  g213
  (
    n235,
    n177,
    n105,
    n181,
    n113
  );


  and
  g214
  (
    n221,
    n84,
    n130,
    n191,
    n141
  );


  and
  g215
  (
    n230,
    n188,
    n161,
    n200,
    n180
  );


  or
  g216
  (
    KeyWire_0_6,
    n144,
    n89,
    n118,
    n142
  );


  xnor
  g217
  (
    n226,
    n112,
    n125,
    n97,
    n164
  );


  nor
  g218
  (
    n233,
    n90,
    n127,
    n189,
    n93
  );


  xor
  g219
  (
    KeyWire_0_25,
    n159,
    n117,
    n80,
    n174
  );


  and
  g220
  (
    n228,
    n201,
    n133,
    n155,
    n205
  );


  xnor
  KeyGate_0_0
  (
    n122,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n105,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n51,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n209,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n93,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n112,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n236,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n107,
    KeyNOTWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n33,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n104,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n136,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n198,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n175,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n25,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n219,
    KeyNOTWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n56,
    keyIn_0_15,
    KeyWire_0_15
  );


  xor
  KeyGate_0_16
  (
    KeyNOTWire_0_16,
    keyIn_0_16,
    KeyWire_0_16
  );


  not
  KeyNOTGate_0_16
  (
    n49,
    KeyNOTWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    KeyNOTWire_0_17,
    keyIn_0_17,
    KeyWire_0_17
  );


  not
  KeyNOTGate_0_17
  (
    n157,
    KeyNOTWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n194,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    KeyNOTWire_0_19,
    keyIn_0_19,
    KeyWire_0_19
  );


  not
  KeyNOTGate_0_19
  (
    n229,
    KeyNOTWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    KeyNOTWire_0_20,
    keyIn_0_20,
    KeyWire_0_20
  );


  not
  KeyNOTGate_0_20
  (
    n184,
    KeyNOTWire_0_20
  );


  xor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n59,
    KeyNOTWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n42,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n137,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n212,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n207,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n92,
    KeyNOTWire_0_26
  );


  xnor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n35,
    KeyNOTWire_0_27
  );


  xor
  KeyGate_0_28
  (
    KeyNOTWire_0_28,
    keyIn_0_28,
    KeyWire_0_28
  );


  not
  KeyNOTGate_0_28
  (
    n123,
    KeyNOTWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n163,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n129,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n133,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    KeyNOTWire_0_32,
    keyIn_0_32,
    KeyWire_0_32
  );


  not
  KeyNOTGate_0_32
  (
    n97,
    KeyNOTWire_0_32
  );


  xor
  KeyGate_0_33
  (
    n159,
    keyIn_0_33,
    KeyWire_0_33
  );


  xnor
  KeyGate_0_34
  (
    n151,
    keyIn_0_34,
    KeyWire_0_34
  );


  xor
  KeyGate_0_35
  (
    n161,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    KeyNOTWire_0_36,
    keyIn_0_36,
    KeyWire_0_36
  );


  not
  KeyNOTGate_0_36
  (
    n146,
    KeyNOTWire_0_36
  );


  xnor
  KeyGate_0_37
  (
    KeyNOTWire_0_37,
    keyIn_0_37,
    KeyWire_0_37
  );


  not
  KeyNOTGate_0_37
  (
    n205,
    KeyNOTWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n216,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    KeyNOTWire_0_39,
    keyIn_0_39,
    KeyWire_0_39
  );


  not
  KeyNOTGate_0_39
  (
    n176,
    KeyNOTWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    KeyNOTWire_0_40,
    keyIn_0_40,
    KeyWire_0_40
  );


  not
  KeyNOTGate_0_40
  (
    n86,
    KeyNOTWire_0_40
  );


  xnor
  KeyGate_0_41
  (
    KeyNOTWire_0_41,
    keyIn_0_41,
    KeyWire_0_41
  );


  not
  KeyNOTGate_0_41
  (
    n69,
    KeyNOTWire_0_41
  );


  xnor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n79,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    KeyNOTWire_0_43,
    keyIn_0_43,
    KeyWire_0_43
  );


  not
  KeyNOTGate_0_43
  (
    n152,
    KeyNOTWire_0_43
  );


  xor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n32,
    KeyNOTWire_0_44
  );


  xor
  KeyGate_0_45
  (
    KeyNOTWire_0_45,
    keyIn_0_45,
    KeyWire_0_45
  );


  not
  KeyNOTGate_0_45
  (
    n180,
    KeyNOTWire_0_45
  );


  xor
  KeyGate_0_46
  (
    n203,
    keyIn_0_46,
    KeyWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    n115,
    keyIn_0_47,
    KeyWire_0_47
  );


  xnor
  KeyGate_0_48
  (
    n29,
    keyIn_0_48,
    KeyWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n70,
    keyIn_0_49,
    KeyWire_0_49
  );


  xnor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n199,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n84,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    n114,
    keyIn_0_52,
    KeyWire_0_52
  );


  xor
  KeyGate_0_53
  (
    n155,
    keyIn_0_53,
    KeyWire_0_53
  );


  xnor
  KeyGate_0_54
  (
    n53,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n166,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    n31,
    keyIn_0_56,
    KeyWire_0_56
  );


  xnor
  KeyGate_0_57
  (
    KeyNOTWire_0_57,
    keyIn_0_57,
    KeyWire_0_57
  );


  not
  KeyNOTGate_0_57
  (
    n21,
    KeyNOTWire_0_57
  );


  xor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n237,
    KeyNOTWire_0_58
  );


  xor
  KeyGate_0_59
  (
    n101,
    keyIn_0_59,
    KeyWire_0_59
  );


  xor
  KeyGate_0_60
  (
    n171,
    keyIn_0_60,
    KeyWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n57,
    KeyNOTWire_0_61
  );


  xnor
  KeyGate_0_62
  (
    KeyNOTWire_0_62,
    keyIn_0_62,
    KeyWire_0_62
  );


  not
  KeyNOTGate_0_62
  (
    n62,
    KeyNOTWire_0_62
  );


  xnor
  KeyGate_0_63
  (
    n37,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

