// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_725_1628 written by SynthGen on 2021/05/24 19:48:29
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_725_1628 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21,
 n655, n652, n667, n666, n662, n669, n653, n665,
 n661, n651, n736, n740, n737, n742, n743, n738,
 n741, n739, n746, n744, n745);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21;

output n655, n652, n667, n666, n662, n669, n653, n665,
 n661, n651, n736, n740, n737, n742, n743, n738,
 n741, n739, n746, n744, n745;

wire n22, n23, n24, n25, n26, n27, n28, n29,
 n30, n31, n32, n33, n34, n35, n36, n37,
 n38, n39, n40, n41, n42, n43, n44, n45,
 n46, n47, n48, n49, n50, n51, n52, n53,
 n54, n55, n56, n57, n58, n59, n60, n61,
 n62, n63, n64, n65, n66, n67, n68, n69,
 n70, n71, n72, n73, n74, n75, n76, n77,
 n78, n79, n80, n81, n82, n83, n84, n85,
 n86, n87, n88, n89, n90, n91, n92, n93,
 n94, n95, n96, n97, n98, n99, n100, n101,
 n102, n103, n104, n105, n106, n107, n108, n109,
 n110, n111, n112, n113, n114, n115, n116, n117,
 n118, n119, n120, n121, n122, n123, n124, n125,
 n126, n127, n128, n129, n130, n131, n132, n133,
 n134, n135, n136, n137, n138, n139, n140, n141,
 n142, n143, n144, n145, n146, n147, n148, n149,
 n150, n151, n152, n153, n154, n155, n156, n157,
 n158, n159, n160, n161, n162, n163, n164, n165,
 n166, n167, n168, n169, n170, n171, n172, n173,
 n174, n175, n176, n177, n178, n179, n180, n181,
 n182, n183, n184, n185, n186, n187, n188, n189,
 n190, n191, n192, n193, n194, n195, n196, n197,
 n198, n199, n200, n201, n202, n203, n204, n205,
 n206, n207, n208, n209, n210, n211, n212, n213,
 n214, n215, n216, n217, n218, n219, n220, n221,
 n222, n223, n224, n225, n226, n227, n228, n229,
 n230, n231, n232, n233, n234, n235, n236, n237,
 n238, n239, n240, n241, n242, n243, n244, n245,
 n246, n247, n248, n249, n250, n251, n252, n253,
 n254, n255, n256, n257, n258, n259, n260, n261,
 n262, n263, n264, n265, n266, n267, n268, n269,
 n270, n271, n272, n273, n274, n275, n276, n277,
 n278, n279, n280, n281, n282, n283, n284, n285,
 n286, n287, n288, n289, n290, n291, n292, n293,
 n294, n295, n296, n297, n298, n299, n300, n301,
 n302, n303, n304, n305, n306, n307, n308, n309,
 n310, n311, n312, n313, n314, n315, n316, n317,
 n318, n319, n320, n321, n322, n323, n324, n325,
 n326, n327, n328, n329, n330, n331, n332, n333,
 n334, n335, n336, n337, n338, n339, n340, n341,
 n342, n343, n344, n345, n346, n347, n348, n349,
 n350, n351, n352, n353, n354, n355, n356, n357,
 n358, n359, n360, n361, n362, n363, n364, n365,
 n366, n367, n368, n369, n370, n371, n372, n373,
 n374, n375, n376, n377, n378, n379, n380, n381,
 n382, n383, n384, n385, n386, n387, n388, n389,
 n390, n391, n392, n393, n394, n395, n396, n397,
 n398, n399, n400, n401, n402, n403, n404, n405,
 n406, n407, n408, n409, n410, n411, n412, n413,
 n414, n415, n416, n417, n418, n419, n420, n421,
 n422, n423, n424, n425, n426, n427, n428, n429,
 n430, n431, n432, n433, n434, n435, n436, n437,
 n438, n439, n440, n441, n442, n443, n444, n445,
 n446, n447, n448, n449, n450, n451, n452, n453,
 n454, n455, n456, n457, n458, n459, n460, n461,
 n462, n463, n464, n465, n466, n467, n468, n469,
 n470, n471, n472, n473, n474, n475, n476, n477,
 n478, n479, n480, n481, n482, n483, n484, n485,
 n486, n487, n488, n489, n490, n491, n492, n493,
 n494, n495, n496, n497, n498, n499, n500, n501,
 n502, n503, n504, n505, n506, n507, n508, n509,
 n510, n511, n512, n513, n514, n515, n516, n517,
 n518, n519, n520, n521, n522, n523, n524, n525,
 n526, n527, n528, n529, n530, n531, n532, n533,
 n534, n535, n536, n537, n538, n539, n540, n541,
 n542, n543, n544, n545, n546, n547, n548, n549,
 n550, n551, n552, n553, n554, n555, n556, n557,
 n558, n559, n560, n561, n562, n563, n564, n565,
 n566, n567, n568, n569, n570, n571, n572, n573,
 n574, n575, n576, n577, n578, n579, n580, n581,
 n582, n583, n584, n585, n586, n587, n588, n589,
 n590, n591, n592, n593, n594, n595, n596, n597,
 n598, n599, n600, n601, n602, n603, n604, n605,
 n606, n607, n608, n609, n610, n611, n612, n613,
 n614, n615, n616, n617, n618, n619, n620, n621,
 n622, n623, n624, n625, n626, n627, n628, n629,
 n630, n631, n632, n633, n634, n635, n636, n637,
 n638, n639, n640, n641, n642, n643, n644, n645,
 n646, n647, n648, n649, n650, n654, n656, n657,
 n658, n659, n660, n663, n664, n668, n670, n671,
 n672, n673, n674, n675, n676, n677, n678, n679,
 n680, n681, n682, n683, n684, n685, n686, n687,
 n688, n689, n690, n691, n692, n693, n694, n695,
 n696, n697, n698, n699, n700, n701, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735;

not  g0 (n83, n15);
buf  g1 (n33, n1);
buf  g2 (n88, n9);
not  g3 (n61, n11);
not  g4 (n73, n1);
buf  g5 (n27, n16);
buf  g6 (n28, n10);
not  g7 (n23, n7);
buf  g8 (n69, n9);
not  g9 (n95, n3);
not  g10 (n25, n2);
not  g11 (n22, n8);
not  g12 (n29, n11);
buf  g13 (n91, n15);
buf  g14 (n85, n19);
buf  g15 (n47, n6);
buf  g16 (n32, n8);
not  g17 (n39, n13);
not  g18 (n36, n11);
not  g19 (n89, n19);
not  g20 (n78, n8);
not  g21 (n55, n19);
buf  g22 (n60, n13);
buf  g23 (n41, n18);
buf  g24 (n96, n5);
buf  g25 (n70, n10);
buf  g26 (n72, n7);
not  g27 (n24, n12);
buf  g28 (n86, n4);
buf  g29 (n74, n14);
buf  g30 (n75, n12);
not  g31 (n77, n6);
buf  g32 (n57, n10);
not  g33 (n43, n11);
buf  g34 (n71, n15);
buf  g35 (n54, n10);
buf  g36 (n53, n7);
buf  g37 (n48, n5);
not  g38 (n44, n1);
buf  g39 (n40, n17);
buf  g40 (n58, n4);
buf  g41 (n67, n2);
buf  g42 (n63, n9);
buf  g43 (n81, n17);
not  g44 (n82, n14);
buf  g45 (n76, n2);
not  g46 (n90, n12);
buf  g47 (n34, n6);
not  g48 (n26, n17);
not  g49 (n31, n15);
buf  g50 (n84, n18);
not  g51 (n62, n14);
not  g52 (n51, n16);
buf  g53 (n94, n13);
not  g54 (n56, n5);
buf  g55 (n59, n8);
buf  g56 (n79, n12);
not  g57 (n80, n3);
buf  g58 (n35, n13);
buf  g59 (n52, n18);
not  g60 (n92, n4);
not  g61 (n50, n16);
not  g62 (n65, n3);
not  g63 (n87, n6);
not  g64 (n37, n4);
not  g65 (n49, n17);
not  g66 (n30, n9);
not  g67 (n45, n14);
buf  g68 (n66, n2);
buf  g69 (n93, n18);
buf  g70 (n38, n1);
buf  g71 (n68, n3);
not  g72 (n42, n7);
buf  g73 (n64, n16);
buf  g74 (n46, n5);
not  g75 (n314, n34);
buf  g76 (n174, n54);
buf  g77 (n225, n62);
buf  g78 (n210, n76);
buf  g79 (n132, n73);
not  g80 (n187, n50);
buf  g81 (n195, n89);
buf  g82 (n276, n76);
not  g83 (n136, n58);
not  g84 (n113, n80);
not  g85 (n162, n27);
not  g86 (n232, n85);
buf  g87 (n266, n29);
buf  g88 (n101, n45);
not  g89 (n285, n28);
buf  g90 (n161, n88);
buf  g91 (n298, n38);
buf  g92 (n323, n27);
buf  g93 (n197, n28);
buf  g94 (n228, n70);
not  g95 (n190, n30);
not  g96 (n185, n80);
buf  g97 (n203, n47);
buf  g98 (n299, n77);
not  g99 (n194, n34);
buf  g100 (n319, n79);
buf  g101 (n175, n56);
not  g102 (n144, n43);
not  g103 (n109, n44);
not  g104 (n155, n55);
buf  g105 (n215, n54);
not  g106 (n333, n36);
buf  g107 (n240, n51);
not  g108 (n116, n82);
buf  g109 (n158, n82);
not  g110 (n335, n47);
not  g111 (n224, n25);
buf  g112 (n238, n86);
not  g113 (n310, n83);
buf  g114 (n153, n32);
not  g115 (n184, n59);
buf  g116 (n246, n78);
buf  g117 (n294, n31);
not  g118 (n181, n41);
not  g119 (n111, n54);
not  g120 (n98, n29);
not  g121 (n103, n75);
buf  g122 (n318, n36);
not  g123 (n202, n74);
buf  g124 (n163, n69);
not  g125 (n325, n83);
buf  g126 (n239, n52);
buf  g127 (n313, n55);
not  g128 (n262, n76);
buf  g129 (n105, n84);
buf  g130 (n265, n65);
buf  g131 (n193, n29);
not  g132 (n229, n81);
not  g133 (n307, n31);
not  g134 (n251, n35);
not  g135 (n236, n88);
not  g136 (n221, n61);
not  g137 (n334, n68);
buf  g138 (n283, n66);
not  g139 (n315, n74);
buf  g140 (n237, n40);
buf  g141 (n308, n64);
not  g142 (n254, n74);
buf  g143 (n128, n43);
buf  g144 (n167, n67);
not  g145 (n281, n56);
buf  g146 (n118, n61);
not  g147 (n189, n37);
not  g148 (n258, n57);
buf  g149 (n231, n57);
buf  g150 (n134, n87);
not  g151 (n164, n28);
buf  g152 (n279, n67);
buf  g153 (n226, n48);
not  g154 (n133, n22);
buf  g155 (n168, n37);
buf  g156 (n178, n24);
buf  g157 (n198, n75);
not  g158 (n119, n44);
not  g159 (n250, n84);
not  g160 (n110, n56);
not  g161 (n192, n69);
buf  g162 (n263, n70);
not  g163 (n150, n62);
buf  g164 (n270, n41);
buf  g165 (n145, n72);
buf  g166 (n141, n72);
buf  g167 (n274, n46);
buf  g168 (n146, n50);
not  g169 (n303, n59);
not  g170 (n324, n63);
buf  g171 (n252, n71);
not  g172 (n289, n57);
buf  g173 (n205, n31);
buf  g174 (n234, n69);
not  g175 (n320, n60);
not  g176 (n242, n41);
not  g177 (n269, n30);
not  g178 (n166, n64);
buf  g179 (n121, n65);
not  g180 (n165, n87);
buf  g181 (n117, n86);
not  g182 (n309, n63);
buf  g183 (n329, n26);
buf  g184 (n212, n38);
buf  g185 (n209, n71);
buf  g186 (n100, n23);
not  g187 (n312, n58);
buf  g188 (n247, n57);
not  g189 (n173, n47);
buf  g190 (n301, n51);
buf  g191 (n260, n52);
not  g192 (n122, n79);
buf  g193 (n152, n50);
buf  g194 (n326, n68);
buf  g195 (n142, n43);
not  g196 (n330, n73);
not  g197 (n104, n39);
not  g198 (n275, n58);
buf  g199 (n256, n50);
not  g200 (n139, n49);
not  g201 (n183, n84);
buf  g202 (n179, n29);
buf  g203 (n293, n61);
not  g204 (n147, n34);
not  g205 (n340, n67);
not  g206 (n255, n30);
buf  g207 (n259, n53);
not  g208 (n126, n39);
buf  g209 (n223, n43);
not  g210 (n108, n79);
not  g211 (n114, n35);
not  g212 (n268, n49);
buf  g213 (n245, n35);
buf  g214 (n339, n47);
not  g215 (n159, n38);
buf  g216 (n273, n80);
not  g217 (n154, n60);
not  g218 (n218, n87);
not  g219 (n125, n42);
buf  g220 (n213, n83);
not  g221 (n135, n26);
buf  g222 (n115, n77);
buf  g223 (n148, n89);
buf  g224 (n287, n30);
buf  g225 (n151, n71);
buf  g226 (n180, n64);
not  g227 (n149, n66);
buf  g228 (n337, n41);
not  g229 (n143, n75);
not  g230 (n284, n81);
buf  g231 (n176, n34);
buf  g232 (n156, n82);
not  g233 (n343, n64);
not  g234 (n131, n51);
not  g235 (n206, n65);
buf  g236 (n169, n66);
not  g237 (n196, n75);
buf  g238 (n140, n25);
buf  g239 (n130, n89);
not  g240 (n177, n48);
buf  g241 (n278, n81);
buf  g242 (n137, n73);
not  g243 (n248, n87);
buf  g244 (n305, n74);
buf  g245 (n297, n36);
not  g246 (n342, n83);
buf  g247 (n97, n82);
not  g248 (n188, n76);
not  g249 (n244, n56);
not  g250 (n295, n42);
not  g251 (n316, n45);
not  g252 (n331, n88);
buf  g253 (n200, n52);
not  g254 (n160, n69);
buf  g255 (n280, n23);
buf  g256 (n272, n49);
not  g257 (n328, n77);
not  g258 (n300, n86);
buf  g259 (n220, n46);
not  g260 (n230, n31);
buf  g261 (n282, n85);
not  g262 (n171, n37);
not  g263 (n204, n45);
not  g264 (n292, n33);
buf  g265 (n107, n48);
not  g266 (n243, n60);
buf  g267 (n214, n52);
not  g268 (n302, n62);
not  g269 (n341, n89);
buf  g270 (n261, n85);
not  g271 (n127, n62);
not  g272 (n112, n55);
not  g273 (n306, n72);
buf  g274 (n102, n53);
not  g275 (n120, n33);
not  g276 (n201, n48);
buf  g277 (n321, n58);
buf  g278 (n277, n70);
buf  g279 (n235, n65);
buf  g280 (n327, n53);
buf  g281 (n317, n68);
not  g282 (n216, n40);
buf  g283 (n172, n39);
buf  g284 (n157, n70);
not  g285 (n191, n63);
not  g286 (n344, n44);
not  g287 (n99, n37);
buf  g288 (n322, n85);
not  g289 (n182, n78);
not  g290 (n124, n35);
not  g291 (n222, n28);
not  g292 (n288, n24);
not  g293 (n249, n60);
not  g294 (n253, n88);
buf  g295 (n336, n46);
not  g296 (n227, n33);
buf  g297 (n286, n81);
not  g298 (n233, n45);
not  g299 (n123, n78);
not  g300 (n311, n38);
buf  g301 (n106, n72);
not  g302 (n291, n84);
buf  g303 (n217, n63);
not  g304 (n219, n55);
not  g305 (n271, n44);
buf  g306 (n186, n54);
not  g307 (n267, n59);
buf  g308 (n199, n46);
not  g309 (n170, n33);
buf  g310 (n264, n61);
buf  g311 (n129, n32);
buf  g312 (n208, n22);
buf  g313 (n290, n73);
not  g314 (n207, n67);
not  g315 (n338, n79);
buf  g316 (n304, n78);
not  g317 (n257, n77);
buf  g318 (n211, n86);
xor  g319 (n138, n66, n59, n51, n40);
nor  g320 (n241, n68, n71, n80, n42);
nand g321 (n332, n49, n42, n40, n32);
xnor g322 (n296, n32, n53, n36, n39);
nor  g323 (n398, n148, n220, n289, n173);
nor  g324 (n349, n237, n157, n281, n211);
xor  g325 (n387, n215, n20, n194, n231);
nand g326 (n361, n299, n306, n122, n201);
nor  g327 (n393, n310, n171, n240, n169);
or   g328 (n382, n307, n185, n142, n241);
or   g329 (n375, n101, n236, n188, n219);
nand g330 (n372, n164, n167, n116, n223);
nand g331 (n383, n277, n229, n301, n121);
nand g332 (n359, n295, n276, n257, n153);
or   g333 (n391, n292, n120, n177, n224);
and  g334 (n351, n287, n114, n228, n245);
xnor g335 (n370, n19, n104, n181, n258);
nand g336 (n397, n172, n217, n238, n191);
xnor g337 (n380, n165, n105, n242, n274);
nand g338 (n368, n260, n108, n226, n133);
and  g339 (n388, n145, n197, n192, n244);
xor  g340 (n399, n221, n235, n267, n204);
nand g341 (n350, n202, n168, n162, n302);
nor  g342 (n371, n175, n268, n225, n273);
nand g343 (n377, n113, n152, n198, n271);
nand g344 (n374, n111, n283, n186, n174);
or   g345 (n355, n20, n208, n146, n115);
or   g346 (n354, n130, n117, n139, n239);
or   g347 (n353, n259, n147, n161, n183);
or   g348 (n348, n97, n288, n230, n280);
or   g349 (n386, n232, n207, n166, n286);
xor  g350 (n362, n284, n123, n218, n250);
nand g351 (n392, n137, n243, n227, n21);
or   g352 (n345, n265, n159, n189, n216);
nor  g353 (n395, n107, n135, n21, n170);
nor  g354 (n363, n253, n300, n119, n297);
nand g355 (n352, n263, n141, n213, n149);
xor  g356 (n385, n180, n196, n247, n200);
nand g357 (n347, n126, n210, n151, n282);
or   g358 (n390, n234, n291, n251, n193);
or   g359 (n389, n311, n304, n278, n285);
xnor g360 (n369, n182, n118, n270, n296);
xnor g361 (n364, n261, n233, n248, n127);
and  g362 (n360, n294, n195, n184, n214);
nand g363 (n384, n102, n178, n99, n179);
and  g364 (n358, n144, n190, n138, n106);
or   g365 (n378, n110, n103, n112, n212);
nand g366 (n365, n209, n21, n269, n132);
xor  g367 (n367, n303, n205, n131, n21);
and  g368 (n394, n155, n143, n279, n203);
and  g369 (n376, n252, n124, n187, n128);
or   g370 (n381, n199, n98, n256, n255);
and  g371 (n373, n298, n266, n129, n160);
or   g372 (n379, n254, n20, n308, n305);
xor  g373 (n396, n154, n264, n158, n100);
nor  g374 (n366, n206, n262, n150, n125);
or   g375 (n400, n272, n249, n109, n290);
nor  g376 (n346, n275, n140, n176, n20);
nor  g377 (n357, n293, n134, n222, n163);
and  g378 (n356, n156, n136, n309, n246);
buf  g379 (n404, n372);
buf  g380 (n403, n360);
not  g381 (n406, n350);
buf  g382 (n416, n363);
not  g383 (n405, n357);
not  g384 (n415, n349);
buf  g385 (n401, n347);
buf  g386 (n408, n90);
buf  g387 (n417, n355);
buf  g388 (n409, n354);
buf  g389 (n412, n345);
buf  g390 (n410, n367);
xor  g391 (n413, n348, n362, n358, n365);
xor  g392 (n411, n90, n90, n353, n359);
xor  g393 (n407, n370, n366, n352, n361);
nor  g394 (n414, n346, n368, n90, n351);
xor  g395 (n402, n371, n369, n356, n364);
not  g396 (n430, n318);
not  g397 (n429, n93);
or   g398 (n424, n324, n91);
and  g399 (n420, n92, n401, n414, n410);
nor  g400 (n422, n321, n404, n406, n91);
or   g401 (n428, n92, n325, n327, n93);
nand g402 (n419, n94, n416, n412, n314);
nand g403 (n421, n409, n402, n91, n94);
or   g404 (n427, n96, n320, n403, n95);
nor  g405 (n426, n91, n319, n405, n93);
xnor g406 (n423, n323, n92, n95, n313);
xnor g407 (n418, n92, n315, n93, n408);
nor  g408 (n431, n411, n94, n415, n326);
and  g409 (n433, n95, n407, n96);
or   g410 (n432, n413, n317, n322, n316);
xor  g411 (n425, n94, n95, n96, n312);
not  g412 (n489, n426);
buf  g413 (n485, n423);
buf  g414 (n475, n422);
buf  g415 (n477, n430);
buf  g416 (n470, n431);
buf  g417 (n480, n422);
buf  g418 (n454, n374);
not  g419 (n436, n427);
not  g420 (n441, n423);
not  g421 (n478, n419);
buf  g422 (n490, n427);
buf  g423 (n450, n420);
buf  g424 (n443, n419);
not  g425 (n474, n421);
not  g426 (n471, n429);
buf  g427 (n469, n418);
buf  g428 (n465, n425);
buf  g429 (n444, n420);
not  g430 (n440, n425);
not  g431 (n484, n418);
buf  g432 (n488, n424);
buf  g433 (n479, n421);
buf  g434 (n461, n418);
buf  g435 (n456, n420);
buf  g436 (n448, n376);
not  g437 (n437, n426);
buf  g438 (n439, n426);
not  g439 (n468, n422);
buf  g440 (n463, n429);
buf  g441 (n457, n424);
buf  g442 (n449, n378);
buf  g443 (n452, n377);
buf  g444 (n473, n431);
buf  g445 (n486, n428);
not  g446 (n434, n431);
buf  g447 (n438, n428);
buf  g448 (n451, n430);
buf  g449 (n482, n424);
not  g450 (n472, n431);
buf  g451 (n447, n430);
buf  g452 (n435, n421);
buf  g453 (n442, n422);
not  g454 (n464, n429);
not  g455 (n467, n432);
buf  g456 (n476, n430);
not  g457 (n462, n373);
not  g458 (n453, n425);
buf  g459 (n455, n424);
not  g460 (n445, n421);
buf  g461 (n466, n420);
not  g462 (n459, n427);
not  g463 (n458, n375);
not  g464 (n487, n428);
and  g465 (n460, n423, n425);
or   g466 (n481, n427, n419);
nor  g467 (n446, n428, n429);
or   g468 (n483, n426, n418, n423, n419);
not  g469 (n513, n436);
buf  g470 (n511, n434);
buf  g471 (n509, n440);
buf  g472 (n514, n438);
buf  g473 (n517, n437);
not  g474 (n499, n437);
not  g475 (n494, n439);
buf  g476 (n498, n438);
not  g477 (n510, n381);
buf  g478 (n502, n439);
not  g479 (n497, n435);
not  g480 (n506, n441);
buf  g481 (n508, n382);
buf  g482 (n515, n439);
buf  g483 (n500, n436);
not  g484 (n491, n434);
not  g485 (n493, n380);
buf  g486 (n504, n435);
buf  g487 (n512, n383);
buf  g488 (n505, n438);
not  g489 (n503, n441);
not  g490 (n495, n440);
not  g491 (n492, n439);
not  g492 (n501, n437);
not  g493 (n516, n436);
nor  g494 (n496, n436, n440);
xnor g495 (n507, n437, n441, n438, n379);
buf  g496 (n519, n495);
buf  g497 (n525, n493);
buf  g498 (n532, n492);
buf  g499 (n526, n492);
not  g500 (n531, n494);
buf  g501 (n528, n495);
buf  g502 (n520, n494);
buf  g503 (n521, n417);
not  g504 (n529, n495);
buf  g505 (n523, n494);
not  g506 (n518, n492);
buf  g507 (n522, n493);
not  g508 (n533, n491);
buf  g509 (n524, n491);
buf  g510 (n527, n492);
buf  g511 (n534, n493);
or   g512 (n530, n494, n493);
or   g513 (n544, n531, n433, n451);
nand g514 (n551, n453, n445, n529);
or   g515 (n541, n443, n432, n523, n518);
or   g516 (n539, n433, n443, n445, n446);
and  g517 (n547, n520, n445, n528, n443);
and  g518 (n535, n446, n450, n447, n525);
xor  g519 (n549, n447, n452, n433, n441);
nor  g520 (n538, n526, n450, n449, n442);
nor  g521 (n546, n524, n442, n533, n453);
and  g522 (n542, n450, n447, n446, n522);
xnor g523 (n552, n527, n446, n534, n449);
nor  g524 (n550, n448, n442, n452, n444);
xnor g525 (n548, n444, n534, n451, n452);
nand g526 (n536, n443, n444, n448, n452);
nand g527 (n537, n449, n521, n432, n448);
nand g528 (n543, n442, n532, n444, n451);
xnor g529 (n545, n432, n448, n530, n453);
or   g530 (n540, n450, n519, n449, n447);
xnor g531 (n563, n461, n465, n502, n547);
and  g532 (n564, n547, n501, n476, n488);
xor  g533 (n583, n474, n498, n487, n536);
xnor g534 (n606, n539, n471, n470, n466);
nor  g535 (n562, n501, n550, n467, n500);
and  g536 (n565, n542, n470, n549, n468);
and  g537 (n582, n501, n488, n480, n546);
or   g538 (n610, n458, n495, n487, n546);
or   g539 (n574, n501, n540, n542, n502);
nor  g540 (n560, n540, n481, n461, n545);
and  g541 (n575, n476, n477, n463, n458);
nand g542 (n601, n478, n543, n467, n474);
or   g543 (n586, n486, n459, n535, n476);
and  g544 (n557, n482, n460, n475, n465);
nand g545 (n594, n458, n483, n478);
nor  g546 (n608, n459, n503, n486, n499);
nand g547 (n568, n504, n475, n482, n544);
nand g548 (n592, n474, n546, n548, n455);
nand g549 (n587, n469, n473, n455, n483);
and  g550 (n578, n488, n473, n543, n468);
or   g551 (n599, n477, n484, n462, n453);
nor  g552 (n554, n464, n485, n470, n478);
nand g553 (n593, n502, n471, n485, n538);
nand g554 (n604, n504, n462, n479, n457);
nor  g555 (n588, n539, n541, n547, n468);
and  g556 (n584, n504, n549, n539, n497);
or   g557 (n571, n484, n464, n465, n474);
or   g558 (n556, n497, n500, n460, n498);
nand g559 (n573, n503, n460, n481, n470);
xnor g560 (n569, n466, n484, n487, n467);
and  g561 (n605, n542, n469, n496);
xnor g562 (n600, n460, n455, n486, n483);
nand g563 (n579, n500, n543, n537, n497);
nor  g564 (n581, n454, n538, n477, n482);
nor  g565 (n555, n536, n548, n462, n472);
nor  g566 (n570, n472, n546, n503, n457);
or   g567 (n566, n463, n475, n464, n476);
xor  g568 (n580, n504, n544, n542, n467);
and  g569 (n602, n539, n502, n536, n484);
and  g570 (n596, n549, n479, n463, n544);
or   g571 (n597, n548, n547, n540, n535);
nand g572 (n577, n498, n454, n545, n536);
xnor g573 (n590, n541, n544, n497, n475);
and  g574 (n567, n537, n471, n480, n473);
and  g575 (n595, n463, n454, n496, n538);
nor  g576 (n576, n454, n498, n485, n469);
or   g577 (n559, n549, n479, n466, n500);
and  g578 (n591, n459, n464, n481, n456);
nand g579 (n609, n543, n461, n499, n473);
xnor g580 (n598, n537, n459, n457, n541);
xnor g581 (n611, n545, n538, n481, n456);
xor  g582 (n561, n478, n485, n462, n461);
nand g583 (n553, n472, n487, n496, n471);
xnor g584 (n585, n457, n480, n458, n472);
nand g585 (n572, n486, n456, n503, n465);
and  g586 (n607, n466, n499, n456, n540);
xnor g587 (n558, n480, n455, n468, n499);
nor  g588 (n589, n479, n545, n541, n548);
xor  g589 (n603, n477, n537, n469, n482);
buf  g590 (n616, n505);
buf  g591 (n617, n507);
buf  g592 (n614, n557);
not  g593 (n621, n556);
not  g594 (n613, n507);
not  g595 (n618, n554);
buf  g596 (n623, n507);
not  g597 (n619, n507);
or   g598 (n612, n558, n506, n557, n505);
or   g599 (n622, n555, n506, n559, n505);
xor  g600 (n615, n553, n555, n559, n506);
xor  g601 (n620, n556, n505, n558, n506);
not  g602 (n647, n392);
buf  g603 (n639, n620);
not  g604 (n643, n619);
not  g605 (n633, n384);
not  g606 (n644, n616);
buf  g607 (n626, n389);
buf  g608 (n641, n612);
not  g609 (n632, n612);
not  g610 (n645, n614);
not  g611 (n629, n617);
not  g612 (n637, n621);
not  g613 (n630, n621);
buf  g614 (n638, n618);
buf  g615 (n634, n621);
not  g616 (n631, n391);
not  g617 (n627, n615);
buf  g618 (n642, n622);
buf  g619 (n624, n613);
not  g620 (n640, n388);
buf  g621 (n625, n620);
nor  g622 (n635, n613, n622);
xnor g623 (n628, n386, n616, n385, n393);
xnor g624 (n636, n387, n615, n617, n618);
nor  g625 (n646, n614, n619, n621, n390);
nand g626 (n665, n625, n552, n561, n572);
xnor g627 (n669, n508, n581, n580, n509);
and  g628 (n664, n509, n566, n395, n574);
nor  g629 (n663, n626, n577, n576, n624);
nor  g630 (n648, n510, n508, n551, n627);
xor  g631 (n672, n394, n564, n561, n584);
nand g632 (n666, n625, n550, n576, n509);
xnor g633 (n670, n396, n579, n624, n573);
nor  g634 (n659, n628, n629, n568, n574);
xnor g635 (n660, n583, n562, n552, n575);
or   g636 (n651, n585, n585, n575, n577);
nor  g637 (n655, n582, n398, n560, n584);
nor  g638 (n654, n509, n400, n569, n571);
and  g639 (n661, n579, n628, n567, n510);
xor  g640 (n652, n626, n563, n551, n630);
nor  g641 (n673, n629, n580, n627, n624);
or   g642 (n650, n550, n508, n628);
xnor g643 (n668, n582, n565, n572, n573);
xor  g644 (n671, n551, n628, n586, n630);
xnor g645 (n656, n570, n578, n624, n625);
nor  g646 (n658, n552, n578, n563, n550);
or   g647 (n649, n560, n629, n569, n551);
nor  g648 (n653, n571, n566, n565, n562);
nand g649 (n657, n625, n568, n570, n626);
and  g650 (n667, n629, n567, n564, n397);
nand g651 (n662, n627, n399, n581, n552);
xnor g652 (n674, n583, n627, n626, n630);
xnor g653 (n689, n596, n659, n605, n660);
or   g654 (n680, n662, n602, n586, n665);
xor  g655 (n682, n610, n611, n600, n668);
or   g656 (n677, n664, n599, n593);
xor  g657 (n684, n606, n597, n666, n607);
or   g658 (n686, n667, n598, n673, n591);
xnor g659 (n685, n594, n588, n605);
xor  g660 (n690, n604, n597, n601, n606);
or   g661 (n691, n590, n604, n589, n603);
nor  g662 (n681, n661, n599, n595, n670);
nand g663 (n679, n601, n663, n609, n600);
and  g664 (n676, n592, n592, n669, n589);
and  g665 (n675, n610, n591, n658, n608);
xnor g666 (n687, n608, n671, n603, n611);
nor  g667 (n678, n609, n595, n587, n596);
nand g668 (n683, n607, n590, n594, n598);
xor  g669 (n688, n602, n674, n587, n672);
xnor g670 (n735, n515, n690, n513, n639);
xor  g671 (n719, n489, n512, n635, n647);
or   g672 (n732, n642, n687, n646, n637);
and  g673 (n714, n513, n513, n636, n640);
and  g674 (n726, n682, n514, n642, n340);
xnor g675 (n696, n640, n635, n623, n684);
or   g676 (n708, n644, n515, n339, n334);
xnor g677 (n724, n490, n676, n516, n517);
xor  g678 (n698, n329, n634, n623, n690);
xor  g679 (n718, n517, n643, n641, n489);
nor  g680 (n720, n622, n515, n335, n642);
nor  g681 (n722, n512, n488, n631, n647);
nand g682 (n715, n632, n511, n644, n678);
xor  g683 (n702, n639, n640, n685, n510);
and  g684 (n734, n637, n639, n678, n644);
xnor g685 (n699, n643, n514, n684, n631);
nand g686 (n700, n646, n676, n517, n644);
and  g687 (n712, n689, n510, n682, n685);
nor  g688 (n733, n635, n641, n638, n684);
xor  g689 (n710, n681, n634, n632, n511);
xor  g690 (n711, n633, n638, n516, n689);
and  g691 (n707, n630, n638, n433, n343);
xor  g692 (n727, n342, n336, n513, n681);
and  g693 (n709, n632, n647, n634, n511);
and  g694 (n695, n636, n633, n689, n517);
xor  g695 (n694, n512, n642, n687, n688);
xnor g696 (n701, n637, n631, n632, n677);
or   g697 (n697, n641, n688, n634, n344);
nand g698 (n713, n685, n489, n516, n643);
nand g699 (n693, n639, n490, n675, n686);
and  g700 (n716, n679, n635, n688, n330);
and  g701 (n731, n623, n691, n328);
xor  g702 (n705, n514, n633, n677, n643);
nor  g703 (n717, n337, n646, n333, n641);
xnor g704 (n704, n647, n515, n638, n623);
nand g705 (n706, n516, n691, n512, n511);
and  g706 (n721, n686, n640, n680, n675);
and  g707 (n729, n646, n680, n686, n683);
or   g708 (n730, n679, n490, n338, n622);
xor  g709 (n703, n636, n690, n489, n645);
nor  g710 (n728, n633, n645, n687, n341);
xnor g711 (n692, n490, n631, n682, n683);
and  g712 (n723, n637, n332, n636, n683);
or   g713 (n725, n331, n645, n514);
nor  g714 (n744, n693, n696, n692, n695);
and  g715 (n739, n721, n723, n701, n709);
nand g716 (n738, n694, n727, n726, n699);
nand g717 (n745, n735, n730, n710, n717);
xor  g718 (n740, n698, n702, n706, n713);
nor  g719 (n746, n719, n708, n724, n700);
xor  g720 (n741, n729, n722, n716, n715);
xor  g721 (n742, n733, n703, n705, n720);
nor  g722 (n736, n728, n732, n711, n734);
xor  g723 (n737, n697, n707, n718, n712);
and  g724 (n743, n725, n714, n731, n704);
endmodule
