

module Stat_1000_153
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n1004,
  n991,
  n988,
  n990,
  n992,
  n995,
  n1005,
  n1010,
  n987,
  n1009,
  n996,
  n1014,
  n994,
  n1012,
  n989,
  n1008,
  n1001,
  n1015,
  n1013,
  n1017,
  n998,
  n1019,
  n1007,
  n993,
  n1011,
  n1018,
  n1020,
  n1022,
  n1024,
  n1025,
  n1032,
  n1031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;input keyIn_0_32;input keyIn_0_33;input keyIn_0_34;input keyIn_0_35;input keyIn_0_36;input keyIn_0_37;input keyIn_0_38;input keyIn_0_39;input keyIn_0_40;input keyIn_0_41;input keyIn_0_42;input keyIn_0_43;input keyIn_0_44;input keyIn_0_45;input keyIn_0_46;input keyIn_0_47;input keyIn_0_48;input keyIn_0_49;input keyIn_0_50;input keyIn_0_51;input keyIn_0_52;input keyIn_0_53;input keyIn_0_54;input keyIn_0_55;input keyIn_0_56;input keyIn_0_57;input keyIn_0_58;input keyIn_0_59;input keyIn_0_60;input keyIn_0_61;input keyIn_0_62;input keyIn_0_63;
  output n1004;output n991;output n988;output n990;output n992;output n995;output n1005;output n1010;output n987;output n1009;output n996;output n1014;output n994;output n1012;output n989;output n1008;output n1001;output n1015;output n1013;output n1017;output n998;output n1019;output n1007;output n993;output n1011;output n1018;output n1020;output n1022;output n1024;output n1025;output n1032;output n1031;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n997;wire n999;wire n1000;wire n1002;wire n1003;wire n1006;wire n1016;wire n1021;wire n1023;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire g_input_0_0;wire gbar_input_0_0;wire g_input_0_1;wire gbar_input_0_1;wire g_input_0_2;wire gbar_input_0_2;wire g_input_0_3;wire gbar_input_0_3;wire g_input_0_4;wire gbar_input_0_4;wire g_input_0_5;wire gbar_input_0_5;wire g_input_0_6;wire gbar_input_0_6;wire g_input_0_7;wire gbar_input_0_7;wire g_input_0_8;wire gbar_input_0_8;wire g_input_0_9;wire gbar_input_0_9;wire g_input_0_10;wire gbar_input_0_10;wire g_input_0_11;wire gbar_input_0_11;wire g_input_0_12;wire gbar_input_0_12;wire g_input_0_13;wire gbar_input_0_13;wire g_input_0_14;wire gbar_input_0_14;wire g_input_0_15;wire gbar_input_0_15;wire g_input_0_16;wire gbar_input_0_16;wire g_input_0_17;wire gbar_input_0_17;wire g_input_0_18;wire gbar_input_0_18;wire g_input_0_19;wire gbar_input_0_19;wire g_input_0_20;wire gbar_input_0_20;wire g_input_0_21;wire gbar_input_0_21;wire g_input_0_22;wire gbar_input_0_22;wire g_input_0_23;wire gbar_input_0_23;wire g_input_0_24;wire gbar_input_0_24;wire g_input_0_25;wire gbar_input_0_25;wire g_input_0_26;wire gbar_input_0_26;wire g_input_0_27;wire gbar_input_0_27;wire g_input_0_28;wire gbar_input_0_28;wire g_input_0_29;wire gbar_input_0_29;wire g_input_0_30;wire gbar_input_0_30;wire g_input_0_31;wire gbar_input_0_31;wire f_g_wire;wire f_gbar_wire;wire AntiSAT_output;

  buf
  g0
  (
    n108,
    n17
  );


  buf
  g1
  (
    n40,
    n23
  );


  buf
  g2
  (
    n139,
    n11
  );


  buf
  g3
  (
    n36,
    n9
  );


  not
  g4
  (
    n126,
    n14
  );


  buf
  g5
  (
    n54,
    n20
  );


  buf
  g6
  (
    n85,
    n3
  );


  not
  g7
  (
    n98,
    n20
  );


  buf
  g8
  (
    n34,
    n4
  );


  not
  g9
  (
    n128,
    n7
  );


  not
  g10
  (
    n41,
    n5
  );


  buf
  g11
  (
    n71,
    n26
  );


  buf
  g12
  (
    n148,
    n10
  );


  buf
  g13
  (
    n152,
    n29
  );


  buf
  g14
  (
    n47,
    n25
  );


  buf
  g15
  (
    n63,
    n24
  );


  buf
  g16
  (
    n94,
    n23
  );


  not
  g17
  (
    n107,
    n30
  );


  not
  g18
  (
    n33,
    n13
  );


  buf
  g19
  (
    n127,
    n14
  );


  not
  g20
  (
    n142,
    n5
  );


  not
  g21
  (
    n84,
    n21
  );


  not
  g22
  (
    n109,
    n21
  );


  buf
  g23
  (
    n104,
    n6
  );


  not
  g24
  (
    n42,
    n21
  );


  buf
  g25
  (
    n61,
    n15
  );


  not
  g26
  (
    n100,
    n9
  );


  not
  g27
  (
    n120,
    n20
  );


  not
  g28
  (
    n66,
    n15
  );


  buf
  g29
  (
    n86,
    n6
  );


  buf
  g30
  (
    n87,
    n12
  );


  not
  g31
  (
    n133,
    n3
  );


  not
  g32
  (
    n93,
    n25
  );


  not
  g33
  (
    n44,
    n19
  );


  buf
  g34
  (
    n48,
    n14
  );


  not
  g35
  (
    n143,
    n16
  );


  buf
  g36
  (
    n39,
    n1
  );


  not
  g37
  (
    n82,
    n19
  );


  buf
  g38
  (
    n130,
    n7
  );


  buf
  g39
  (
    n81,
    n17
  );


  not
  g40
  (
    n96,
    n31
  );


  buf
  g41
  (
    n146,
    n9
  );


  buf
  g42
  (
    n149,
    n16
  );


  buf
  g43
  (
    n125,
    n14
  );


  not
  g44
  (
    n45,
    n9
  );


  not
  g45
  (
    n80,
    n16
  );


  buf
  g46
  (
    n118,
    n5
  );


  not
  g47
  (
    n60,
    n7
  );


  buf
  g48
  (
    n52,
    n2
  );


  not
  g49
  (
    n132,
    n16
  );


  not
  g50
  (
    n70,
    n15
  );


  buf
  g51
  (
    n90,
    n10
  );


  buf
  g52
  (
    n105,
    n29
  );


  not
  g53
  (
    n151,
    n27
  );


  buf
  g54
  (
    n123,
    n31
  );


  buf
  g55
  (
    n131,
    n22
  );


  buf
  g56
  (
    n53,
    n1
  );


  buf
  g57
  (
    n67,
    n19
  );


  buf
  g58
  (
    n88,
    n17
  );


  not
  g59
  (
    n141,
    n29
  );


  not
  g60
  (
    n113,
    n11
  );


  not
  g61
  (
    n116,
    n13
  );


  not
  g62
  (
    n137,
    n24
  );


  buf
  g63
  (
    n62,
    n26
  );


  buf
  g64
  (
    n49,
    n19
  );


  buf
  g65
  (
    n124,
    n30
  );


  not
  g66
  (
    n57,
    n22
  );


  buf
  g67
  (
    n144,
    n23
  );


  buf
  g68
  (
    n35,
    n30
  );


  not
  g69
  (
    n46,
    n4
  );


  buf
  g70
  (
    n112,
    n8
  );


  buf
  g71
  (
    n77,
    n12
  );


  not
  g72
  (
    n64,
    n28
  );


  not
  g73
  (
    n83,
    n18
  );


  not
  g74
  (
    n135,
    n8
  );


  buf
  g75
  (
    n145,
    n13
  );


  buf
  g76
  (
    n99,
    n18
  );


  not
  g77
  (
    n37,
    n4
  );


  not
  g78
  (
    n69,
    n20
  );


  buf
  g79
  (
    n68,
    n31
  );


  buf
  g80
  (
    n122,
    n22
  );


  buf
  g81
  (
    n89,
    n7
  );


  buf
  g82
  (
    n138,
    n6
  );


  buf
  g83
  (
    n72,
    n8
  );


  buf
  g84
  (
    n121,
    n30
  );


  not
  g85
  (
    n91,
    n4
  );


  not
  g86
  (
    n140,
    n21
  );


  not
  g87
  (
    n101,
    n26
  );


  not
  g88
  (
    n103,
    n3
  );


  not
  g89
  (
    n58,
    n1
  );


  buf
  g90
  (
    n43,
    n18
  );


  buf
  g91
  (
    n136,
    n25
  );


  buf
  g92
  (
    n97,
    n11
  );


  buf
  g93
  (
    n129,
    n12
  );


  buf
  g94
  (
    n117,
    n26
  );


  buf
  g95
  (
    n55,
    n11
  );


  not
  g96
  (
    n38,
    n8
  );


  not
  g97
  (
    n119,
    n2
  );


  buf
  g98
  (
    n92,
    n5
  );


  buf
  g99
  (
    n65,
    n23
  );


  not
  g100
  (
    n147,
    n24
  );


  not
  g101
  (
    n111,
    n6
  );


  buf
  g102
  (
    n56,
    n10
  );


  not
  g103
  (
    n74,
    n15
  );


  buf
  g104
  (
    n51,
    n28
  );


  not
  g105
  (
    n114,
    n27
  );


  not
  g106
  (
    n106,
    n18
  );


  buf
  g107
  (
    n102,
    n10
  );


  not
  g108
  (
    n110,
    n28
  );


  buf
  g109
  (
    n73,
    n29
  );


  buf
  g110
  (
    n79,
    n12
  );


  buf
  g111
  (
    n150,
    n17
  );


  buf
  g112
  (
    n59,
    n28
  );


  not
  g113
  (
    n134,
    n27
  );


  not
  g114
  (
    n115,
    n24
  );


  not
  g115
  (
    n75,
    n13
  );


  not
  g116
  (
    n95,
    n22
  );


  buf
  g117
  (
    n76,
    n25
  );


  buf
  g118
  (
    n78,
    n27
  );


  not
  g119
  (
    n50,
    n2
  );


  not
  g120
  (
    n291,
    n56
  );


  not
  g121
  (
    n327,
    n33
  );


  buf
  g122
  (
    n233,
    n40
  );


  buf
  g123
  (
    n303,
    n34
  );


  buf
  g124
  (
    n219,
    n63
  );


  buf
  g125
  (
    n260,
    n37
  );


  buf
  g126
  (
    n302,
    n56
  );


  buf
  g127
  (
    n316,
    n46
  );


  not
  g128
  (
    n189,
    n35
  );


  buf
  g129
  (
    n325,
    n52
  );


  buf
  g130
  (
    n211,
    n73
  );


  not
  g131
  (
    n156,
    n73
  );


  buf
  g132
  (
    n162,
    n46
  );


  not
  g133
  (
    n193,
    n62
  );


  buf
  g134
  (
    n235,
    n38
  );


  buf
  g135
  (
    n241,
    n70
  );


  not
  g136
  (
    n209,
    n47
  );


  buf
  g137
  (
    n246,
    n56
  );


  not
  g138
  (
    n312,
    n40
  );


  buf
  g139
  (
    n252,
    n56
  );


  not
  g140
  (
    n282,
    n69
  );


  not
  g141
  (
    n185,
    n76
  );


  buf
  g142
  (
    n247,
    n54
  );


  not
  g143
  (
    n216,
    n42
  );


  buf
  g144
  (
    n323,
    n64
  );


  not
  g145
  (
    n250,
    n50
  );


  not
  g146
  (
    n321,
    n65
  );


  not
  g147
  (
    n191,
    n45
  );


  not
  g148
  (
    n256,
    n50
  );


  buf
  g149
  (
    n217,
    n71
  );


  not
  g150
  (
    n164,
    n47
  );


  not
  g151
  (
    n244,
    n51
  );


  buf
  g152
  (
    n227,
    n53
  );


  not
  g153
  (
    n163,
    n57
  );


  not
  g154
  (
    n290,
    n75
  );


  not
  g155
  (
    n236,
    n59
  );


  not
  g156
  (
    n218,
    n72
  );


  not
  g157
  (
    n175,
    n51
  );


  not
  g158
  (
    n172,
    n37
  );


  not
  g159
  (
    n157,
    n68
  );


  buf
  g160
  (
    n258,
    n67
  );


  buf
  g161
  (
    n155,
    n36
  );


  buf
  g162
  (
    n311,
    n50
  );


  buf
  g163
  (
    n269,
    n53
  );


  buf
  g164
  (
    n285,
    n48
  );


  buf
  g165
  (
    n314,
    n52
  );


  buf
  g166
  (
    n309,
    n68
  );


  not
  g167
  (
    n170,
    n62
  );


  buf
  g168
  (
    n226,
    n48
  );


  buf
  g169
  (
    n153,
    n37
  );


  not
  g170
  (
    n243,
    n49
  );


  not
  g171
  (
    n300,
    n35
  );


  not
  g172
  (
    n166,
    n63
  );


  buf
  g173
  (
    n293,
    n55
  );


  buf
  g174
  (
    n232,
    n41
  );


  buf
  g175
  (
    n313,
    n76
  );


  not
  g176
  (
    n305,
    n38
  );


  not
  g177
  (
    n186,
    n73
  );


  not
  g178
  (
    n284,
    n36
  );


  buf
  g179
  (
    n304,
    n68
  );


  buf
  g180
  (
    n322,
    n75
  );


  buf
  g181
  (
    n263,
    n74
  );


  buf
  g182
  (
    n173,
    n52
  );


  not
  g183
  (
    n165,
    n49
  );


  not
  g184
  (
    n265,
    n53
  );


  not
  g185
  (
    n274,
    n61
  );


  not
  g186
  (
    n308,
    n48
  );


  not
  g187
  (
    n229,
    n58
  );


  buf
  g188
  (
    n295,
    n66
  );


  not
  g189
  (
    n206,
    n74
  );


  buf
  g190
  (
    n286,
    n51
  );


  not
  g191
  (
    n188,
    n35
  );


  not
  g192
  (
    n329,
    n63
  );


  buf
  g193
  (
    n196,
    n63
  );


  buf
  g194
  (
    n179,
    n45
  );


  buf
  g195
  (
    n177,
    n33
  );


  buf
  g196
  (
    n223,
    n41
  );


  not
  g197
  (
    n181,
    n46
  );


  buf
  g198
  (
    n264,
    n75
  );


  buf
  g199
  (
    n254,
    n36
  );


  buf
  g200
  (
    n310,
    n35
  );


  buf
  g201
  (
    n301,
    n70
  );


  buf
  g202
  (
    n326,
    n55
  );


  not
  g203
  (
    n272,
    n62
  );


  not
  g204
  (
    n294,
    n57
  );


  not
  g205
  (
    n180,
    n61
  );


  buf
  g206
  (
    n242,
    n61
  );


  buf
  g207
  (
    n195,
    n37
  );


  not
  g208
  (
    n281,
    n34
  );


  not
  g209
  (
    n324,
    n36
  );


  not
  g210
  (
    n200,
    n44
  );


  not
  g211
  (
    n187,
    n42
  );


  buf
  g212
  (
    n296,
    n38
  );


  not
  g213
  (
    n237,
    n38
  );


  buf
  g214
  (
    n292,
    n54
  );


  buf
  g215
  (
    n255,
    n76
  );


  not
  g216
  (
    n280,
    n66
  );


  buf
  g217
  (
    n205,
    n45
  );


  not
  g218
  (
    n299,
    n43
  );


  buf
  g219
  (
    n184,
    n57
  );


  not
  g220
  (
    n202,
    n71
  );


  buf
  g221
  (
    n198,
    n48
  );


  buf
  g222
  (
    n262,
    n65
  );


  not
  g223
  (
    n270,
    n44
  );


  not
  g224
  (
    n306,
    n46
  );


  buf
  g225
  (
    n214,
    n70
  );


  not
  g226
  (
    n231,
    n72
  );


  not
  g227
  (
    n251,
    n39
  );


  buf
  g228
  (
    n288,
    n42
  );


  buf
  g229
  (
    n176,
    n77
  );


  buf
  g230
  (
    n277,
    n53
  );


  buf
  g231
  (
    n230,
    n62
  );


  not
  g232
  (
    n275,
    n64
  );


  buf
  g233
  (
    n317,
    n33
  );


  not
  g234
  (
    n192,
    n59
  );


  not
  g235
  (
    n276,
    n58
  );


  buf
  g236
  (
    n319,
    n42
  );


  not
  g237
  (
    n183,
    n45
  );


  not
  g238
  (
    n215,
    n68
  );


  buf
  g239
  (
    n154,
    n73
  );


  buf
  g240
  (
    n210,
    n41
  );


  buf
  g241
  (
    n182,
    n52
  );


  buf
  g242
  (
    n289,
    n41
  );


  not
  g243
  (
    n208,
    n71
  );


  not
  g244
  (
    n160,
    n69
  );


  buf
  g245
  (
    n174,
    n44
  );


  not
  g246
  (
    n261,
    n71
  );


  buf
  g247
  (
    n167,
    n43
  );


  not
  g248
  (
    n224,
    n47
  );


  not
  g249
  (
    n178,
    n49
  );


  buf
  g250
  (
    n245,
    n47
  );


  buf
  g251
  (
    n161,
    n39
  );


  not
  g252
  (
    n328,
    n65
  );


  buf
  g253
  (
    n213,
    n61
  );


  not
  g254
  (
    n225,
    n39
  );


  buf
  g255
  (
    n234,
    n39
  );


  buf
  g256
  (
    n283,
    n74
  );


  buf
  g257
  (
    n253,
    n34
  );


  not
  g258
  (
    n279,
    n72
  );


  buf
  g259
  (
    n320,
    n51
  );


  buf
  g260
  (
    n257,
    n57
  );


  buf
  g261
  (
    n239,
    n34
  );


  buf
  g262
  (
    n228,
    n65
  );


  buf
  g263
  (
    n220,
    n59
  );


  buf
  g264
  (
    n287,
    n43
  );


  not
  g265
  (
    n197,
    n58
  );


  not
  g266
  (
    n240,
    n70
  );


  buf
  g267
  (
    n297,
    n60
  );


  not
  g268
  (
    n271,
    n66
  );


  buf
  g269
  (
    n199,
    n64
  );


  buf
  g270
  (
    n273,
    n49
  );


  not
  g271
  (
    n158,
    n50
  );


  buf
  g272
  (
    n318,
    n66
  );


  buf
  g273
  (
    n278,
    n69
  );


  buf
  g274
  (
    n204,
    n76
  );


  buf
  g275
  (
    n203,
    n58
  );


  not
  g276
  (
    n159,
    n75
  );


  buf
  g277
  (
    n267,
    n55
  );


  buf
  g278
  (
    n268,
    n72
  );


  buf
  g279
  (
    n307,
    n69
  );


  not
  g280
  (
    n201,
    n59
  );


  not
  g281
  (
    n207,
    n55
  );


  not
  g282
  (
    n222,
    n74
  );


  not
  g283
  (
    n315,
    n40
  );


  buf
  g284
  (
    n194,
    n33
  );


  buf
  g285
  (
    n190,
    n60
  );


  buf
  g286
  (
    n238,
    n67
  );


  buf
  g287
  (
    n248,
    n60
  );


  not
  g288
  (
    n249,
    n54
  );


  not
  g289
  (
    n259,
    n67
  );


  buf
  g290
  (
    n221,
    n67
  );


  not
  g291
  (
    n212,
    n43
  );


  buf
  g292
  (
    n298,
    n40
  );


  buf
  g293
  (
    n168,
    n60
  );


  buf
  g294
  (
    n266,
    n54
  );


  buf
  g295
  (
    n171,
    n64
  );


  buf
  g296
  (
    n169,
    n44
  );


  not
  g297
  (
    n519,
    n220
  );


  buf
  g298
  (
    n476,
    n322
  );


  not
  g299
  (
    n345,
    n227
  );


  not
  g300
  (
    n516,
    n189
  );


  buf
  g301
  (
    n405,
    n290
  );


  buf
  g302
  (
    n397,
    n307
  );


  not
  g303
  (
    n420,
    n303
  );


  not
  g304
  (
    n391,
    n265
  );


  buf
  g305
  (
    n571,
    n262
  );


  not
  g306
  (
    n555,
    n266
  );


  buf
  g307
  (
    n562,
    n279
  );


  buf
  g308
  (
    n483,
    n274
  );


  buf
  g309
  (
    n374,
    n183
  );


  buf
  g310
  (
    n347,
    n160
  );


  not
  g311
  (
    n379,
    n254
  );


  buf
  g312
  (
    n518,
    n286
  );


  buf
  g313
  (
    n498,
    n164
  );


  buf
  g314
  (
    n487,
    n191
  );


  not
  g315
  (
    n552,
    n203
  );


  buf
  g316
  (
    n439,
    n82
  );


  buf
  g317
  (
    n400,
    n313
  );


  not
  g318
  (
    n526,
    n235
  );


  buf
  g319
  (
    n393,
    n313
  );


  buf
  g320
  (
    n425,
    n168
  );


  not
  g321
  (
    n448,
    n288
  );


  not
  g322
  (
    n422,
    n274
  );


  buf
  g323
  (
    n511,
    n199
  );


  not
  g324
  (
    n560,
    n169
  );


  buf
  g325
  (
    n394,
    n252
  );


  buf
  g326
  (
    n433,
    n292
  );


  buf
  g327
  (
    n482,
    n247
  );


  buf
  g328
  (
    n428,
    n200
  );


  not
  g329
  (
    n427,
    n154
  );


  not
  g330
  (
    n356,
    n234
  );


  not
  g331
  (
    n340,
    n218
  );


  not
  g332
  (
    n419,
    n318
  );


  buf
  g333
  (
    n387,
    n266
  );


  buf
  g334
  (
    n543,
    n325
  );


  buf
  g335
  (
    n554,
    n79
  );


  not
  g336
  (
    n401,
    n306
  );


  buf
  g337
  (
    n495,
    n296
  );


  not
  g338
  (
    n556,
    n300
  );


  buf
  g339
  (
    n354,
    n222
  );


  not
  g340
  (
    n375,
    n261
  );


  buf
  g341
  (
    n463,
    n294
  );


  not
  g342
  (
    n440,
    n154
  );


  buf
  g343
  (
    n453,
    n301
  );


  not
  g344
  (
    n462,
    n189
  );


  buf
  g345
  (
    n536,
    n291
  );


  not
  g346
  (
    n538,
    n267
  );


  not
  g347
  (
    n565,
    n168
  );


  buf
  g348
  (
    n456,
    n232
  );


  not
  g349
  (
    n540,
    n82
  );


  not
  g350
  (
    n435,
    n298
  );


  not
  g351
  (
    n352,
    n295
  );


  buf
  g352
  (
    n344,
    n277
  );


  buf
  g353
  (
    n521,
    n276
  );


  buf
  g354
  (
    n541,
    n304
  );


  not
  g355
  (
    n572,
    n223
  );


  buf
  g356
  (
    n468,
    n320
  );


  not
  g357
  (
    n331,
    n299
  );


  not
  g358
  (
    n548,
    n260
  );


  not
  g359
  (
    n492,
    n264
  );


  not
  g360
  (
    n535,
    n239
  );


  not
  g361
  (
    n349,
    n296
  );


  not
  g362
  (
    n359,
    n218
  );


  not
  g363
  (
    n389,
    n210
  );


  not
  g364
  (
    n549,
    n188
  );


  buf
  g365
  (
    n564,
    n317
  );


  not
  g366
  (
    n402,
    n246
  );


  not
  g367
  (
    n355,
    n77
  );


  buf
  g368
  (
    n348,
    n214
  );


  not
  g369
  (
    n525,
    n294
  );


  buf
  g370
  (
    n574,
    n204
  );


  buf
  g371
  (
    n496,
    n282
  );


  buf
  g372
  (
    n413,
    n316
  );


  not
  g373
  (
    n534,
    n299
  );


  buf
  g374
  (
    n503,
    n296
  );


  not
  g375
  (
    n467,
    n239
  );


  not
  g376
  (
    n418,
    n209
  );


  buf
  g377
  (
    n371,
    n166
  );


  buf
  g378
  (
    n406,
    n288
  );


  buf
  g379
  (
    n442,
    n177
  );


  not
  g380
  (
    n411,
    n267
  );


  not
  g381
  (
    n542,
    n302
  );


  not
  g382
  (
    n522,
    n272
  );


  buf
  g383
  (
    n444,
    n271
  );


  buf
  g384
  (
    n415,
    n303
  );


  not
  g385
  (
    n514,
    n324
  );


  not
  g386
  (
    n508,
    n277
  );


  not
  g387
  (
    n458,
    n255
  );


  not
  g388
  (
    n491,
    n292
  );


  buf
  g389
  (
    n424,
    n228
  );


  not
  g390
  (
    n373,
    n187
  );


  not
  g391
  (
    n333,
    n195
  );


  not
  g392
  (
    n421,
    n273
  );


  buf
  g393
  (
    n545,
    n325
  );


  buf
  g394
  (
    n550,
    n309
  );


  buf
  g395
  (
    n377,
    n300
  );


  buf
  g396
  (
    n409,
    n78
  );


  buf
  g397
  (
    n489,
    n246
  );


  not
  g398
  (
    n475,
    n207
  );


  not
  g399
  (
    n523,
    n259
  );


  not
  g400
  (
    n396,
    n315
  );


  not
  g401
  (
    n416,
    n298
  );


  not
  g402
  (
    n384,
    n236
  );


  not
  g403
  (
    n392,
    n322
  );


  buf
  g404
  (
    n423,
    n309
  );


  not
  g405
  (
    n484,
    n291
  );


  not
  g406
  (
    n513,
    n221
  );


  buf
  g407
  (
    n461,
    n219
  );


  not
  g408
  (
    n412,
    n193
  );


  buf
  g409
  (
    n343,
    n271
  );


  not
  g410
  (
    n459,
    n165
  );


  not
  g411
  (
    n460,
    n305
  );


  buf
  g412
  (
    n517,
    n170
  );


  not
  g413
  (
    n330,
    n157
  );


  not
  g414
  (
    n366,
    n264
  );


  not
  g415
  (
    n553,
    n268
  );


  not
  g416
  (
    n529,
    n318
  );


  not
  g417
  (
    n378,
    n323
  );


  not
  g418
  (
    n507,
    n81
  );


  not
  g419
  (
    n465,
    n187
  );


  buf
  g420
  (
    n395,
    n160
  );


  buf
  g421
  (
    n334,
    n259
  );


  buf
  g422
  (
    n474,
    n257
  );


  not
  g423
  (
    n557,
    n246
  );


  not
  g424
  (
    n342,
    n269
  );


  buf
  g425
  (
    n382,
    n224
  );


  not
  g426
  (
    n490,
    n194
  );


  buf
  g427
  (
    n341,
    n170
  );


  buf
  g428
  (
    n486,
    n190
  );


  not
  g429
  (
    n500,
    n78
  );


  not
  g430
  (
    n504,
    n242
  );


  buf
  g431
  (
    n501,
    n202
  );


  buf
  g432
  (
    n417,
    n242
  );


  buf
  g433
  (
    n469,
    n310
  );


  not
  g434
  (
    n568,
    n299
  );


  buf
  g435
  (
    n376,
    n198
  );


  not
  g436
  (
    n351,
    n223
  );


  buf
  g437
  (
    n505,
    n240
  );


  not
  g438
  (
    n558,
    n248
  );


  not
  g439
  (
    n403,
    n196
  );


  not
  g440
  (
    n383,
    n311
  );


  not
  g441
  (
    n559,
    n317
  );


  buf
  g442
  (
    n499,
    n272
  );


  not
  g443
  (
    n451,
    n270
  );


  buf
  g444
  (
    n528,
    n286
  );


  xor
  g445
  (
    n436,
    n295,
    n282
  );


  and
  g446
  (
    n502,
    n290,
    n263,
    n302,
    n307
  );


  nand
  g447
  (
    n365,
    n181,
    n153,
    n278,
    n155
  );


  nor
  g448
  (
    n477,
    n83,
    n245,
    n215,
    n180
  );


  and
  g449
  (
    n539,
    n297,
    n283,
    n313,
    n236
  );


  nor
  g450
  (
    n357,
    n277,
    n202,
    n249,
    n78
  );


  nor
  g451
  (
    n480,
    n316,
    n305,
    n297,
    n269
  );


  or
  g452
  (
    n446,
    n208,
    n214,
    n273,
    n321
  );


  or
  g453
  (
    n399,
    n323,
    n285,
    n312,
    n294
  );


  xor
  g454
  (
    n338,
    n283,
    n295,
    n176,
    n196
  );


  nor
  g455
  (
    n404,
    n269,
    n226,
    n186,
    n212
  );


  or
  g456
  (
    n488,
    n288,
    n296,
    n317,
    n251
  );


  or
  g457
  (
    n443,
    n216,
    n324,
    n182,
    n79
  );


  nor
  g458
  (
    n367,
    n321,
    n173,
    n279,
    n250
  );


  xnor
  g459
  (
    n429,
    n260,
    n285,
    n175,
    n259
  );


  or
  g460
  (
    n370,
    n306,
    n181,
    n158,
    n263
  );


  and
  g461
  (
    n431,
    n258,
    n291,
    n203,
    n235
  );


  nand
  g462
  (
    n390,
    n311,
    n219,
    n251,
    n276
  );


  nand
  g463
  (
    n533,
    n247,
    n184,
    n193,
    n228
  );


  or
  g464
  (
    n547,
    n294,
    n284,
    n314,
    n216
  );


  or
  g465
  (
    n524,
    n254,
    n307,
    n268,
    n303
  );


  xor
  g466
  (
    n455,
    n276,
    n178,
    n255,
    n308
  );


  and
  g467
  (
    n509,
    n258,
    n210,
    n261,
    n243
  );


  or
  g468
  (
    n479,
    n270,
    n81,
    n293,
    n302
  );


  and
  g469
  (
    n454,
    n318,
    n317,
    n319,
    n284
  );


  and
  g470
  (
    n407,
    n275,
    n211,
    n174,
    n213
  );


  xnor
  g471
  (
    n364,
    n234,
    n322,
    n199,
    n251
  );


  xor
  g472
  (
    n358,
    n310,
    n323,
    n250,
    n185
  );


  nand
  g473
  (
    n532,
    n229,
    n278,
    n287,
    n163
  );


  nand
  g474
  (
    n493,
    n311,
    n265,
    n263,
    n171
  );


  xnor
  g475
  (
    n449,
    n319,
    n320,
    n162,
    n293
  );


  nor
  g476
  (
    n481,
    n293,
    n309,
    n180,
    n253
  );


  or
  g477
  (
    n437,
    n325,
    n245,
    n237,
    n82
  );


  nor
  g478
  (
    n438,
    n271,
    n287,
    n300,
    n265
  );


  xor
  g479
  (
    n464,
    n278,
    n253,
    n262,
    n306
  );


  and
  g480
  (
    n512,
    n191,
    n291,
    n255,
    n252
  );


  nand
  g481
  (
    n339,
    n184,
    n221,
    n268,
    n204
  );


  and
  g482
  (
    n473,
    n194,
    n78,
    n289,
    n224
  );


  nand
  g483
  (
    n527,
    n307,
    n249,
    n217,
    n175
  );


  nor
  g484
  (
    n494,
    n232,
    n246,
    n308,
    n230
  );


  xor
  g485
  (
    n472,
    n258,
    n325,
    n312,
    n226
  );


  or
  g486
  (
    n398,
    n179,
    n249,
    n188,
    n222
  );


  nor
  g487
  (
    n369,
    n82,
    n273,
    n304,
    n233
  );


  nor
  g488
  (
    n537,
    n192,
    n164,
    n79,
    n283
  );


  nor
  g489
  (
    n381,
    n310,
    n304,
    n270,
    n79
  );


  or
  g490
  (
    n506,
    n281,
    n297,
    n306,
    n282
  );


  or
  g491
  (
    n388,
    n314,
    n285,
    n161,
    n230
  );


  nor
  g492
  (
    n368,
    n295,
    n81,
    n257,
    n270
  );


  xor
  g493
  (
    n569,
    n272,
    n323,
    n250,
    n286
  );


  or
  g494
  (
    n441,
    n261,
    n83,
    n256,
    n299
  );


  and
  g495
  (
    n361,
    n266,
    n280,
    n319,
    n315
  );


  or
  g496
  (
    n497,
    n269,
    n243,
    n183,
    n309
  );


  and
  g497
  (
    n567,
    n217,
    n192,
    n279,
    n247
  );


  and
  g498
  (
    n386,
    n312,
    n254,
    n206,
    n205
  );


  xnor
  g499
  (
    n573,
    n162,
    n205,
    n267,
    n238
  );


  or
  g500
  (
    n466,
    n318,
    n182,
    n215,
    n167
  );


  xor
  g501
  (
    n337,
    n247,
    n157,
    n301,
    n195
  );


  nor
  g502
  (
    n563,
    n253,
    n271,
    n206,
    n283
  );


  nand
  g503
  (
    n531,
    n281,
    n256,
    n166,
    n304
  );


  or
  g504
  (
    n510,
    n158,
    n301,
    n163,
    n197
  );


  or
  g505
  (
    n372,
    n240,
    n264,
    n248,
    n281
  );


  xor
  g506
  (
    n434,
    n263,
    n171,
    n290,
    n314
  );


  xnor
  g507
  (
    n350,
    n298,
    n80,
    n177,
    n268
  );


  or
  g508
  (
    n362,
    n256,
    n179,
    n305,
    n253
  );


  xor
  g509
  (
    n546,
    n77,
    n297,
    n290,
    n316
  );


  and
  g510
  (
    n457,
    n282,
    n261,
    n185,
    n280
  );


  nand
  g511
  (
    n426,
    n190,
    n287,
    n314,
    n264
  );


  or
  g512
  (
    n385,
    n213,
    n267,
    n159,
    n81
  );


  and
  g513
  (
    n478,
    n178,
    n275,
    n249,
    n197
  );


  nor
  g514
  (
    n551,
    n244,
    n324,
    n308,
    n156
  );


  xnor
  g515
  (
    n408,
    n227,
    n259,
    n319,
    n153
  );


  and
  g516
  (
    n335,
    n172,
    n159,
    n280,
    n208
  );


  nor
  g517
  (
    n353,
    n167,
    n200,
    n315,
    n322
  );


  xor
  g518
  (
    n515,
    n279,
    n275,
    n265,
    n284
  );


  or
  g519
  (
    n450,
    n320,
    n252,
    n241,
    n251
  );


  and
  g520
  (
    n380,
    n315,
    n165,
    n161,
    n237
  );


  and
  g521
  (
    n430,
    n198,
    n155,
    n241,
    n245
  );


  or
  g522
  (
    n544,
    n281,
    n209,
    n248,
    n257
  );


  nor
  g523
  (
    n447,
    n320,
    n258,
    n186,
    n248
  );


  nand
  g524
  (
    n346,
    n276,
    n274,
    n289,
    n312
  );


  or
  g525
  (
    n410,
    n176,
    n316,
    n284,
    n254
  );


  nand
  g526
  (
    n470,
    n308,
    n300,
    n288,
    n231
  );


  xor
  g527
  (
    n414,
    n262,
    n156,
    n321,
    n225
  );


  and
  g528
  (
    n432,
    n313,
    n238,
    n273,
    n174
  );


  and
  g529
  (
    n520,
    n292,
    n278,
    n262,
    n287
  );


  xnor
  g530
  (
    n452,
    n289,
    n274,
    n303,
    n201
  );


  nor
  g531
  (
    n530,
    n77,
    n266,
    n301,
    n260
  );


  xor
  g532
  (
    n336,
    n244,
    n83,
    n321,
    n277
  );


  or
  g533
  (
    n360,
    n293,
    n220,
    n280,
    n286
  );


  and
  g534
  (
    n471,
    n311,
    n80,
    n298,
    n229
  );


  xnor
  g535
  (
    n445,
    n289,
    n256,
    n207,
    n250
  );


  or
  g536
  (
    n561,
    n275,
    n272,
    n305,
    n245
  );


  nand
  g537
  (
    n485,
    n173,
    n302,
    n255,
    n80
  );


  nor
  g538
  (
    n566,
    n324,
    n201,
    n260,
    n80
  );


  nand
  g539
  (
    n570,
    n169,
    n225,
    n285,
    n257
  );


  or
  g540
  (
    n332,
    n233,
    n252,
    n172,
    n231
  );


  nor
  g541
  (
    n363,
    n212,
    n211,
    n310,
    n292
  );


  buf
  g542
  (
    n635,
    n360
  );


  buf
  g543
  (
    n584,
    n384
  );


  buf
  g544
  (
    n620,
    n380
  );


  not
  g545
  (
    n631,
    n389
  );


  buf
  g546
  (
    n597,
    n346
  );


  buf
  g547
  (
    n610,
    n377
  );


  not
  g548
  (
    n578,
    n393
  );


  not
  g549
  (
    n608,
    n333
  );


  buf
  g550
  (
    n590,
    n368
  );


  not
  g551
  (
    n607,
    n334
  );


  not
  g552
  (
    n602,
    n379
  );


  buf
  g553
  (
    n595,
    n330
  );


  not
  g554
  (
    n592,
    n371
  );


  buf
  g555
  (
    n589,
    n349
  );


  not
  g556
  (
    n626,
    n359
  );


  not
  g557
  (
    n624,
    n372
  );


  buf
  g558
  (
    n616,
    n373
  );


  not
  g559
  (
    n579,
    n352
  );


  not
  g560
  (
    n600,
    n358
  );


  buf
  g561
  (
    n614,
    n344
  );


  buf
  g562
  (
    n606,
    n388
  );


  not
  g563
  (
    n588,
    n347
  );


  not
  g564
  (
    n605,
    n362
  );


  buf
  g565
  (
    n632,
    n331
  );


  not
  g566
  (
    n638,
    n361
  );


  not
  g567
  (
    n599,
    n375
  );


  buf
  g568
  (
    n612,
    n381
  );


  not
  g569
  (
    n630,
    n338
  );


  not
  g570
  (
    n634,
    n351
  );


  buf
  g571
  (
    n586,
    n365
  );


  not
  g572
  (
    n625,
    n386
  );


  not
  g573
  (
    n576,
    n363
  );


  buf
  g574
  (
    n598,
    n383
  );


  not
  g575
  (
    n617,
    n336
  );


  buf
  g576
  (
    n596,
    n376
  );


  buf
  g577
  (
    n637,
    n355
  );


  buf
  g578
  (
    n583,
    n335
  );


  not
  g579
  (
    n636,
    n369
  );


  not
  g580
  (
    n581,
    n392
  );


  not
  g581
  (
    n613,
    n366
  );


  buf
  g582
  (
    n619,
    n354
  );


  not
  g583
  (
    n627,
    n345
  );


  buf
  g584
  (
    n615,
    n337
  );


  buf
  g585
  (
    n580,
    n356
  );


  buf
  g586
  (
    n601,
    n350
  );


  buf
  g587
  (
    n633,
    n348
  );


  not
  g588
  (
    n594,
    n364
  );


  buf
  g589
  (
    n593,
    n339
  );


  buf
  g590
  (
    n621,
    n341
  );


  not
  g591
  (
    n587,
    n374
  );


  not
  g592
  (
    n628,
    n343
  );


  buf
  g593
  (
    n577,
    n370
  );


  buf
  g594
  (
    n591,
    n357
  );


  buf
  g595
  (
    n604,
    n387
  );


  not
  g596
  (
    n575,
    n340
  );


  buf
  g597
  (
    n618,
    n353
  );


  buf
  g598
  (
    n609,
    n378
  );


  buf
  g599
  (
    n603,
    n391
  );


  buf
  g600
  (
    n611,
    n390
  );


  buf
  g601
  (
    n582,
    n382
  );


  not
  g602
  (
    n585,
    n342
  );


  buf
  g603
  (
    n622,
    n367
  );


  not
  g604
  (
    n629,
    n385
  );


  buf
  g605
  (
    n623,
    n332
  );


  or
  g606
  (
    n643,
    n469,
    n584
  );


  and
  g607
  (
    n662,
    n467,
    n406,
    n499,
    n416
  );


  xor
  g608
  (
    n677,
    n577,
    n585,
    n578,
    n441
  );


  xor
  g609
  (
    n651,
    n517,
    n408,
    n581,
    n491
  );


  or
  g610
  (
    n676,
    n493,
    n395,
    n494,
    n409
  );


  xor
  g611
  (
    n639,
    n421,
    n453,
    n470,
    n579
  );


  nand
  g612
  (
    n647,
    n457,
    n412,
    n446,
    n497
  );


  and
  g613
  (
    n640,
    n584,
    n437,
    n580,
    n521
  );


  xnor
  g614
  (
    n660,
    n503,
    n581,
    n508,
    n468
  );


  xor
  g615
  (
    n671,
    n501,
    n496,
    n460,
    n576
  );


  and
  g616
  (
    n667,
    n450,
    n403,
    n415,
    n397
  );


  and
  g617
  (
    n670,
    n523,
    n433,
    n476,
    n413
  );


  nor
  g618
  (
    n658,
    n514,
    n522,
    n473,
    n455
  );


  xor
  g619
  (
    n650,
    n502,
    n480,
    n579,
    n581
  );


  or
  g620
  (
    n661,
    n575,
    n513,
    n492,
    n444
  );


  or
  g621
  (
    n656,
    n472,
    n509,
    n580,
    n479
  );


  nand
  g622
  (
    n675,
    n424,
    n405,
    n442,
    n581
  );


  nor
  g623
  (
    n668,
    n586,
    n434,
    n454,
    n578
  );


  and
  g624
  (
    n665,
    n448,
    n486,
    n582,
    n427
  );


  xnor
  g625
  (
    n646,
    n440,
    n422,
    n520,
    n585
  );


  xor
  g626
  (
    n681,
    n498,
    n584,
    n426,
    n474
  );


  xor
  g627
  (
    n652,
    n483,
    n585,
    n582,
    n402
  );


  nand
  g628
  (
    n655,
    n583,
    n425,
    n580,
    n459
  );


  nand
  g629
  (
    n679,
    n414,
    n515,
    n394,
    n429
  );


  xnor
  g630
  (
    n644,
    n586,
    n464,
    n435,
    n452
  );


  nor
  g631
  (
    n678,
    n505,
    n458,
    n439,
    n478
  );


  nand
  g632
  (
    n663,
    n461,
    n506,
    n485,
    n579
  );


  nor
  g633
  (
    n674,
    n420,
    n451,
    n575,
    n510
  );


  or
  g634
  (
    n664,
    n576,
    n511,
    n518,
    n577
  );


  xnor
  g635
  (
    n645,
    n585,
    n430,
    n436,
    n431
  );


  xnor
  g636
  (
    n654,
    n418,
    n404,
    n399,
    n456
  );


  nand
  g637
  (
    n682,
    n417,
    n583,
    n481,
    n423
  );


  and
  g638
  (
    n669,
    n471,
    n487,
    n443,
    n578
  );


  xnor
  g639
  (
    n672,
    n577,
    n512,
    n576,
    n438
  );


  or
  g640
  (
    n680,
    n407,
    n462,
    n584,
    n477
  );


  nand
  g641
  (
    n659,
    n504,
    n400,
    n580,
    n583
  );


  nor
  g642
  (
    n653,
    n495,
    n582,
    n445,
    n432
  );


  or
  g643
  (
    n649,
    n419,
    n447,
    n582,
    n583
  );


  nand
  g644
  (
    n642,
    n484,
    n475,
    n579,
    n428
  );


  and
  g645
  (
    n666,
    n488,
    n578,
    n482,
    n489
  );


  nor
  g646
  (
    n648,
    n396,
    n500,
    n516,
    n465
  );


  nand
  g647
  (
    n657,
    n519,
    n449,
    n401,
    n411
  );


  xor
  g648
  (
    n673,
    n463,
    n466,
    n507,
    n490
  );


  xnor
  g649
  (
    n641,
    n575,
    n410,
    n398,
    n577
  );


  xnor
  g650
  (
    n693,
    n629,
    n621,
    n627,
    n607
  );


  xnor
  g651
  (
    n690,
    n88,
    n588,
    n631,
    n93
  );


  nor
  g652
  (
    n725,
    n587,
    n603,
    n681,
    n628
  );


  xor
  g653
  (
    n685,
    n657,
    n624,
    n609,
    n663
  );


  nor
  g654
  (
    n747,
    n670,
    n587,
    n88,
    n86
  );


  or
  g655
  (
    n717,
    n596,
    n613,
    n622,
    n611
  );


  and
  g656
  (
    n754,
    n525,
    n617,
    n603,
    n622
  );


  and
  g657
  (
    n759,
    n605,
    n637,
    n675,
    n594
  );


  xor
  g658
  (
    n756,
    n604,
    n96,
    n631,
    n635
  );


  or
  g659
  (
    n692,
    n604,
    n593,
    n587,
    n616
  );


  xnor
  g660
  (
    n694,
    n592,
    n594,
    n85
  );


  nand
  g661
  (
    n689,
    n606,
    n679,
    n603,
    n93
  );


  and
  g662
  (
    n684,
    n644,
    n653,
    n595,
    n651
  );


  nand
  g663
  (
    n738,
    n598,
    n93,
    n607,
    n591
  );


  or
  g664
  (
    n696,
    n606,
    n591,
    n94,
    n587
  );


  nand
  g665
  (
    n723,
    n592,
    n643,
    n636,
    n590
  );


  xnor
  g666
  (
    n757,
    n619,
    n615,
    n654,
    n86
  );


  xnor
  g667
  (
    n760,
    n660,
    n590,
    n602,
    n623
  );


  or
  g668
  (
    n710,
    n593,
    n629,
    n661,
    n588
  );


  nor
  g669
  (
    n709,
    n93,
    n91,
    n597
  );


  nor
  g670
  (
    n708,
    n679,
    n92,
    n88,
    n610
  );


  and
  g671
  (
    n722,
    n660,
    n634,
    n90,
    n627
  );


  and
  g672
  (
    n711,
    n599,
    n624,
    n597,
    n623
  );


  or
  g673
  (
    n700,
    n662,
    n597,
    n97,
    n589
  );


  nor
  g674
  (
    n719,
    n671,
    n681,
    n632,
    n611
  );


  xnor
  g675
  (
    n765,
    n674,
    n640,
    n614,
    n88
  );


  nand
  g676
  (
    n727,
    n649,
    n601,
    n592,
    n607
  );


  xor
  g677
  (
    n745,
    n594,
    n618,
    n605
  );


  and
  g678
  (
    n713,
    n608,
    n600,
    n603,
    n590
  );


  nor
  g679
  (
    n712,
    n608,
    n621,
    n596,
    n84
  );


  xnor
  g680
  (
    n720,
    n592,
    n90,
    n658,
    n87
  );


  nand
  g681
  (
    n763,
    n616,
    n624,
    n595,
    n610
  );


  xnor
  g682
  (
    n751,
    n677,
    n90,
    n675,
    n602
  );


  or
  g683
  (
    n715,
    n682,
    n84,
    n646,
    n680
  );


  nor
  g684
  (
    n691,
    n613,
    n666,
    n655,
    n625
  );


  or
  g685
  (
    n770,
    n640,
    n662,
    n86,
    n621
  );


  and
  g686
  (
    n766,
    n89,
    n614,
    n672,
    n616
  );


  xnor
  g687
  (
    n737,
    n664,
    n87,
    n639,
    n629
  );


  and
  g688
  (
    n698,
    n665,
    n615,
    n668,
    n651
  );


  nor
  g689
  (
    n743,
    n586,
    n635,
    n598,
    n605
  );


  xnor
  g690
  (
    n721,
    n666,
    n682,
    n627,
    n626
  );


  and
  g691
  (
    n686,
    n669,
    n671,
    n524,
    n599
  );


  or
  g692
  (
    n697,
    n604,
    n596,
    n622,
    n94
  );


  nand
  g693
  (
    n705,
    n602,
    n673,
    n664,
    n649
  );


  or
  g694
  (
    n687,
    n613,
    n634,
    n657,
    n648
  );


  and
  g695
  (
    n731,
    n620,
    n627,
    n631,
    n594
  );


  xnor
  g696
  (
    n706,
    n614,
    n623,
    n631,
    n630
  );


  xnor
  g697
  (
    n724,
    n605,
    n680,
    n616,
    n619
  );


  xor
  g698
  (
    n702,
    n85,
    n95,
    n87,
    n633
  );


  nor
  g699
  (
    n740,
    n635,
    n91,
    n673,
    n90
  );


  xor
  g700
  (
    n703,
    n621,
    n644,
    n628,
    n611
  );


  nand
  g701
  (
    n750,
    n632,
    n614,
    n647,
    n600
  );


  nand
  g702
  (
    n729,
    n95,
    n628,
    n647,
    n615
  );


  or
  g703
  (
    n758,
    n637,
    n593,
    n591,
    n588
  );


  nand
  g704
  (
    n714,
    n643,
    n609,
    n650,
    n639
  );


  nand
  g705
  (
    n716,
    n630,
    n674,
    n611,
    n89
  );


  xor
  g706
  (
    n739,
    n648,
    n658,
    n94,
    n625
  );


  xnor
  g707
  (
    n707,
    n628,
    n676,
    n608,
    n597
  );


  and
  g708
  (
    n768,
    n615,
    n610,
    n677,
    n618
  );


  nand
  g709
  (
    n683,
    n642,
    n91,
    n676,
    n89
  );


  and
  g710
  (
    n762,
    n604,
    n656,
    n601,
    n620
  );


  nor
  g711
  (
    n755,
    n590,
    n617,
    n596,
    n645
  );


  xor
  g712
  (
    n733,
    n595,
    n625,
    n600,
    n652
  );


  and
  g713
  (
    n732,
    n618,
    n667,
    n665,
    n642
  );


  xor
  g714
  (
    n726,
    n85,
    n96,
    n669,
    n617
  );


  xor
  g715
  (
    n704,
    n613,
    n632,
    n593,
    n620
  );


  or
  g716
  (
    n753,
    n622,
    n624,
    n84,
    n87
  );


  nand
  g717
  (
    n748,
    n600,
    n650,
    n92,
    n653
  );


  nor
  g718
  (
    n695,
    n89,
    n645,
    n670,
    n598
  );


  or
  g719
  (
    n761,
    n608,
    n678,
    n652,
    n667
  );


  and
  g720
  (
    n746,
    n94,
    n96,
    n609,
    n655
  );


  and
  g721
  (
    n764,
    n599,
    n626,
    n659,
    n617
  );


  nand
  g722
  (
    n742,
    n610,
    n663,
    n620,
    n601
  );


  and
  g723
  (
    n718,
    n634,
    n635,
    n612,
    n591
  );


  xor
  g724
  (
    n688,
    n606,
    n661,
    n612,
    n630
  );


  nand
  g725
  (
    n730,
    n659,
    n589,
    n92,
    n602
  );


  nor
  g726
  (
    n734,
    n95,
    n84,
    n619,
    n641
  );


  or
  g727
  (
    n741,
    n633,
    n601,
    n632,
    n612
  );


  nand
  g728
  (
    n767,
    n625,
    n656,
    n86,
    n646
  );


  xnor
  g729
  (
    n744,
    n678,
    n641,
    n607,
    n634
  );


  xor
  g730
  (
    n728,
    n629,
    n619,
    n96,
    n83
  );


  or
  g731
  (
    n769,
    n95,
    n92,
    n588,
    n595
  );


  xor
  g732
  (
    n699,
    n626,
    n589,
    n668,
    n609
  );


  or
  g733
  (
    n736,
    n636,
    n598,
    n599,
    n672
  );


  xnor
  g734
  (
    n752,
    n589,
    n633,
    n637
  );


  or
  g735
  (
    n749,
    n606,
    n626,
    n97,
    n612
  );


  xnor
  g736
  (
    n701,
    n636,
    n586,
    n633,
    n630
  );


  xnor
  g737
  (
    n735,
    n623,
    n97,
    n654,
    n636
  );


  and
  g738
  (
    n849,
    n720,
    n735,
    n756,
    n721
  );


  xnor
  g739
  (
    n773,
    n124,
    n739,
    n106,
    n756
  );


  and
  g740
  (
    n861,
    n733,
    n108,
    n140,
    n750
  );


  nand
  g741
  (
    n800,
    n138,
    n754,
    n740,
    n103
  );


  xnor
  g742
  (
    n822,
    n707,
    n730,
    n755,
    n749
  );


  xnor
  g743
  (
    n825,
    n121,
    n140,
    n128,
    n722
  );


  nor
  g744
  (
    n821,
    n692,
    n105,
    n757,
    n117
  );


  xnor
  g745
  (
    n791,
    n101,
    n709,
    n737,
    n722
  );


  xor
  g746
  (
    n854,
    n715,
    n98,
    n104,
    n118
  );


  or
  g747
  (
    n788,
    n683,
    n107,
    n726,
    n757
  );


  and
  g748
  (
    n840,
    n120,
    n693,
    n140,
    n133
  );


  xor
  g749
  (
    n864,
    n704,
    n749,
    n119,
    n103
  );


  or
  g750
  (
    n806,
    n705,
    n121,
    n130,
    n748
  );


  xor
  g751
  (
    n789,
    n103,
    n106,
    n132,
    n700
  );


  and
  g752
  (
    n792,
    n704,
    n145,
    n111,
    n703
  );


  nor
  g753
  (
    n834,
    n119,
    n735,
    n716,
    n743
  );


  and
  g754
  (
    n809,
    n123,
    n762,
    n711,
    n769
  );


  xnor
  g755
  (
    n829,
    n752,
    n762,
    n694,
    n120
  );


  and
  g756
  (
    n855,
    n110,
    n738,
    n142,
    n766
  );


  xor
  g757
  (
    n823,
    n114,
    n683,
    n142,
    n689
  );


  nor
  g758
  (
    n814,
    n133,
    n746,
    n144,
    n103
  );


  xor
  g759
  (
    n799,
    n131,
    n709,
    n729,
    n759
  );


  and
  g760
  (
    n803,
    n730,
    n765,
    n713,
    n685
  );


  or
  g761
  (
    n815,
    n134,
    n133,
    n110,
    n144
  );


  xor
  g762
  (
    n862,
    n747,
    n723,
    n99,
    n126
  );


  xor
  g763
  (
    n782,
    n723,
    n718,
    n748,
    n125
  );


  and
  g764
  (
    n816,
    n100,
    n135,
    n766,
    n687
  );


  xor
  g765
  (
    n836,
    n131,
    n144,
    n696,
    n684
  );


  and
  g766
  (
    n824,
    n695,
    n143,
    n741
  );


  xor
  g767
  (
    n796,
    n770,
    n761,
    n727,
    n714
  );


  xor
  g768
  (
    n798,
    n684,
    n768,
    n132,
    n114
  );


  xor
  g769
  (
    n801,
    n108,
    n726,
    n146,
    n757
  );


  xor
  g770
  (
    n843,
    n690,
    n736,
    n105,
    n145
  );


  xnor
  g771
  (
    n784,
    n689,
    n692,
    n98,
    n115
  );


  and
  g772
  (
    n802,
    n764,
    n99,
    n751,
    n118
  );


  nor
  g773
  (
    n812,
    n135,
    n128,
    n143,
    n132
  );


  or
  g774
  (
    n851,
    n715,
    n751,
    n97,
    n755
  );


  nor
  g775
  (
    n804,
    n729,
    n113,
    n765,
    n731
  );


  xor
  g776
  (
    n847,
    n740,
    n117,
    n697,
    n758
  );


  or
  g777
  (
    n790,
    n123,
    n731,
    n145,
    n702
  );


  or
  g778
  (
    n805,
    n104,
    n750,
    n130,
    n121
  );


  or
  g779
  (
    n837,
    n767,
    n121,
    n763
  );


  nand
  g780
  (
    n839,
    n697,
    n770,
    n129,
    n139
  );


  nor
  g781
  (
    n841,
    n714,
    n125,
    n713,
    n129
  );


  or
  g782
  (
    n863,
    n701,
    n768,
    n116,
    n98
  );


  and
  g783
  (
    n771,
    n109,
    n753,
    n754,
    n744
  );


  nor
  g784
  (
    n781,
    n100,
    n105,
    n762,
    n131
  );


  xor
  g785
  (
    n830,
    n759,
    n760,
    n104,
    n758
  );


  nor
  g786
  (
    n795,
    n142,
    n686,
    n102,
    n756
  );


  nand
  g787
  (
    n844,
    n702,
    n769,
    n742,
    n112
  );


  or
  g788
  (
    n860,
    n101,
    n712,
    n741,
    n761
  );


  or
  g789
  (
    n820,
    n122,
    n701,
    n111,
    n127
  );


  or
  g790
  (
    n777,
    n750,
    n109,
    n703,
    n717
  );


  xnor
  g791
  (
    n867,
    n752,
    n136,
    n127,
    n690
  );


  nor
  g792
  (
    n794,
    n101,
    n767,
    n128,
    n122
  );


  xor
  g793
  (
    n865,
    n119,
    n124,
    n753,
    n734
  );


  xor
  g794
  (
    n858,
    n685,
    n122,
    n746,
    n753
  );


  nor
  g795
  (
    n783,
    n707,
    n698,
    n114,
    n691
  );


  nand
  g796
  (
    n866,
    n137,
    n136,
    n724,
    n130
  );


  and
  g797
  (
    n852,
    n134,
    n124,
    n705,
    n107
  );


  or
  g798
  (
    n832,
    n108,
    n770,
    n110,
    n112
  );


  xor
  g799
  (
    n828,
    n126,
    n135,
    n109,
    n100
  );


  nor
  g800
  (
    n817,
    n719,
    n141,
    n105,
    n694
  );


  nor
  g801
  (
    n835,
    n126,
    n687,
    n717,
    n99
  );


  and
  g802
  (
    n780,
    n113,
    n139,
    n131,
    n695
  );


  xnor
  g803
  (
    n786,
    n123,
    n732,
    n725,
    n126
  );


  nand
  g804
  (
    n811,
    n127,
    n768,
    n102,
    n112
  );


  nor
  g805
  (
    n859,
    n754,
    n696,
    n738,
    n708
  );


  or
  g806
  (
    n838,
    n130,
    n111,
    n109
  );


  nor
  g807
  (
    n797,
    n767,
    n120,
    n133,
    n747
  );


  xnor
  g808
  (
    n857,
    n129,
    n108,
    n132,
    n102
  );


  and
  g809
  (
    n776,
    n765,
    n710,
    n693,
    n739
  );


  xnor
  g810
  (
    n833,
    n728,
    n724,
    n118,
    n113
  );


  nor
  g811
  (
    n842,
    n137,
    n107,
    n706,
    n699
  );


  nor
  g812
  (
    n810,
    n769,
    n140,
    n137,
    n764
  );


  and
  g813
  (
    n819,
    n708,
    n110,
    n101,
    n760
  );


  nor
  g814
  (
    n779,
    n755,
    n141,
    n142,
    n734
  );


  nor
  g815
  (
    n807,
    n124,
    n115,
    n135,
    n112
  );


  nor
  g816
  (
    n827,
    n706,
    n116,
    n691,
    n136
  );


  or
  g817
  (
    n785,
    n733,
    n764,
    n727,
    n106
  );


  and
  g818
  (
    n774,
    n99,
    n766,
    n123,
    n719
  );


  xor
  g819
  (
    n787,
    n710,
    n125,
    n744,
    n698
  );


  xnor
  g820
  (
    n775,
    n146,
    n138,
    n117,
    n120
  );


  or
  g821
  (
    n831,
    n114,
    n116,
    n134,
    n145
  );


  nand
  g822
  (
    n818,
    n721,
    n115,
    n116,
    n104
  );


  or
  g823
  (
    n772,
    n737,
    n712,
    n763,
    n761
  );


  or
  g824
  (
    n868,
    n751,
    n138,
    n127,
    n102
  );


  or
  g825
  (
    n850,
    n143,
    n128,
    n745,
    n139
  );


  nand
  g826
  (
    n845,
    n758,
    n736,
    n106,
    n699
  );


  nor
  g827
  (
    n808,
    n141,
    n688,
    n686,
    n752
  );


  and
  g828
  (
    n793,
    n98,
    n136,
    n100,
    n759
  );


  nor
  g829
  (
    n846,
    n745,
    n134,
    n688,
    n760
  );


  xnor
  g830
  (
    n856,
    n138,
    n139,
    n725,
    n144
  );


  and
  g831
  (
    n778,
    n742,
    n129,
    n118,
    n107
  );


  xor
  g832
  (
    n853,
    n117,
    n720,
    n728,
    n732
  );


  xnor
  g833
  (
    n848,
    n716,
    n125,
    n113,
    n137
  );


  xor
  g834
  (
    n826,
    n115,
    n141,
    n122,
    n743
  );


  nor
  g835
  (
    n813,
    n718,
    n711,
    n700,
    n119
  );


  buf
  g836
  (
    n878,
    n816
  );


  buf
  g837
  (
    n887,
    n821
  );


  not
  g838
  (
    n884,
    n781
  );


  not
  g839
  (
    n879,
    n771
  );


  buf
  g840
  (
    n896,
    n812
  );


  not
  g841
  (
    n882,
    n845
  );


  nand
  g842
  (
    n892,
    n789,
    n834
  );


  and
  g843
  (
    n886,
    n798,
    n783,
    n785
  );


  nor
  g844
  (
    n885,
    n833,
    n807,
    n830
  );


  nand
  g845
  (
    n895,
    n844,
    n815,
    n786
  );


  and
  g846
  (
    n899,
    n776,
    n843,
    n838
  );


  and
  g847
  (
    n893,
    n823,
    n809,
    n795
  );


  xor
  g848
  (
    n874,
    n841,
    n832,
    n819
  );


  or
  g849
  (
    n880,
    n835,
    n784,
    n808
  );


  or
  g850
  (
    n877,
    n849,
    n790,
    n846
  );


  or
  g851
  (
    n870,
    n824,
    n774,
    n836
  );


  nand
  g852
  (
    n890,
    n829,
    n817,
    n788
  );


  nor
  g853
  (
    n871,
    n782,
    n794,
    n837
  );


  xor
  g854
  (
    n875,
    n803,
    n806,
    n822
  );


  and
  g855
  (
    n891,
    n802,
    n792,
    n825
  );


  xnor
  g856
  (
    n883,
    n775,
    n791,
    n813
  );


  nand
  g857
  (
    n888,
    n811,
    n820,
    n800
  );


  or
  g858
  (
    n869,
    n810,
    n827,
    n840
  );


  xnor
  g859
  (
    n881,
    n772,
    n826,
    n793
  );


  or
  g860
  (
    n898,
    n778,
    n796,
    n805
  );


  nand
  g861
  (
    n876,
    n799,
    n847,
    n839
  );


  or
  g862
  (
    n894,
    n801,
    n842,
    n797
  );


  nand
  g863
  (
    n889,
    n831,
    n787,
    n804
  );


  or
  g864
  (
    n872,
    n773,
    n818,
    n828
  );


  nand
  g865
  (
    n897,
    n850,
    n814,
    n780
  );


  or
  g866
  (
    n873,
    n779,
    n777,
    n848
  );


  not
  g867
  (
    n926,
    n534
  );


  not
  g868
  (
    n916,
    n563
  );


  buf
  g869
  (
    n919,
    n537
  );


  buf
  g870
  (
    n924,
    n874
  );


  or
  g871
  (
    n901,
    n875,
    n874
  );


  nand
  g872
  (
    n911,
    n558,
    n549,
    n876
  );


  xor
  g873
  (
    n928,
    n556,
    n540,
    n560,
    n527
  );


  xnor
  g874
  (
    n922,
    n552,
    n535,
    n871
  );


  nor
  g875
  (
    n909,
    n872,
    n562,
    n877,
    n873
  );


  xnor
  g876
  (
    n927,
    n876,
    n528,
    n547,
    n533
  );


  nor
  g877
  (
    n920,
    n872,
    n872,
    n551,
    n545
  );


  nand
  g878
  (
    n915,
    n877,
    n877,
    n557,
    n560
  );


  xor
  g879
  (
    n929,
    n878,
    n536,
    n877,
    n561
  );


  nand
  g880
  (
    n900,
    n547,
    n564,
    n542,
    n875
  );


  or
  g881
  (
    n910,
    n536,
    n878,
    n546,
    n540
  );


  and
  g882
  (
    n925,
    n550,
    n875,
    n873,
    n871
  );


  xnor
  g883
  (
    n921,
    n870,
    n869,
    n533,
    n553
  );


  nand
  g884
  (
    n914,
    n874,
    n556,
    n550,
    n554
  );


  xor
  g885
  (
    n907,
    n544,
    n538,
    n548,
    n534
  );


  and
  g886
  (
    n903,
    n554,
    n555,
    n875,
    n537
  );


  nor
  g887
  (
    n904,
    n553,
    n543,
    n546,
    n530
  );


  nand
  g888
  (
    n906,
    n543,
    n538,
    n870
  );


  nand
  g889
  (
    n902,
    n545,
    n869,
    n871,
    n559
  );


  nand
  g890
  (
    n913,
    n562,
    n539,
    n549
  );


  xnor
  g891
  (
    n908,
    n872,
    n558,
    n557,
    n559
  );


  xor
  g892
  (
    n912,
    n870,
    n873,
    n561,
    n876
  );


  nor
  g893
  (
    n905,
    n542,
    n548,
    n544,
    n529
  );


  xnor
  g894
  (
    n923,
    n532,
    n552,
    n871,
    n551
  );


  and
  g895
  (
    n917,
    n541,
    n555,
    n563,
    n526
  );


  nor
  g896
  (
    n918,
    n873,
    n531,
    n874,
    n541
  );


  and
  g897
  (
    n937,
    n896,
    n892,
    n908
  );


  or
  g898
  (
    n946,
    n882,
    n893,
    n884
  );


  xor
  g899
  (
    n931,
    n895,
    n919,
    n906,
    n917
  );


  nand
  g900
  (
    n935,
    n881,
    n897,
    n879
  );


  nor
  g901
  (
    n955,
    n883,
    n925,
    n886,
    n920
  );


  or
  g902
  (
    n934,
    n891,
    n915,
    n884,
    n898
  );


  nor
  g903
  (
    n939,
    n912,
    n896,
    n905
  );


  xor
  g904
  (
    n938,
    n894,
    n897,
    n890
  );


  xor
  g905
  (
    n930,
    n889,
    n893,
    n926,
    n887
  );


  nand
  g906
  (
    n945,
    n888,
    n911,
    n887,
    n890
  );


  xnor
  g907
  (
    n957,
    n898,
    n891,
    n893,
    n887
  );


  xor
  g908
  (
    n952,
    n904,
    n903,
    n881,
    n922
  );


  and
  g909
  (
    n949,
    n880,
    n890,
    n900,
    n894
  );


  xor
  g910
  (
    n951,
    n882,
    n879,
    n902,
    n884
  );


  xnor
  g911
  (
    n942,
    n878,
    n885,
    n881,
    n910
  );


  and
  g912
  (
    n940,
    n909,
    n884,
    n888,
    n881
  );


  and
  g913
  (
    n941,
    n880,
    n898,
    n887,
    n899
  );


  nand
  g914
  (
    n953,
    n886,
    n878,
    n899,
    n885
  );


  nand
  g915
  (
    n936,
    n892,
    n927,
    n897,
    n889
  );


  nand
  g916
  (
    n947,
    n895,
    n883,
    n898,
    n888
  );


  and
  g917
  (
    n950,
    n901,
    n883,
    n907,
    n914
  );


  nand
  g918
  (
    n948,
    n880,
    n894,
    n921,
    n886
  );


  xor
  g919
  (
    n933,
    n879,
    n883,
    n889,
    n888
  );


  xnor
  g920
  (
    n944,
    n924,
    n880,
    n923,
    n885
  );


  nand
  g921
  (
    n956,
    n894,
    n916,
    n882,
    n886
  );


  xor
  g922
  (
    n932,
    n891,
    n913,
    n896,
    n889
  );


  nor
  g923
  (
    n954,
    n885,
    n895,
    n918
  );


  xor
  g924
  (
    n943,
    n892,
    n891,
    n882,
    n890
  );


  buf
  g925
  (
    n978,
    n32
  );


  buf
  g926
  (
    n958,
    n328
  );


  not
  g927
  (
    n967,
    n929
  );


  buf
  g928
  (
    n969,
    n148
  );


  buf
  g929
  (
    n964,
    n942
  );


  buf
  g930
  (
    n972,
    n933
  );


  buf
  g931
  (
    n979,
    n329
  );


  buf
  g932
  (
    n984,
    n329
  );


  buf
  g933
  (
    n966,
    n566
  );


  buf
  g934
  (
    n973,
    n936
  );


  buf
  g935
  (
    n975,
    n326
  );


  not
  g936
  (
    n959,
    n928
  );


  nand
  g937
  (
    n976,
    n32,
    n147,
    n940,
    n567
  );


  xnor
  g938
  (
    n981,
    n944,
    n954,
    n949,
    n568
  );


  or
  g939
  (
    n971,
    n327,
    n570,
    n569,
    n957
  );


  or
  g940
  (
    n983,
    n326,
    n932,
    n328,
    n568
  );


  or
  g941
  (
    n962,
    n148,
    n931,
    n947,
    n570
  );


  nand
  g942
  (
    n980,
    n572,
    n950,
    n957,
    n945
  );


  and
  g943
  (
    n982,
    n930,
    n326,
    n147
  );


  nor
  g944
  (
    n965,
    n327,
    n328,
    n571,
    n565
  );


  xor
  g945
  (
    n970,
    n569,
    n327,
    n934,
    n938
  );


  xnor
  g946
  (
    n977,
    n943,
    n147,
    n939,
    n927
  );


  or
  g947
  (
    n985,
    n929,
    n146,
    n564
  );


  nand
  g948
  (
    n963,
    n948,
    n956,
    n327,
    n851
  );


  nor
  g949
  (
    n986,
    n937,
    n329,
    n566,
    n953
  );


  or
  g950
  (
    n974,
    n565,
    n571,
    n32,
    n328
  );


  nand
  g951
  (
    n968,
    n946,
    n32,
    n951,
    n928
  );


  and
  g952
  (
    n960,
    n147,
    n567,
    n935,
    n952
  );


  xnor
  g953
  (
    n961,
    n329,
    n955,
    n941,
    n31
  );


  xnor
  g954
  (
    n993,
    n149,
    n974,
    n982,
    n980
  );


  xnor
  g955
  (
    n995,
    n150,
    n150,
    n972,
    n966
  );


  and
  g956
  (
    n1011,
    n976,
    n976,
    n979,
    n983
  );


  or
  g957
  (
    n1003,
    n970,
    n151,
    n961,
    n959
  );


  xnor
  g958
  (
    n1018,
    n985,
    n960,
    n979,
    n965
  );


  xor
  g959
  (
    n1006,
    n984,
    n148,
    n968,
    n151
  );


  and
  g960
  (
    n1005,
    n983,
    n971,
    n977,
    n980
  );


  or
  g961
  (
    n1004,
    n964,
    n978,
    n573,
    n965
  );


  xnor
  g962
  (
    n1010,
    n958,
    n981,
    n971,
    n974
  );


  nor
  g963
  (
    n999,
    n972,
    n971,
    n961,
    n964
  );


  xnor
  g964
  (
    n997,
    n978,
    n982,
    n974,
    n852
  );


  and
  g965
  (
    n1016,
    n973,
    n985,
    n983,
    n969
  );


  xnor
  g966
  (
    n1008,
    n973,
    n981,
    n977,
    n980
  );


  and
  g967
  (
    n992,
    n965,
    n958,
    n969,
    n964
  );


  and
  g968
  (
    n991,
    n974,
    n149,
    n975,
    n960
  );


  xnor
  g969
  (
    n1020,
    n964,
    n959,
    n152,
    n961
  );


  nor
  g970
  (
    n1013,
    n572,
    n573,
    n971,
    n960
  );


  nand
  g971
  (
    n990,
    n968,
    n958,
    n970,
    n980
  );


  and
  g972
  (
    n1012,
    n970,
    n961,
    n149,
    n152
  );


  xor
  g973
  (
    n994,
    n976,
    n982,
    n963
  );


  nor
  g974
  (
    n1014,
    n981,
    n977,
    n976,
    n966
  );


  xnor
  g975
  (
    n989,
    n959,
    n985,
    n969
  );


  nand
  g976
  (
    n1000,
    n962,
    n978,
    n152,
    n975
  );


  nor
  g977
  (
    n1017,
    n966,
    n977,
    n149,
    n968
  );


  xnor
  g978
  (
    n1009,
    n981,
    n150,
    n984,
    n962
  );


  nand
  g979
  (
    n1007,
    n963,
    n968,
    n967,
    n972
  );


  nand
  g980
  (
    n1015,
    n962,
    n967,
    n152,
    n969
  );


  xnor
  g981
  (
    n1019,
    n975,
    n962,
    n963,
    n979
  );


  xnor
  g982
  (
    n1001,
    n150,
    n983,
    n973,
    n574
  );


  nor
  g983
  (
    AntiSAT_key_wire,
    n986,
    n967,
    n970,
    n973
  );


  or
  g984
  (
    n1002,
    n984,
    n967,
    n151,
    n965
  );


  or
  g985
  (
    n987,
    n984,
    n151,
    n972,
    n978
  );


  xnor
  g986
  (
    n996,
    n958,
    n975,
    n959,
    n960
  );


  xor
  g987
  (
    n988,
    n982,
    n966,
    n148,
    n979
  );


  xnor
  g988
  (
    n1027,
    n854,
    n1018,
    n986,
    n1019
  );


  xor
  g989
  (
    n1026,
    n861,
    n1016,
    n856,
    n860
  );


  nand
  g990
  (
    n1022,
    n1014,
    n867,
    n868,
    n857
  );


  nor
  g991
  (
    n1025,
    n864,
    n899,
    n866,
    n859
  );


  and
  g992
  (
    n1023,
    n1015,
    n858,
    n863,
    n862
  );


  xor
  g993
  (
    n1021,
    n853,
    n1020,
    n865,
    n855
  );


  nand
  g994
  (
    n1024,
    n1017,
    n986,
    n899
  );


  buf
  g995
  (
    n1030,
    n574
  );


  not
  g996
  (
    n1028,
    n1025
  );


  nand
  g997
  (
    n1029,
    n1024,
    n1026
  );


  and
  g998
  (
    n1032,
    n1027,
    n1028,
    n638
  );


  xnor
  g999
  (
    n1031,
    n1029,
    n638,
    n1030
  );


  xor
  KeyPIGate_0_0
  (
    g_input_0_0,
    keyIn_0_0,
    n1
  );


  xor
  KeyPIGate_0_32
  (
    gbar_input_0_0,
    keyIn_0_32,
    n1
  );


  xor
  KeyPIGate_0_1
  (
    g_input_0_1,
    keyIn_0_1,
    n2
  );


  xor
  KeyPIGate_0_33
  (
    gbar_input_0_1,
    keyIn_0_33,
    n2
  );


  xor
  KeyPIGate_0_2
  (
    g_input_0_2,
    keyIn_0_2,
    n3
  );


  xor
  KeyPIGate_0_34
  (
    gbar_input_0_2,
    keyIn_0_34,
    n3
  );


  xor
  KeyPIGate_0_3
  (
    g_input_0_3,
    keyIn_0_3,
    n4
  );


  xor
  KeyPIGate_0_35
  (
    gbar_input_0_3,
    keyIn_0_35,
    n4
  );


  xor
  KeyPIGate_0_4
  (
    g_input_0_4,
    keyIn_0_4,
    n5
  );


  xor
  KeyPIGate_0_36
  (
    gbar_input_0_4,
    keyIn_0_36,
    n5
  );


  xor
  KeyPIGate_0_5
  (
    g_input_0_5,
    keyIn_0_5,
    n6
  );


  xor
  KeyPIGate_0_37
  (
    gbar_input_0_5,
    keyIn_0_37,
    n6
  );


  xor
  KeyPIGate_0_6
  (
    g_input_0_6,
    keyIn_0_6,
    n7
  );


  xor
  KeyPIGate_0_38
  (
    gbar_input_0_6,
    keyIn_0_38,
    n7
  );


  xor
  KeyPIGate_0_7
  (
    g_input_0_7,
    keyIn_0_7,
    n8
  );


  xor
  KeyPIGate_0_39
  (
    gbar_input_0_7,
    keyIn_0_39,
    n8
  );


  xor
  KeyPIGate_0_8
  (
    g_input_0_8,
    keyIn_0_8,
    n9
  );


  xor
  KeyPIGate_0_40
  (
    gbar_input_0_8,
    keyIn_0_40,
    n9
  );


  xor
  KeyPIGate_0_9
  (
    g_input_0_9,
    keyIn_0_9,
    n10
  );


  xor
  KeyPIGate_0_41
  (
    gbar_input_0_9,
    keyIn_0_41,
    n10
  );


  xor
  KeyPIGate_0_10
  (
    g_input_0_10,
    keyIn_0_10,
    n11
  );


  xor
  KeyPIGate_0_42
  (
    gbar_input_0_10,
    keyIn_0_42,
    n11
  );


  xor
  KeyPIGate_0_11
  (
    g_input_0_11,
    keyIn_0_11,
    n12
  );


  xor
  KeyPIGate_0_43
  (
    gbar_input_0_11,
    keyIn_0_43,
    n12
  );


  xor
  KeyPIGate_0_12
  (
    g_input_0_12,
    keyIn_0_12,
    n13
  );


  xor
  KeyPIGate_0_44
  (
    gbar_input_0_12,
    keyIn_0_44,
    n13
  );


  xor
  KeyPIGate_0_13
  (
    g_input_0_13,
    keyIn_0_13,
    n14
  );


  xor
  KeyPIGate_0_45
  (
    gbar_input_0_13,
    keyIn_0_45,
    n14
  );


  xor
  KeyPIGate_0_14
  (
    g_input_0_14,
    keyIn_0_14,
    n15
  );


  xor
  KeyPIGate_0_46
  (
    gbar_input_0_14,
    keyIn_0_46,
    n15
  );


  xor
  KeyPIGate_0_15
  (
    g_input_0_15,
    keyIn_0_15,
    n16
  );


  xor
  KeyPIGate_0_47
  (
    gbar_input_0_15,
    keyIn_0_47,
    n16
  );


  xor
  KeyPIGate_0_16
  (
    g_input_0_16,
    keyIn_0_16,
    n17
  );


  xor
  KeyPIGate_0_48
  (
    gbar_input_0_16,
    keyIn_0_48,
    n17
  );


  xor
  KeyPIGate_0_17
  (
    g_input_0_17,
    keyIn_0_17,
    n18
  );


  xor
  KeyPIGate_0_49
  (
    gbar_input_0_17,
    keyIn_0_49,
    n18
  );


  xor
  KeyPIGate_0_18
  (
    g_input_0_18,
    keyIn_0_18,
    n19
  );


  xor
  KeyPIGate_0_50
  (
    gbar_input_0_18,
    keyIn_0_50,
    n19
  );


  xor
  KeyPIGate_0_19
  (
    g_input_0_19,
    keyIn_0_19,
    n20
  );


  xor
  KeyPIGate_0_51
  (
    gbar_input_0_19,
    keyIn_0_51,
    n20
  );


  xor
  KeyPIGate_0_20
  (
    g_input_0_20,
    keyIn_0_20,
    n21
  );


  xor
  KeyPIGate_0_52
  (
    gbar_input_0_20,
    keyIn_0_52,
    n21
  );


  xor
  KeyPIGate_0_21
  (
    g_input_0_21,
    keyIn_0_21,
    n22
  );


  xor
  KeyPIGate_0_53
  (
    gbar_input_0_21,
    keyIn_0_53,
    n22
  );


  xor
  KeyPIGate_0_22
  (
    g_input_0_22,
    keyIn_0_22,
    n23
  );


  xor
  KeyPIGate_0_54
  (
    gbar_input_0_22,
    keyIn_0_54,
    n23
  );


  xor
  KeyPIGate_0_23
  (
    g_input_0_23,
    keyIn_0_23,
    n24
  );


  xor
  KeyPIGate_0_55
  (
    gbar_input_0_23,
    keyIn_0_55,
    n24
  );


  xor
  KeyPIGate_0_24
  (
    g_input_0_24,
    keyIn_0_24,
    n25
  );


  xor
  KeyPIGate_0_56
  (
    gbar_input_0_24,
    keyIn_0_56,
    n25
  );


  xor
  KeyPIGate_0_25
  (
    g_input_0_25,
    keyIn_0_25,
    n26
  );


  xor
  KeyPIGate_0_57
  (
    gbar_input_0_25,
    keyIn_0_57,
    n26
  );


  xor
  KeyPIGate_0_26
  (
    g_input_0_26,
    keyIn_0_26,
    n27
  );


  xor
  KeyPIGate_0_58
  (
    gbar_input_0_26,
    keyIn_0_58,
    n27
  );


  xor
  KeyPIGate_0_27
  (
    g_input_0_27,
    keyIn_0_27,
    n28
  );


  xor
  KeyPIGate_0_59
  (
    gbar_input_0_27,
    keyIn_0_59,
    n28
  );


  xor
  KeyPIGate_0_28
  (
    g_input_0_28,
    keyIn_0_28,
    n29
  );


  xor
  KeyPIGate_0_60
  (
    gbar_input_0_28,
    keyIn_0_60,
    n29
  );


  xor
  KeyPIGate_0_29
  (
    g_input_0_29,
    keyIn_0_29,
    n30
  );


  xor
  KeyPIGate_0_61
  (
    gbar_input_0_29,
    keyIn_0_61,
    n30
  );


  xor
  KeyPIGate_0_30
  (
    g_input_0_30,
    keyIn_0_30,
    n31
  );


  xor
  KeyPIGate_0_62
  (
    gbar_input_0_30,
    keyIn_0_62,
    n31
  );


  xor
  KeyPIGate_0_31
  (
    g_input_0_31,
    keyIn_0_31,
    n32
  );


  xor
  KeyPIGate_0_63
  (
    gbar_input_0_31,
    keyIn_0_63,
    n32
  );


  and
  f_g
  (
    f_g_wire,
    g_input_0_0,
    g_input_0_1,
    g_input_0_2,
    g_input_0_3,
    g_input_0_4,
    g_input_0_5,
    g_input_0_6,
    g_input_0_7,
    g_input_0_8,
    g_input_0_9,
    g_input_0_10,
    g_input_0_11,
    g_input_0_12,
    g_input_0_13,
    g_input_0_14,
    g_input_0_15,
    g_input_0_16,
    g_input_0_17,
    g_input_0_18,
    g_input_0_19,
    g_input_0_20,
    g_input_0_21,
    g_input_0_22,
    g_input_0_23,
    g_input_0_24,
    g_input_0_25,
    g_input_0_26,
    g_input_0_27,
    g_input_0_28,
    g_input_0_29,
    g_input_0_30,
    g_input_0_31
  );


  nand
  f_gbar
  (
    f_gbar_wire,
    gbar_input_0_0,
    gbar_input_0_1,
    gbar_input_0_2,
    gbar_input_0_3,
    gbar_input_0_4,
    gbar_input_0_5,
    gbar_input_0_6,
    gbar_input_0_7,
    gbar_input_0_8,
    gbar_input_0_9,
    gbar_input_0_10,
    gbar_input_0_11,
    gbar_input_0_12,
    gbar_input_0_13,
    gbar_input_0_14,
    gbar_input_0_15,
    gbar_input_0_16,
    gbar_input_0_17,
    gbar_input_0_18,
    gbar_input_0_19,
    gbar_input_0_20,
    gbar_input_0_21,
    gbar_input_0_22,
    gbar_input_0_23,
    gbar_input_0_24,
    gbar_input_0_25,
    gbar_input_0_26,
    gbar_input_0_27,
    gbar_input_0_28,
    gbar_input_0_29,
    gbar_input_0_30,
    gbar_input_0_31
  );


  and
  G
  (
    AntiSAT_output,
    f_g_wire,
    f_gbar_wire
  );


  xor
  flip_it
  (
    n998,
    AntiSAT_output,
    AntiSAT_key_wire
  );


endmodule

