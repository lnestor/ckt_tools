// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1197_31_10 written by SynthGen on 2021/05/24 19:42:17
module Stat_1197_31_10( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23,
 n989, n996, n990, n1013, n1017, n993, n981, n1014,
 n994, n991, n1008, n1001, n999, n992, n1005, n987,
 n997, n985, n982, n1004, n988, n1028, n1026, n1031,
 n1023, n1029, n1025, n1022, n1027, n1181, n1197, n1220);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23;

output n989, n996, n990, n1013, n1017, n993, n981, n1014,
 n994, n991, n1008, n1001, n999, n992, n1005, n987,
 n997, n985, n982, n1004, n988, n1028, n1026, n1031,
 n1023, n1029, n1025, n1022, n1027, n1181, n1197, n1220;

wire n24, n25, n26, n27, n28, n29, n30, n31,
 n32, n33, n34, n35, n36, n37, n38, n39,
 n40, n41, n42, n43, n44, n45, n46, n47,
 n48, n49, n50, n51, n52, n53, n54, n55,
 n56, n57, n58, n59, n60, n61, n62, n63,
 n64, n65, n66, n67, n68, n69, n70, n71,
 n72, n73, n74, n75, n76, n77, n78, n79,
 n80, n81, n82, n83, n84, n85, n86, n87,
 n88, n89, n90, n91, n92, n93, n94, n95,
 n96, n97, n98, n99, n100, n101, n102, n103,
 n104, n105, n106, n107, n108, n109, n110, n111,
 n112, n113, n114, n115, n116, n117, n118, n119,
 n120, n121, n122, n123, n124, n125, n126, n127,
 n128, n129, n130, n131, n132, n133, n134, n135,
 n136, n137, n138, n139, n140, n141, n142, n143,
 n144, n145, n146, n147, n148, n149, n150, n151,
 n152, n153, n154, n155, n156, n157, n158, n159,
 n160, n161, n162, n163, n164, n165, n166, n167,
 n168, n169, n170, n171, n172, n173, n174, n175,
 n176, n177, n178, n179, n180, n181, n182, n183,
 n184, n185, n186, n187, n188, n189, n190, n191,
 n192, n193, n194, n195, n196, n197, n198, n199,
 n200, n201, n202, n203, n204, n205, n206, n207,
 n208, n209, n210, n211, n212, n213, n214, n215,
 n216, n217, n218, n219, n220, n221, n222, n223,
 n224, n225, n226, n227, n228, n229, n230, n231,
 n232, n233, n234, n235, n236, n237, n238, n239,
 n240, n241, n242, n243, n244, n245, n246, n247,
 n248, n249, n250, n251, n252, n253, n254, n255,
 n256, n257, n258, n259, n260, n261, n262, n263,
 n264, n265, n266, n267, n268, n269, n270, n271,
 n272, n273, n274, n275, n276, n277, n278, n279,
 n280, n281, n282, n283, n284, n285, n286, n287,
 n288, n289, n290, n291, n292, n293, n294, n295,
 n296, n297, n298, n299, n300, n301, n302, n303,
 n304, n305, n306, n307, n308, n309, n310, n311,
 n312, n313, n314, n315, n316, n317, n318, n319,
 n320, n321, n322, n323, n324, n325, n326, n327,
 n328, n329, n330, n331, n332, n333, n334, n335,
 n336, n337, n338, n339, n340, n341, n342, n343,
 n344, n345, n346, n347, n348, n349, n350, n351,
 n352, n353, n354, n355, n356, n357, n358, n359,
 n360, n361, n362, n363, n364, n365, n366, n367,
 n368, n369, n370, n371, n372, n373, n374, n375,
 n376, n377, n378, n379, n380, n381, n382, n383,
 n384, n385, n386, n387, n388, n389, n390, n391,
 n392, n393, n394, n395, n396, n397, n398, n399,
 n400, n401, n402, n403, n404, n405, n406, n407,
 n408, n409, n410, n411, n412, n413, n414, n415,
 n416, n417, n418, n419, n420, n421, n422, n423,
 n424, n425, n426, n427, n428, n429, n430, n431,
 n432, n433, n434, n435, n436, n437, n438, n439,
 n440, n441, n442, n443, n444, n445, n446, n447,
 n448, n449, n450, n451, n452, n453, n454, n455,
 n456, n457, n458, n459, n460, n461, n462, n463,
 n464, n465, n466, n467, n468, n469, n470, n471,
 n472, n473, n474, n475, n476, n477, n478, n479,
 n480, n481, n482, n483, n484, n485, n486, n487,
 n488, n489, n490, n491, n492, n493, n494, n495,
 n496, n497, n498, n499, n500, n501, n502, n503,
 n504, n505, n506, n507, n508, n509, n510, n511,
 n512, n513, n514, n515, n516, n517, n518, n519,
 n520, n521, n522, n523, n524, n525, n526, n527,
 n528, n529, n530, n531, n532, n533, n534, n535,
 n536, n537, n538, n539, n540, n541, n542, n543,
 n544, n545, n546, n547, n548, n549, n550, n551,
 n552, n553, n554, n555, n556, n557, n558, n559,
 n560, n561, n562, n563, n564, n565, n566, n567,
 n568, n569, n570, n571, n572, n573, n574, n575,
 n576, n577, n578, n579, n580, n581, n582, n583,
 n584, n585, n586, n587, n588, n589, n590, n591,
 n592, n593, n594, n595, n596, n597, n598, n599,
 n600, n601, n602, n603, n604, n605, n606, n607,
 n608, n609, n610, n611, n612, n613, n614, n615,
 n616, n617, n618, n619, n620, n621, n622, n623,
 n624, n625, n626, n627, n628, n629, n630, n631,
 n632, n633, n634, n635, n636, n637, n638, n639,
 n640, n641, n642, n643, n644, n645, n646, n647,
 n648, n649, n650, n651, n652, n653, n654, n655,
 n656, n657, n658, n659, n660, n661, n662, n663,
 n664, n665, n666, n667, n668, n669, n670, n671,
 n672, n673, n674, n675, n676, n677, n678, n679,
 n680, n681, n682, n683, n684, n685, n686, n687,
 n688, n689, n690, n691, n692, n693, n694, n695,
 n696, n697, n698, n699, n700, n701, n702, n703,
 n704, n705, n706, n707, n708, n709, n710, n711,
 n712, n713, n714, n715, n716, n717, n718, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n731, n732, n733, n734, n735,
 n736, n737, n738, n739, n740, n741, n742, n743,
 n744, n745, n746, n747, n748, n749, n750, n751,
 n752, n753, n754, n755, n756, n757, n758, n759,
 n760, n761, n762, n763, n764, n765, n766, n767,
 n768, n769, n770, n771, n772, n773, n774, n775,
 n776, n777, n778, n779, n780, n781, n782, n783,
 n784, n785, n786, n787, n788, n789, n790, n791,
 n792, n793, n794, n795, n796, n797, n798, n799,
 n800, n801, n802, n803, n804, n805, n806, n807,
 n808, n809, n810, n811, n812, n813, n814, n815,
 n816, n817, n818, n819, n820, n821, n822, n823,
 n824, n825, n826, n827, n828, n829, n830, n831,
 n832, n833, n834, n835, n836, n837, n838, n839,
 n840, n841, n842, n843, n844, n845, n846, n847,
 n848, n849, n850, n851, n852, n853, n854, n855,
 n856, n857, n858, n859, n860, n861, n862, n863,
 n864, n865, n866, n867, n868, n869, n870, n871,
 n872, n873, n874, n875, n876, n877, n878, n879,
 n880, n881, n882, n883, n884, n885, n886, n887,
 n888, n889, n890, n891, n892, n893, n894, n895,
 n896, n897, n898, n899, n900, n901, n902, n903,
 n904, n905, n906, n907, n908, n909, n910, n911,
 n912, n913, n914, n915, n916, n917, n918, n919,
 n920, n921, n922, n923, n924, n925, n926, n927,
 n928, n929, n930, n931, n932, n933, n934, n935,
 n936, n937, n938, n939, n940, n941, n942, n943,
 n944, n945, n946, n947, n948, n949, n950, n951,
 n952, n953, n954, n955, n956, n957, n958, n959,
 n960, n961, n962, n963, n964, n965, n966, n967,
 n968, n969, n970, n971, n972, n973, n974, n975,
 n976, n977, n978, n979, n980, n983, n984, n986,
 n995, n998, n1000, n1002, n1003, n1006, n1007, n1009,
 n1010, n1011, n1012, n1015, n1016, n1018, n1019, n1020,
 n1021, n1024, n1030, n1032, n1033, n1034, n1035, n1036,
 n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
 n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
 n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
 n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
 n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
 n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
 n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
 n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
 n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
 n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
 n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
 n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
 n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
 n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
 n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
 n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
 n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
 n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
 n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
 n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1198,
 n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
 n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
 n1215, n1216, n1217, n1218, n1219;

buf  g0 (n78, n7);
buf  g1 (n82, n13);
not  g2 (n71, n6);
not  g3 (n36, n8);
not  g4 (n26, n6);
not  g5 (n113, n11);
not  g6 (n91, n23);
not  g7 (n114, n6);
not  g8 (n112, n16);
buf  g9 (n81, n21);
buf  g10 (n84, n6);
not  g11 (n70, n23);
buf  g12 (n25, n11);
not  g13 (n85, n18);
buf  g14 (n33, n21);
not  g15 (n34, n13);
buf  g16 (n99, n18);
not  g17 (n64, n4);
not  g18 (n56, n8);
not  g19 (n67, n16);
buf  g20 (n59, n10);
not  g21 (n57, n14);
not  g22 (n51, n4);
not  g23 (n89, n15);
not  g24 (n100, n19);
not  g25 (n106, n20);
not  g26 (n76, n13);
not  g27 (n29, n18);
not  g28 (n44, n1);
buf  g29 (n115, n20);
buf  g30 (n88, n16);
buf  g31 (n94, n19);
buf  g32 (n48, n1);
not  g33 (n80, n22);
buf  g34 (n75, n23);
not  g35 (n43, n19);
buf  g36 (n32, n3);
not  g37 (n60, n9);
buf  g38 (n53, n9);
not  g39 (n45, n3);
buf  g40 (n95, n17);
not  g41 (n68, n12);
not  g42 (n27, n16);
buf  g43 (n101, n2);
buf  g44 (n55, n1);
buf  g45 (n58, n11);
buf  g46 (n105, n17);
not  g47 (n65, n21);
not  g48 (n49, n4);
buf  g49 (n103, n15);
buf  g50 (n31, n17);
buf  g51 (n111, n20);
not  g52 (n83, n12);
not  g53 (n52, n10);
buf  g54 (n73, n8);
not  g55 (n97, n7);
not  g56 (n28, n23);
not  g57 (n24, n10);
not  g58 (n61, n14);
not  g59 (n92, n2);
buf  g60 (n30, n4);
buf  g61 (n47, n12);
buf  g62 (n86, n15);
not  g63 (n69, n12);
not  g64 (n40, n9);
buf  g65 (n63, n10);
buf  g66 (n93, n1);
not  g67 (n98, n3);
buf  g68 (n108, n14);
not  g69 (n109, n19);
not  g70 (n66, n5);
buf  g71 (n79, n3);
not  g72 (n104, n15);
buf  g73 (n39, n14);
not  g74 (n107, n18);
buf  g75 (n102, n21);
not  g76 (n110, n22);
buf  g77 (n90, n13);
buf  g78 (n74, n7);
not  g79 (n54, n2);
not  g80 (n50, n22);
not  g81 (n87, n22);
not  g82 (n96, n5);
not  g83 (n77, n11);
not  g84 (n72, n17);
not  g85 (n35, n2);
not  g86 (n38, n5);
not  g87 (n42, n7);
buf  g88 (n62, n8);
not  g89 (n37, n5);
not  g90 (n41, n20);
buf  g91 (n46, n9);
not  g92 (n355, n77);
buf  g93 (n343, n111);
not  g94 (n246, n112);
not  g95 (n414, n42);
buf  g96 (n283, n31);
buf  g97 (n444, n71);
not  g98 (n135, n30);
buf  g99 (n367, n25);
not  g100 (n155, n85);
buf  g101 (n124, n38);
buf  g102 (n420, n37);
buf  g103 (n276, n108);
not  g104 (n482, n57);
not  g105 (n456, n34);
not  g106 (n223, n45);
not  g107 (n141, n46);
buf  g108 (n221, n102);
not  g109 (n396, n42);
buf  g110 (n169, n103);
buf  g111 (n303, n110);
not  g112 (n455, n95);
buf  g113 (n332, n93);
not  g114 (n237, n47);
not  g115 (n173, n80);
buf  g116 (n277, n104);
buf  g117 (n401, n40);
not  g118 (n405, n49);
buf  g119 (n447, n62);
not  g120 (n333, n27);
not  g121 (n361, n76);
not  g122 (n296, n70);
buf  g123 (n418, n50);
not  g124 (n366, n54);
buf  g125 (n218, n59);
not  g126 (n119, n54);
buf  g127 (n442, n67);
not  g128 (n352, n75);
not  g129 (n369, n97);
not  g130 (n229, n107);
buf  g131 (n335, n77);
buf  g132 (n269, n69);
not  g133 (n408, n73);
buf  g134 (n323, n56);
not  g135 (n454, n79);
buf  g136 (n469, n49);
buf  g137 (n285, n44);
buf  g138 (n353, n98);
not  g139 (n232, n108);
buf  g140 (n429, n42);
buf  g141 (n432, n102);
not  g142 (n397, n34);
not  g143 (n172, n85);
buf  g144 (n437, n112);
not  g145 (n165, n75);
buf  g146 (n300, n110);
not  g147 (n449, n75);
buf  g148 (n242, n33);
not  g149 (n189, n89);
not  g150 (n194, n94);
not  g151 (n208, n61);
buf  g152 (n306, n82);
buf  g153 (n328, n85);
buf  g154 (n346, n27);
not  g155 (n130, n84);
not  g156 (n268, n82);
buf  g157 (n294, n111);
not  g158 (n251, n91);
buf  g159 (n249, n101);
not  g160 (n211, n97);
not  g161 (n382, n41);
buf  g162 (n468, n106);
not  g163 (n471, n48);
not  g164 (n185, n30);
not  g165 (n458, n71);
buf  g166 (n406, n99);
buf  g167 (n433, n38);
buf  g168 (n383, n65);
not  g169 (n461, n92);
buf  g170 (n290, n107);
not  g171 (n282, n46);
not  g172 (n476, n81);
not  g173 (n215, n48);
not  g174 (n395, n61);
not  g175 (n257, n104);
buf  g176 (n373, n38);
buf  g177 (n180, n58);
not  g178 (n327, n114);
not  g179 (n326, n68);
not  g180 (n273, n113);
buf  g181 (n117, n68);
buf  g182 (n133, n28);
buf  g183 (n375, n98);
not  g184 (n402, n70);
not  g185 (n310, n28);
buf  g186 (n329, n72);
not  g187 (n219, n68);
not  g188 (n260, n35);
not  g189 (n261, n51);
not  g190 (n190, n50);
buf  g191 (n132, n62);
not  g192 (n201, n109);
not  g193 (n336, n44);
not  g194 (n407, n70);
buf  g195 (n467, n76);
not  g196 (n378, n46);
not  g197 (n118, n66);
buf  g198 (n143, n115);
buf  g199 (n388, n52);
buf  g200 (n274, n100);
not  g201 (n216, n49);
buf  g202 (n145, n109);
not  g203 (n195, n50);
not  g204 (n236, n75);
buf  g205 (n439, n67);
not  g206 (n428, n43);
buf  g207 (n252, n57);
not  g208 (n364, n40);
not  g209 (n160, n100);
not  g210 (n295, n92);
buf  g211 (n142, n36);
not  g212 (n341, n83);
not  g213 (n234, n39);
buf  g214 (n187, n71);
buf  g215 (n386, n27);
buf  g216 (n146, n103);
not  g217 (n230, n84);
not  g218 (n435, n41);
buf  g219 (n253, n61);
buf  g220 (n284, n101);
not  g221 (n411, n51);
not  g222 (n241, n91);
not  g223 (n156, n76);
not  g224 (n421, n53);
not  g225 (n213, n110);
buf  g226 (n379, n69);
buf  g227 (n280, n47);
buf  g228 (n123, n26);
buf  g229 (n391, n55);
buf  g230 (n116, n65);
not  g231 (n417, n57);
not  g232 (n462, n29);
buf  g233 (n440, n51);
buf  g234 (n199, n104);
buf  g235 (n314, n72);
not  g236 (n394, n69);
not  g237 (n392, n30);
not  g238 (n272, n76);
not  g239 (n245, n80);
buf  g240 (n321, n113);
buf  g241 (n360, n32);
buf  g242 (n424, n43);
not  g243 (n288, n64);
not  g244 (n174, n24);
not  g245 (n316, n29);
not  g246 (n409, n79);
buf  g247 (n349, n109);
not  g248 (n224, n100);
not  g249 (n178, n36);
not  g250 (n466, n24);
buf  g251 (n415, n106);
not  g252 (n176, n31);
not  g253 (n149, n33);
not  g254 (n450, n105);
not  g255 (n473, n55);
not  g256 (n151, n33);
not  g257 (n270, n55);
not  g258 (n319, n26);
not  g259 (n254, n98);
not  g260 (n400, n47);
buf  g261 (n431, n68);
buf  g262 (n197, n82);
buf  g263 (n287, n41);
buf  g264 (n203, n77);
not  g265 (n315, n114);
not  g266 (n330, n54);
buf  g267 (n480, n113);
not  g268 (n264, n102);
buf  g269 (n479, n86);
not  g270 (n265, n45);
not  g271 (n168, n115);
buf  g272 (n472, n43);
not  g273 (n144, n34);
buf  g274 (n183, n52);
not  g275 (n318, n59);
buf  g276 (n292, n91);
buf  g277 (n210, n56);
not  g278 (n298, n48);
not  g279 (n281, n101);
buf  g280 (n351, n93);
not  g281 (n381, n59);
not  g282 (n275, n83);
buf  g283 (n259, n24);
not  g284 (n419, n107);
buf  g285 (n175, n53);
buf  g286 (n436, n92);
buf  g287 (n416, n90);
buf  g288 (n475, n115);
not  g289 (n302, n94);
buf  g290 (n404, n105);
buf  g291 (n164, n81);
buf  g292 (n181, n67);
not  g293 (n297, n73);
buf  g294 (n425, n106);
buf  g295 (n412, n59);
buf  g296 (n247, n63);
buf  g297 (n387, n83);
not  g298 (n138, n72);
not  g299 (n363, n115);
not  g300 (n122, n53);
buf  g301 (n374, n31);
buf  g302 (n368, n107);
not  g303 (n289, n24);
buf  g304 (n121, n48);
not  g305 (n293, n64);
not  g306 (n163, n58);
not  g307 (n186, n37);
buf  g308 (n129, n96);
not  g309 (n147, n96);
buf  g310 (n354, n85);
not  g311 (n474, n93);
not  g312 (n206, n32);
not  g313 (n477, n73);
buf  g314 (n339, n66);
not  g315 (n128, n78);
buf  g316 (n350, n79);
not  g317 (n157, n86);
buf  g318 (n430, n65);
buf  g319 (n322, n81);
buf  g320 (n154, n102);
buf  g321 (n403, n35);
not  g322 (n120, n114);
buf  g323 (n198, n39);
not  g324 (n207, n97);
not  g325 (n158, n43);
buf  g326 (n214, n113);
not  g327 (n342, n36);
buf  g328 (n389, n89);
buf  g329 (n271, n94);
buf  g330 (n131, n90);
buf  g331 (n324, n33);
not  g332 (n347, n66);
not  g333 (n423, n49);
not  g334 (n313, n84);
buf  g335 (n126, n82);
buf  g336 (n209, n64);
not  g337 (n483, n87);
buf  g338 (n243, n103);
buf  g339 (n240, n94);
not  g340 (n202, n37);
not  g341 (n307, n30);
not  g342 (n309, n69);
buf  g343 (n345, n112);
buf  g344 (n212, n70);
not  g345 (n365, n95);
buf  g346 (n153, n88);
not  g347 (n348, n42);
not  g348 (n312, n109);
buf  g349 (n334, n46);
buf  g350 (n399, n90);
buf  g351 (n279, n96);
not  g352 (n377, n52);
buf  g353 (n459, n31);
not  g354 (n443, n78);
buf  g355 (n337, n87);
not  g356 (n311, n83);
buf  g357 (n325, n60);
buf  g358 (n193, n40);
buf  g359 (n262, n56);
buf  g360 (n255, n91);
buf  g361 (n136, n105);
buf  g362 (n179, n64);
buf  g363 (n205, n44);
not  g364 (n320, n87);
buf  g365 (n463, n114);
buf  g366 (n278, n86);
buf  g367 (n286, n95);
buf  g368 (n384, n74);
not  g369 (n304, n89);
not  g370 (n267, n28);
buf  g371 (n413, n101);
not  g372 (n222, n73);
buf  g373 (n427, n74);
not  g374 (n170, n62);
buf  g375 (n362, n104);
not  g376 (n250, n99);
buf  g377 (n305, n81);
buf  g378 (n344, n98);
buf  g379 (n438, n51);
buf  g380 (n248, n87);
not  g381 (n340, n50);
buf  g382 (n227, n62);
not  g383 (n448, n77);
not  g384 (n191, n44);
buf  g385 (n238, n108);
not  g386 (n457, n99);
buf  g387 (n148, n80);
not  g388 (n372, n61);
not  g389 (n239, n97);
not  g390 (n452, n29);
not  g391 (n139, n63);
not  g392 (n184, n45);
not  g393 (n226, n111);
buf  g394 (n171, n78);
not  g395 (n235, n88);
buf  g396 (n233, n74);
not  g397 (n200, n39);
not  g398 (n451, n36);
not  g399 (n358, n112);
not  g400 (n478, n54);
buf  g401 (n359, n92);
buf  g402 (n263, n58);
buf  g403 (n152, n65);
buf  g404 (n140, n41);
not  g405 (n150, n38);
buf  g406 (n371, n32);
buf  g407 (n162, n57);
not  g408 (n182, n84);
buf  g409 (n390, n86);
not  g410 (n299, n89);
buf  g411 (n177, n34);
buf  g412 (n244, n35);
not  g413 (n422, n37);
buf  g414 (n445, n25);
buf  g415 (n393, n47);
buf  g416 (n446, n88);
buf  g417 (n464, n111);
not  g418 (n166, n25);
buf  g419 (n385, n29);
buf  g420 (n125, n103);
not  g421 (n376, n45);
not  g422 (n204, n110);
not  g423 (n481, n60);
not  g424 (n370, n105);
buf  g425 (n127, n28);
buf  g426 (n357, n106);
not  g427 (n228, n60);
not  g428 (n338, n39);
buf  g429 (n137, n78);
buf  g430 (n220, n80);
buf  g431 (n301, n27);
buf  g432 (n410, n26);
buf  g433 (n161, n55);
not  g434 (n134, n52);
not  g435 (n317, n56);
not  g436 (n453, n25);
not  g437 (n398, n53);
not  g438 (n308, n58);
buf  g439 (n441, n66);
not  g440 (n460, n60);
not  g441 (n231, n40);
buf  g442 (n434, n32);
not  g443 (n291, n71);
buf  g444 (n380, n99);
not  g445 (n167, n96);
not  g446 (n470, n93);
not  g447 (n465, n26);
buf  g448 (n192, n108);
buf  g449 (n258, n74);
buf  g450 (n426, n63);
not  g451 (n217, n67);
buf  g452 (n159, n72);
not  g453 (n256, n63);
buf  g454 (n331, n90);
not  g455 (n356, n35);
buf  g456 (n225, n95);
not  g457 (n188, n79);
buf  g458 (n196, n100);
buf  g459 (n266, n88);
nand g460 (n671, n381, n379, n325, n332);
and  g461 (n591, n411, n331, n281, n409);
and  g462 (n701, n239, n331, n232, n367);
nor  g463 (n533, n412, n276, n309, n248);
nor  g464 (n517, n371, n420, n269, n397);
nor  g465 (n546, n317, n330, n334, n400);
and  g466 (n495, n385, n397, n434, n353);
xnor g467 (n624, n386, n426, n320, n409);
and  g468 (n710, n336, n404, n291, n416);
and  g469 (n650, n436, n357, n318, n245);
nand g470 (n513, n386, n345, n346, n348);
nand g471 (n580, n401, n199, n309, n362);
nand g472 (n519, n343, n408, n416, n310);
and  g473 (n581, n322, n445, n382, n347);
nand g474 (n699, n315, n381, n228, n281);
nand g475 (n574, n344, n374, n417, n429);
xor  g476 (n697, n447, n427, n245, n337);
or   g477 (n582, n272, n378, n306, n349);
and  g478 (n622, n166, n312, n376, n165);
or   g479 (n493, n259, n403, n424, n435);
nor  g480 (n616, n424, n267, n238, n252);
xnor g481 (n549, n251, n418, n425, n436);
xnor g482 (n615, n313, n326, n442, n443);
xnor g483 (n526, n277, n421, n381, n375);
xnor g484 (n562, n319, n301, n248, n293);
xnor g485 (n684, n296, n384, n441, n403);
xnor g486 (n536, n344, n338, n286, n194);
xnor g487 (n644, n361, n283, n119, n253);
or   g488 (n523, n197, n355, n432, n363);
or   g489 (n649, n255, n378, n148, n327);
and  g490 (n494, n310, n279, n126, n180);
xnor g491 (n648, n396, n408, n325, n404);
nor  g492 (n576, n379, n285, n236, n334);
or   g493 (n658, n294, n297, n365, n332);
or   g494 (n610, n383, n258, n213, n127);
and  g495 (n510, n392, n273, n343, n121);
xnor g496 (n599, n395, n142, n431, n151);
and  g497 (n543, n307, n370, n316, n225);
xnor g498 (n572, n153, n422, n313, n284);
nor  g499 (n695, n304, n206, n239, n358);
nor  g500 (n503, n150, n315, n221, n262);
or   g501 (n601, n271, n441, n412, n269);
xor  g502 (n652, n363, n161, n277, n359);
xnor g503 (n587, n227, n415, n308, n407);
or   g504 (n609, n386, n124, n334, n341);
xor  g505 (n507, n420, n278, n287, n139);
or   g506 (n542, n144, n287, n292, n316);
nor  g507 (n702, n242, n445, n177, n364);
or   g508 (n515, n274, n303, n192, n332);
and  g509 (n566, n274, n313, n307, n342);
xor  g510 (n537, n435, n405, n446, n372);
and  g511 (n489, n363, n339, n391, n223);
nor  g512 (n682, n391, n414, n179, n247);
and  g513 (n556, n211, n212, n130, n372);
xor  g514 (n643, n438, n306, n333, n277);
or   g515 (n598, n434, n388, n314, n353);
and  g516 (n578, n406, n254, n277, n286);
nand g517 (n501, n422, n305, n356, n386);
and  g518 (n540, n203, n198, n219, n325);
xnor g519 (n676, n351, n378, n385, n347);
xor  g520 (n498, n350, n300, n327, n360);
xor  g521 (n508, n355, n281, n217, n395);
and  g522 (n618, n309, n276, n335, n387);
nor  g523 (n569, n390, n176, n145, n288);
nand g524 (n612, n427, n371, n293);
xnor g525 (n657, n331, n400, n357, n375);
xor  g526 (n647, n275, n433, n292, n346);
nor  g527 (n584, n403, n341, n417, n345);
nand g528 (n535, n364, n424, n254, n274);
xnor g529 (n593, n349, n437, n377, n322);
nor  g530 (n573, n282, n445, n188, n131);
nor  g531 (n512, n394, n430, n134, n332);
or   g532 (n558, n258, n321, n259, n352);
xnor g533 (n655, n261, n380, n310, n238);
xnor g534 (n511, n225, n329, n439, n376);
and  g535 (n674, n135, n421, n412, n379);
xor  g536 (n588, n296, n343, n366, n270);
xnor g537 (n527, n383, n442, n210, n347);
nor  g538 (n575, n314, n340, n370, n392);
xnor g539 (n504, n324, n389, n443, n339);
xnor g540 (n662, n302, n162, n289, n421);
nor  g541 (n564, n393, n395, n381, n389);
and  g542 (n653, n249, n222, n229, n272);
and  g543 (n525, n326, n243, n337, n368);
and  g544 (n611, n428, n356, n349, n233);
xnor g545 (n613, n444, n328, n207, n301);
nand g546 (n669, n428, n328, n402, n255);
nor  g547 (n524, n307, n306, n123, n168);
nor  g548 (n626, n413, n440, n367, n283);
xor  g549 (n675, n435, n322, n374, n302);
nand g550 (n547, n388, n389, n440, n428);
xor  g551 (n659, n402, n242, n427, n366);
xnor g552 (n565, n340, n415, n326, n311);
xnor g553 (n681, n380, n289, n337, n327);
or   g554 (n641, n214, n323, n348, n293);
nor  g555 (n585, n396, n270, n359, n330);
xor  g556 (n663, n430, n411, n429, n351);
xor  g557 (n545, n333, n320, n442, n291);
xor  g558 (n607, n352, n424, n292, n319);
nand g559 (n531, n312, n396, n390, n374);
xnor g560 (n595, n404, n329, n439, n167);
xnor g561 (n686, n364, n300, n388, n414);
nand g562 (n520, n299, n445, n169, n409);
nor  g563 (n634, n384, n250, n183, n361);
xor  g564 (n500, n260, n227, n328, n208);
xnor g565 (n698, n337, n361, n132, n419);
and  g566 (n560, n354, n285, n289, n423);
xnor g567 (n706, n122, n283, n346, n300);
nor  g568 (n561, n304, n338, n250, n195);
and  g569 (n567, n420, n425, n307, n380);
and  g570 (n552, n437, n251, n233, n305);
nand g571 (n705, n321, n412, n402, n365);
or   g572 (n665, n201, n433, n368, n181);
or   g573 (n656, n387, n432, n252, n312);
nor  g574 (n538, n338, n241, n370, n284);
xor  g575 (n621, n367, n247, n117, n295);
nand g576 (n497, n156, n279, n447, n370);
nand g577 (n630, n393, n446, n348, n118);
xor  g578 (n603, n446, n345, n292, n191);
nand g579 (n687, n116, n322, n400, n444);
and  g580 (n534, n387, n431, n354, n443);
nand g581 (n484, n275, n414, n383, n447);
xnor g582 (n492, n363, n342, n280, n244);
or   g583 (n579, n308, n413, n320, n303);
xor  g584 (n666, n407, n422, n434, n185);
and  g585 (n677, n421, n398, n432, n265);
xnor g586 (n596, n289, n375, n282, n202);
and  g587 (n553, n266, n417, n138, n431);
nor  g588 (n619, n186, n415, n273, n305);
nor  g589 (n683, n297, n164, n278, n369);
or   g590 (n532, n311, n272, n120, n315);
xnor g591 (n590, n246, n129, n330, n268);
nor  g592 (n548, n340, n299, n403, n311);
nor  g593 (n506, n405, n280, n297, n373);
and  g594 (n638, n368, n371, n344, n352);
xor  g595 (n586, n228, n359, n360, n351);
nand g596 (n680, n410, n418, n340, n444);
nand g597 (n694, n390, n368, n365, n393);
nand g598 (n668, n323, n408, n246, n425);
and  g599 (n505, n286, n355, n299, n205);
or   g600 (n544, n358, n439, n318, n175);
xnor g601 (n516, n394, n336, n149, n288);
and  g602 (n673, n282, n317, n434, n236);
and  g603 (n592, n273, n290, n379, n429);
xor  g604 (n707, n137, n441, n329, n360);
xor  g605 (n530, n281, n172, n410, n357);
nand g606 (n559, n418, n257, n317, n350);
and  g607 (n509, n373, n325, n282, n280);
and  g608 (n696, n285, n304, n209, n283);
nand g609 (n642, n285, n356, n423, n157);
or   g610 (n690, n226, n319, n298, n312);
xor  g611 (n577, n290, n173, n366, n369);
xor  g612 (n528, n243, n399, n384, n244);
and  g613 (n486, n354, n399, n406, n408);
or   g614 (n594, n398, n441, n402, n397);
nor  g615 (n496, n339, n336, n367, n416);
and  g616 (n633, n229, n348, n345, n240);
nor  g617 (n488, n400, n356, n140, n411);
xnor g618 (n709, n392, n433, n437, n141);
and  g619 (n554, n342, n394, n261, n335);
xnor g620 (n514, n216, n297, n317, n133);
or   g621 (n667, n383, n318, n218, n329);
nand g622 (n623, n284, n387, n362, n406);
nand g623 (n637, n342, n237, n382, n302);
or   g624 (n518, n361, n391, n235, n275);
and  g625 (n555, n351, n313, n365, n440);
nand g626 (n678, n384, n328, n274, n419);
xor  g627 (n708, n298, n350, n234, n413);
and  g628 (n654, n136, n350, n300, n398);
xnor g629 (n522, n196, n291, n253, n323);
and  g630 (n490, n318, n373, n413, n125);
nand g631 (n693, n303, n295, n237, n308);
xnor g632 (n632, n264, n163, n369, n260);
xor  g633 (n491, n158, n366, n330, n436);
nor  g634 (n664, n407, n423, n401, n428);
xor  g635 (n589, n286, n439, n419, n231);
xnor g636 (n640, n436, n407, n257, n326);
xnor g637 (n600, n224, n200, n349, n397);
and  g638 (n521, n298, n391, n429, n288);
xor  g639 (n627, n220, n288, n338, n316);
nand g640 (n606, n395, n426, n182, n343);
and  g641 (n685, n190, n389, n392, n414);
xor  g642 (n604, n334, n287, n159, n353);
nand g643 (n570, n310, n290, n422, n152);
nand g644 (n691, n360, n147, n278, n401);
or   g645 (n672, n438, n303, n390, n341);
nand g646 (n703, n265, n331, n426, n315);
nand g647 (n563, n278, n396, n410, n321);
and  g648 (n539, n324, n226, n287, n430);
xor  g649 (n617, n352, n170, n435, n420);
nand g650 (n704, n442, n279, n437, n362);
nand g651 (n485, n256, n333, n404, n262);
xor  g652 (n614, n373, n440, n240, n146);
xor  g653 (n636, n230, n358, n362, n380);
and  g654 (n635, n372, n296, n294, n447);
xnor g655 (n487, n319, n143, n336, n364);
xnor g656 (n692, n256, n369, n446, n398);
xnor g657 (n550, n335, n346, n433, n423);
xor  g658 (n700, n154, n430, n306, n296);
nor  g659 (n639, n302, n372, n301, n275);
nand g660 (n568, n301, n241, n393, n266);
and  g661 (n646, n432, n399, n377, n298);
nand g662 (n571, n264, n189, n410, n347);
or   g663 (n661, n267, n359, n427, n280);
xnor g664 (n608, n279, n415, n378, n394);
or   g665 (n557, n385, n294, n295, n409);
or   g666 (n602, n295, n284, n401, n438);
and  g667 (n597, n324, n333, n377, n271);
and  g668 (n502, n425, n263, n234, n375);
or   g669 (n620, n187, n128, n341, n444);
nand g670 (n541, n418, n388, n399, n323);
and  g671 (n645, n417, n276, n155, n263);
xor  g672 (n689, n204, n377, n160, n406);
nor  g673 (n651, n321, n193, n405, n358);
nor  g674 (n605, n316, n273, n431, n290);
or   g675 (n499, n308, n231, n294, n299);
nand g676 (n625, n327, n215, n224, n355);
nor  g677 (n629, n232, n382, n311, n374);
xor  g678 (n529, n272, n304, n339, n411);
or   g679 (n660, n353, n419, n314, n438);
or   g680 (n583, n178, n371, n174, n249);
nor  g681 (n628, n171, n268, n309, n235);
and  g682 (n670, n184, n324, n385, n357);
xnor g683 (n688, n443, n405, n376, n230);
xor  g684 (n679, n426, n320, n416, n376);
or   g685 (n551, n354, n382, n314, n291);
or   g686 (n631, n335, n305, n344, n276);
not  g687 (n736, n513);
not  g688 (n728, n507);
not  g689 (n713, n497);
buf  g690 (n723, n506);
not  g691 (n739, n509);
buf  g692 (n711, n511);
not  g693 (n741, n515);
not  g694 (n735, n505);
not  g695 (n715, n503);
buf  g696 (n731, n489);
buf  g697 (n714, n514);
not  g698 (n726, n508);
not  g699 (n733, n491);
buf  g700 (n730, n502);
not  g701 (n721, n500);
not  g702 (n719, n490);
not  g703 (n724, n486);
not  g704 (n729, n492);
buf  g705 (n738, n487);
buf  g706 (n712, n493);
buf  g707 (n727, n501);
not  g708 (n722, n512);
buf  g709 (n717, n485);
not  g710 (n737, n498);
not  g711 (n716, n510);
buf  g712 (n725, n494);
not  g713 (n740, n499);
not  g714 (n720, n484);
not  g715 (n742, n496);
not  g716 (n734, n488);
not  g717 (n718, n495);
not  g718 (n732, n504);
buf  g719 (n757, n719);
not  g720 (n762, n729);
buf  g721 (n754, n713);
buf  g722 (n761, n723);
buf  g723 (n746, n727);
buf  g724 (n750, n725);
buf  g725 (n744, n730);
not  g726 (n752, n721);
buf  g727 (n743, n715);
buf  g728 (n751, n717);
not  g729 (n745, n728);
not  g730 (n755, n716);
not  g731 (n756, n718);
not  g732 (n749, n722);
not  g733 (n747, n720);
not  g734 (n748, n711);
not  g735 (n759, n714);
not  g736 (n758, n726);
not  g737 (n753, n724);
not  g738 (n760, n712);
not  g739 (n801, n744);
buf  g740 (n818, n538);
not  g741 (n810, n745);
not  g742 (n808, n520);
not  g743 (n814, n734);
buf  g744 (n821, n756);
not  g745 (n816, n541);
buf  g746 (n786, n751);
buf  g747 (n823, n548);
not  g748 (n765, n753);
not  g749 (n773, n745);
not  g750 (n794, n751);
not  g751 (n793, n750);
not  g752 (n770, n751);
buf  g753 (n817, n741);
buf  g754 (n798, n543);
not  g755 (n781, n753);
not  g756 (n788, n741);
buf  g757 (n800, n552);
buf  g758 (n766, n524);
not  g759 (n779, n523);
not  g760 (n802, n750);
not  g761 (n796, n742);
not  g762 (n790, n521);
buf  g763 (n769, n749);
buf  g764 (n775, n747);
not  g765 (n764, n528);
not  g766 (n797, n540);
not  g767 (n812, n756);
not  g768 (n782, n745);
buf  g769 (n776, n747);
buf  g770 (n763, n752);
not  g771 (n771, n743);
buf  g772 (n807, n549);
not  g773 (n813, n547);
not  g774 (n787, n741);
buf  g775 (n806, n533);
not  g776 (n811, n530);
buf  g777 (n809, n738);
not  g778 (n767, n518);
buf  g779 (n819, n516);
not  g780 (n804, n527);
and  g781 (n792, n746, n551, n757, n748);
nor  g782 (n778, n739, n744, n748, n732);
xor  g783 (n805, n537, n755, n546, n522);
nand g784 (n820, n536, n753, n757, n745);
or   g785 (n789, n755, n735, n535, n743);
nand g786 (n783, n754, n733, n532, n517);
and  g787 (n815, n751, n756, n746, n748);
and  g788 (n822, n748, n553, n747, n529);
xor  g789 (n774, n550, n757, n746, n754);
xnor g790 (n768, n555, n525, n526, n531);
xor  g791 (n780, n746, n752, n754, n554);
nand g792 (n777, n740, n545, n534, n736);
or   g793 (n784, n756, n755, n753, n750);
xnor g794 (n785, n749, n749, n737, n731);
nand g795 (n795, n752, n758, n744, n743);
nor  g796 (n791, n757, n519, n743, n539);
nor  g797 (n803, n747, n742, n752, n542);
xor  g798 (n799, n741, n744, n740, n754);
xnor g799 (n772, n749, n750, n544, n755);
buf  g800 (n867, n570);
buf  g801 (n837, n458);
not  g802 (n858, n454);
not  g803 (n856, n598);
buf  g804 (n834, n467);
not  g805 (n859, n473);
xor  g806 (n833, n784, n592, n794, n476);
xor  g807 (n826, n450, n472, n772, n580);
nor  g808 (n868, n785, n768, n808, n562);
nor  g809 (n882, n449, n461, n472, n465);
or   g810 (n852, n579, n469, n468);
xnor g811 (n869, n472, n587, n810, n556);
and  g812 (n831, n822, n593, n468, n795);
nand g813 (n848, n475, n460, n456);
nand g814 (n847, n455, n458, n758, n804);
and  g815 (n832, n459, n817, n816, n796);
xnor g816 (n830, n465, n459, n470, n809);
xnor g817 (n884, n563, n451, n813, n452);
xor  g818 (n866, n814, n823, n818, n450);
nor  g819 (n865, n449, n597, n461, n805);
nand g820 (n861, n448, n797, n771, n578);
nor  g821 (n829, n758, n455, n470, n557);
nor  g822 (n851, n450, n464, n759, n448);
nor  g823 (n843, n590, n585, n467);
xnor g824 (n881, n476, n571, n802, n798);
xor  g825 (n879, n453, n451, n474, n788);
nor  g826 (n877, n470, n591, n473, n451);
nand g827 (n842, n589, n764, n453, n807);
nand g828 (n876, n779, n469, n477, n594);
and  g829 (n840, n786, n577, n584, n462);
xor  g830 (n878, n799, n778, n475, n561);
and  g831 (n870, n811, n458, n776, n473);
or   g832 (n874, n783, n758, n450, n567);
nand g833 (n863, n449, n466, n789, n456);
nor  g834 (n827, n457, n454, n467, n560);
xor  g835 (n846, n472, n466, n474, n458);
nand g836 (n845, n806, n581, n568, n462);
or   g837 (n854, n576, n582, n463, n787);
xor  g838 (n883, n466, n452, n460, n453);
nor  g839 (n862, n558, n766, n469, n765);
nor  g840 (n875, n574, n453, n575, n463);
and  g841 (n872, n572, n759, n457, n821);
xnor g842 (n864, n460, n763, n566, n803);
and  g843 (n839, n464, n596, n792, n461);
xor  g844 (n838, n464, n449, n473, n476);
or   g845 (n849, n815, n455, n793);
xnor g846 (n825, n586, n463, n475, n460);
xor  g847 (n841, n583, n565, n465, n595);
nor  g848 (n873, n559, n448, n474, n465);
and  g849 (n828, n790, n461, n454, n777);
nand g850 (n836, n463, n471, n800, n464);
or   g851 (n835, n781, n474, n471, n564);
nor  g852 (n880, n770, n791, n780, n469);
xor  g853 (n853, n773, n451, n782, n452);
xnor g854 (n857, n819, n459, n573, n569);
or   g855 (n871, n470, n774, n466, n459);
xnor g856 (n850, n769, n476, n452, n448);
nor  g857 (n860, n471, n457, n767, n462);
or   g858 (n855, n462, n801, n454, n468);
nand g859 (n824, n471, n588, n820, n475);
xor  g860 (n844, n457, n775, n456, n812);
buf  g861 (n953, n610);
buf  g862 (n888, n826);
buf  g863 (n915, n857);
buf  g864 (n949, n617);
not  g865 (n933, n833);
not  g866 (n889, n634);
not  g867 (n922, n846);
buf  g868 (n967, n841);
buf  g869 (n886, n843);
buf  g870 (n904, n850);
not  g871 (n961, n846);
buf  g872 (n979, n826);
buf  g873 (n891, n833);
not  g874 (n958, n853);
buf  g875 (n962, n843);
not  g876 (n893, n841);
buf  g877 (n902, n854);
buf  g878 (n931, n845);
not  g879 (n927, n850);
buf  g880 (n963, n847);
not  g881 (n978, n852);
not  g882 (n945, n834);
buf  g883 (n950, n621);
not  g884 (n926, n840);
not  g885 (n914, n825);
buf  g886 (n955, n632);
buf  g887 (n912, n633);
not  g888 (n906, n825);
buf  g889 (n952, n853);
not  g890 (n939, n625);
not  g891 (n923, n840);
buf  g892 (n897, n840);
not  g893 (n918, n836);
buf  g894 (n930, n842);
buf  g895 (n917, n606);
not  g896 (n894, n603);
not  g897 (n916, n840);
buf  g898 (n934, n852);
not  g899 (n970, n854);
buf  g900 (n890, n851);
not  g901 (n959, n824);
buf  g902 (n980, n837);
buf  g903 (n972, n847);
not  g904 (n948, n612);
not  g905 (n907, n844);
buf  g906 (n947, n827);
buf  g907 (n909, n848);
not  g908 (n957, n827);
not  g909 (n941, n834);
not  g910 (n946, n627);
not  g911 (n975, n849);
not  g912 (n966, n611);
not  g913 (n954, n858);
not  g914 (n938, n835);
not  g915 (n977, n830);
not  g916 (n956, n845);
not  g917 (n895, n623);
buf  g918 (n885, n624);
not  g919 (n965, n851);
buf  g920 (n896, n619);
not  g921 (n900, n839);
not  g922 (n937, n857);
not  g923 (n942, n834);
buf  g924 (n932, n852);
not  g925 (n944, n853);
buf  g926 (n976, n841);
buf  g927 (n943, n855);
buf  g928 (n969, n836);
buf  g929 (n921, n850);
buf  g930 (n973, n608);
xor  g931 (n935, n832, n838, n849, n847);
and  g932 (n892, n626, n829, n844, n848);
and  g933 (n903, n839, n828, n629, n615);
nand g934 (n920, n857, n829, n601, n841);
nor  g935 (n928, n829, n829, n852, n855);
xor  g936 (n929, n837, n602, n635, n827);
or   g937 (n887, n836, n848, n824, n856);
xor  g938 (n968, n834, n599, n849, n836);
or   g939 (n924, n830, n848, n628, n838);
or   g940 (n901, n837, n844, n846, n616);
xor  g941 (n936, n849, n855, n842, n828);
nor  g942 (n899, n622, n607, n831, n609);
and  g943 (n911, n828, n832, n855, n833);
xnor g944 (n964, n856, n839, n832, n631);
xnor g945 (n951, n828, n856, n843, n857);
nor  g946 (n925, n853, n825, n835, n854);
xnor g947 (n960, n605, n838, n845, n614);
and  g948 (n974, n826, n838, n851, n831);
or   g949 (n898, n839, n604, n835, n850);
xnor g950 (n940, n600, n824, n831, n613);
and  g951 (n905, n844, n842, n830, n833);
xor  g952 (n971, n826, n847, n835, n832);
and  g953 (n919, n618, n842, n825, n831);
or   g954 (n913, n854, n851, n824, n830);
and  g955 (n910, n846, n843, n837, n827);
xor  g956 (n908, n630, n856, n845, n620);
xnor g957 (n1012, n872, n865, n860, n893);
xor  g958 (n1008, n933, n944, n874, n909);
nand g959 (n997, n919, n927, n876, n898);
nand g960 (n1003, n899, n877, n872, n878);
xor  g961 (n1013, n861, n859, n945, n873);
nor  g962 (n986, n875, n866, n938);
xor  g963 (n1015, n871, n895, n929, n940);
xor  g964 (n1009, n879, n874, n942, n941);
xnor g965 (n990, n905, n863, n930, n888);
nand g966 (n982, n932, n870, n879, n892);
and  g967 (n995, n865, n858, n866, n876);
nor  g968 (n1016, n939, n860, n934, n859);
or   g969 (n981, n868, n870, n931, n860);
nand g970 (n1004, n928, n862, n911, n858);
xor  g971 (n1011, n907, n863, n947, n918);
xor  g972 (n993, n878, n877, n923, n912);
xnor g973 (n984, n894, n878, n868, n900);
nand g974 (n999, n914, n946, n876, n864);
and  g975 (n1002, n902, n861, n863, n876);
and  g976 (n988, n875, n878, n877, n915);
nor  g977 (n1006, n867, n859, n887, n910);
nor  g978 (n983, n874, n862, n864, n872);
xnor g979 (n998, n903, n867, n859);
nor  g980 (n991, n871, n864, n913, n890);
or   g981 (n992, n937, n858, n901, n868);
nor  g982 (n985, n922, n866, n874, n873);
xor  g983 (n989, n925, n935, n870, n865);
nor  g984 (n1005, n875, n896, n865, n908);
or   g985 (n1001, n861, n862, n916, n870);
nor  g986 (n1014, n871, n943, n869, n936);
or   g987 (n994, n906, n863, n868, n872);
xor  g988 (n1000, n924, n904, n889, n886);
nand g989 (n987, n862, n917, n873, n867);
nand g990 (n996, n869, n869, n877, n920);
nor  g991 (n1017, n875, n926, n873, n864);
nor  g992 (n1010, n921, n885, n869, n860);
xor  g993 (n1007, n861, n891, n897, n871);
not  g994 (n1021, n1002);
buf  g995 (n1018, n1003);
buf  g996 (n1019, n1004);
buf  g997 (n1020, n1005);
nor  g998 (n1030, n644, n1012, n641, n646);
and  g999 (n1022, n1018, n639, n647, n1013);
xnor g1000 (n1027, n645, n652, n648, n1019);
nor  g1001 (n1028, n1007, n636, n1011, n651);
nor  g1002 (n1031, n1020, n948, n1009, n642);
xnor g1003 (n1024, n1015, n649, n650, n637);
xor  g1004 (n1023, n643, n1010, n1018, n1019);
or   g1005 (n1026, n1018, n638, n1014, n640);
and  g1006 (n1029, n1020, n1016, n1017, n1019);
nand g1007 (n1025, n1019, n1006, n1018, n1008);
or   g1008 (n1032, n1031, n478, n1030);
xnor g1009 (n1033, n478, n477);
buf  g1010 (n1039, n1033);
buf  g1011 (n1034, n1033);
not  g1012 (n1037, n1033);
buf  g1013 (n1040, n1032);
buf  g1014 (n1036, n1032);
buf  g1015 (n1038, n1032);
not  g1016 (n1035, n1032);
xor  g1017 (n1041, n951, n653);
xor  g1018 (n1047, n953, n655, n956);
nor  g1019 (n1043, n742, n1037, n1036);
nand g1020 (n1048, n1038, n656, n1040);
xnor g1021 (n1042, n654, n949, n1039);
nor  g1022 (n1046, n1035, n957, n1033);
or   g1023 (n1049, n1034, n954, n958);
nand g1024 (n1045, n1039, n952, n1038);
xor  g1025 (n1044, n478, n950, n955);
not  g1026 (n1055, n479);
xnor g1027 (n1054, n1049, n961, n959);
nand g1028 (n1058, n962, n1049, n1044);
or   g1029 (n1056, n479, n657, n1040);
or   g1030 (n1052, n1047, n1040);
and  g1031 (n1050, n1045, n963, n879);
xor  g1032 (n1053, n965, n880, n964);
xnor g1033 (n1059, n1042, n1041, n1046);
xnor g1034 (n1051, n1048, n960, n879);
nor  g1035 (n1057, n966, n479, n1043);
not  g1036 (n1064, n1050);
buf  g1037 (n1063, n1052);
not  g1038 (n1061, n1053);
buf  g1039 (n1062, n968);
buf  g1040 (n1067, n1051);
not  g1041 (n1066, n967);
not  g1042 (n1060, n1050);
and  g1043 (n1065, n1051, n1053, n1052);
not  g1044 (n1082, n1056);
buf  g1045 (n1076, n658);
not  g1046 (n1084, n1055);
not  g1047 (n1080, n1057);
buf  g1048 (n1078, n481);
not  g1049 (n1081, n659);
not  g1050 (n1072, n1061);
and  g1051 (n1069, n1064, n1063, n1062, n1061);
nand g1052 (n1083, n1063, n480, n1060, n665);
and  g1053 (n1074, n1063, n668, n667, n1056);
or   g1054 (n1070, n1062, n1062, n662, n661);
nand g1055 (n1079, n1062, n480, n1057, n1054);
nand g1056 (n1073, n1059, n479, n480, n1060);
nand g1057 (n1068, n660, n1064, n1054, n1058);
xnor g1058 (n1075, n663, n1059, n1063, n1061);
nand g1059 (n1071, n666, n1058, n664, n1061);
xor  g1060 (n1077, n481, n1060, n1055, n480);
not  g1061 (n1091, n1064);
not  g1062 (n1096, n1072);
buf  g1063 (n1093, n481);
not  g1064 (n1095, n1070);
not  g1065 (n1085, n669);
not  g1066 (n1100, n1080);
buf  g1067 (n1097, n1067);
not  g1068 (n1092, n1066);
and  g1069 (n1087, n1075, n1065);
nor  g1070 (n1086, n1067, n1084, n1065);
nand g1071 (n1088, n1069, n1082, n670);
nand g1072 (n1094, n1068, n1065, n1071);
nor  g1073 (n1089, n1079, n1066, n1078);
or   g1074 (n1099, n1066, n1073, n1074);
xor  g1075 (n1098, n671, n1064, n1076);
or   g1076 (n1090, n1067, n1066, n969);
and  g1077 (n1101, n1077, n1083, n1067, n1081);
not  g1078 (n1104, n1086);
buf  g1079 (n1105, n1088);
buf  g1080 (n1103, n1087);
buf  g1081 (n1102, n1085);
xnor g1082 (n1116, n683, n1102, n686, n687);
nand g1083 (n1118, n1095, n698, n1104, n695);
xnor g1084 (n1119, n709, n674, n676, n1090);
nor  g1085 (n1112, n1094, n689, n707, n1104);
nand g1086 (n1117, n694, n708, n1105, n1093);
nor  g1087 (n1107, n682, n1089, n696, n1103);
nor  g1088 (n1115, n1105, n675, n1103, n702);
xnor g1089 (n1111, n692, n701, n677, n679);
or   g1090 (n1108, n680, n681, n1102, n1105);
or   g1091 (n1106, n699, n700, n688, n1105);
nand g1092 (n1121, n684, n1097, n691, n1091);
xnor g1093 (n1120, n1104, n697, n690, n1092);
nor  g1094 (n1109, n703, n672, n693, n705);
and  g1095 (n1113, n685, n1102, n1096, n1104);
nor  g1096 (n1114, n1102, n704, n1098, n706);
nand g1097 (n1110, n673, n1103, n678);
buf  g1098 (n1146, n1120);
buf  g1099 (n1132, n1113);
buf  g1100 (n1125, n1117);
buf  g1101 (n1138, n1117);
buf  g1102 (n1124, n1120);
buf  g1103 (n1135, n1119);
buf  g1104 (n1129, n1119);
buf  g1105 (n1144, n1116);
not  g1106 (n1128, n1106);
buf  g1107 (n1139, n1118);
not  g1108 (n1133, n1108);
not  g1109 (n1142, n1119);
not  g1110 (n1131, n1117);
buf  g1111 (n1151, n1109);
buf  g1112 (n1123, n1118);
not  g1113 (n1147, n1120);
not  g1114 (n1141, n1118);
buf  g1115 (n1140, n1117);
not  g1116 (n1136, n1121);
not  g1117 (n1126, n1121);
buf  g1118 (n1145, n1118);
buf  g1119 (n1149, n1119);
not  g1120 (n1134, n1114);
buf  g1121 (n1122, n1121);
not  g1122 (n1137, n1111);
not  g1123 (n1127, n1120);
not  g1124 (n1130, n1115);
buf  g1125 (n1143, n1107);
buf  g1126 (n1148, n1112);
buf  g1127 (n1150, n1110);
not  g1128 (n1152, n1122);
not  g1129 (n1153, n1123);
buf  g1130 (n1156, n1153);
xor  g1131 (n1160, n1153, n1126, n1129);
and  g1132 (n1154, n1152, n1133, n1128, n1134);
nand g1133 (n1157, n1135, n1141, n1132, n1130);
nor  g1134 (n1155, n1139, n1143, n1138, n1153);
xor  g1135 (n1158, n1152, n1131, n1136, n1127);
nor  g1136 (n1159, n1124, n1137, n1152);
nor  g1137 (n1161, n1125, n1142, n1140, n1153);
and  g1138 (n1164, n482, n482, n1155, n483);
or   g1139 (n1163, n1154, n482, n483);
and  g1140 (n1162, n481, n1154, n483);
and  g1141 (n1169, n1164, n1163, n1158, n1155);
or   g1142 (n1167, n1158, n972, n1159, n1163);
xor  g1143 (n1166, n1156, n970, n973, n1160);
or   g1144 (n1168, n971, n1156, n1164, n1162);
nand g1145 (n1165, n1159, n1157, n974);
not  g1146 (n1173, n1166);
not  g1147 (n1176, n1165);
buf  g1148 (n1172, n1166);
not  g1149 (n1174, n1165);
buf  g1150 (n1170, n1165);
not  g1151 (n1171, n1166);
not  g1152 (n1175, n1165);
nand g1153 (n1197, n1020, n1168, n1172);
and  g1154 (n1186, n975, n977, n1176, n761);
or   g1155 (n1183, n1172, n1161, n762, n1167);
nor  g1156 (n1195, n1021, n1161, n1175, n1160);
xor  g1157 (n1177, n1170, n759, n1166, n760);
nor  g1158 (n1187, n1173, n978, n1167);
nor  g1159 (n1180, n1168, n882, n1171, n1173);
and  g1160 (n1196, n761, n1021, n1175, n1169);
nand g1161 (n1188, n1175, n1169, n1168, n1176);
and  g1162 (n1191, n976, n880, n760);
and  g1163 (n1189, n1101, n1021, n762, n1100);
xnor g1164 (n1182, n1172, n1174, n1169, n1170);
xor  g1165 (n1178, n761, n759, n1170);
and  g1166 (n1193, n881, n1099, n1171, n762);
xor  g1167 (n1184, n1174, n1121, n881);
xnor g1168 (n1185, n1176, n742, n1100, n979);
xnor g1169 (n1190, n1169, n762, n1172, n1171);
or   g1170 (n1181, n1173, n881, n1171, n761);
or   g1171 (n1194, n1176, n1101, n1173, n1021);
or   g1172 (n1179, n880, n1174, n760, n1020);
nor  g1173 (n1192, n1167, n880, n1174, n1175);
buf  g1174 (n1198, n1179);
buf  g1175 (n1202, n1181);
buf  g1176 (n1201, n1180);
buf  g1177 (n1199, n1182);
not  g1178 (n1200, n1183);
nor  g1179 (n1213, n883, n980, n882, n1201);
nand g1180 (n1204, n1191, n882, n1199, n710);
and  g1181 (n1203, n1201, n1190, n1146, n1150);
xor  g1182 (n1206, n1200, n883);
and  g1183 (n1211, n1193, n1200, n1201, n1198);
xnor g1184 (n1210, n1147, n1148, n884, n1201);
xnor g1185 (n1209, n1145, n1149, n1198, n882);
xnor g1186 (n1205, n1199, n1198, n1188, n1189);
xor  g1187 (n1214, n1192, n884, n1202, n1199);
or   g1188 (n1208, n884, n1194, n1197, n1198);
xnor g1189 (n1212, n1185, n884, n1199, n1184);
nor  g1190 (n1215, n1187, n1196, n883, n1186);
or   g1191 (n1207, n1200, n1195, n1144, n1151);
xnor g1192 (n1219, n1215, n1212, n1202);
or   g1193 (n1217, n1210, n1208, n1207, n1214);
xor  g1194 (n1216, n1211, n1213, n1205, n1203);
and  g1195 (n1218, n1204, n1202, n1206, n1209);
xnor g1196 (n1220, n1219, n1218, n1217, n1216);
endmodule
