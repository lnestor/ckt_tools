

module Stat_100_510
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n86,
  n96,
  n117,
  n111,
  n81,
  n80,
  n108,
  n97,
  n92,
  n85,
  n94,
  n93,
  n106,
  n114,
  n107,
  n104,
  n95,
  n113,
  n102,
  n110,
  n90,
  n84,
  n82,
  n91,
  n88,
  n83,
  n118,
  n101,
  n105,
  n100,
  n132,
  n131,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n86;
  output n96;
  output n117;
  output n111;
  output n81;
  output n80;
  output n108;
  output n97;
  output n92;
  output n85;
  output n94;
  output n93;
  output n106;
  output n114;
  output n107;
  output n104;
  output n95;
  output n113;
  output n102;
  output n110;
  output n90;
  output n84;
  output n82;
  output n91;
  output n88;
  output n83;
  output n118;
  output n101;
  output n105;
  output n100;
  output n132;
  output n131;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n87;
  wire n89;
  wire n98;
  wire n99;
  wire n103;
  wire n109;
  wire n112;
  wire n115;
  wire n116;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire KeyWire_0_0;
  wire KeyNOTWire_0_0;
  wire KeyWire_0_1;
  wire KeyNOTWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyNOTWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;

  not
  g0
  (
    n38,
    n13
  );


  not
  g1
  (
    n48,
    n13
  );


  buf
  g2
  (
    n37,
    n25
  );


  not
  g3
  (
    n52,
    n27
  );


  not
  g4
  (
    n71,
    n25
  );


  buf
  g5
  (
    n54,
    n14
  );


  buf
  g6
  (
    n50,
    n8
  );


  buf
  g7
  (
    n55,
    n14
  );


  buf
  g8
  (
    n56,
    n20
  );


  buf
  g9
  (
    KeyWire_0_11,
    n1
  );


  not
  g10
  (
    KeyWire_0_15,
    n10
  );


  buf
  g11
  (
    n74,
    n17
  );


  not
  g12
  (
    n40,
    n19
  );


  not
  g13
  (
    n53,
    n30
  );


  not
  g14
  (
    n75,
    n25
  );


  not
  g15
  (
    n68,
    n18
  );


  buf
  g16
  (
    n76,
    n30
  );


  buf
  g17
  (
    n42,
    n31
  );


  not
  g18
  (
    n61,
    n10
  );


  buf
  g19
  (
    n77,
    n4
  );


  buf
  g20
  (
    n46,
    n16
  );


  or
  g21
  (
    n59,
    n10,
    n3,
    n23
  );


  and
  g22
  (
    n36,
    n23,
    n1,
    n20,
    n30
  );


  and
  g23
  (
    n66,
    n29,
    n26,
    n14,
    n13
  );


  xor
  g24
  (
    KeyWire_0_3,
    n17,
    n2,
    n23,
    n24
  );


  and
  g25
  (
    n57,
    n19,
    n31,
    n28,
    n7
  );


  xor
  g26
  (
    n79,
    n17,
    n26,
    n31,
    n3
  );


  and
  g27
  (
    n62,
    n9,
    n11,
    n22,
    n3
  );


  xnor
  g28
  (
    KeyWire_0_1,
    n6,
    n15,
    n28,
    n16
  );


  nor
  g29
  (
    n45,
    n6,
    n19,
    n18,
    n1
  );


  xor
  g30
  (
    KeyWire_0_2,
    n10,
    n4,
    n8,
    n16
  );


  xnor
  g31
  (
    n43,
    n18,
    n9,
    n22,
    n14
  );


  nand
  g32
  (
    n67,
    n24,
    n12,
    n23,
    n29
  );


  xor
  g33
  (
    n33,
    n11,
    n5,
    n25
  );


  xor
  g34
  (
    n41,
    n24,
    n11,
    n12,
    n5
  );


  and
  g35
  (
    KeyWire_0_9,
    n21,
    n29,
    n18,
    n7
  );


  nand
  g36
  (
    n51,
    n9,
    n6
  );


  and
  g37
  (
    n72,
    n12,
    n21,
    n19
  );


  nand
  g38
  (
    n70,
    n5,
    n20,
    n17,
    n1
  );


  nand
  g39
  (
    KeyWire_0_5,
    n22,
    n2,
    n16,
    n24
  );


  and
  g40
  (
    n73,
    n27,
    n28,
    n11,
    n13
  );


  nand
  g41
  (
    n60,
    n29,
    n3,
    n8
  );


  nand
  g42
  (
    n39,
    n15,
    n22,
    n7,
    n27
  );


  nand
  g43
  (
    n58,
    n4,
    n30,
    n28,
    n31
  );


  nor
  g44
  (
    n78,
    n12,
    n20,
    n15
  );


  nand
  g45
  (
    KeyWire_0_8,
    n4,
    n2,
    n27,
    n21
  );


  nand
  g46
  (
    n49,
    n2,
    n26,
    n7
  );


  nor
  g47
  (
    n94,
    n53,
    n58,
    n51,
    n52
  );


  or
  g48
  (
    KeyWire_0_0,
    n50,
    n67,
    n45,
    n59
  );


  nor
  g49
  (
    n97,
    n63,
    n53,
    n59,
    n70
  );


  nand
  g50
  (
    n114,
    n41,
    n64,
    n38,
    n74
  );


  nor
  g51
  (
    n81,
    n69,
    n68,
    n66,
    n48
  );


  or
  g52
  (
    n117,
    n46,
    n58,
    n52,
    n65
  );


  or
  g53
  (
    n116,
    n39,
    n36,
    n75,
    n43
  );


  xnor
  g54
  (
    n104,
    n73,
    n52,
    n57,
    n60
  );


  xnor
  g55
  (
    n110,
    n71,
    n65,
    n60,
    n77
  );


  or
  g56
  (
    n86,
    n78,
    n54,
    n43,
    n53
  );


  or
  g57
  (
    n109,
    n48,
    n78,
    n47,
    n67
  );


  xnor
  g58
  (
    n102,
    n48,
    n56,
    n50,
    n78
  );


  xnor
  g59
  (
    n83,
    n55,
    n47,
    n70,
    n74
  );


  xor
  g60
  (
    KeyWire_0_10,
    n54,
    n77,
    n62,
    n47
  );


  nand
  g61
  (
    KeyWire_0_4,
    n62,
    n67,
    n76,
    n42
  );


  nor
  g62
  (
    n118,
    n61,
    n75,
    n76,
    n34
  );


  xor
  g63
  (
    n100,
    n38,
    n56,
    n55,
    n68
  );


  and
  g64
  (
    n101,
    n41,
    n76,
    n64,
    n75
  );


  or
  g65
  (
    n88,
    n61,
    n66,
    n37,
    n73
  );


  xnor
  g66
  (
    n113,
    n45,
    n46,
    n56,
    n77
  );


  nor
  g67
  (
    n92,
    n58,
    n73,
    n51
  );


  or
  g68
  (
    n87,
    n79,
    n60,
    n66,
    n40
  );


  nor
  g69
  (
    n90,
    n57,
    n50,
    n73,
    n48
  );


  xor
  g70
  (
    n106,
    n64,
    n59,
    n39,
    n57
  );


  xnor
  g71
  (
    n103,
    n60,
    n63,
    n55,
    n36
  );


  nand
  g72
  (
    KeyWire_0_13,
    n51,
    n69,
    n74,
    n59
  );


  xnor
  g73
  (
    n89,
    n68,
    n37,
    n54,
    n50
  );


  or
  g74
  (
    n95,
    n49,
    n74,
    n79,
    n75
  );


  nand
  g75
  (
    n84,
    n78,
    n64,
    n61,
    n70
  );


  nor
  g76
  (
    n119,
    n35,
    n72,
    n79,
    n52
  );


  or
  g77
  (
    n91,
    n57,
    n35,
    n49,
    n71
  );


  nand
  g78
  (
    n108,
    n58,
    n33,
    n44,
    n62
  );


  nand
  g79
  (
    KeyWire_0_14,
    n44,
    n61,
    n33,
    n65
  );


  xnor
  g80
  (
    n93,
    n66,
    n67,
    n53,
    n49
  );


  nand
  g81
  (
    n82,
    n69,
    n55,
    n72,
    n70
  );


  nand
  g82
  (
    n105,
    n77,
    n68,
    n40,
    n65
  );


  and
  g83
  (
    n96,
    n62,
    n71,
    n34,
    n49
  );


  nor
  g84
  (
    n99,
    n47,
    n79,
    n69,
    n71
  );


  nor
  g85
  (
    n112,
    n72,
    n63,
    n76,
    n54
  );


  and
  g86
  (
    n98,
    n56,
    n72,
    n42,
    n63
  );


  buf
  g87
  (
    n122,
    n111
  );


  not
  g88
  (
    KeyWire_0_7,
    n114
  );


  buf
  g89
  (
    n124,
    n113
  );


  not
  g90
  (
    KeyWire_0_12,
    n112
  );


  not
  g91
  (
    n120,
    n110
  );


  nor
  g92
  (
    n129,
    n121,
    n123,
    n117
  );


  or
  g93
  (
    n130,
    n124,
    n32,
    n122,
    n115
  );


  xnor
  g94
  (
    n127,
    n121,
    n119,
    n32,
    n120
  );


  or
  g95
  (
    n128,
    n124,
    n32
  );


  xor
  g96
  (
    n126,
    n121,
    n120,
    n124,
    n118
  );


  and
  g97
  (
    n125,
    n116,
    n123,
    n122
  );


  xor
  g98
  (
    KeyWire_0_6,
    n128,
    n130,
    n129,
    n126
  );


  xnor
  g99
  (
    n131,
    n127,
    n130,
    n129,
    n125
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n80,
    KeyNOTWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n63,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n35,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n34,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n107,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n44,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    KeyNOTWire_0_6,
    keyIn_0_6,
    KeyWire_0_6
  );


  not
  KeyNOTGate_0_6
  (
    n132,
    KeyNOTWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n121,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n47,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n64,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n111,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n65,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n123,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n85,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n115,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n69,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule

