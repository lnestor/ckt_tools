// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\5_24_randomized_params\Stat_1336_14_6 written by SynthGen on 2021/05/24 19:42:18
module Stat_1336_14_6( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17,
 n1341, n1337, n1336, n1346, n1345, n1351, n1342, n1347,
 n1350, n1334, n1353, n1343, n1335, n1352, n1331, n1330,
 n1338, n1332, n1333, n1339, n1348, n1340, n1349, n1344);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17;

output n1341, n1337, n1336, n1346, n1345, n1351, n1342, n1347,
 n1350, n1334, n1353, n1343, n1335, n1352, n1331, n1330,
 n1338, n1332, n1333, n1339, n1348, n1340, n1349, n1344;

wire n18, n19, n20, n21, n22, n23, n24, n25,
 n26, n27, n28, n29, n30, n31, n32, n33,
 n34, n35, n36, n37, n38, n39, n40, n41,
 n42, n43, n44, n45, n46, n47, n48, n49,
 n50, n51, n52, n53, n54, n55, n56, n57,
 n58, n59, n60, n61, n62, n63, n64, n65,
 n66, n67, n68, n69, n70, n71, n72, n73,
 n74, n75, n76, n77, n78, n79, n80, n81,
 n82, n83, n84, n85, n86, n87, n88, n89,
 n90, n91, n92, n93, n94, n95, n96, n97,
 n98, n99, n100, n101, n102, n103, n104, n105,
 n106, n107, n108, n109, n110, n111, n112, n113,
 n114, n115, n116, n117, n118, n119, n120, n121,
 n122, n123, n124, n125, n126, n127, n128, n129,
 n130, n131, n132, n133, n134, n135, n136, n137,
 n138, n139, n140, n141, n142, n143, n144, n145,
 n146, n147, n148, n149, n150, n151, n152, n153,
 n154, n155, n156, n157, n158, n159, n160, n161,
 n162, n163, n164, n165, n166, n167, n168, n169,
 n170, n171, n172, n173, n174, n175, n176, n177,
 n178, n179, n180, n181, n182, n183, n184, n185,
 n186, n187, n188, n189, n190, n191, n192, n193,
 n194, n195, n196, n197, n198, n199, n200, n201,
 n202, n203, n204, n205, n206, n207, n208, n209,
 n210, n211, n212, n213, n214, n215, n216, n217,
 n218, n219, n220, n221, n222, n223, n224, n225,
 n226, n227, n228, n229, n230, n231, n232, n233,
 n234, n235, n236, n237, n238, n239, n240, n241,
 n242, n243, n244, n245, n246, n247, n248, n249,
 n250, n251, n252, n253, n254, n255, n256, n257,
 n258, n259, n260, n261, n262, n263, n264, n265,
 n266, n267, n268, n269, n270, n271, n272, n273,
 n274, n275, n276, n277, n278, n279, n280, n281,
 n282, n283, n284, n285, n286, n287, n288, n289,
 n290, n291, n292, n293, n294, n295, n296, n297,
 n298, n299, n300, n301, n302, n303, n304, n305,
 n306, n307, n308, n309, n310, n311, n312, n313,
 n314, n315, n316, n317, n318, n319, n320, n321,
 n322, n323, n324, n325, n326, n327, n328, n329,
 n330, n331, n332, n333, n334, n335, n336, n337,
 n338, n339, n340, n341, n342, n343, n344, n345,
 n346, n347, n348, n349, n350, n351, n352, n353,
 n354, n355, n356, n357, n358, n359, n360, n361,
 n362, n363, n364, n365, n366, n367, n368, n369,
 n370, n371, n372, n373, n374, n375, n376, n377,
 n378, n379, n380, n381, n382, n383, n384, n385,
 n386, n387, n388, n389, n390, n391, n392, n393,
 n394, n395, n396, n397, n398, n399, n400, n401,
 n402, n403, n404, n405, n406, n407, n408, n409,
 n410, n411, n412, n413, n414, n415, n416, n417,
 n418, n419, n420, n421, n422, n423, n424, n425,
 n426, n427, n428, n429, n430, n431, n432, n433,
 n434, n435, n436, n437, n438, n439, n440, n441,
 n442, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n608, n609,
 n610, n611, n612, n613, n614, n615, n616, n617,
 n618, n619, n620, n621, n622, n623, n624, n625,
 n626, n627, n628, n629, n630, n631, n632, n633,
 n634, n635, n636, n637, n638, n639, n640, n641,
 n642, n643, n644, n645, n646, n647, n648, n649,
 n650, n651, n652, n653, n654, n655, n656, n657,
 n658, n659, n660, n661, n662, n663, n664, n665,
 n666, n667, n668, n669, n670, n671, n672, n673,
 n674, n675, n676, n677, n678, n679, n680, n681,
 n682, n683, n684, n685, n686, n687, n688, n689,
 n690, n691, n692, n693, n694, n695, n696, n697,
 n698, n699, n700, n701, n702, n703, n704, n705,
 n706, n707, n708, n709, n710, n711, n712, n713,
 n714, n715, n716, n717, n718, n719, n720, n721,
 n722, n723, n724, n725, n726, n727, n728, n729,
 n730, n731, n732, n733, n734, n735, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
 n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
 n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
 n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
 n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
 n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
 n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
 n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
 n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
 n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
 n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
 n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
 n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
 n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
 n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
 n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
 n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
 n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
 n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
 n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
 n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
 n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
 n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
 n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
 n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
 n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
 n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
 n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
 n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
 n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
 n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
 n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
 n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
 n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
 n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
 n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
 n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
 n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
 n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
 n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329;

not  g0 (n66, n11);
not  g1 (n40, n16);
buf  g2 (n18, n2);
not  g3 (n34, n14);
buf  g4 (n53, n7);
buf  g5 (n76, n16);
buf  g6 (n63, n16);
buf  g7 (n72, n2);
not  g8 (n50, n15);
not  g9 (n25, n1);
buf  g10 (n78, n14);
not  g11 (n35, n17);
not  g12 (n20, n10);
not  g13 (n68, n13);
not  g14 (n80, n11);
not  g15 (n48, n3);
not  g16 (n43, n17);
not  g17 (n55, n12);
buf  g18 (n27, n15);
not  g19 (n81, n4);
buf  g20 (n51, n12);
not  g21 (n60, n10);
not  g22 (n77, n11);
not  g23 (n58, n9);
not  g24 (n42, n14);
not  g25 (n73, n10);
buf  g26 (n29, n17);
not  g27 (n49, n6);
buf  g28 (n65, n4);
buf  g29 (n62, n3);
buf  g30 (n47, n12);
not  g31 (n32, n6);
buf  g32 (n31, n2);
not  g33 (n56, n8);
not  g34 (n23, n3);
buf  g35 (n83, n9);
buf  g36 (n52, n1);
buf  g37 (n44, n13);
not  g38 (n30, n16);
buf  g39 (n82, n12);
buf  g40 (n46, n9);
not  g41 (n54, n13);
buf  g42 (n24, n5);
buf  g43 (n19, n6);
buf  g44 (n70, n9);
buf  g45 (n84, n1);
buf  g46 (n75, n15);
buf  g47 (n71, n17);
buf  g48 (n39, n4);
buf  g49 (n79, n5);
not  g50 (n64, n3);
not  g51 (n41, n1);
buf  g52 (n59, n2);
buf  g53 (n45, n6);
buf  g54 (n57, n8);
not  g55 (n61, n8);
not  g56 (n69, n7);
not  g57 (n38, n11);
buf  g58 (n36, n5);
not  g59 (n22, n5);
not  g60 (n85, n7);
not  g61 (n26, n15);
not  g62 (n67, n7);
buf  g63 (n33, n13);
buf  g64 (n21, n14);
not  g65 (n28, n10);
not  g66 (n74, n8);
not  g67 (n37, n4);
buf  g68 (n123, n33);
buf  g69 (n102, n59);
not  g70 (n233, n80);
not  g71 (n106, n19);
buf  g72 (n169, n63);
not  g73 (n322, n80);
buf  g74 (n177, n60);
not  g75 (n315, n38);
buf  g76 (n202, n26);
not  g77 (n171, n85);
buf  g78 (n264, n24);
not  g79 (n303, n36);
not  g80 (n97, n55);
buf  g81 (n138, n23);
buf  g82 (n304, n50);
buf  g83 (n231, n77);
not  g84 (n154, n30);
not  g85 (n333, n84);
buf  g86 (n272, n46);
buf  g87 (n190, n37);
not  g88 (n318, n34);
buf  g89 (n161, n67);
not  g90 (n105, n44);
buf  g91 (n288, n61);
not  g92 (n227, n83);
not  g93 (n168, n27);
buf  g94 (n175, n29);
buf  g95 (n115, n49);
buf  g96 (n212, n81);
buf  g97 (n343, n68);
buf  g98 (n158, n48);
not  g99 (n95, n70);
not  g100 (n179, n66);
not  g101 (n305, n63);
not  g102 (n142, n67);
buf  g103 (n307, n41);
buf  g104 (n252, n80);
not  g105 (n324, n49);
not  g106 (n193, n76);
buf  g107 (n290, n73);
buf  g108 (n133, n65);
not  g109 (n357, n48);
buf  g110 (n98, n19);
buf  g111 (n165, n46);
buf  g112 (n295, n68);
not  g113 (n215, n50);
not  g114 (n88, n82);
not  g115 (n244, n44);
buf  g116 (n116, n34);
buf  g117 (n146, n30);
not  g118 (n336, n67);
not  g119 (n281, n71);
buf  g120 (n176, n85);
buf  g121 (n240, n41);
not  g122 (n300, n81);
buf  g123 (n124, n66);
buf  g124 (n335, n31);
not  g125 (n241, n42);
buf  g126 (n145, n69);
buf  g127 (n232, n43);
buf  g128 (n152, n41);
buf  g129 (n130, n33);
not  g130 (n329, n54);
buf  g131 (n132, n35);
not  g132 (n253, n40);
buf  g133 (n234, n56);
buf  g134 (n205, n55);
buf  g135 (n164, n75);
not  g136 (n317, n25);
not  g137 (n188, n28);
not  g138 (n274, n53);
buf  g139 (n348, n51);
not  g140 (n314, n82);
buf  g141 (n122, n35);
not  g142 (n259, n79);
buf  g143 (n269, n32);
not  g144 (n126, n83);
not  g145 (n237, n52);
not  g146 (n214, n42);
not  g147 (n277, n76);
buf  g148 (n285, n85);
not  g149 (n198, n29);
buf  g150 (n163, n19);
buf  g151 (n119, n28);
buf  g152 (n211, n65);
buf  g153 (n120, n45);
buf  g154 (n134, n64);
not  g155 (n230, n81);
buf  g156 (n207, n24);
buf  g157 (n260, n53);
not  g158 (n256, n71);
not  g159 (n181, n73);
not  g160 (n262, n50);
not  g161 (n331, n56);
buf  g162 (n249, n68);
buf  g163 (n157, n78);
buf  g164 (n287, n60);
buf  g165 (n292, n70);
buf  g166 (n127, n36);
buf  g167 (n208, n56);
not  g168 (n286, n45);
buf  g169 (n206, n84);
not  g170 (n89, n25);
buf  g171 (n121, n61);
buf  g172 (n276, n64);
not  g173 (n320, n59);
not  g174 (n239, n67);
not  g175 (n265, n83);
not  g176 (n137, n23);
not  g177 (n155, n74);
not  g178 (n312, n79);
buf  g179 (n297, n51);
buf  g180 (n342, n69);
buf  g181 (n254, n28);
buf  g182 (n337, n60);
not  g183 (n167, n66);
buf  g184 (n136, n22);
buf  g185 (n268, n82);
buf  g186 (n144, n51);
not  g187 (n345, n53);
not  g188 (n306, n39);
buf  g189 (n131, n84);
not  g190 (n243, n57);
buf  g191 (n141, n45);
not  g192 (n258, n42);
buf  g193 (n325, n64);
buf  g194 (n299, n47);
buf  g195 (n282, n65);
not  g196 (n112, n64);
not  g197 (n310, n62);
not  g198 (n294, n71);
buf  g199 (n108, n26);
buf  g200 (n151, n31);
not  g201 (n180, n24);
not  g202 (n289, n43);
not  g203 (n184, n21);
buf  g204 (n117, n47);
buf  g205 (n94, n35);
buf  g206 (n330, n21);
buf  g207 (n173, n36);
not  g208 (n327, n31);
buf  g209 (n114, n25);
buf  g210 (n223, n58);
buf  g211 (n153, n84);
not  g212 (n182, n66);
not  g213 (n356, n29);
not  g214 (n313, n24);
buf  g215 (n323, n48);
not  g216 (n326, n18);
buf  g217 (n280, n19);
not  g218 (n218, n74);
buf  g219 (n332, n30);
not  g220 (n346, n49);
buf  g221 (n220, n70);
buf  g222 (n174, n51);
buf  g223 (n156, n45);
not  g224 (n263, n39);
buf  g225 (n189, n58);
buf  g226 (n245, n30);
not  g227 (n143, n55);
not  g228 (n203, n21);
not  g229 (n226, n37);
buf  g230 (n99, n18);
not  g231 (n224, n62);
buf  g232 (n91, n75);
buf  g233 (n349, n78);
buf  g234 (n352, n39);
not  g235 (n90, n27);
buf  g236 (n311, n80);
buf  g237 (n316, n85);
buf  g238 (n135, n77);
buf  g239 (n270, n38);
not  g240 (n340, n54);
buf  g241 (n172, n33);
not  g242 (n147, n46);
not  g243 (n275, n78);
not  g244 (n103, n39);
not  g245 (n110, n29);
buf  g246 (n328, n75);
not  g247 (n187, n83);
not  g248 (n238, n63);
not  g249 (n200, n52);
buf  g250 (n266, n57);
not  g251 (n107, n20);
not  g252 (n225, n79);
not  g253 (n350, n38);
buf  g254 (n194, n49);
not  g255 (n216, n27);
not  g256 (n204, n46);
not  g257 (n92, n58);
buf  g258 (n192, n71);
buf  g259 (n93, n34);
buf  g260 (n334, n50);
not  g261 (n321, n76);
not  g262 (n104, n18);
buf  g263 (n235, n72);
not  g264 (n298, n62);
buf  g265 (n159, n52);
buf  g266 (n101, n38);
not  g267 (n278, n47);
buf  g268 (n341, n77);
not  g269 (n186, n60);
buf  g270 (n209, n54);
buf  g271 (n291, n21);
buf  g272 (n199, n33);
buf  g273 (n178, n59);
not  g274 (n148, n70);
not  g275 (n309, n69);
buf  g276 (n302, n78);
not  g277 (n109, n31);
not  g278 (n246, n44);
buf  g279 (n267, n43);
not  g280 (n221, n48);
not  g281 (n242, n55);
not  g282 (n338, n28);
buf  g283 (n354, n22);
buf  g284 (n344, n27);
buf  g285 (n255, n20);
buf  g286 (n301, n54);
buf  g287 (n283, n20);
not  g288 (n129, n59);
buf  g289 (n308, n72);
buf  g290 (n87, n52);
buf  g291 (n347, n32);
buf  g292 (n183, n43);
buf  g293 (n196, n74);
not  g294 (n273, n32);
buf  g295 (n149, n36);
buf  g296 (n296, n57);
buf  g297 (n351, n18);
not  g298 (n191, n69);
not  g299 (n247, n25);
not  g300 (n257, n53);
not  g301 (n139, n22);
buf  g302 (n217, n40);
not  g303 (n150, n68);
buf  g304 (n279, n42);
not  g305 (n355, n74);
buf  g306 (n160, n62);
not  g307 (n236, n35);
not  g308 (n128, n65);
not  g309 (n100, n20);
not  g310 (n210, n23);
buf  g311 (n166, n58);
not  g312 (n219, n63);
not  g313 (n162, n26);
not  g314 (n195, n79);
not  g315 (n319, n23);
buf  g316 (n170, n26);
not  g317 (n271, n47);
buf  g318 (n118, n37);
buf  g319 (n111, n73);
buf  g320 (n261, n77);
buf  g321 (n86, n82);
buf  g322 (n96, n40);
not  g323 (n293, n61);
buf  g324 (n229, n32);
buf  g325 (n248, n44);
buf  g326 (n201, n34);
buf  g327 (n213, n37);
not  g328 (n140, n75);
not  g329 (n250, n73);
not  g330 (n339, n22);
not  g331 (n113, n72);
buf  g332 (n185, n56);
buf  g333 (n125, n81);
not  g334 (n197, n76);
not  g335 (n284, n72);
not  g336 (n222, n57);
not  g337 (n353, n61);
buf  g338 (n251, n40);
not  g339 (n228, n41);
buf  g340 (n830, n117);
buf  g341 (n430, n86);
buf  g342 (n868, n235);
not  g343 (n861, n246);
buf  g344 (n834, n148);
not  g345 (n447, n274);
not  g346 (n681, n102);
not  g347 (n775, n139);
buf  g348 (n822, n345);
buf  g349 (n882, n351);
buf  g350 (n513, n274);
buf  g351 (n664, n292);
buf  g352 (n803, n251);
not  g353 (n812, n230);
not  g354 (n712, n111);
not  g355 (n710, n203);
buf  g356 (n836, n189);
buf  g357 (n793, n349);
buf  g358 (n888, n246);
buf  g359 (n561, n332);
buf  g360 (n363, n290);
buf  g361 (n599, n265);
not  g362 (n691, n293);
buf  g363 (n399, n331);
not  g364 (n772, n304);
buf  g365 (n508, n298);
not  g366 (n394, n190);
buf  g367 (n554, n262);
not  g368 (n719, n293);
not  g369 (n385, n163);
not  g370 (n887, n249);
buf  g371 (n751, n308);
buf  g372 (n547, n320);
not  g373 (n536, n202);
buf  g374 (n864, n92);
not  g375 (n723, n353);
buf  g376 (n413, n241);
not  g377 (n824, n261);
buf  g378 (n419, n154);
not  g379 (n813, n93);
not  g380 (n828, n244);
not  g381 (n798, n278);
buf  g382 (n627, n97);
buf  g383 (n455, n343);
buf  g384 (n382, n228);
not  g385 (n359, n158);
not  g386 (n741, n91);
buf  g387 (n545, n107);
buf  g388 (n833, n104);
not  g389 (n422, n303);
buf  g390 (n483, n350);
buf  g391 (n758, n118);
buf  g392 (n528, n224);
buf  g393 (n555, n345);
buf  g394 (n853, n143);
not  g395 (n441, n124);
not  g396 (n452, n156);
not  g397 (n552, n234);
not  g398 (n485, n302);
buf  g399 (n476, n215);
buf  g400 (n589, n313);
not  g401 (n587, n200);
not  g402 (n629, n296);
not  g403 (n506, n177);
not  g404 (n383, n231);
not  g405 (n635, n226);
buf  g406 (n880, n309);
not  g407 (n360, n254);
not  g408 (n366, n238);
not  g409 (n729, n270);
buf  g410 (n526, n246);
not  g411 (n659, n307);
not  g412 (n451, n114);
not  g413 (n425, n259);
not  g414 (n865, n234);
buf  g415 (n529, n121);
buf  g416 (n605, n195);
buf  g417 (n610, n346);
not  g418 (n489, n224);
not  g419 (n432, n106);
buf  g420 (n740, n352);
buf  g421 (n597, n341);
not  g422 (n546, n182);
not  g423 (n390, n88);
not  g424 (n661, n272);
not  g425 (n794, n270);
not  g426 (n639, n280);
not  g427 (n580, n96);
buf  g428 (n820, n335);
buf  g429 (n431, n109);
buf  g430 (n439, n142);
buf  g431 (n846, n143);
not  g432 (n746, n327);
not  g433 (n510, n166);
not  g434 (n693, n286);
not  g435 (n645, n189);
buf  g436 (n749, n312);
not  g437 (n782, n345);
buf  g438 (n512, n292);
buf  g439 (n875, n346);
not  g440 (n467, n172);
not  g441 (n755, n247);
not  g442 (n698, n146);
buf  g443 (n595, n227);
buf  g444 (n504, n226);
not  g445 (n825, n174);
buf  g446 (n827, n153);
not  g447 (n789, n257);
not  g448 (n548, n275);
not  g449 (n374, n98);
not  g450 (n896, n135);
buf  g451 (n884, n281);
buf  g452 (n801, n176);
buf  g453 (n449, n238);
buf  g454 (n396, n220);
not  g455 (n668, n354);
buf  g456 (n524, n296);
not  g457 (n666, n303);
not  g458 (n538, n228);
buf  g459 (n611, n244);
buf  g460 (n700, n236);
buf  g461 (n622, n178);
buf  g462 (n810, n227);
not  g463 (n550, n203);
not  g464 (n800, n338);
not  g465 (n401, n300);
not  g466 (n637, n141);
buf  g467 (n486, n144);
buf  g468 (n638, n178);
not  g469 (n418, n230);
not  g470 (n881, n267);
not  g471 (n500, n211);
buf  g472 (n457, n179);
buf  g473 (n609, n199);
buf  g474 (n750, n314);
not  g475 (n613, n167);
buf  g476 (n724, n186);
buf  g477 (n395, n207);
buf  g478 (n487, n140);
buf  g479 (n785, n258);
not  g480 (n721, n180);
buf  g481 (n591, n137);
not  g482 (n764, n264);
buf  g483 (n462, n133);
not  g484 (n886, n125);
buf  g485 (n835, n103);
buf  g486 (n871, n308);
buf  g487 (n615, n275);
buf  g488 (n761, n125);
buf  g489 (n706, n194);
buf  g490 (n753, n137);
buf  g491 (n603, n280);
not  g492 (n616, n137);
buf  g493 (n628, n327);
buf  g494 (n727, n230);
buf  g495 (n588, n321);
not  g496 (n762, n186);
buf  g497 (n651, n139);
buf  g498 (n665, n228);
buf  g499 (n774, n132);
buf  g500 (n598, n133);
buf  g501 (n371, n302);
not  g502 (n844, n345);
buf  g503 (n380, n101);
not  g504 (n448, n150);
not  g505 (n474, n347);
not  g506 (n873, n200);
buf  g507 (n734, n201);
buf  g508 (n477, n214);
buf  g509 (n389, n238);
not  g510 (n696, n356);
buf  g511 (n392, n259);
not  g512 (n362, n237);
buf  g513 (n454, n203);
not  g514 (n663, n339);
not  g515 (n876, n201);
buf  g516 (n444, n247);
not  g517 (n542, n254);
not  g518 (n643, n279);
buf  g519 (n565, n165);
not  g520 (n799, n307);
buf  g521 (n579, n120);
not  g522 (n652, n174);
not  g523 (n450, n169);
buf  g524 (n501, n211);
buf  g525 (n445, n269);
buf  g526 (n514, n114);
not  g527 (n517, n342);
buf  g528 (n669, n234);
buf  g529 (n409, n353);
not  g530 (n891, n338);
not  g531 (n807, n189);
not  g532 (n578, n198);
buf  g533 (n358, n209);
not  g534 (n583, n296);
not  g535 (n496, n237);
not  g536 (n373, n281);
buf  g537 (n641, n92);
buf  g538 (n688, n132);
not  g539 (n414, n275);
not  g540 (n894, n317);
not  g541 (n468, n102);
not  g542 (n657, n173);
not  g543 (n730, n279);
buf  g544 (n421, n248);
not  g545 (n567, n161);
not  g546 (n658, n252);
buf  g547 (n644, n250);
buf  g548 (n708, n318);
buf  g549 (n368, n216);
buf  g550 (n446, n271);
not  g551 (n437, n182);
buf  g552 (n671, n256);
not  g553 (n424, n274);
not  g554 (n747, n331);
not  g555 (n826, n311);
not  g556 (n403, n91);
not  g557 (n842, n208);
buf  g558 (n889, n218);
buf  g559 (n614, n225);
buf  g560 (n654, n282);
not  g561 (n662, n334);
not  g562 (n745, n268);
not  g563 (n544, n161);
not  g564 (n515, n199);
not  g565 (n686, n319);
not  g566 (n792, n242);
buf  g567 (n559, n204);
buf  g568 (n776, n342);
not  g569 (n811, n356);
buf  g570 (n640, n352);
not  g571 (n502, n240);
buf  g572 (n715, n266);
not  g573 (n535, n235);
not  g574 (n471, n325);
buf  g575 (n505, n323);
not  g576 (n849, n232);
not  g577 (n773, n128);
buf  g578 (n594, n138);
not  g579 (n634, n266);
not  g580 (n885, n171);
not  g581 (n716, n353);
buf  g582 (n707, n225);
not  g583 (n509, n173);
not  g584 (n470, n236);
not  g585 (n379, n323);
buf  g586 (n584, n282);
not  g587 (n725, n142);
not  g588 (n636, n192);
not  g589 (n530, n242);
buf  g590 (n768, n134);
not  g591 (n843, n272);
buf  g592 (n420, n170);
not  g593 (n795, n243);
not  g594 (n582, n279);
buf  g595 (n642, n349);
buf  g596 (n375, n274);
buf  g597 (n694, n300);
not  g598 (n858, n271);
not  g599 (n797, n258);
not  g600 (n893, n113);
buf  g601 (n784, n140);
not  g602 (n684, n277);
not  g603 (n819, n130);
not  g604 (n466, n168);
buf  g605 (n463, n185);
buf  g606 (n543, n256);
buf  g607 (n456, n215);
not  g608 (n402, n160);
not  g609 (n845, n136);
buf  g610 (n702, n262);
not  g611 (n631, n280);
not  g612 (n870, n203);
not  g613 (n570, n299);
buf  g614 (n673, n120);
buf  g615 (n541, n297);
buf  g616 (n831, n173);
not  g617 (n711, n252);
buf  g618 (n408, n191);
buf  g619 (n498, n229);
buf  g620 (n581, n233);
buf  g621 (n387, n350);
not  g622 (n670, n287);
buf  g623 (n577, n288);
not  g624 (n783, n172);
not  g625 (n847, n346);
not  g626 (n743, n162);
buf  g627 (n722, n221);
buf  g628 (n593, n349);
buf  g629 (n805, n222);
not  g630 (n461, n221);
not  g631 (n575, n264);
not  g632 (n416, n295);
not  g633 (n562, n324);
buf  g634 (n796, n301);
not  g635 (n623, n155);
buf  g636 (n838, n291);
not  g637 (n675, n310);
buf  g638 (n840, n273);
not  g639 (n632, n182);
buf  g640 (n484, n151);
buf  g641 (n370, n151);
not  g642 (n539, n315);
not  g643 (n841, n147);
not  g644 (n621, n192);
not  g645 (n832, n133);
buf  g646 (n464, n94);
buf  g647 (n503, n260);
buf  g648 (n735, n181);
not  g649 (n626, n211);
not  g650 (n520, n181);
buf  g651 (n771, n112);
buf  g652 (n780, n335);
buf  g653 (n697, n167);
buf  g654 (n685, n337);
buf  g655 (n458, n347);
buf  g656 (n683, n309);
buf  g657 (n619, n205);
not  g658 (n617, n169);
buf  g659 (n679, n256);
not  g660 (n839, n262);
not  g661 (n742, n237);
not  g662 (n608, n288);
not  g663 (n647, n225);
buf  g664 (n364, n200);
buf  g665 (n625, n178);
buf  g666 (n653, n244);
buf  g667 (n407, n215);
buf  g668 (n563, n295);
not  g669 (n817, n286);
buf  g670 (n862, n261);
buf  g671 (n872, n212);
not  g672 (n410, n355);
not  g673 (n411, n108);
buf  g674 (n655, n94);
buf  g675 (n633, n209);
buf  g676 (n551, n348);
not  g677 (n781, n139);
not  g678 (n600, n326);
not  g679 (n556, n248);
buf  g680 (n714, n316);
not  g681 (n415, n152);
not  g682 (n854, n170);
not  g683 (n677, n158);
not  g684 (n699, n144);
not  g685 (n571, n333);
buf  g686 (n705, n175);
not  g687 (n511, n146);
buf  g688 (n406, n213);
not  g689 (n689, n305);
not  g690 (n527, n166);
buf  g691 (n815, n201);
not  g692 (n818, n247);
not  g693 (n493, n323);
not  g694 (n660, n164);
buf  g695 (n434, n217);
buf  g696 (n404, n177);
not  g697 (n473, n204);
not  g698 (n377, n284);
buf  g699 (n537, n335);
not  g700 (n863, n332);
buf  g701 (n460, n314);
buf  g702 (n495, n153);
buf  g703 (n488, n299);
buf  g704 (n592, n210);
not  g705 (n672, n263);
buf  g706 (n786, n253);
buf  g707 (n744, n148);
buf  g708 (n895, n159);
buf  g709 (n427, n201);
not  g710 (n829, n119);
buf  g711 (n667, n311);
not  g712 (n397, n136);
buf  g713 (n808, n137);
not  g714 (n733, n273);
not  g715 (n494, n255);
not  g716 (n569, n104);
not  g717 (n850, n155);
buf  g718 (n438, n246);
buf  g719 (n766, n149);
not  g720 (n478, n299);
not  g721 (n393, n324);
not  g722 (n624, n119);
buf  g723 (n429, n213);
buf  g724 (n436, n257);
not  g725 (n472, n304);
buf  g726 (n674, n272);
buf  g727 (n890, n206);
nand g728 (n770, n166, n330, n264, n328);
or   g729 (n391, n310, n171, n276, n295);
and  g730 (n620, n127, n300, n138, n89);
nor  g731 (n823, n194, n354, n299, n164);
xor  g732 (n480, n251, n346, n204, n343);
or   g733 (n779, n170, n320, n266, n338);
xor  g734 (n720, n193, n191, n330, n339);
nand g735 (n534, n207, n160, n176);
xnor g736 (n837, n231, n231, n314, n340);
or   g737 (n748, n318, n276, n218, n161);
xnor g738 (n709, n172, n113, n252, n131);
xor  g739 (n736, n226, n217, n264, n123);
xnor g740 (n648, n301, n297, n196, n205);
xor  g741 (n869, n330, n325, n350, n188);
nor  g742 (n398, n283, n298, n145, n184);
nand g743 (n566, n318, n325, n202, n290);
and  g744 (n759, n152, n135, n134, n212);
or   g745 (n867, n239, n250, n148, n340);
or   g746 (n479, n232, n178, n224, n342);
nor  g747 (n778, n227, n129, n315, n93);
and  g748 (n372, n143, n217, n243, n322);
xnor g749 (n378, n337, n352, n143, n110);
xor  g750 (n531, n340, n168, n170, n243);
or   g751 (n442, n255, n127, n157, n138);
nor  g752 (n690, n150, n230, n219, n273);
or   g753 (n435, n279, n245, n313, n288);
xor  g754 (n423, n254, n291, n214, n144);
or   g755 (n540, n306, n255, n185, n117);
or   g756 (n767, n256, n267, n232, n263);
nor  g757 (n453, n193, n242, n332, n88);
nor  g758 (n676, n238, n206, n195, n315);
nand g759 (n852, n163, n180, n343, n90);
nand g760 (n728, n208, n89, n240, n233);
nor  g761 (n491, n187, n240, n305, n325);
nor  g762 (n656, n332, n190, n327, n340);
nor  g763 (n469, n157, n300, n255, n164);
and  g764 (n752, n316, n196, n289, n294);
nor  g765 (n465, n217, n322, n351, n301);
nor  g766 (n756, n261, n165, n301, n268);
xor  g767 (n874, n199, n283, n128, n145);
and  g768 (n630, n188, n141, n306, n261);
and  g769 (n713, n154, n146, n336, n294);
xnor g770 (n851, n105, n122, n222, n228);
nor  g771 (n618, n344, n239, n292, n229);
or   g772 (n533, n197, n309, n355, n287);
xor  g773 (n572, n186, n190, n193, n336);
xnor g774 (n585, n177, n283, n196, n349);
nor  g775 (n692, n322, n167, n224, n298);
xor  g776 (n704, n146, n329, n257, n212);
nand g777 (n440, n223, n354, n220, n251);
and  g778 (n549, n245, n152, n308);
nand g779 (n522, n151, n286, n282, n154);
or   g780 (n757, n315, n247, n269, n226);
xor  g781 (n859, n195, n248, n214);
and  g782 (n737, n294, n265, n287, n147);
or   g783 (n601, n341, n147, n312, n90);
or   g784 (n760, n150, n334, n181, n249);
and  g785 (n739, n96, n145, n188, n241);
nor  g786 (n726, n289, n284, n303, n157);
xnor g787 (n497, n164, n339, n347, n206);
xnor g788 (n765, n97, n306, n191, n221);
nand g789 (n519, n157, n179, n229, n353);
xnor g790 (n703, n133, n337, n87, n334);
and  g791 (n769, n179, n142, n182, n271);
xnor g792 (n856, n262, n210, n187, n200);
nand g793 (n384, n328, n356, n138, n305);
or   g794 (n481, n199, n292, n129, n352);
nand g795 (n754, n348, n336, n197, n195);
xnor g796 (n586, n188, n223, n326, n169);
and  g797 (n695, n136, n282, n343, n194);
xnor g798 (n731, n311, n313, n339, n268);
or   g799 (n791, n99, n276, n260, n278);
or   g800 (n806, n277, n320, n337, n272);
xnor g801 (n848, n253, n183, n169, n163);
and  g802 (n388, n273, n136, n297, n174);
xor  g803 (n680, n156, n265, n231, n271);
or   g804 (n400, n258, n210, n316, n347);
xnor g805 (n788, n260, n174, n148, n122);
nand g806 (n574, n263, n180, n348, n185);
and  g807 (n821, n115, n177, n233, n95);
xnor g808 (n568, n121, n162, n260, n151);
or   g809 (n433, n152, n317, n305, n123);
and  g810 (n809, n259, n356, n258, n236);
or   g811 (n492, n191, n317, n290, n158);
xnor g812 (n763, n329, n141, n294);
or   g813 (n650, n312, n269, n263, n350);
nor  g814 (n573, n227, n285, n184, n115);
and  g815 (n790, n190, n319, n259, n202);
or   g816 (n814, n223, n307, n351, n150);
xnor g817 (n518, n186, n245, n298, n225);
or   g818 (n777, n341, n289, n253, n326);
nand g819 (n523, n235, n131, n314, n205);
and  g820 (n557, n313, n180, n197, n333);
and  g821 (n883, n335, n344, n316, n155);
and  g822 (n576, n193, n318, n331, n253);
nor  g823 (n604, n307, n216, n192, n179);
or   g824 (n602, n218, n86, n310, n112);
nand g825 (n701, n194, n250, n175, n323);
or   g826 (n507, n257, n241, n211, n183);
xor  g827 (n860, n166, n176, n302, n134);
or   g828 (n687, n160, n209, n285, n159);
nand g829 (n855, n205, n218, n116, n269);
nand g830 (n428, n132, n111, n184, n311);
xor  g831 (n866, n293, n134, n142, n334);
nand g832 (n381, n139, n162, n338, n341);
and  g833 (n443, n196, n319, n106, n306);
nor  g834 (n564, n324, n354, n250, n175);
xnor g835 (n361, n181, n321, n324, n241);
or   g836 (n738, n130, n155, n189, n198);
xnor g837 (n386, n159, n207, n229, n348);
xnor g838 (n532, n320, n243, n249, n296);
and  g839 (n367, n233, n270, n208, n197);
xnor g840 (n590, n333, n184, n278, n355);
and  g841 (n596, n222, n149, n303, n173);
and  g842 (n459, n185, n187, n153);
and  g843 (n607, n222, n175, n344, n124);
xor  g844 (n417, n212, n159, n281, n132);
nand g845 (n877, n267, n336, n232, n183);
xor  g846 (n482, n285, n145, n144, n321);
nand g847 (n612, n265, n277, n220, n245);
or   g848 (n516, n202, n277, n156, n216);
or   g849 (n682, n289, n219, n330, n331);
nand g850 (n376, n237, n321, n209, n344);
xor  g851 (n857, n198, n291, n286, n244);
and  g852 (n787, n116, n103, n156, n118);
xnor g853 (n405, n278, n287, n252, n219);
nor  g854 (n525, n280, n351, n223, n291);
xor  g855 (n490, n240, n149, n108, n206);
and  g856 (n646, n153, n284, n239, n215);
and  g857 (n558, n100, n165, n107, n309);
or   g858 (n412, n317, n268, n333, n147);
nor  g859 (n879, n295, n126, n158, n167);
and  g860 (n553, n254, n221, n176, n95);
nor  g861 (n606, n168, n312, n207, n302);
xnor g862 (n499, n239, n326, n328, n281);
xor  g863 (n878, n135, n171, n183, n192);
xor  g864 (n892, n149, n98, n216, n210);
nor  g865 (n717, n327, n214, n267, n162);
and  g866 (n678, n171, n284, n161, n204);
xnor g867 (n804, n304, n140, n220, n219);
xor  g868 (n649, n109, n101, n297, n266);
nor  g869 (n365, n293, n105, n110, n283);
or   g870 (n369, n213, n329, n140, n322);
nand g871 (n732, n310, n304, n208, n270);
nand g872 (n816, n288, n319, n135, n213);
xor  g873 (n475, n242, n355, n168, n87);
and  g874 (n521, n236, n99, n126, n249);
xnor g875 (n426, n163, n328, n235, n290);
xnor g876 (n560, n276, n165, n251, n275);
and  g877 (n718, n198, n100, n234, n342);
xnor g878 (n802, n329, n285, n172, n154);
and  g879 (n904, n441, n369, n407, n412);
nor  g880 (n910, n394, n465, n457, n512);
and  g881 (n933, n497, n380, n452, n505);
xnor g882 (n920, n444, n496, n360, n447);
and  g883 (n916, n498, n459, n473, n420);
nor  g884 (n932, n479, n373, n397, n379);
xnor g885 (n897, n414, n361, n416, n430);
or   g886 (n917, n437, n364, n391, n466);
or   g887 (n907, n408, n393, n453, n508);
and  g888 (n913, n388, n456, n382, n385);
xor  g889 (n924, n377, n383, n448, n418);
nor  g890 (n906, n427, n492, n455, n477);
nor  g891 (n899, n451, n432, n413, n384);
nand g892 (n909, n474, n446, n398, n366);
nor  g893 (n912, n480, n402, n359, n502);
and  g894 (n900, n499, n485, n370, n365);
xor  g895 (n905, n481, n450, n490, n494);
or   g896 (n931, n468, n460, n511, n392);
xor  g897 (n903, n510, n426, n443, n399);
or   g898 (n922, n417, n440, n475, n396);
and  g899 (n919, n431, n495, n469, n454);
nand g900 (n935, n406, n462, n400, n442);
nand g901 (n898, n429, n363, n439, n395);
nand g902 (n921, n509, n483, n371, n405);
nand g903 (n914, n367, n428, n381, n467);
xnor g904 (n929, n449, n491, n438, n484);
xnor g905 (n925, n368, n422, n389, n436);
xor  g906 (n926, n500, n513, n435, n425);
xor  g907 (n934, n507, n470, n434, n488);
nor  g908 (n928, n504, n372, n410, n501);
xor  g909 (n918, n463, n411, n374, n387);
nand g910 (n927, n482, n489, n424, n423);
xor  g911 (n908, n375, n478, n461, n362);
or   g912 (n930, n419, n390, n472, n404);
xnor g913 (n901, n409, n464, n471, n403);
or   g914 (n915, n503, n415, n506, n378);
and  g915 (n902, n476, n376, n487, n458);
xor  g916 (n923, n493, n401, n486, n386);
xor  g917 (n911, n358, n421, n433, n445);
not  g918 (n943, n521);
buf  g919 (n938, n514);
not  g920 (n944, n905);
buf  g921 (n941, n523);
buf  g922 (n940, n520);
nor  g923 (n945, n904, n902, n519);
nand g924 (n936, n898, n516, n900);
or   g925 (n942, n903, n901, n897);
xnor g926 (n937, n906, n522, n517);
nand g927 (n939, n515, n899, n518);
buf  g928 (n979, n912);
not  g929 (n973, n936);
not  g930 (n977, n940);
not  g931 (n966, n914);
not  g932 (n953, n938);
not  g933 (n983, n943);
buf  g934 (n956, n939);
buf  g935 (n962, n563);
not  g936 (n957, n559);
buf  g937 (n951, n928);
not  g938 (n972, n937);
buf  g939 (n980, n945);
not  g940 (n981, n560);
buf  g941 (n970, n556);
not  g942 (n969, n547);
not  g943 (n963, n943);
buf  g944 (n950, n921);
buf  g945 (n961, n936);
or   g946 (n960, n543, n939, n937);
and  g947 (n982, n927, n357, n941, n919);
xnor g948 (n984, n944, n915, n940);
xnor g949 (n974, n937, n911, n530, n943);
or   g950 (n948, n940, n937, n941, n909);
xnor g951 (n959, n943, n918, n544, n923);
nor  g952 (n955, n910, n944, n532);
and  g953 (n978, n553, n527, n533, n526);
or   g954 (n976, n938, n555, n924, n541);
xnor g955 (n975, n538, n551, n550, n536);
or   g956 (n958, n534, n920, n942, n554);
nor  g957 (n946, n561, n944, n936, n945);
nor  g958 (n971, n942, n925, n548, n941);
and  g959 (n954, n528, n916, n917, n524);
xor  g960 (n965, n537, n558, n939, n545);
nor  g961 (n968, n529, n913, n535, n938);
nand g962 (n952, n557, n941, n540, n542);
xor  g963 (n967, n549, n908, n531, n907);
or   g964 (n964, n552, n562, n922, n539);
and  g965 (n947, n942, n945, n525, n938);
nand g966 (n949, n936, n942, n546, n926);
not  g967 (n1001, n950);
not  g968 (n995, n953);
not  g969 (n985, n952);
buf  g970 (n997, n953);
not  g971 (n991, n952);
not  g972 (n990, n947);
buf  g973 (n988, n949);
not  g974 (n1000, n951);
not  g975 (n987, n950);
not  g976 (n999, n947);
buf  g977 (n1002, n951);
buf  g978 (n986, n949);
not  g979 (n998, n948);
not  g980 (n992, n951);
not  g981 (n989, n952);
not  g982 (n993, n952);
not  g983 (n1004, n946);
buf  g984 (n996, n946);
buf  g985 (n1003, n948);
not  g986 (n994, n951);
not  g987 (n1063, n973);
not  g988 (n1038, n1001);
buf  g989 (n1007, n977);
buf  g990 (n1058, n971);
not  g991 (n1056, n1000);
buf  g992 (n1019, n979);
buf  g993 (n1061, n954);
buf  g994 (n1009, n1003);
buf  g995 (n1067, n967);
buf  g996 (n1062, n1000);
not  g997 (n1042, n995);
buf  g998 (n1026, n985);
not  g999 (n1021, n579);
not  g1000 (n1068, n573);
buf  g1001 (n1064, n961);
buf  g1002 (n1057, n991);
not  g1003 (n1011, n961);
buf  g1004 (n1072, n983);
not  g1005 (n1050, n983);
buf  g1006 (n1051, n970);
not  g1007 (n1082, n1002);
buf  g1008 (n1054, n980);
not  g1009 (n1078, n995);
not  g1010 (n1076, n994);
not  g1011 (n1037, n993);
buf  g1012 (n1028, n989);
not  g1013 (n1074, n1004);
buf  g1014 (n1020, n957);
buf  g1015 (n1006, n958);
not  g1016 (n1073, n992);
not  g1017 (n1043, n973);
buf  g1018 (n1033, n570);
xor  g1019 (n1036, n1004, n980);
or   g1020 (n1047, n970, n959, n984, n978);
nand g1021 (n1005, n955, n977, n962, n989);
and  g1022 (n1066, n978, n969, n956, n955);
nand g1023 (n1027, n964, n960, n976, n963);
nand g1024 (n1035, n976, n960, n970, n985);
nor  g1025 (n1031, n988, n999, n972, n978);
xor  g1026 (n1081, n993, n1002, n954, n982);
nor  g1027 (n1017, n958, n984, n1001, n974);
and  g1028 (n1013, n973, n992, n979, n986);
xnor g1029 (n1034, n958, n1003, n1002, n961);
xor  g1030 (n1080, n974, n956, n987, n991);
nor  g1031 (n1055, n975, n953, n988, n972);
and  g1032 (n1010, n995, n997, n955, n978);
xnor g1033 (n1065, n966, n965, n569, n972);
xor  g1034 (n1029, n977, n960, n971, n966);
xnor g1035 (n1022, n998, n996, n981, n963);
or   g1036 (n1049, n971, n997, n975, n979);
nand g1037 (n1084, n576, n1003, n976, n998);
nor  g1038 (n1083, n1000, n967, n963);
nand g1039 (n1015, n957, n980, n566, n985);
and  g1040 (n1024, n959, n966, n985, n968);
xnor g1041 (n1023, n962, n968, n999, n989);
xor  g1042 (n1039, n567, n1004, n991, n970);
xor  g1043 (n1018, n994, n572, n990, n968);
xnor g1044 (n1044, n969, n962, n957, n577);
nor  g1045 (n1052, n991, n977, n565, n966);
nand g1046 (n1075, n956, n564, n968, n996);
nand g1047 (n1012, n962, n969, n986, n983);
and  g1048 (n1014, n982, n993, n574, n992);
nor  g1049 (n1059, n955, n964, n983, n969);
nor  g1050 (n1048, n971, n1001, n999, n578);
xnor g1051 (n1030, n992, n980, n960, n967);
nand g1052 (n1032, n957, n997, n981, n953);
xor  g1053 (n1060, n956, n571, n988, n965);
nand g1054 (n1008, n987, n1001, n982, n975);
xnor g1055 (n1046, n1003, n987, n975, n984);
xnor g1056 (n1071, n995, n998, n575, n959);
nand g1057 (n1040, n993, n996, n963, n961);
xor  g1058 (n1053, n999, n994, n984, n981);
nor  g1059 (n1016, n990, n987, n994, n964);
and  g1060 (n1025, n979, n974, n976, n988);
nand g1061 (n1045, n981, n954, n982, n958);
or   g1062 (n1077, n990, n973, n954, n974);
nor  g1063 (n1070, n965, n998, n986);
and  g1064 (n1079, n990, n1002, n568, n1000);
and  g1065 (n1041, n989, n996, n964, n1004);
and  g1066 (n1069, n965, n972, n997, n959);
xor  g1067 (n1093, n357, n1010, n580);
nor  g1068 (n1089, n1020, n1019, n581);
and  g1069 (n1092, n1015, n1018, n1008);
xor  g1070 (n1090, n1016, n1008, n1006);
or   g1071 (n1087, n1016, n1012, n1005, n1011);
or   g1072 (n1095, n582, n1007, n1020);
or   g1073 (n1097, n1019, n1013, n1016, n1005);
nand g1074 (n1086, n1016, n357, n1011, n1013);
xnor g1075 (n1094, n1014, n1017, n1012, n1006);
nor  g1076 (n1099, n585, n1009, n1017, n945);
or   g1077 (n1088, n583, n1017, n1015);
nor  g1078 (n1096, n1009, n1013, n1012, n1018);
nand g1079 (n1091, n1014, n1012, n1019);
xnor g1080 (n1085, n1011, n1014, n1010, n1018);
xor  g1081 (n1100, n1017, n1013, n1014, n584);
nand g1082 (n1098, n1018, n357, n1011, n1015);
not  g1083 (n1103, n587);
buf  g1084 (n1107, n1094);
buf  g1085 (n1104, n1097);
buf  g1086 (n1111, n586);
buf  g1087 (n1110, n1088);
buf  g1088 (n1112, n592);
not  g1089 (n1106, n1092);
not  g1090 (n1101, n588);
buf  g1091 (n1105, n600);
buf  g1092 (n1109, n597);
and  g1093 (n1113, n1093, n1098, n593, n1096);
and  g1094 (n1114, n1091, n1090, n1087, n598);
nor  g1095 (n1108, n590, n591, n1095, n1086);
and  g1096 (n1115, n1089, n594, n1099, n599);
nand g1097 (n1102, n1085, n596, n595, n589);
not  g1098 (n1121, n1109);
not  g1099 (n1118, n1101);
not  g1100 (n1137, n1105);
not  g1101 (n1126, n1108);
not  g1102 (n1119, n1110);
not  g1103 (n1124, n1102);
not  g1104 (n1117, n1111);
buf  g1105 (n1129, n1111);
not  g1106 (n1128, n1108);
not  g1107 (n1127, n1104);
not  g1108 (n1134, n1103);
not  g1109 (n1130, n1102);
buf  g1110 (n1133, n1106);
buf  g1111 (n1136, n1112);
buf  g1112 (n1131, n1112);
not  g1113 (n1138, n1103);
buf  g1114 (n1139, n1104);
buf  g1115 (n1135, n1107);
not  g1116 (n1123, n1110);
not  g1117 (n1132, n1101);
buf  g1118 (n1116, n1105);
buf  g1119 (n1122, n1109);
not  g1120 (n1125, n1106);
not  g1121 (n1120, n1107);
and  g1122 (n1168, n1073, n1032, n1077, n1042);
nand g1123 (n1183, n1122, n1071, n1031, n1084);
nor  g1124 (n1193, n1049, n1119, n1138, n1054);
xor  g1125 (n1176, n1058, n1127, n1047, n1125);
nand g1126 (n1219, n1061, n1137, n1130, n1136);
nor  g1127 (n1206, n1078, n1135, n1070, n1137);
xnor g1128 (n1144, n1126, n1078, n1042, n1116);
nand g1129 (n1162, n1119, n1045, n1139, n1083);
or   g1130 (n1150, n1027, n1061, n1038, n1134);
nor  g1131 (n1169, n1044, n1059, n1036, n1131);
xnor g1132 (n1231, n1116, n1075, n1123, n1073);
nor  g1133 (n1222, n1135, n1137, n933, n1047);
nand g1134 (n1181, n605, n1023, n1029, n1021);
and  g1135 (n1189, n1127, n1046, n1059, n1044);
xnor g1136 (n1156, n1117, n1127, n1060, n1069);
xnor g1137 (n1212, n1033, n1139, n1120, n1056);
xor  g1138 (n1175, n1068, n1070, n1117, n1028);
xnor g1139 (n1196, n932, n1082, n1072, n1079);
and  g1140 (n1164, n1121, n1080, n1037, n1050);
nor  g1141 (n1228, n1058, n1022, n1082, n1076);
xnor g1142 (n1204, n1138, n1123, n1050, n1034);
or   g1143 (n1201, n1040, n1124, n1051, n1055);
and  g1144 (n1140, n1045, n1119, n1034, n1026);
xnor g1145 (n1226, n934, n1026, n1077, n1124);
nor  g1146 (n1191, n1035, n1135, n1074, n1123);
or   g1147 (n1172, n1118, n1137, n1076, n931);
or   g1148 (n1227, n1030, n929, n1130, n1079);
nor  g1149 (n1163, n1020, n1048, n1079, n1139);
nor  g1150 (n1192, n1065, n1121, n1035, n1072);
xor  g1151 (n1171, n1035, n1113, n1134, n1028);
xnor g1152 (n1151, n1036, n1064, n1025, n1138);
xnor g1153 (n1207, n1069, n1075, n1021, n604);
and  g1154 (n1147, n1057, n1132, n1041, n1029);
or   g1155 (n1154, n1027, n1130, n1084, n1122);
xor  g1156 (n1232, n1057, n1052, n1036);
xnor g1157 (n1186, n1037, n1027, n1118, n1080);
nand g1158 (n1180, n1044, n1068, n1031, n1072);
xor  g1159 (n1173, n1074, n1119, n1082, n1062);
nor  g1160 (n1190, n1061, n1025, n1122, n1128);
or   g1161 (n1194, n1067, n1062, n1068, n1028);
xnor g1162 (n1233, n1029, n1049, n1046, n1120);
xor  g1163 (n1203, n601, n1053, n1042, n1041);
xnor g1164 (n1197, n1069, n1052, n1067, n1058);
or   g1165 (n1215, n1066, n1032, n1056, n1038);
or   g1166 (n1220, n1045, n1131, n1121, n1054);
xnor g1167 (n1187, n1078, n1048, n1026, n1021);
xnor g1168 (n1148, n1123, n1113, n1057, n1083);
nand g1169 (n1221, n1125, n1034, n1032, n1068);
and  g1170 (n1166, n1038, n1053, n1075, n1071);
and  g1171 (n1142, n1033, n606, n1039, n1125);
nand g1172 (n1185, n1070, n1082, n1056, n1115);
nand g1173 (n1141, n1083, n1062, n1065, n1028);
xnor g1174 (n1208, n1037, n1041, n1023, n1133);
and  g1175 (n1165, n1054, n1132, n1115, n1065);
and  g1176 (n1225, n1039, n1124, n1041, n1024);
xor  g1177 (n1178, n1077, n607, n1080, n1050);
or   g1178 (n1214, n1081, n1040, n1044, n1021);
xnor g1179 (n1213, n1043, n1071, n1059);
and  g1180 (n1146, n1053, n930, n1076, n1070);
nor  g1181 (n1143, n1040, n1057, n1129, n1055);
nor  g1182 (n1179, n1053, n1022, n1061, n1081);
and  g1183 (n1229, n1115, n1046, n1051, n1081);
xnor g1184 (n1218, n1025, n1074, n1023, n1126);
and  g1185 (n1155, n1139, n1129, n1022, n1073);
or   g1186 (n1158, n1129, n1128, n608, n1100);
nor  g1187 (n1216, n1032, n1114, n1079, n1128);
xor  g1188 (n1209, n1067, n1027, n1066, n1074);
xnor g1189 (n1182, n1133, n1029, n1066, n1040);
xnor g1190 (n1149, n1076, n1080, n1063, n1064);
and  g1191 (n1210, n1048, n1034, n1133, n1120);
nand g1192 (n1167, n1064, n1039, n1117, n1047);
xor  g1193 (n1157, n1035, n1045, n1135, n1129);
nand g1194 (n1177, n1055, n1033, n1066, n1063);
or   g1195 (n1195, n1136, n1024, n1031, n1131);
and  g1196 (n1217, n1132, n603, n1054, n1078);
nand g1197 (n1198, n1043, n1063, n1024, n1049);
or   g1198 (n1145, n1067, n1042, n1126, n1048);
or   g1199 (n1161, n1136, n1024, n1134, n1050);
or   g1200 (n1174, n1071, n1052, n602, n1072);
xnor g1201 (n1200, n1052, n1030, n1026, n1077);
nor  g1202 (n1230, n1022, n1030, n1037, n1118);
xor  g1203 (n1224, n1046, n1063, n1131, n1065);
xor  g1204 (n1153, n1043, n1047, n1130, n1083);
xor  g1205 (n1223, n1023, n1039, n1081, n1127);
xor  g1206 (n1202, n1120, n1134, n1058, n1064);
nand g1207 (n1188, n1084, n1075, n1038, n1138);
and  g1208 (n1199, n1030, n1060, n1115);
and  g1209 (n1205, n1049, n1051, n935, n1025);
or   g1210 (n1160, n1069, n1051, n1132, n1033);
xnor g1211 (n1211, n1126, n1124, n1055, n1060);
nor  g1212 (n1152, n1133, n1136, n1020, n1084);
and  g1213 (n1159, n1122, n1056, n1121, n1118);
xnor g1214 (n1170, n1125, n1073, n1062, n1128);
nand g1215 (n1184, n1043, n1031, n1117, n1114);
nor  g1216 (n1290, n712, n753, n749, n726);
nor  g1217 (n1288, n617, n781, n783, n629);
nor  g1218 (n1322, n627, n785, n896, n872);
nand g1219 (n1260, n729, n757, n648, n624);
nor  g1220 (n1300, n1188, n774, n855, n1155);
and  g1221 (n1301, n642, n730, n782, n640);
nand g1222 (n1264, n867, n646, n739, n1173);
xnor g1223 (n1279, n1229, n1159, n701, n611);
nor  g1224 (n1303, n615, n862, n639, n771);
and  g1225 (n1271, n653, n799, n690, n1181);
xor  g1226 (n1255, n1197, n664, n843, n873);
nand g1227 (n1311, n770, n836, n800, n860);
nor  g1228 (n1263, n673, n831, n850, n669);
xor  g1229 (n1316, n1195, n676, n792, n813);
nand g1230 (n1310, n722, n609, n789, n895);
nand g1231 (n1305, n1147, n1166, n735, n1171);
nor  g1232 (n1258, n635, n623, n1158, n696);
and  g1233 (n1320, n746, n821, n824, n732);
xor  g1234 (n1307, n1194, n681, n1168, n661);
or   g1235 (n1250, n744, n830, n765, n761);
and  g1236 (n1324, n864, n882, n691, n734);
or   g1237 (n1273, n1223, n755, n892, n779);
nor  g1238 (n1249, n694, n894, n875, n1164);
and  g1239 (n1253, n1172, n1193, n1143, n689);
nand g1240 (n1268, n1161, n854, n798, n1210);
xnor g1241 (n1325, n794, n876, n657, n1214);
nor  g1242 (n1244, n1221, n743, n1233, n742);
nand g1243 (n1329, n758, n803, n636, n637);
xor  g1244 (n1297, n849, n846, n674, n820);
or   g1245 (n1315, n647, n1231, n886, n769);
or   g1246 (n1319, n877, n1205, n1191, n801);
xnor g1247 (n1321, n662, n812, n773, n638);
nand g1248 (n1272, n1227, n890, n1233, n767);
nor  g1249 (n1302, n1232, n861, n740, n764);
nand g1250 (n1293, n1209, n718, n1180, n818);
nand g1251 (n1287, n795, n802, n645, n724);
nor  g1252 (n1306, n612, n698, n871, n808);
xor  g1253 (n1242, n679, n660, n870, n677);
nor  g1254 (n1327, n869, n707, n832, n1212);
nand g1255 (n1257, n1176, n695, n848, n1175);
or   g1256 (n1270, n1167, n706, n614, n1226);
nor  g1257 (n1323, n641, n1179, n804, n716);
nor  g1258 (n1266, n790, n1224, n1202, n1145);
and  g1259 (n1294, n827, n834, n1151, n685);
xor  g1260 (n1240, n833, n858, n786, n1183);
xnor g1261 (n1298, n1141, n1160, n737, n634);
xor  g1262 (n1304, n720, n885, n811, n823);
xnor g1263 (n1277, n619, n1169, n654, n888);
xor  g1264 (n1235, n1186, n667, n709, n704);
and  g1265 (n1247, n1200, n1217, n793, n699);
xnor g1266 (n1241, n845, n878, n1178, n747);
nand g1267 (n1291, n1228, n745, n1196, n625);
or   g1268 (n1285, n656, n879, n814, n784);
or   g1269 (n1256, n766, n859, n693, n1177);
nand g1270 (n1262, n631, n678, n675, n828);
and  g1271 (n1234, n633, n655, n768, n1156);
nand g1272 (n1278, n1152, n668, n751, n1140);
nand g1273 (n1246, n1182, n711, n838, n719);
or   g1274 (n1274, n644, n1207, n759, n727);
xor  g1275 (n1317, n687, n630, n1192, n760);
nand g1276 (n1282, n1190, n1211, n725, n1220);
or   g1277 (n1283, n756, n1199, n650, n702);
nor  g1278 (n1251, n738, n874, n622, n1232);
xnor g1279 (n1265, n1157, n663, n868, n825);
nand g1280 (n1254, n1170, n723, n1198, n717);
nand g1281 (n1289, n822, n620, n710, n893);
xnor g1282 (n1243, n844, n810, n780, n672);
xor  g1283 (n1259, n778, n682, n817, n649);
xor  g1284 (n1275, n697, n1162, n705, n1174);
and  g1285 (n1292, n852, n1149, n775, n680);
and  g1286 (n1237, n1153, n1165, n715, n816);
nor  g1287 (n1252, n643, n713, n658, n652);
or   g1288 (n1267, n1215, n703, n1154, n621);
xnor g1289 (n1314, n1230, n847, n700, n1208);
or   g1290 (n1236, n807, n1218, n787, n728);
or   g1291 (n1286, n651, n1216, n754, n1203);
or   g1292 (n1299, n610, n826, n819, n671);
nand g1293 (n1261, n1144, n887, n797, n1184);
and  g1294 (n1238, n884, n1206, n670, n626);
or   g1295 (n1280, n1150, n1219, n665, n809);
xnor g1296 (n1312, n851, n1146, n1187, n776);
xor  g1297 (n1245, n883, n632, n1163, n840);
xnor g1298 (n1276, n889, n815, n684, n865);
or   g1299 (n1239, n863, n618, n841, n777);
nor  g1300 (n1269, n829, n866, n748, n881);
or   g1301 (n1328, n688, n805, n857, n791);
nor  g1302 (n1309, n613, n683, n1213, n659);
xor  g1303 (n1326, n1225, n788, n721, n1201);
xnor g1304 (n1296, n741, n835, n880, n842);
xor  g1305 (n1308, n763, n733, n772, n692);
or   g1306 (n1248, n839, n837, n736, n853);
xnor g1307 (n1313, n1222, n1185, n616, n752);
xnor g1308 (n1318, n1189, n1204, n731, n666);
and  g1309 (n1284, n856, n750, n686, n796);
and  g1310 (n1295, n628, n762, n891, n714);
nand g1311 (n1281, n708, n806, n1142, n1148);
or   g1312 (n1342, n1305, n1257, n1315, n1263);
and  g1313 (n1332, n1302, n1280, n1304, n1277);
and  g1314 (n1352, n1313, n1317, n1329, n1252);
xor  g1315 (n1344, n1244, n1235, n1300, n1261);
or   g1316 (n1333, n1286, n1320, n1264, n1316);
nand g1317 (n1346, n1275, n1276, n1326, n1245);
or   g1318 (n1341, n1272, n1236, n1292, n1262);
xor  g1319 (n1339, n1249, n1321, n1295, n1234);
and  g1320 (n1350, n1255, n1296, n1242, n1299);
nand g1321 (n1351, n1291, n1238, n1279, n1324);
and  g1322 (n1337, n1269, n1325, n1237, n1240);
xnor g1323 (n1330, n1294, n1284, n1314, n1270);
nand g1324 (n1343, n1248, n1268, n1323, n1289);
nor  g1325 (n1353, n1293, n1251, n1246, n1274);
and  g1326 (n1348, n1301, n1281, n1266, n1287);
and  g1327 (n1331, n1308, n1241, n1318, n1311);
nand g1328 (n1340, n1247, n1273, n1322, n1319);
xnor g1329 (n1349, n1285, n1260, n1303, n1253);
nand g1330 (n1336, n1307, n1298, n1265, n1306);
xor  g1331 (n1345, n1328, n1256, n1312, n1259);
and  g1332 (n1335, n1288, n1290, n1282, n1267);
nor  g1333 (n1334, n1243, n1278, n1239, n1310);
xor  g1334 (n1347, n1283, n1250, n1297, n1327);
xor  g1335 (n1338, n1271, n1254, n1309, n1258);
endmodule
