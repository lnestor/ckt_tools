

module Stat_3000_306
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n323,
  n356,
  n3020,
  n3022,
  n3032,
  n3005,
  n3011,
  n3017,
  n3003,
  n3008,
  n3031,
  n3021,
  n3009,
  n3026,
  n3004,
  n3023,
  n3010,
  n3014,
  n3016,
  n3025,
  n3024,
  n3013,
  n3027,
  n3019,
  n3029,
  n3007,
  n3028,
  n3030,
  n3015,
  n3018,
  n3012,
  n3006
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n323;output n356;output n3020;output n3022;output n3032;output n3005;output n3011;output n3017;output n3003;output n3008;output n3031;output n3021;output n3009;output n3026;output n3004;output n3023;output n3010;output n3014;output n3016;output n3025;output n3024;output n3013;output n3027;output n3019;output n3029;output n3007;output n3028;output n3030;output n3015;output n3018;output n3012;output n3006;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2795;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2844;wire n2845;wire n2846;wire n2847;wire n2848;wire n2849;wire n2850;wire n2851;wire n2852;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n68,
    n8
  );


  buf
  g1
  (
    n46,
    n8
  );


  buf
  g2
  (
    n86,
    n6
  );


  buf
  g3
  (
    n38,
    n13
  );


  not
  g4
  (
    n77,
    n7
  );


  not
  g5
  (
    n82,
    n11
  );


  buf
  g6
  (
    n75,
    n6
  );


  not
  g7
  (
    n51,
    n10
  );


  buf
  g8
  (
    n87,
    n12
  );


  buf
  g9
  (
    n63,
    n9
  );


  not
  g10
  (
    n45,
    n10
  );


  not
  g11
  (
    n44,
    n9
  );


  buf
  g12
  (
    n55,
    n12
  );


  buf
  g13
  (
    n54,
    n6
  );


  buf
  g14
  (
    n67,
    n12
  );


  not
  g15
  (
    n79,
    n2
  );


  buf
  g16
  (
    n48,
    n5
  );


  buf
  g17
  (
    n50,
    n3
  );


  buf
  g18
  (
    n36,
    n14
  );


  not
  g19
  (
    n49,
    n4
  );


  not
  g20
  (
    n65,
    n7
  );


  buf
  g21
  (
    n81,
    n3
  );


  buf
  g22
  (
    n78,
    n13
  );


  not
  g23
  (
    n76,
    n5
  );


  buf
  g24
  (
    n34,
    n8
  );


  buf
  g25
  (
    n80,
    n7
  );


  not
  g26
  (
    n47,
    n3
  );


  buf
  g27
  (
    n85,
    n13
  );


  buf
  g28
  (
    n83,
    n9
  );


  not
  g29
  (
    n59,
    n2
  );


  buf
  g30
  (
    n61,
    n2
  );


  not
  g31
  (
    n35,
    n2
  );


  buf
  g32
  (
    n74,
    n12
  );


  buf
  g33
  (
    n64,
    n3
  );


  buf
  g34
  (
    n41,
    n8
  );


  buf
  g35
  (
    n84,
    n15
  );


  not
  g36
  (
    n70,
    n1
  );


  buf
  g37
  (
    n53,
    n5
  );


  buf
  g38
  (
    n72,
    n9
  );


  buf
  g39
  (
    n73,
    n14
  );


  buf
  g40
  (
    n66,
    n15
  );


  buf
  g41
  (
    n58,
    n4
  );


  not
  g42
  (
    n69,
    n7
  );


  not
  g43
  (
    n71,
    n14
  );


  buf
  g44
  (
    n88,
    n10
  );


  not
  g45
  (
    n60,
    n13
  );


  not
  g46
  (
    n39,
    n4
  );


  buf
  g47
  (
    n33,
    n10
  );


  buf
  g48
  (
    n52,
    n1
  );


  not
  g49
  (
    n42,
    n5
  );


  not
  g50
  (
    n62,
    n11
  );


  buf
  g51
  (
    n37,
    n11
  );


  buf
  g52
  (
    n57,
    n11
  );


  buf
  g53
  (
    n43,
    n14
  );


  buf
  g54
  (
    n56,
    n4
  );


  buf
  g55
  (
    n40,
    n6
  );


  not
  g56
  (
    n98,
    n54
  );


  not
  g57
  (
    n279,
    n39
  );


  buf
  g58
  (
    n176,
    n48
  );


  not
  g59
  (
    n135,
    n58
  );


  not
  g60
  (
    n198,
    n62
  );


  not
  g61
  (
    n123,
    n34
  );


  buf
  g62
  (
    n154,
    n53
  );


  buf
  g63
  (
    n246,
    n81
  );


  buf
  g64
  (
    n142,
    n59
  );


  buf
  g65
  (
    n97,
    n61
  );


  not
  g66
  (
    n170,
    n69
  );


  not
  g67
  (
    n149,
    n33
  );


  not
  g68
  (
    n116,
    n83
  );


  not
  g69
  (
    n182,
    n53
  );


  buf
  g70
  (
    n157,
    n78
  );


  not
  g71
  (
    n228,
    n59
  );


  buf
  g72
  (
    n188,
    n74
  );


  not
  g73
  (
    n236,
    n79
  );


  not
  g74
  (
    n100,
    n44
  );


  buf
  g75
  (
    n265,
    n36
  );


  buf
  g76
  (
    n112,
    n40
  );


  not
  g77
  (
    n220,
    n64
  );


  buf
  g78
  (
    n167,
    n67
  );


  buf
  g79
  (
    n238,
    n56
  );


  not
  g80
  (
    n259,
    n73
  );


  buf
  g81
  (
    n150,
    n82
  );


  buf
  g82
  (
    n127,
    n79
  );


  not
  g83
  (
    n200,
    n47
  );


  buf
  g84
  (
    n284,
    n75
  );


  not
  g85
  (
    n229,
    n67
  );


  not
  g86
  (
    n204,
    n49
  );


  buf
  g87
  (
    n146,
    n73
  );


  buf
  g88
  (
    n264,
    n42
  );


  buf
  g89
  (
    n222,
    n38
  );


  buf
  g90
  (
    n275,
    n48
  );


  not
  g91
  (
    n129,
    n74
  );


  not
  g92
  (
    n90,
    n45
  );


  buf
  g93
  (
    n174,
    n57
  );


  buf
  g94
  (
    n155,
    n39
  );


  buf
  g95
  (
    n282,
    n72
  );


  not
  g96
  (
    n255,
    n50
  );


  buf
  g97
  (
    n166,
    n62
  );


  not
  g98
  (
    n201,
    n40
  );


  not
  g99
  (
    n253,
    n79
  );


  not
  g100
  (
    n216,
    n55
  );


  not
  g101
  (
    n148,
    n35
  );


  not
  g102
  (
    n191,
    n82
  );


  buf
  g103
  (
    n271,
    n47
  );


  not
  g104
  (
    n226,
    n57
  );


  not
  g105
  (
    n256,
    n41
  );


  buf
  g106
  (
    n141,
    n37
  );


  not
  g107
  (
    n99,
    n34
  );


  not
  g108
  (
    n156,
    n43
  );


  buf
  g109
  (
    n104,
    n60
  );


  buf
  g110
  (
    n108,
    n72
  );


  not
  g111
  (
    n239,
    n59
  );


  not
  g112
  (
    n213,
    n54
  );


  buf
  g113
  (
    n117,
    n43
  );


  not
  g114
  (
    n272,
    n57
  );


  not
  g115
  (
    n210,
    n75
  );


  not
  g116
  (
    n107,
    n83
  );


  buf
  g117
  (
    n126,
    n69
  );


  buf
  g118
  (
    n207,
    n33
  );


  not
  g119
  (
    n241,
    n61
  );


  not
  g120
  (
    n134,
    n35
  );


  buf
  g121
  (
    n163,
    n47
  );


  buf
  g122
  (
    n287,
    n63
  );


  not
  g123
  (
    n267,
    n62
  );


  buf
  g124
  (
    n161,
    n52
  );


  buf
  g125
  (
    n119,
    n75
  );


  buf
  g126
  (
    n189,
    n71
  );


  not
  g127
  (
    n249,
    n37
  );


  buf
  g128
  (
    n292,
    n77
  );


  not
  g129
  (
    n197,
    n55
  );


  not
  g130
  (
    n92,
    n53
  );


  buf
  g131
  (
    n288,
    n56
  );


  not
  g132
  (
    n274,
    n65
  );


  buf
  g133
  (
    n203,
    n64
  );


  not
  g134
  (
    n181,
    n40
  );


  not
  g135
  (
    n247,
    n65
  );


  buf
  g136
  (
    n192,
    n78
  );


  not
  g137
  (
    n175,
    n79
  );


  buf
  g138
  (
    n130,
    n35
  );


  not
  g139
  (
    n223,
    n34
  );


  buf
  g140
  (
    n140,
    n60
  );


  not
  g141
  (
    n250,
    n71
  );


  buf
  g142
  (
    n102,
    n76
  );


  not
  g143
  (
    n180,
    n36
  );


  buf
  g144
  (
    n93,
    n70
  );


  not
  g145
  (
    n251,
    n61
  );


  not
  g146
  (
    n269,
    n52
  );


  not
  g147
  (
    n96,
    n41
  );


  not
  g148
  (
    n277,
    n38
  );


  buf
  g149
  (
    n280,
    n50
  );


  buf
  g150
  (
    n202,
    n67
  );


  not
  g151
  (
    n131,
    n52
  );


  buf
  g152
  (
    n122,
    n46
  );


  not
  g153
  (
    n270,
    n42
  );


  buf
  g154
  (
    n244,
    n58
  );


  buf
  g155
  (
    n206,
    n51
  );


  buf
  g156
  (
    n111,
    n56
  );


  buf
  g157
  (
    n245,
    n77
  );


  buf
  g158
  (
    n194,
    n38
  );


  not
  g159
  (
    n232,
    n81
  );


  buf
  g160
  (
    n138,
    n45
  );


  not
  g161
  (
    n144,
    n65
  );


  not
  g162
  (
    n212,
    n45
  );


  buf
  g163
  (
    n243,
    n62
  );


  not
  g164
  (
    n266,
    n80
  );


  buf
  g165
  (
    n214,
    n67
  );


  buf
  g166
  (
    n235,
    n73
  );


  not
  g167
  (
    n125,
    n34
  );


  not
  g168
  (
    n132,
    n75
  );


  not
  g169
  (
    n151,
    n43
  );


  not
  g170
  (
    n106,
    n63
  );


  not
  g171
  (
    n173,
    n74
  );


  buf
  g172
  (
    n120,
    n76
  );


  buf
  g173
  (
    n291,
    n59
  );


  buf
  g174
  (
    n273,
    n80
  );


  not
  g175
  (
    n128,
    n83
  );


  not
  g176
  (
    n224,
    n58
  );


  not
  g177
  (
    n281,
    n44
  );


  not
  g178
  (
    n168,
    n71
  );


  buf
  g179
  (
    n233,
    n37
  );


  buf
  g180
  (
    n258,
    n66
  );


  not
  g181
  (
    n242,
    n77
  );


  not
  g182
  (
    n113,
    n63
  );


  buf
  g183
  (
    n268,
    n51
  );


  buf
  g184
  (
    n219,
    n76
  );


  buf
  g185
  (
    n195,
    n64
  );


  buf
  g186
  (
    n105,
    n43
  );


  buf
  g187
  (
    n221,
    n49
  );


  not
  g188
  (
    n152,
    n66
  );


  buf
  g189
  (
    n205,
    n61
  );


  buf
  g190
  (
    n95,
    n65
  );


  buf
  g191
  (
    n262,
    n55
  );


  buf
  g192
  (
    n121,
    n76
  );


  not
  g193
  (
    n225,
    n39
  );


  not
  g194
  (
    n136,
    n56
  );


  not
  g195
  (
    n109,
    n80
  );


  not
  g196
  (
    KeyWire_0_14,
    n39
  );


  buf
  g197
  (
    n285,
    n63
  );


  buf
  g198
  (
    n257,
    n82
  );


  not
  g199
  (
    n103,
    n66
  );


  not
  g200
  (
    n162,
    n41
  );


  buf
  g201
  (
    n115,
    n66
  );


  not
  g202
  (
    n183,
    n45
  );


  buf
  g203
  (
    n215,
    n36
  );


  buf
  g204
  (
    n289,
    n46
  );


  not
  g205
  (
    n158,
    n33
  );


  buf
  g206
  (
    n254,
    n81
  );


  not
  g207
  (
    n230,
    n83
  );


  buf
  g208
  (
    n276,
    n69
  );


  buf
  g209
  (
    n91,
    n37
  );


  not
  g210
  (
    n199,
    n60
  );


  not
  g211
  (
    n139,
    n44
  );


  buf
  g212
  (
    n209,
    n70
  );


  buf
  g213
  (
    n186,
    n35
  );


  not
  g214
  (
    n237,
    n36
  );


  not
  g215
  (
    n290,
    n46
  );


  not
  g216
  (
    n240,
    n82
  );


  buf
  g217
  (
    n234,
    n48
  );


  not
  g218
  (
    n177,
    n40
  );


  not
  g219
  (
    n263,
    n53
  );


  not
  g220
  (
    n89,
    n78
  );


  buf
  g221
  (
    n172,
    n68
  );


  not
  g222
  (
    n101,
    n70
  );


  not
  g223
  (
    n164,
    n74
  );


  not
  g224
  (
    n143,
    n78
  );


  buf
  g225
  (
    n178,
    n47
  );


  not
  g226
  (
    n218,
    n50
  );


  not
  g227
  (
    n165,
    n70
  );


  not
  g228
  (
    n278,
    n80
  );


  buf
  g229
  (
    n211,
    n38
  );


  buf
  g230
  (
    n110,
    n68
  );


  not
  g231
  (
    n184,
    n50
  );


  buf
  g232
  (
    n283,
    n51
  );


  buf
  g233
  (
    n124,
    n44
  );


  buf
  g234
  (
    n94,
    n42
  );


  not
  g235
  (
    n231,
    n58
  );


  not
  g236
  (
    n153,
    n49
  );


  buf
  g237
  (
    n193,
    n46
  );


  not
  g238
  (
    n145,
    n69
  );


  buf
  g239
  (
    n114,
    n81
  );


  buf
  g240
  (
    n190,
    n57
  );


  not
  g241
  (
    n171,
    n49
  );


  buf
  g242
  (
    n208,
    n55
  );


  buf
  g243
  (
    n217,
    n60
  );


  buf
  g244
  (
    n252,
    n64
  );


  buf
  g245
  (
    n160,
    n48
  );


  buf
  g246
  (
    n159,
    n72
  );


  not
  g247
  (
    n169,
    n51
  );


  not
  g248
  (
    n133,
    n52
  );


  buf
  g249
  (
    n118,
    n68
  );


  buf
  g250
  (
    n187,
    n68
  );


  not
  g251
  (
    n286,
    n72
  );


  not
  g252
  (
    n179,
    n54
  );


  buf
  g253
  (
    n248,
    n71
  );


  not
  g254
  (
    n196,
    n33
  );


  buf
  g255
  (
    n261,
    n73
  );


  not
  g256
  (
    n227,
    n77
  );


  not
  g257
  (
    n137,
    n54
  );


  not
  g258
  (
    n260,
    n41
  );


  not
  g259
  (
    n147,
    n42
  );


  not
  g260
  (
    n315,
    n90
  );


  not
  g261
  (
    n298,
    n92
  );


  not
  g262
  (
    n294,
    n96
  );


  buf
  g263
  (
    n308,
    n91
  );


  buf
  g264
  (
    n305,
    n94
  );


  not
  g265
  (
    n311,
    n94
  );


  not
  g266
  (
    n301,
    n90
  );


  buf
  g267
  (
    n306,
    n91
  );


  not
  g268
  (
    n300,
    n89
  );


  not
  g269
  (
    n313,
    n94
  );


  not
  g270
  (
    n314,
    n92
  );


  not
  g271
  (
    n321,
    n91
  );


  not
  g272
  (
    n293,
    n89
  );


  not
  g273
  (
    n299,
    n95
  );


  not
  g274
  (
    n309,
    n92
  );


  buf
  g275
  (
    n320,
    n95
  );


  buf
  g276
  (
    n319,
    n91
  );


  buf
  g277
  (
    n297,
    n93
  );


  buf
  g278
  (
    n317,
    n89
  );


  buf
  g279
  (
    n316,
    n90
  );


  not
  g280
  (
    n307,
    n89
  );


  not
  g281
  (
    KeyWire_0_11,
    n96
  );


  not
  g282
  (
    n295,
    n92
  );


  buf
  g283
  (
    n310,
    n93
  );


  buf
  g284
  (
    n304,
    n90
  );


  not
  g285
  (
    n303,
    n95
  );


  buf
  g286
  (
    n302,
    n94
  );


  buf
  g287
  (
    n318,
    n93
  );


  nand
  g288
  (
    n296,
    n95,
    n93
  );


  buf
  g289
  (
    n322,
    n294
  );


  not
  g290
  (
    n323,
    n293
  );


  and
  g291
  (
    n324,
    n323,
    n84
  );


  xor
  g292
  (
    n326,
    n324,
    n96
  );


  nor
  g293
  (
    n327,
    n97,
    n98,
    n324
  );


  or
  g294
  (
    n325,
    n324,
    n97
  );


  nand
  g295
  (
    n329,
    n327,
    n298,
    n316,
    n301
  );


  or
  g296
  (
    n330,
    n304,
    n299,
    n302,
    n319
  );


  nor
  g297
  (
    n335,
    n316,
    n296,
    n315,
    n326
  );


  and
  g298
  (
    n328,
    n312,
    n305,
    n295,
    n326
  );


  nor
  g299
  (
    n334,
    n325,
    n311,
    n318,
    n315
  );


  nor
  g300
  (
    n337,
    n327,
    n325,
    n297,
    n318
  );


  xnor
  g301
  (
    n333,
    n326,
    n327,
    n310
  );


  nand
  g302
  (
    n332,
    n326,
    n300,
    n309,
    n313
  );


  xnor
  g303
  (
    n336,
    n307,
    n319,
    n317,
    n308
  );


  xor
  g304
  (
    n331,
    n314,
    n317,
    n306,
    n303
  );


  buf
  g305
  (
    n341,
    n328
  );


  buf
  g306
  (
    n339,
    n16
  );


  xor
  g307
  (
    n340,
    n15,
    n16,
    n328
  );


  nor
  g308
  (
    n338,
    n16,
    n328,
    n15
  );


  buf
  g309
  (
    n342,
    n338
  );


  and
  g310
  (
    n343,
    n342,
    n98
  );


  xnor
  g311
  (
    n345,
    n330,
    n329,
    n343
  );


  and
  g312
  (
    n344,
    n330,
    n329
  );


  or
  g313
  (
    n349,
    n344,
    n340,
    n345
  );


  or
  g314
  (
    n350,
    n340,
    n341,
    n344
  );


  xor
  g315
  (
    n347,
    n341,
    n344,
    n338
  );


  xor
  g316
  (
    n348,
    n340,
    n339,
    n338,
    n344
  );


  or
  g317
  (
    n346,
    n341,
    n339
  );


  nand
  g318
  (
    n358,
    n84,
    n348
  );


  nand
  g319
  (
    n355,
    n346,
    n350,
    n320,
    n321
  );


  xor
  g320
  (
    n354,
    n99,
    n86,
    n350,
    n347
  );


  and
  g321
  (
    n356,
    n350,
    n85,
    n320,
    n346
  );


  xnor
  g322
  (
    n353,
    n348,
    n342,
    n99,
    n330
  );


  and
  g323
  (
    n357,
    n85,
    n349,
    n320,
    n350
  );


  nor
  g324
  (
    n351,
    n84,
    n86,
    n85
  );


  xnor
  g325
  (
    n359,
    n349,
    n347,
    n84,
    n85
  );


  nor
  g326
  (
    n352,
    n345,
    n345,
    n320,
    n342
  );


  buf
  g327
  (
    n365,
    n17
  );


  buf
  g328
  (
    n363,
    n355
  );


  not
  g329
  (
    n361,
    n17
  );


  buf
  g330
  (
    n364,
    n356
  );


  buf
  g331
  (
    n362,
    n353
  );


  nor
  g332
  (
    n360,
    n357,
    n354,
    n352
  );


  not
  g333
  (
    n369,
    n87
  );


  buf
  g334
  (
    n370,
    n362
  );


  xnor
  g335
  (
    n367,
    n360,
    n361
  );


  xnor
  g336
  (
    n366,
    n17,
    n364
  );


  xor
  g337
  (
    n368,
    n86,
    n363
  );


  not
  g338
  (
    n376,
    n366
  );


  not
  g339
  (
    n373,
    n367
  );


  buf
  g340
  (
    n375,
    n367
  );


  buf
  g341
  (
    n371,
    n367
  );


  not
  g342
  (
    n374,
    n366
  );


  not
  g343
  (
    n377,
    n366
  );


  xor
  g344
  (
    n372,
    n99,
    n366
  );


  buf
  g345
  (
    n401,
    n101
  );


  buf
  g346
  (
    n400,
    n374
  );


  buf
  g347
  (
    n396,
    n99
  );


  not
  g348
  (
    n382,
    n375
  );


  buf
  g349
  (
    n385,
    n377
  );


  buf
  g350
  (
    n402,
    n376
  );


  buf
  g351
  (
    n397,
    n371
  );


  buf
  g352
  (
    n405,
    n375
  );


  not
  g353
  (
    n383,
    n377
  );


  not
  g354
  (
    n389,
    n100
  );


  buf
  g355
  (
    n404,
    n359
  );


  not
  g356
  (
    n381,
    n100
  );


  buf
  g357
  (
    n379,
    n376
  );


  not
  g358
  (
    n388,
    n374
  );


  buf
  g359
  (
    n392,
    n373
  );


  buf
  g360
  (
    n394,
    n373
  );


  buf
  g361
  (
    n390,
    n375
  );


  not
  g362
  (
    n391,
    n101
  );


  buf
  g363
  (
    n398,
    n373
  );


  buf
  g364
  (
    n387,
    n372
  );


  not
  g365
  (
    n378,
    n374
  );


  buf
  g366
  (
    n399,
    n375
  );


  not
  g367
  (
    n384,
    n371
  );


  not
  g368
  (
    n403,
    n358
  );


  not
  g369
  (
    n386,
    n376
  );


  nor
  g370
  (
    n395,
    n377,
    n100,
    n372,
    n376
  );


  xor
  g371
  (
    n380,
    n373,
    n372,
    n371
  );


  xor
  g372
  (
    n393,
    n374,
    n377,
    n100,
    n371
  );


  or
  g373
  (
    n406,
    n378,
    n365
  );


  not
  g374
  (
    n407,
    n406
  );


  not
  g375
  (
    n408,
    n406
  );


  not
  g376
  (
    n409,
    n408
  );


  buf
  g377
  (
    n412,
    n408
  );


  buf
  g378
  (
    n411,
    n408
  );


  buf
  g379
  (
    n415,
    n407
  );


  not
  g380
  (
    n410,
    n408
  );


  not
  g381
  (
    n413,
    n407
  );


  buf
  g382
  (
    n414,
    n407
  );


  not
  g383
  (
    n416,
    n407
  );


  or
  g384
  (
    n434,
    n389,
    n382,
    n410,
    n380
  );


  nand
  g385
  (
    KeyWire_0_12,
    n382,
    n385,
    n386,
    n412
  );


  nand
  g386
  (
    n420,
    n379,
    n411,
    n381,
    n385
  );


  xnor
  g387
  (
    n430,
    n385,
    n380,
    n378,
    n390
  );


  xor
  g388
  (
    n423,
    n387,
    n391,
    n388,
    n384
  );


  nor
  g389
  (
    n421,
    n409,
    n383,
    n390
  );


  nand
  g390
  (
    n427,
    n383,
    n412,
    n381
  );


  xor
  g391
  (
    n428,
    n389,
    n381,
    n379,
    n384
  );


  xnor
  g392
  (
    n422,
    n391,
    n386,
    n410
  );


  xnor
  g393
  (
    n429,
    n379,
    n378,
    n380,
    n391
  );


  nand
  g394
  (
    n419,
    n409,
    n382,
    n390,
    n411
  );


  xor
  g395
  (
    n418,
    n385,
    n382,
    n411,
    n390
  );


  or
  g396
  (
    n424,
    n379,
    n388,
    n380,
    n412
  );


  xor
  g397
  (
    n417,
    n409,
    n413,
    n384,
    n387
  );


  nand
  g398
  (
    n425,
    n409,
    n386,
    n411,
    n383
  );


  nand
  g399
  (
    n426,
    n381,
    n378,
    n387,
    n410
  );


  xnor
  g400
  (
    n432,
    n387,
    n389,
    n388,
    n413
  );


  nand
  g401
  (
    n431,
    n389,
    n388,
    n410,
    n384
  );


  buf
  g402
  (
    n435,
    n87
  );


  not
  g403
  (
    n443,
    n419
  );


  buf
  g404
  (
    n436,
    n368
  );


  xnor
  g405
  (
    n439,
    n422,
    n321,
    n88,
    n369
  );


  nand
  g406
  (
    n438,
    n423,
    n369,
    n392,
    n87
  );


  xnor
  g407
  (
    n440,
    n88,
    n369,
    n420,
    n406
  );


  xor
  g408
  (
    n441,
    n426,
    n427,
    n392,
    n391
  );


  xnor
  g409
  (
    n444,
    n417,
    n406,
    n321,
    n368
  );


  and
  g410
  (
    n445,
    n369,
    n424,
    n87,
    n425
  );


  xor
  g411
  (
    n442,
    n421,
    n321,
    n418,
    n88
  );


  nor
  g412
  (
    n437,
    n368,
    n368,
    n367,
    n88
  );


  not
  g413
  (
    n448,
    n438
  );


  buf
  g414
  (
    n450,
    n439
  );


  buf
  g415
  (
    n467,
    n439
  );


  not
  g416
  (
    n464,
    n436
  );


  buf
  g417
  (
    n469,
    n435
  );


  not
  g418
  (
    n466,
    n440
  );


  buf
  g419
  (
    n447,
    n440
  );


  buf
  g420
  (
    n454,
    n438
  );


  not
  g421
  (
    n468,
    n440
  );


  buf
  g422
  (
    n462,
    n437
  );


  not
  g423
  (
    n460,
    n437
  );


  buf
  g424
  (
    n456,
    n439
  );


  not
  g425
  (
    n457,
    n437
  );


  not
  g426
  (
    n452,
    n436
  );


  not
  g427
  (
    n453,
    n437
  );


  buf
  g428
  (
    n458,
    n435
  );


  not
  g429
  (
    n446,
    n440
  );


  buf
  g430
  (
    n465,
    n438
  );


  buf
  g431
  (
    n459,
    n436
  );


  buf
  g432
  (
    n455,
    n438
  );


  buf
  g433
  (
    n461,
    n435
  );


  buf
  g434
  (
    n451,
    n435
  );


  buf
  g435
  (
    n449,
    n439
  );


  buf
  g436
  (
    n463,
    n436
  );


  buf
  g437
  (
    n531,
    n393
  );


  not
  g438
  (
    n481,
    n102
  );


  buf
  g439
  (
    n532,
    n451
  );


  buf
  g440
  (
    n533,
    n448
  );


  not
  g441
  (
    n487,
    n416
  );


  buf
  g442
  (
    n564,
    n401
  );


  not
  g443
  (
    n493,
    n447
  );


  buf
  g444
  (
    n512,
    n400
  );


  buf
  g445
  (
    n485,
    n399
  );


  not
  g446
  (
    n476,
    n451
  );


  not
  g447
  (
    n489,
    n399
  );


  not
  g448
  (
    n504,
    n452
  );


  buf
  g449
  (
    n474,
    n468
  );


  buf
  g450
  (
    n497,
    n463
  );


  not
  g451
  (
    n560,
    n467
  );


  buf
  g452
  (
    n541,
    n401
  );


  not
  g453
  (
    n470,
    n468
  );


  buf
  g454
  (
    n501,
    n450
  );


  not
  g455
  (
    n516,
    n397
  );


  buf
  g456
  (
    n500,
    n397
  );


  buf
  g457
  (
    n494,
    n451
  );


  buf
  g458
  (
    n549,
    n456
  );


  not
  g459
  (
    n505,
    n103
  );


  not
  g460
  (
    n561,
    n454
  );


  buf
  g461
  (
    n551,
    n18
  );


  not
  g462
  (
    n546,
    n450
  );


  buf
  g463
  (
    n514,
    n103
  );


  not
  g464
  (
    n499,
    n447
  );


  buf
  g465
  (
    n511,
    n402
  );


  not
  g466
  (
    n507,
    n465
  );


  buf
  g467
  (
    n491,
    n415
  );


  not
  g468
  (
    n556,
    n469
  );


  not
  g469
  (
    n563,
    n459
  );


  not
  g470
  (
    n530,
    n365
  );


  buf
  g471
  (
    n539,
    n396
  );


  buf
  g472
  (
    n517,
    n448
  );


  buf
  g473
  (
    n525,
    n453
  );


  buf
  g474
  (
    n550,
    n392
  );


  buf
  g475
  (
    n527,
    n463
  );


  not
  g476
  (
    n515,
    n459
  );


  buf
  g477
  (
    n498,
    n398
  );


  not
  g478
  (
    n557,
    n18
  );


  buf
  g479
  (
    n554,
    n453
  );


  not
  g480
  (
    n534,
    n459
  );


  not
  g481
  (
    n486,
    n466
  );


  buf
  g482
  (
    n529,
    n17
  );


  not
  g483
  (
    n536,
    n103
  );


  buf
  g484
  (
    n490,
    n458
  );


  buf
  g485
  (
    n537,
    n464
  );


  not
  g486
  (
    n492,
    n469
  );


  buf
  g487
  (
    n508,
    n456
  );


  not
  g488
  (
    n479,
    n394
  );


  not
  g489
  (
    n503,
    n466
  );


  buf
  g490
  (
    n535,
    n462
  );


  xnor
  g491
  (
    n472,
    n467,
    n453,
    n459
  );


  or
  g492
  (
    n544,
    n324,
    n394,
    n446
  );


  nor
  g493
  (
    n510,
    n452,
    n395,
    n101
  );


  nor
  g494
  (
    n526,
    n402,
    n399,
    n398
  );


  nor
  g495
  (
    n545,
    n456,
    n467,
    n465
  );


  nor
  g496
  (
    n518,
    n450,
    n464,
    n455
  );


  and
  g497
  (
    n484,
    n457,
    n446,
    n396
  );


  xnor
  g498
  (
    n559,
    n458,
    n393,
    n395
  );


  nor
  g499
  (
    n548,
    n415,
    n398,
    n468
  );


  xor
  g500
  (
    n471,
    n467,
    n403,
    n396
  );


  xor
  g501
  (
    n480,
    n102,
    n466,
    n463
  );


  xor
  g502
  (
    n519,
    n464,
    n451,
    n461
  );


  and
  g503
  (
    n478,
    n397,
    n400,
    n452
  );


  xor
  g504
  (
    n520,
    n460,
    n404,
    n416
  );


  or
  g505
  (
    n523,
    n447,
    n403,
    n458
  );


  and
  g506
  (
    n552,
    n102,
    n413,
    n453
  );


  nand
  g507
  (
    n553,
    n393,
    n104,
    n413
  );


  xor
  g508
  (
    n562,
    n461,
    n462,
    n450
  );


  xor
  g509
  (
    n540,
    n392,
    n446,
    n393
  );


  nor
  g510
  (
    n502,
    n449,
    n458,
    n104
  );


  nand
  g511
  (
    n542,
    n402,
    n395,
    n416
  );


  and
  g512
  (
    n475,
    n399,
    n400,
    n446
  );


  nor
  g513
  (
    n555,
    n401,
    n462,
    n102
  );


  and
  g514
  (
    n473,
    n461,
    n101,
    n414
  );


  xor
  g515
  (
    n483,
    n414,
    n415,
    n395
  );


  xor
  g516
  (
    n522,
    n398,
    n452,
    n457
  );


  xnor
  g517
  (
    n524,
    n449,
    n465,
    n455
  );


  or
  g518
  (
    n513,
    n414,
    n400,
    n456
  );


  or
  g519
  (
    n528,
    n402,
    n394,
    n454
  );


  xor
  g520
  (
    n521,
    n447,
    n455,
    n457
  );


  xor
  g521
  (
    n477,
    n396,
    n404
  );


  or
  g522
  (
    n543,
    n449,
    n455,
    n461
  );


  nand
  g523
  (
    n558,
    n414,
    n460,
    n469
  );


  nand
  g524
  (
    n496,
    n415,
    n466,
    n449
  );


  or
  g525
  (
    n482,
    n464,
    n403,
    n401
  );


  xnor
  g526
  (
    n509,
    n416,
    n454
  );


  xor
  g527
  (
    n547,
    n460,
    n463,
    n457
  );


  xor
  g528
  (
    n488,
    n462,
    n394,
    n448
  );


  and
  g529
  (
    n495,
    n468,
    n448,
    n397
  );


  nand
  g530
  (
    n538,
    n460,
    n18,
    n404
  );


  and
  g531
  (
    n506,
    n465,
    n403,
    n103
  );


  or
  g532
  (
    n738,
    n495,
    n476,
    n225,
    n173
  );


  or
  g533
  (
    n625,
    n144,
    n182,
    n196,
    n104
  );


  xor
  g534
  (
    n635,
    n121,
    n206,
    n133,
    n221
  );


  nor
  g535
  (
    n644,
    n133,
    n491,
    n514,
    n486
  );


  xor
  g536
  (
    n803,
    n220,
    n217,
    n479,
    n473
  );


  and
  g537
  (
    n655,
    n166,
    n515,
    n480,
    n107
  );


  xor
  g538
  (
    n742,
    n116,
    n237,
    n494,
    n234
  );


  xor
  g539
  (
    n748,
    n254,
    n486,
    n513,
    n184
  );


  xor
  g540
  (
    n676,
    n276,
    n470,
    n266,
    n278
  );


  nor
  g541
  (
    n791,
    n199,
    n432,
    n147,
    n477
  );


  nor
  g542
  (
    n628,
    n173,
    n224,
    n115,
    n201
  );


  and
  g543
  (
    n609,
    n162,
    n274,
    n146,
    n520
  );


  nand
  g544
  (
    n566,
    n254,
    n471,
    n507,
    n128
  );


  xor
  g545
  (
    n781,
    n236,
    n121,
    n252,
    n166
  );


  xor
  g546
  (
    n769,
    n196,
    n526,
    n529,
    n165
  );


  nor
  g547
  (
    n712,
    n174,
    n481,
    n259,
    n154
  );


  xor
  g548
  (
    n577,
    n206,
    n239,
    n247,
    n117
  );


  and
  g549
  (
    n706,
    n516,
    n499,
    n479,
    n510
  );


  xor
  g550
  (
    n693,
    n277,
    n161,
    n494,
    n137
  );


  xnor
  g551
  (
    n787,
    n270,
    n231,
    n108,
    n222
  );


  xor
  g552
  (
    n740,
    n271,
    n137,
    n135,
    n142
  );


  nand
  g553
  (
    n623,
    n210,
    n160,
    n510,
    n405
  );


  nor
  g554
  (
    n802,
    n154,
    n144,
    n248,
    n512
  );


  and
  g555
  (
    n749,
    n493,
    n131,
    n127,
    n429
  );


  nor
  g556
  (
    n689,
    n267,
    n220,
    n138,
    n122
  );


  xor
  g557
  (
    n801,
    n250,
    n488,
    n122,
    n269
  );


  xor
  g558
  (
    n729,
    n203,
    n478,
    n508,
    n135
  );


  xnor
  g559
  (
    n745,
    n230,
    n264,
    n485,
    n184
  );


  and
  g560
  (
    n732,
    n148,
    n154,
    n482,
    n211
  );


  and
  g561
  (
    n670,
    n157,
    n272,
    n405,
    n522
  );


  nor
  g562
  (
    n698,
    n405,
    n153,
    n228,
    n520
  );


  and
  g563
  (
    n647,
    n153,
    n147,
    n197,
    n485
  );


  and
  g564
  (
    n649,
    n111,
    n158,
    n185,
    n524
  );


  xor
  g565
  (
    n757,
    n152,
    n110,
    n174,
    n519
  );


  xnor
  g566
  (
    n643,
    n497,
    n528,
    n525,
    n195
  );


  nand
  g567
  (
    n597,
    n131,
    n489,
    n238,
    n244
  );


  nand
  g568
  (
    n768,
    n175,
    n171,
    n114,
    n111
  );


  xor
  g569
  (
    n719,
    n430,
    n185,
    n194,
    n271
  );


  xnor
  g570
  (
    n614,
    n269,
    n503,
    n481,
    n166
  );


  nor
  g571
  (
    n630,
    n151,
    n145,
    n184,
    n256
  );


  or
  g572
  (
    n733,
    n172,
    n152,
    n236,
    n139
  );


  nand
  g573
  (
    n793,
    n118,
    n259,
    n169,
    n127
  );


  nand
  g574
  (
    n708,
    n219,
    n178,
    n110,
    n180
  );


  and
  g575
  (
    n619,
    n276,
    n498,
    n120,
    n251
  );


  nand
  g576
  (
    n761,
    n480,
    n183,
    n251,
    n509
  );


  xor
  g577
  (
    n578,
    n273,
    n105,
    n109,
    n202
  );


  and
  g578
  (
    n794,
    n124,
    n480,
    n526,
    n266
  );


  or
  g579
  (
    n595,
    n208,
    n156,
    n152,
    n240
  );


  or
  g580
  (
    n701,
    n475,
    n189,
    n478,
    n473
  );


  nor
  g581
  (
    n717,
    n209,
    n139,
    n202,
    n106
  );


  xnor
  g582
  (
    n603,
    n279,
    n491,
    n131,
    n212
  );


  nand
  g583
  (
    n798,
    n274,
    n116,
    n205,
    n494
  );


  or
  g584
  (
    n568,
    n526,
    n253,
    n120,
    n251
  );


  xor
  g585
  (
    n796,
    n218,
    n159,
    n496,
    n206
  );


  nand
  g586
  (
    n621,
    n513,
    n144,
    n234,
    n203
  );


  nand
  g587
  (
    n610,
    n268,
    n471,
    n256,
    n119
  );


  and
  g588
  (
    n661,
    n482,
    n242,
    n183,
    n212
  );


  nand
  g589
  (
    n799,
    n253,
    n221,
    n268,
    n111
  );


  or
  g590
  (
    n611,
    n164,
    n518,
    n172,
    n499
  );


  nor
  g591
  (
    n687,
    n265,
    n228,
    n138,
    n497
  );


  nand
  g592
  (
    n574,
    n109,
    n501,
    n505,
    n157
  );


  or
  g593
  (
    n778,
    n248,
    n488,
    n268,
    n505
  );


  nor
  g594
  (
    n713,
    n370,
    n263,
    n132,
    n495
  );


  nor
  g595
  (
    n772,
    n171,
    n506,
    n242,
    n524
  );


  xnor
  g596
  (
    n572,
    n235,
    n192,
    n263,
    n527
  );


  nand
  g597
  (
    n800,
    n221,
    n107,
    n246,
    n182
  );


  nand
  g598
  (
    n764,
    n235,
    n274,
    n213,
    n241
  );


  nand
  g599
  (
    n656,
    n493,
    n519,
    n470,
    n142
  );


  nand
  g600
  (
    n645,
    n161,
    n226,
    n109,
    n241
  );


  or
  g601
  (
    n722,
    n479,
    n474,
    n250,
    n153
  );


  nor
  g602
  (
    n771,
    n515,
    n274,
    n140
  );


  xnor
  g603
  (
    n770,
    n485,
    n245,
    n145,
    n181
  );


  nand
  g604
  (
    n784,
    n474,
    n160,
    n216,
    n229
  );


  or
  g605
  (
    n581,
    n124,
    n228,
    n475,
    n496
  );


  and
  g606
  (
    n721,
    n499,
    n232,
    n210,
    n162
  );


  or
  g607
  (
    n631,
    n204,
    n181,
    n115,
    n270
  );


  xnor
  g608
  (
    n684,
    n161,
    n197,
    n225,
    n230
  );


  nand
  g609
  (
    n753,
    n504,
    n496,
    n176,
    n173
  );


  xnor
  g610
  (
    n598,
    n235,
    n260,
    n504,
    n229
  );


  nor
  g611
  (
    n620,
    n175,
    n240,
    n262,
    n511
  );


  nand
  g612
  (
    n567,
    n500,
    n126,
    n187,
    n512
  );


  or
  g613
  (
    n695,
    n185,
    n162,
    n263,
    n249
  );


  or
  g614
  (
    n589,
    n428,
    n128,
    n239
  );


  nand
  g615
  (
    n629,
    n147,
    n474,
    n517,
    n271
  );


  nor
  g616
  (
    n606,
    n233,
    n169,
    n242,
    n155
  );


  xnor
  g617
  (
    n667,
    n206,
    n254,
    n227,
    n224
  );


  xor
  g618
  (
    n780,
    n471,
    n498,
    n132,
    n275
  );


  and
  g619
  (
    n744,
    n499,
    n151,
    n106,
    n167
  );


  nor
  g620
  (
    n680,
    n495,
    n515,
    n106,
    n268
  );


  or
  g621
  (
    n677,
    n180,
    n278,
    n264,
    n218
  );


  nor
  g622
  (
    n710,
    n232,
    n178,
    n158,
    n249
  );


  xor
  g623
  (
    n754,
    n510,
    n148,
    n504,
    n521
  );


  xnor
  g624
  (
    n590,
    n528,
    n130,
    n258,
    n139
  );


  nand
  g625
  (
    n736,
    n209,
    n477,
    n520,
    n252
  );


  or
  g626
  (
    KeyWire_0_5,
    n140,
    n266,
    n134,
    n216
  );


  and
  g627
  (
    n636,
    n107,
    n112,
    n248,
    n260
  );


  nand
  g628
  (
    n613,
    n489,
    n502,
    n132,
    n246
  );


  xnor
  g629
  (
    n776,
    n136,
    n201,
    n203,
    n212
  );


  xor
  g630
  (
    n783,
    n172,
    n175,
    n181,
    n177
  );


  nand
  g631
  (
    n594,
    n182,
    n179,
    n118,
    n260
  );


  xnor
  g632
  (
    n569,
    n514,
    n214,
    n141,
    n243
  );


  nand
  g633
  (
    n755,
    n209,
    n472,
    n490,
    n186
  );


  xor
  g634
  (
    n583,
    n523,
    n199,
    n119,
    n156
  );


  xnor
  g635
  (
    n660,
    n245,
    n161,
    n124,
    n191
  );


  xnor
  g636
  (
    n585,
    n168,
    n142,
    n140,
    n506
  );


  xnor
  g637
  (
    n751,
    n258,
    n473,
    n475,
    n511
  );


  xor
  g638
  (
    n599,
    n197,
    n168,
    n509,
    n234
  );


  and
  g639
  (
    n612,
    n507,
    n487,
    n488,
    n264
  );


  xor
  g640
  (
    n675,
    n245,
    n511,
    n150,
    n255
  );


  nor
  g641
  (
    n699,
    n149,
    n198,
    n492,
    n522
  );


  nor
  g642
  (
    n663,
    n265,
    n257,
    n126,
    n237
  );


  xnor
  g643
  (
    n724,
    n180,
    n147,
    n126,
    n186
  );


  nor
  g644
  (
    n705,
    n164,
    n160,
    n123,
    n195
  );


  xnor
  g645
  (
    n746,
    n500,
    n512,
    n227,
    n171
  );


  or
  g646
  (
    n664,
    n144,
    n522,
    n370,
    n278
  );


  nand
  g647
  (
    n634,
    n497,
    n256,
    n128,
    n189
  );


  xnor
  g648
  (
    n653,
    n519,
    n502,
    n214,
    n252
  );


  nand
  g649
  (
    n765,
    n258,
    n175,
    n476,
    n220
  );


  nor
  g650
  (
    n718,
    n223,
    n487,
    n278,
    n481
  );


  and
  g651
  (
    n694,
    n195,
    n261,
    n129,
    n484
  );


  xor
  g652
  (
    n767,
    n514,
    n240,
    n221,
    n210
  );


  and
  g653
  (
    n786,
    n254,
    n500,
    n244,
    n527
  );


  nand
  g654
  (
    n624,
    n202,
    n489,
    n154,
    n119
  );


  nand
  g655
  (
    n602,
    n115,
    n188,
    n143,
    n170
  );


  nor
  g656
  (
    n573,
    n222,
    n200,
    n226,
    n176
  );


  xor
  g657
  (
    n575,
    n213,
    n190,
    n492,
    n330
  );


  xnor
  g658
  (
    n674,
    n518,
    n493,
    n198,
    n523
  );


  nand
  g659
  (
    n703,
    n169,
    n227,
    n259,
    n272
  );


  nor
  g660
  (
    n604,
    n267,
    n130,
    n483,
    n179
  );


  nor
  g661
  (
    n692,
    n135,
    n112,
    n242,
    n157
  );


  xnor
  g662
  (
    KeyWire_0_9,
    n198,
    n196,
    n529,
    n238
  );


  xor
  g663
  (
    n659,
    n152,
    n518,
    n502,
    n150
  );


  and
  g664
  (
    n587,
    n243,
    n163,
    n149
  );


  nand
  g665
  (
    n788,
    n191,
    n215,
    n108,
    n273
  );


  nor
  g666
  (
    n766,
    n119,
    n247,
    n513,
    n507
  );


  and
  g667
  (
    n608,
    n190,
    n277,
    n145,
    n192
  );


  xor
  g668
  (
    n571,
    n250,
    n233,
    n483,
    n179
  );


  xor
  g669
  (
    n691,
    n488,
    n136,
    n146,
    n195
  );


  or
  g670
  (
    n642,
    n222,
    n483,
    n137,
    n113
  );


  or
  g671
  (
    n743,
    n527,
    n187,
    n157,
    n138
  );


  nor
  g672
  (
    n633,
    n115,
    n143,
    n208
  );


  and
  g673
  (
    n707,
    n170,
    n217,
    n508,
    n126
  );


  nor
  g674
  (
    n641,
    n159,
    n517,
    n165,
    n194
  );


  and
  g675
  (
    n618,
    n150,
    n502,
    n136,
    n487
  );


  xor
  g676
  (
    n709,
    n262,
    n190,
    n198,
    n113
  );


  xor
  g677
  (
    n741,
    n112,
    n486,
    n472,
    n160
  );


  xor
  g678
  (
    n711,
    n470,
    n273,
    n519,
    n370
  );


  nor
  g679
  (
    n605,
    n516,
    n229,
    n141,
    n247
  );


  nand
  g680
  (
    n622,
    n130,
    n110,
    n480,
    n262
  );


  xor
  g681
  (
    n762,
    n507,
    n238,
    n225,
    n210
  );


  nor
  g682
  (
    n596,
    n216,
    n528,
    n200,
    n231
  );


  nor
  g683
  (
    n588,
    n505,
    n476,
    n188,
    n146
  );


  and
  g684
  (
    n627,
    n267,
    n259,
    n264,
    n182
  );


  xnor
  g685
  (
    n720,
    n163,
    n118,
    n233,
    n204
  );


  xnor
  g686
  (
    n580,
    n271,
    n508,
    n263,
    n155
  );


  nor
  g687
  (
    n731,
    n269,
    n174,
    n169,
    n168
  );


  xor
  g688
  (
    n593,
    n201,
    n223,
    n473,
    n162
  );


  or
  g689
  (
    n678,
    n257,
    n471,
    n125,
    n501
  );


  or
  g690
  (
    n730,
    n474,
    n127,
    n483,
    n170
  );


  nor
  g691
  (
    n739,
    n166,
    n193,
    n176,
    n248
  );


  and
  g692
  (
    n752,
    n214,
    n477,
    n494,
    n120
  );


  and
  g693
  (
    n782,
    n500,
    n112,
    n183,
    n232
  );


  nor
  g694
  (
    n673,
    n191,
    n219,
    n232,
    n164
  );


  xnor
  g695
  (
    n640,
    n238,
    n186,
    n170,
    n224
  );


  xor
  g696
  (
    n747,
    n224,
    n158,
    n218,
    n129
  );


  or
  g697
  (
    n756,
    n496,
    n521,
    n241,
    n272
  );


  xor
  g698
  (
    n734,
    n236,
    n176,
    n189,
    n244
  );


  nor
  g699
  (
    n658,
    n201,
    n516,
    n117,
    n218
  );


  xor
  g700
  (
    n626,
    n484,
    n514,
    n117,
    n125
  );


  xnor
  g701
  (
    n576,
    n159,
    n521,
    n527,
    n233
  );


  xor
  g702
  (
    n688,
    n177,
    n433,
    n482,
    n491
  );


  xnor
  g703
  (
    n637,
    n197,
    n146,
    n155,
    n105
  );


  or
  g704
  (
    n760,
    n205,
    n114,
    n526,
    n156
  );


  and
  g705
  (
    n570,
    n192,
    n199,
    n128,
    n275
  );


  nand
  g706
  (
    n639,
    n167,
    n490,
    n117,
    n183
  );


  xnor
  g707
  (
    n671,
    n501,
    n246,
    n164,
    n107
  );


  nand
  g708
  (
    n617,
    n165,
    n106,
    n225,
    n243
  );


  or
  g709
  (
    n727,
    n217,
    n226,
    n475,
    n213
  );


  and
  g710
  (
    n775,
    n498,
    n267,
    n260,
    n129
  );


  and
  g711
  (
    n565,
    n511,
    n143,
    n145,
    n345
  );


  xnor
  g712
  (
    n790,
    n118,
    n528,
    n153,
    n151
  );


  xnor
  g713
  (
    n792,
    n524,
    n205,
    n165,
    n196
  );


  xnor
  g714
  (
    n696,
    n212,
    n249,
    n132,
    n523
  );


  nand
  g715
  (
    n763,
    n134,
    n220,
    n192,
    n188
  );


  xor
  g716
  (
    n615,
    n184,
    n215,
    n275,
    n187
  );


  xor
  g717
  (
    n579,
    n227,
    n481,
    n123,
    n251
  );


  or
  g718
  (
    n607,
    n174,
    n492,
    n148,
    n155
  );


  nor
  g719
  (
    n672,
    n492,
    n114,
    n130,
    n270
  );


  nor
  g720
  (
    n591,
    n234,
    n205,
    n250,
    n215
  );


  or
  g721
  (
    n686,
    n127,
    n110,
    n185,
    n133
  );


  xor
  g722
  (
    n714,
    n487,
    n194,
    n108,
    n252
  );


  nand
  g723
  (
    n704,
    n525,
    n269,
    n270,
    n524
  );


  nand
  g724
  (
    n669,
    n490,
    n482,
    n529,
    n240
  );


  or
  g725
  (
    n726,
    n199,
    n256,
    n262,
    n219
  );


  or
  g726
  (
    n654,
    n178,
    n261,
    n190,
    n504
  );


  nand
  g727
  (
    n584,
    n266,
    n523,
    n211,
    n136
  );


  nor
  g728
  (
    n690,
    n116,
    n223,
    n204,
    n173
  );


  xor
  g729
  (
    n582,
    n503,
    n405,
    n207,
    n521
  );


  xnor
  g730
  (
    n648,
    n172,
    n211,
    n123,
    n134
  );


  nand
  g731
  (
    n668,
    n141,
    n188,
    n193,
    n213
  );


  xnor
  g732
  (
    n681,
    n472,
    n167,
    n277,
    n237
  );


  nand
  g733
  (
    n666,
    n207,
    n503,
    n191,
    n479
  );


  or
  g734
  (
    n702,
    n509,
    n484,
    n125,
    n209
  );


  xnor
  g735
  (
    n592,
    n498,
    n104,
    n223,
    n508
  );


  or
  g736
  (
    n662,
    n503,
    n253,
    n133,
    n151
  );


  xnor
  g737
  (
    n728,
    n178,
    n520,
    n163,
    n109
  );


  nor
  g738
  (
    n773,
    n275,
    n241,
    n505,
    n276
  );


  xnor
  g739
  (
    n586,
    n189,
    n485,
    n129,
    n497
  );


  and
  g740
  (
    n665,
    n517,
    n489,
    n207,
    n491
  );


  and
  g741
  (
    n758,
    n230,
    n139,
    n200,
    n219
  );


  nand
  g742
  (
    n683,
    n510,
    n186,
    n237,
    n258
  );


  xnor
  g743
  (
    n774,
    n194,
    n214,
    n167,
    n249
  );


  or
  g744
  (
    n716,
    n141,
    n493,
    n484,
    n114
  );


  nor
  g745
  (
    n652,
    n478,
    n203,
    n231,
    n193
  );


  nor
  g746
  (
    n759,
    n517,
    n228,
    n168,
    n265
  );


  and
  g747
  (
    n601,
    n229,
    n486,
    n277,
    n113
  );


  nand
  g748
  (
    n638,
    n120,
    n134,
    n222,
    n142
  );


  nand
  g749
  (
    n700,
    n159,
    n180,
    n121,
    n193
  );


  xnor
  g750
  (
    n735,
    n501,
    n207,
    n243,
    n226
  );


  and
  g751
  (
    n785,
    n113,
    n512,
    n434,
    n490
  );


  nand
  g752
  (
    n650,
    n495,
    n122,
    n135,
    n272
  );


  and
  g753
  (
    n795,
    n478,
    n516,
    n137,
    n122
  );


  and
  g754
  (
    n685,
    n200,
    n208,
    n171,
    n177
  );


  nand
  g755
  (
    n723,
    n131,
    n181,
    n111,
    n245
  );


  xnor
  g756
  (
    n646,
    n211,
    n253,
    n509,
    n235
  );


  nor
  g757
  (
    n616,
    n149,
    n476,
    n231,
    n116
  );


  xnor
  g758
  (
    n682,
    n525,
    n124,
    n470,
    n247
  );


  nand
  g759
  (
    n715,
    n255,
    n156,
    n216,
    n257
  );


  nand
  g760
  (
    KeyWire_0_18,
    n177,
    n204,
    n506,
    n158
  );


  and
  g761
  (
    n777,
    n265,
    n255,
    n261,
    n506
  );


  and
  g762
  (
    n750,
    n513,
    n431,
    n125,
    n108
  );


  nand
  g763
  (
    n797,
    n244,
    n257,
    n525,
    n150
  );


  nor
  g764
  (
    n789,
    n515,
    n121,
    n217,
    n105
  );


  nor
  g765
  (
    n657,
    n143,
    n261,
    n518,
    n123
  );


  or
  g766
  (
    n632,
    n105,
    n255,
    n276,
    n163
  );


  nand
  g767
  (
    n600,
    n472,
    n522,
    n239,
    n279
  );


  and
  g768
  (
    KeyWire_0_31,
    n215,
    n273,
    n187,
    n148
  );


  and
  g769
  (
    n651,
    n477,
    n179,
    n246,
    n370
  );


  or
  g770
  (
    n679,
    n202,
    n230,
    n236,
    n138
  );


  not
  g771
  (
    n998,
    n741
  );


  buf
  g772
  (
    n1116,
    n694
  );


  not
  g773
  (
    n1518,
    n702
  );


  buf
  g774
  (
    n1388,
    n585
  );


  not
  g775
  (
    n1090,
    n720
  );


  buf
  g776
  (
    n937,
    n581
  );


  buf
  g777
  (
    n1265,
    n732
  );


  buf
  g778
  (
    n1063,
    n794
  );


  not
  g779
  (
    n1638,
    n750
  );


  buf
  g780
  (
    n973,
    n676
  );


  buf
  g781
  (
    n1375,
    n788
  );


  buf
  g782
  (
    n975,
    n759
  );


  buf
  g783
  (
    n1315,
    n587
  );


  buf
  g784
  (
    n1425,
    n752
  );


  not
  g785
  (
    n1312,
    n627
  );


  not
  g786
  (
    n1166,
    n640
  );


  buf
  g787
  (
    n1724,
    n331
  );


  not
  g788
  (
    n905,
    n770
  );


  not
  g789
  (
    n807,
    n707
  );


  not
  g790
  (
    n1377,
    n791
  );


  buf
  g791
  (
    n1629,
    n653
  );


  not
  g792
  (
    n1616,
    n676
  );


  buf
  g793
  (
    n1172,
    n656
  );


  buf
  g794
  (
    n865,
    n663
  );


  not
  g795
  (
    n1115,
    n791
  );


  not
  g796
  (
    n892,
    n653
  );


  buf
  g797
  (
    n1209,
    n710
  );


  not
  g798
  (
    n1514,
    n682
  );


  buf
  g799
  (
    n1142,
    n789
  );


  not
  g800
  (
    n1089,
    n753
  );


  not
  g801
  (
    n1319,
    n598
  );


  not
  g802
  (
    n1485,
    n631
  );


  not
  g803
  (
    n1646,
    n708
  );


  not
  g804
  (
    n1422,
    n782
  );


  buf
  g805
  (
    n1126,
    n685
  );


  not
  g806
  (
    n1134,
    n768
  );


  not
  g807
  (
    n1570,
    n794
  );


  not
  g808
  (
    n1573,
    n700
  );


  not
  g809
  (
    n972,
    n566
  );


  not
  g810
  (
    n854,
    n643
  );


  buf
  g811
  (
    n1269,
    n773
  );


  not
  g812
  (
    KeyWire_0_10,
    n585
  );


  buf
  g813
  (
    n1510,
    n444
  );


  not
  g814
  (
    n1230,
    n629
  );


  buf
  g815
  (
    n1176,
    n594
  );


  not
  g816
  (
    n899,
    n776
  );


  not
  g817
  (
    n1586,
    n604
  );


  not
  g818
  (
    n1179,
    n766
  );


  buf
  g819
  (
    n826,
    n795
  );


  buf
  g820
  (
    n1195,
    n287
  );


  buf
  g821
  (
    n871,
    n716
  );


  not
  g822
  (
    n1049,
    n569
  );


  buf
  g823
  (
    n1019,
    n694
  );


  not
  g824
  (
    n1363,
    n335
  );


  buf
  g825
  (
    n894,
    n731
  );


  buf
  g826
  (
    n1196,
    n736
  );


  buf
  g827
  (
    n1007,
    n782
  );


  buf
  g828
  (
    n1017,
    n751
  );


  not
  g829
  (
    n1520,
    n608
  );


  not
  g830
  (
    KeyWire_0_27,
    n664
  );


  buf
  g831
  (
    n1270,
    n740
  );


  not
  g832
  (
    n1060,
    n743
  );


  buf
  g833
  (
    n1608,
    n598
  );


  not
  g834
  (
    n1087,
    n644
  );


  not
  g835
  (
    n1550,
    n672
  );


  buf
  g836
  (
    n1306,
    n719
  );


  not
  g837
  (
    n1342,
    n781
  );


  buf
  g838
  (
    n1181,
    n292
  );


  not
  g839
  (
    n1512,
    n661
  );


  buf
  g840
  (
    n1393,
    n786
  );


  not
  g841
  (
    n1033,
    n787
  );


  not
  g842
  (
    n1591,
    n716
  );


  buf
  g843
  (
    n1385,
    n713
  );


  not
  g844
  (
    n1748,
    n751
  );


  not
  g845
  (
    n1036,
    n658
  );


  not
  g846
  (
    n1291,
    n572
  );


  not
  g847
  (
    n1031,
    n753
  );


  buf
  g848
  (
    n939,
    n784
  );


  buf
  g849
  (
    n1352,
    n675
  );


  buf
  g850
  (
    n1530,
    n689
  );


  buf
  g851
  (
    n1233,
    n713
  );


  not
  g852
  (
    n1649,
    n672
  );


  not
  g853
  (
    n1636,
    n573
  );


  not
  g854
  (
    n1073,
    n593
  );


  buf
  g855
  (
    n1424,
    n286
  );


  not
  g856
  (
    n847,
    n444
  );


  not
  g857
  (
    n1466,
    n611
  );


  not
  g858
  (
    n919,
    n673
  );


  not
  g859
  (
    n1370,
    n284
  );


  buf
  g860
  (
    n1286,
    n579
  );


  buf
  g861
  (
    n853,
    n623
  );


  not
  g862
  (
    n1117,
    n685
  );


  buf
  g863
  (
    n1039,
    n630
  );


  buf
  g864
  (
    n1340,
    n783
  );


  not
  g865
  (
    n1524,
    n769
  );


  not
  g866
  (
    n1605,
    n708
  );


  buf
  g867
  (
    n1462,
    n794
  );


  buf
  g868
  (
    n1202,
    n776
  );


  buf
  g869
  (
    n1307,
    n282
  );


  not
  g870
  (
    n1034,
    n620
  );


  not
  g871
  (
    n1584,
    n653
  );


  not
  g872
  (
    n1075,
    n578
  );


  buf
  g873
  (
    n1184,
    n678
  );


  not
  g874
  (
    n886,
    n596
  );


  buf
  g875
  (
    n1238,
    n756
  );


  not
  g876
  (
    n1305,
    n769
  );


  buf
  g877
  (
    n1679,
    n761
  );


  not
  g878
  (
    n1441,
    n569
  );


  not
  g879
  (
    n952,
    n729
  );


  not
  g880
  (
    n1384,
    n722
  );


  buf
  g881
  (
    n1250,
    n623
  );


  not
  g882
  (
    n947,
    n632
  );


  buf
  g883
  (
    n1062,
    n679
  );


  not
  g884
  (
    n815,
    n686
  );


  buf
  g885
  (
    n1501,
    n696
  );


  buf
  g886
  (
    n1430,
    n582
  );


  buf
  g887
  (
    n1664,
    n603
  );


  not
  g888
  (
    n1735,
    n788
  );


  buf
  g889
  (
    n1506,
    n605
  );


  not
  g890
  (
    n1741,
    n702
  );


  not
  g891
  (
    n1752,
    n799
  );


  not
  g892
  (
    n1137,
    n603
  );


  not
  g893
  (
    n1277,
    n597
  );


  buf
  g894
  (
    n1403,
    n691
  );


  not
  g895
  (
    n839,
    n671
  );


  not
  g896
  (
    n1658,
    n714
  );


  not
  g897
  (
    n1394,
    n752
  );


  buf
  g898
  (
    n1251,
    n650
  );


  not
  g899
  (
    n1604,
    n621
  );


  not
  g900
  (
    n1589,
    n639
  );


  buf
  g901
  (
    n1734,
    n684
  );


  buf
  g902
  (
    n1634,
    n604
  );


  buf
  g903
  (
    n1279,
    n633
  );


  not
  g904
  (
    n1171,
    n666
  );


  not
  g905
  (
    n1438,
    n717
  );


  buf
  g906
  (
    n834,
    n284
  );


  buf
  g907
  (
    n946,
    n589
  );


  buf
  g908
  (
    n860,
    n763
  );


  buf
  g909
  (
    n1022,
    n701
  );


  not
  g910
  (
    n1200,
    n331
  );


  buf
  g911
  (
    n1402,
    n583
  );


  not
  g912
  (
    n1443,
    n674
  );


  buf
  g913
  (
    n1526,
    n724
  );


  not
  g914
  (
    n1472,
    n680
  );


  not
  g915
  (
    n1127,
    n662
  );


  not
  g916
  (
    n902,
    n634
  );


  buf
  g917
  (
    n1220,
    n738
  );


  buf
  g918
  (
    n1482,
    n734
  );


  buf
  g919
  (
    n1560,
    n659
  );


  buf
  g920
  (
    n1387,
    n608
  );


  not
  g921
  (
    n1552,
    n780
  );


  buf
  g922
  (
    n1667,
    n287
  );


  buf
  g923
  (
    n1397,
    n684
  );


  buf
  g924
  (
    n862,
    n747
  );


  not
  g925
  (
    n938,
    n710
  );


  not
  g926
  (
    n909,
    n595
  );


  buf
  g927
  (
    n1427,
    n592
  );


  not
  g928
  (
    n1657,
    n618
  );


  not
  g929
  (
    n1678,
    n728
  );


  not
  g930
  (
    n1040,
    n689
  );


  not
  g931
  (
    n933,
    n675
  );


  buf
  g932
  (
    n1298,
    n670
  );


  buf
  g933
  (
    n995,
    n625
  );


  not
  g934
  (
    n1476,
    n765
  );


  buf
  g935
  (
    n1350,
    n802
  );


  buf
  g936
  (
    n829,
    n656
  );


  not
  g937
  (
    n968,
    n688
  );


  not
  g938
  (
    n1600,
    n748
  );


  not
  g939
  (
    KeyWire_0_29,
    n633
  );


  not
  g940
  (
    n1177,
    n746
  );


  not
  g941
  (
    n1288,
    n645
  );


  not
  g942
  (
    n1732,
    n627
  );


  not
  g943
  (
    n1050,
    n783
  );


  buf
  g944
  (
    n949,
    n626
  );


  not
  g945
  (
    n1626,
    n625
  );


  not
  g946
  (
    n1351,
    n727
  );


  buf
  g947
  (
    n1241,
    n612
  );


  not
  g948
  (
    n1395,
    n333
  );


  buf
  g949
  (
    n816,
    n335
  );


  not
  g950
  (
    n1738,
    n669
  );


  buf
  g951
  (
    n1318,
    n281
  );


  buf
  g952
  (
    n1149,
    n773
  );


  buf
  g953
  (
    n1416,
    n580
  );


  buf
  g954
  (
    n1454,
    n756
  );


  buf
  g955
  (
    n1631,
    n585
  );


  buf
  g956
  (
    n1122,
    n683
  );


  not
  g957
  (
    n1689,
    n744
  );


  buf
  g958
  (
    n1446,
    n332
  );


  not
  g959
  (
    n1577,
    n777
  );


  buf
  g960
  (
    n1301,
    n802
  );


  buf
  g961
  (
    n1190,
    n587
  );


  not
  g962
  (
    n948,
    n753
  );


  buf
  g963
  (
    n1376,
    n288
  );


  not
  g964
  (
    n1615,
    n759
  );


  buf
  g965
  (
    n1541,
    n654
  );


  not
  g966
  (
    n1575,
    n694
  );


  buf
  g967
  (
    n1228,
    n772
  );


  not
  g968
  (
    n817,
    n715
  );


  not
  g969
  (
    n1107,
    n760
  );


  not
  g970
  (
    n1408,
    n705
  );


  not
  g971
  (
    n1165,
    n606
  );


  buf
  g972
  (
    n1725,
    n568
  );


  buf
  g973
  (
    n1313,
    n592
  );


  not
  g974
  (
    n858,
    n725
  );


  not
  g975
  (
    n1145,
    n601
  );


  not
  g976
  (
    n1272,
    n748
  );


  not
  g977
  (
    n923,
    n622
  );


  buf
  g978
  (
    n1110,
    n751
  );


  not
  g979
  (
    n1215,
    n758
  );


  buf
  g980
  (
    n1358,
    n607
  );


  not
  g981
  (
    n883,
    n734
  );


  not
  g982
  (
    n1094,
    n692
  );


  buf
  g983
  (
    n1392,
    n682
  );


  not
  g984
  (
    n962,
    n443
  );


  buf
  g985
  (
    n893,
    n789
  );


  buf
  g986
  (
    n1688,
    n693
  );


  not
  g987
  (
    n1225,
    n589
  );


  not
  g988
  (
    n1364,
    n690
  );


  not
  g989
  (
    n1593,
    n734
  );


  not
  g990
  (
    n1002,
    n660
  );


  buf
  g991
  (
    n1681,
    n776
  );


  buf
  g992
  (
    n1295,
    n605
  );


  buf
  g993
  (
    n1661,
    n610
  );


  not
  g994
  (
    n852,
    n570
  );


  not
  g995
  (
    n980,
    n598
  );


  buf
  g996
  (
    n1044,
    n656
  );


  not
  g997
  (
    n875,
    n599
  );


  not
  g998
  (
    n969,
    n763
  );


  not
  g999
  (
    n1515,
    n624
  );


  buf
  g1000
  (
    n1452,
    n654
  );


  buf
  g1001
  (
    n1598,
    n622
  );


  buf
  g1002
  (
    n1739,
    n579
  );


  buf
  g1003
  (
    n1458,
    n580
  );


  buf
  g1004
  (
    n812,
    n600
  );


  buf
  g1005
  (
    n1339,
    n788
  );


  buf
  g1006
  (
    n1474,
    n576
  );


  buf
  g1007
  (
    n1133,
    n678
  );


  buf
  g1008
  (
    n895,
    n721
  );


  not
  g1009
  (
    n943,
    n626
  );


  not
  g1010
  (
    n976,
    n620
  );


  not
  g1011
  (
    n934,
    n285
  );


  not
  g1012
  (
    n920,
    n731
  );


  buf
  g1013
  (
    n1096,
    n644
  );


  buf
  g1014
  (
    n1255,
    n758
  );


  not
  g1015
  (
    n1420,
    n789
  );


  buf
  g1016
  (
    n1614,
    n688
  );


  not
  g1017
  (
    n907,
    n730
  );


  not
  g1018
  (
    n1609,
    n610
  );


  buf
  g1019
  (
    n1456,
    n594
  );


  buf
  g1020
  (
    n906,
    n679
  );


  not
  g1021
  (
    n1348,
    n725
  );


  not
  g1022
  (
    n1354,
    n718
  );


  buf
  g1023
  (
    n1652,
    n444
  );


  not
  g1024
  (
    n1193,
    n654
  );


  not
  g1025
  (
    n1459,
    n331
  );


  buf
  g1026
  (
    n842,
    n683
  );


  not
  g1027
  (
    n1123,
    n721
  );


  buf
  g1028
  (
    n1449,
    n597
  );


  not
  g1029
  (
    n1302,
    n616
  );


  buf
  g1030
  (
    n1199,
    n723
  );


  not
  g1031
  (
    n874,
    n654
  );


  buf
  g1032
  (
    KeyWire_0_26,
    n598
  );


  buf
  g1033
  (
    n818,
    n692
  );


  not
  g1034
  (
    n1071,
    n779
  );


  not
  g1035
  (
    n846,
    n803
  );


  not
  g1036
  (
    n1296,
    n630
  );


  buf
  g1037
  (
    n1747,
    n737
  );


  buf
  g1038
  (
    n1677,
    n667
  );


  not
  g1039
  (
    n925,
    n735
  );


  not
  g1040
  (
    n1189,
    n290
  );


  not
  g1041
  (
    n1009,
    n713
  );


  not
  g1042
  (
    n1246,
    n684
  );


  buf
  g1043
  (
    n960,
    n782
  );


  not
  g1044
  (
    n915,
    n736
  );


  not
  g1045
  (
    n970,
    n727
  );


  not
  g1046
  (
    n1360,
    n721
  );


  buf
  g1047
  (
    n1730,
    n575
  );


  not
  g1048
  (
    n1637,
    n762
  );


  buf
  g1049
  (
    n819,
    n592
  );


  buf
  g1050
  (
    n832,
    n597
  );


  buf
  g1051
  (
    n1599,
    n682
  );


  not
  g1052
  (
    n1610,
    n717
  );


  buf
  g1053
  (
    n1281,
    n641
  );


  not
  g1054
  (
    n1755,
    n605
  );


  not
  g1055
  (
    n1536,
    n784
  );


  not
  g1056
  (
    n977,
    n653
  );


  buf
  g1057
  (
    n1559,
    n803
  );


  buf
  g1058
  (
    n877,
    n800
  );


  buf
  g1059
  (
    n1240,
    n590
  );


  buf
  g1060
  (
    n896,
    n442
  );


  buf
  g1061
  (
    n1128,
    n665
  );


  buf
  g1062
  (
    n1381,
    n668
  );


  not
  g1063
  (
    n1700,
    n672
  );


  not
  g1064
  (
    n1380,
    n606
  );


  buf
  g1065
  (
    n1194,
    n745
  );


  not
  g1066
  (
    n1065,
    n660
  );


  buf
  g1067
  (
    n979,
    n741
  );


  not
  g1068
  (
    n965,
    n712
  );


  buf
  g1069
  (
    n1164,
    n569
  );


  buf
  g1070
  (
    n1205,
    n768
  );


  buf
  g1071
  (
    n1201,
    n285
  );


  not
  g1072
  (
    n1345,
    n740
  );


  buf
  g1073
  (
    n1275,
    n671
  );


  not
  g1074
  (
    n1051,
    n787
  );


  buf
  g1075
  (
    n974,
    n716
  );


  not
  g1076
  (
    n876,
    n702
  );


  buf
  g1077
  (
    n1743,
    n286
  );


  not
  g1078
  (
    n1426,
    n770
  );


  not
  g1079
  (
    n1157,
    n607
  );


  not
  g1080
  (
    n1447,
    n599
  );


  not
  g1081
  (
    n1642,
    n335
  );


  buf
  g1082
  (
    n1135,
    n754
  );


  buf
  g1083
  (
    n929,
    n733
  );


  buf
  g1084
  (
    n917,
    n617
  );


  not
  g1085
  (
    n1278,
    n724
  );


  buf
  g1086
  (
    n1571,
    n785
  );


  not
  g1087
  (
    n1576,
    n767
  );


  buf
  g1088
  (
    n1254,
    n681
  );


  not
  g1089
  (
    n1655,
    n675
  );


  buf
  g1090
  (
    n1486,
    n577
  );


  not
  g1091
  (
    n1706,
    n790
  );


  buf
  g1092
  (
    n1746,
    n771
  );


  not
  g1093
  (
    n1043,
    n674
  );


  not
  g1094
  (
    n1156,
    n590
  );


  not
  g1095
  (
    n1182,
    n686
  );


  buf
  g1096
  (
    n1758,
    n602
  );


  buf
  g1097
  (
    n1736,
    n737
  );


  buf
  g1098
  (
    n1226,
    n715
  );


  buf
  g1099
  (
    n1492,
    n597
  );


  not
  g1100
  (
    n1692,
    n649
  );


  not
  g1101
  (
    n1332,
    n334
  );


  not
  g1102
  (
    n994,
    n614
  );


  buf
  g1103
  (
    n1085,
    n679
  );


  not
  g1104
  (
    n811,
    n589
  );


  buf
  g1105
  (
    n1558,
    n789
  );


  not
  g1106
  (
    n1026,
    n778
  );


  buf
  g1107
  (
    n1542,
    n763
  );


  not
  g1108
  (
    n857,
    n737
  );


  buf
  g1109
  (
    n1588,
    n801
  );


  not
  g1110
  (
    KeyWire_0_2,
    n577
  );


  buf
  g1111
  (
    n809,
    n588
  );


  not
  g1112
  (
    n1231,
    n676
  );


  buf
  g1113
  (
    n1622,
    n750
  );


  not
  g1114
  (
    n870,
    n638
  );


  buf
  g1115
  (
    n1054,
    n573
  );


  not
  g1116
  (
    n1670,
    n680
  );


  buf
  g1117
  (
    n1058,
    n703
  );


  buf
  g1118
  (
    n1084,
    n762
  );


  not
  g1119
  (
    n1068,
    n657
  );


  buf
  g1120
  (
    n990,
    n780
  );


  not
  g1121
  (
    n913,
    n646
  );


  not
  g1122
  (
    n935,
    n665
  );


  buf
  g1123
  (
    n1432,
    n609
  );


  buf
  g1124
  (
    n982,
    n599
  );


  buf
  g1125
  (
    n898,
    n745
  );


  buf
  g1126
  (
    n1021,
    n691
  );


  buf
  g1127
  (
    n1322,
    n652
  );


  not
  g1128
  (
    n903,
    n699
  );


  buf
  g1129
  (
    n955,
    n750
  );


  buf
  g1130
  (
    n901,
    n621
  );


  not
  g1131
  (
    n1701,
    n707
  );


  not
  g1132
  (
    n971,
    n750
  );


  buf
  g1133
  (
    n1038,
    n734
  );


  not
  g1134
  (
    n1263,
    n601
  );


  not
  g1135
  (
    n837,
    n740
  );


  not
  g1136
  (
    n1330,
    n740
  );


  not
  g1137
  (
    n1258,
    n793
  );


  buf
  g1138
  (
    n1168,
    n749
  );


  not
  g1139
  (
    n1715,
    n757
  );


  buf
  g1140
  (
    n1079,
    n775
  );


  buf
  g1141
  (
    n1704,
    n764
  );


  buf
  g1142
  (
    n1709,
    n615
  );


  buf
  g1143
  (
    n880,
    n571
  );


  not
  g1144
  (
    n1641,
    n768
  );


  buf
  g1145
  (
    n823,
    n793
  );


  not
  g1146
  (
    n991,
    n797
  );


  not
  g1147
  (
    n1434,
    n593
  );


  buf
  g1148
  (
    n1186,
    n665
  );


  not
  g1149
  (
    n1047,
    n707
  );


  not
  g1150
  (
    n1544,
    n786
  );


  buf
  g1151
  (
    n1372,
    n571
  );


  buf
  g1152
  (
    n1523,
    n690
  );


  not
  g1153
  (
    n1656,
    n634
  );


  buf
  g1154
  (
    n1460,
    n650
  );


  buf
  g1155
  (
    n1208,
    n793
  );


  buf
  g1156
  (
    n1378,
    n331
  );


  not
  g1157
  (
    n957,
    n291
  );


  not
  g1158
  (
    n1653,
    n784
  );


  buf
  g1159
  (
    n1003,
    n738
  );


  not
  g1160
  (
    n1522,
    n677
  );


  buf
  g1161
  (
    n1273,
    n634
  );


  not
  g1162
  (
    n1143,
    n591
  );


  buf
  g1163
  (
    n1662,
    n772
  );


  not
  g1164
  (
    n1628,
    n636
  );


  not
  g1165
  (
    n1369,
    n798
  );


  buf
  g1166
  (
    n981,
    n333
  );


  not
  g1167
  (
    n1669,
    n720
  );


  buf
  g1168
  (
    n1750,
    n641
  );


  buf
  g1169
  (
    n1727,
    n678
  );


  not
  g1170
  (
    n1401,
    n668
  );


  buf
  g1171
  (
    n1547,
    n659
  );


  not
  g1172
  (
    n1495,
    n781
  );


  not
  g1173
  (
    n1180,
    n642
  );


  buf
  g1174
  (
    n1578,
    n741
  );


  buf
  g1175
  (
    n1723,
    n748
  );


  not
  g1176
  (
    n1102,
    n778
  );


  not
  g1177
  (
    n1448,
    n747
  );


  not
  g1178
  (
    n1083,
    n762
  );


  buf
  g1179
  (
    n1491,
    n755
  );


  buf
  g1180
  (
    n1070,
    n612
  );


  buf
  g1181
  (
    n1644,
    n723
  );


  buf
  g1182
  (
    n986,
    n568
  );


  not
  g1183
  (
    n1611,
    n751
  );


  buf
  g1184
  (
    n864,
    n777
  );


  not
  g1185
  (
    n1519,
    n619
  );


  buf
  g1186
  (
    n1707,
    n733
  );


  buf
  g1187
  (
    n1030,
    n643
  );


  not
  g1188
  (
    KeyWire_0_28,
    n747
  );


  not
  g1189
  (
    n1632,
    n712
  );


  not
  g1190
  (
    n1645,
    n565
  );


  buf
  g1191
  (
    n1234,
    n685
  );


  buf
  g1192
  (
    n940,
    n681
  );


  not
  g1193
  (
    n1243,
    n602
  );


  buf
  g1194
  (
    n944,
    n644
  );


  buf
  g1195
  (
    n890,
    n656
  );


  buf
  g1196
  (
    n1696,
    n698
  );


  not
  g1197
  (
    n1546,
    n689
  );


  not
  g1198
  (
    n1502,
    n629
  );


  buf
  g1199
  (
    n1311,
    n761
  );


  not
  g1200
  (
    n824,
    n645
  );


  not
  g1201
  (
    n1170,
    n775
  );


  buf
  g1202
  (
    n827,
    n611
  );


  not
  g1203
  (
    n1721,
    n671
  );


  not
  g1204
  (
    n951,
    n697
  );


  not
  g1205
  (
    n1192,
    n717
  );


  buf
  g1206
  (
    n1647,
    n442
  );


  not
  g1207
  (
    n1555,
    n673
  );


  not
  g1208
  (
    n1290,
    n575
  );


  not
  g1209
  (
    n1297,
    n636
  );


  not
  g1210
  (
    n1093,
    n288
  );


  not
  g1211
  (
    n921,
    n573
  );


  not
  g1212
  (
    n1672,
    n617
  );


  buf
  g1213
  (
    n887,
    n726
  );


  not
  g1214
  (
    n1141,
    n801
  );


  buf
  g1215
  (
    n1590,
    n739
  );


  buf
  g1216
  (
    n1211,
    n582
  );


  buf
  g1217
  (
    n1504,
    n766
  );


  not
  g1218
  (
    n1595,
    n336
  );


  not
  g1219
  (
    n1057,
    n575
  );


  buf
  g1220
  (
    n1483,
    n759
  );


  buf
  g1221
  (
    n1334,
    n770
  );


  not
  g1222
  (
    n1248,
    n730
  );


  buf
  g1223
  (
    n1371,
    n670
  );


  not
  g1224
  (
    n1139,
    n742
  );


  not
  g1225
  (
    n1722,
    n744
  );


  not
  g1226
  (
    n1053,
    n703
  );


  buf
  g1227
  (
    n1415,
    n767
  );


  not
  g1228
  (
    n999,
    n677
  );


  buf
  g1229
  (
    n1437,
    n637
  );


  not
  g1230
  (
    n1130,
    n291
  );


  buf
  g1231
  (
    n1496,
    n687
  );


  not
  g1232
  (
    n1262,
    n593
  );


  buf
  g1233
  (
    n1567,
    n631
  );


  buf
  g1234
  (
    n1292,
    n291
  );


  buf
  g1235
  (
    n1316,
    n756
  );


  buf
  g1236
  (
    n855,
    n664
  );


  not
  g1237
  (
    n950,
    n652
  );


  buf
  g1238
  (
    n1239,
    n618
  );


  buf
  g1239
  (
    n1016,
    n643
  );


  not
  g1240
  (
    n931,
    n284
  );


  buf
  g1241
  (
    n996,
    n602
  );


  not
  g1242
  (
    n873,
    n729
  );


  buf
  g1243
  (
    n1191,
    n632
  );


  buf
  g1244
  (
    n1745,
    n630
  );


  buf
  g1245
  (
    n966,
    n651
  );


  buf
  g1246
  (
    n1630,
    n695
  );


  buf
  g1247
  (
    n1751,
    n764
  );


  buf
  g1248
  (
    n1445,
    n719
  );


  not
  g1249
  (
    n848,
    n761
  );


  not
  g1250
  (
    n1582,
    n626
  );


  not
  g1251
  (
    n964,
    n732
  );


  not
  g1252
  (
    n1303,
    n594
  );


  buf
  g1253
  (
    n1359,
    n649
  );


  buf
  g1254
  (
    n861,
    n661
  );


  buf
  g1255
  (
    n1411,
    n719
  );


  not
  g1256
  (
    n1687,
    n736
  );


  not
  g1257
  (
    n1042,
    n688
  );


  not
  g1258
  (
    n1711,
    n668
  );


  not
  g1259
  (
    n918,
    n642
  );


  not
  g1260
  (
    n1601,
    n691
  );


  buf
  g1261
  (
    n1635,
    n650
  );


  not
  g1262
  (
    n1285,
    n670
  );


  not
  g1263
  (
    n1431,
    n679
  );


  buf
  g1264
  (
    n1185,
    n678
  );


  buf
  g1265
  (
    n1710,
    n796
  );


  buf
  g1266
  (
    n1321,
    n700
  );


  not
  g1267
  (
    n841,
    n692
  );


  not
  g1268
  (
    n1158,
    n626
  );


  buf
  g1269
  (
    n1235,
    n665
  );


  not
  g1270
  (
    n1001,
    n600
  );


  buf
  g1271
  (
    n1581,
    n611
  );


  buf
  g1272
  (
    n1338,
    n674
  );


  not
  g1273
  (
    n1543,
    n281
  );


  buf
  g1274
  (
    n1607,
    n289
  );


  not
  g1275
  (
    n1173,
    n615
  );


  buf
  g1276
  (
    n1175,
    n760
  );


  not
  g1277
  (
    n1357,
    n783
  );


  not
  g1278
  (
    n1695,
    n619
  );


  buf
  g1279
  (
    n1624,
    n579
  );


  buf
  g1280
  (
    n1423,
    n633
  );


  not
  g1281
  (
    n1569,
    n565
  );


  not
  g1282
  (
    n1497,
    n568
  );


  buf
  g1283
  (
    n1507,
    n614
  );


  not
  g1284
  (
    n958,
    n687
  );


  buf
  g1285
  (
    n814,
    n767
  );


  buf
  g1286
  (
    n1680,
    n798
  );


  not
  g1287
  (
    n1245,
    n798
  );


  not
  g1288
  (
    n1405,
    n601
  );


  buf
  g1289
  (
    n1602,
    n285
  );


  not
  g1290
  (
    n1685,
    n753
  );


  buf
  g1291
  (
    n1064,
    n586
  );


  buf
  g1292
  (
    n1503,
    n640
  );


  not
  g1293
  (
    n1355,
    n744
  );


  not
  g1294
  (
    n926,
    n647
  );


  buf
  g1295
  (
    n912,
    n584
  );


  not
  g1296
  (
    n1744,
    n774
  );


  buf
  g1297
  (
    n1549,
    n625
  );


  not
  g1298
  (
    n1341,
    n683
  );


  buf
  g1299
  (
    n1095,
    n655
  );


  buf
  g1300
  (
    n821,
    n332
  );


  not
  g1301
  (
    n1525,
    n667
  );


  not
  g1302
  (
    n1451,
    n591
  );


  not
  g1303
  (
    n1082,
    n715
  );


  buf
  g1304
  (
    n1106,
    n771
  );


  not
  g1305
  (
    n1187,
    n737
  );


  not
  g1306
  (
    n1236,
    n680
  );


  not
  g1307
  (
    n1621,
    n667
  );


  not
  g1308
  (
    n1478,
    n663
  );


  not
  g1309
  (
    n1344,
    n780
  );


  buf
  g1310
  (
    n1216,
    n778
  );


  buf
  g1311
  (
    n1294,
    n661
  );


  not
  g1312
  (
    KeyWire_0_19,
    n624
  );


  not
  g1313
  (
    n1343,
    n582
  );


  not
  g1314
  (
    n1274,
    n754
  );


  not
  g1315
  (
    n930,
    n792
  );


  buf
  g1316
  (
    n1457,
    n635
  );


  not
  g1317
  (
    n1557,
    n773
  );


  not
  g1318
  (
    n1147,
    n603
  );


  buf
  g1319
  (
    n1024,
    n698
  );


  buf
  g1320
  (
    n1464,
    n721
  );


  not
  g1321
  (
    n1517,
    n607
  );


  not
  g1322
  (
    n1406,
    n775
  );


  buf
  g1323
  (
    n1153,
    n613
  );


  not
  g1324
  (
    n1583,
    n659
  );


  not
  g1325
  (
    n1154,
    n767
  );


  not
  g1326
  (
    n1639,
    n586
  );


  buf
  g1327
  (
    n1268,
    n627
  );


  not
  g1328
  (
    n888,
    n723
  );


  not
  g1329
  (
    n1465,
    n744
  );


  not
  g1330
  (
    n1072,
    n669
  );


  not
  g1331
  (
    n1121,
    n799
  );


  not
  g1332
  (
    n1613,
    n695
  );


  not
  g1333
  (
    n1148,
    n666
  );


  not
  g1334
  (
    n1708,
    n720
  );


  not
  g1335
  (
    n1487,
    n337
  );


  not
  g1336
  (
    n1623,
    n710
  );


  buf
  g1337
  (
    n916,
    n752
  );


  buf
  g1338
  (
    n1328,
    n607
  );


  not
  g1339
  (
    n1204,
    n279
  );


  buf
  g1340
  (
    n932,
    n631
  );


  buf
  g1341
  (
    n1553,
    n604
  );


  buf
  g1342
  (
    n820,
    n655
  );


  buf
  g1343
  (
    n1561,
    n443
  );


  not
  g1344
  (
    n1280,
    n795
  );


  not
  g1345
  (
    n1717,
    n775
  );


  not
  g1346
  (
    n1712,
    n583
  );


  not
  g1347
  (
    n1222,
    n727
  );


  buf
  g1348
  (
    n1221,
    n619
  );


  not
  g1349
  (
    n1442,
    n596
  );


  buf
  g1350
  (
    n810,
    n773
  );


  not
  g1351
  (
    n1564,
    n660
  );


  not
  g1352
  (
    n1421,
    n567
  );


  buf
  g1353
  (
    n1264,
    n442
  );


  buf
  g1354
  (
    n1067,
    n581
  );


  buf
  g1355
  (
    n1011,
    n798
  );


  buf
  g1356
  (
    n1702,
    n699
  );


  buf
  g1357
  (
    n1594,
    n735
  );


  buf
  g1358
  (
    n1556,
    n577
  );


  not
  g1359
  (
    n1046,
    n615
  );


  buf
  g1360
  (
    KeyWire_0_13,
    n780
  );


  buf
  g1361
  (
    n1206,
    n729
  );


  buf
  g1362
  (
    n1138,
    n803
  );


  buf
  g1363
  (
    n1467,
    n614
  );


  buf
  g1364
  (
    n808,
    n688
  );


  not
  g1365
  (
    n1548,
    n285
  );


  buf
  g1366
  (
    n1320,
    n570
  );


  buf
  g1367
  (
    n1155,
    n648
  );


  not
  g1368
  (
    n1373,
    n445
  );


  buf
  g1369
  (
    n1488,
    n620
  );


  buf
  g1370
  (
    n1618,
    n693
  );


  not
  g1371
  (
    n1580,
    n797
  );


  buf
  g1372
  (
    n1109,
    n754
  );


  not
  g1373
  (
    n885,
    n728
  );


  not
  g1374
  (
    n1534,
    n445
  );


  buf
  g1375
  (
    n1284,
    n612
  );


  not
  g1376
  (
    n1150,
    n795
  );


  buf
  g1377
  (
    n825,
    n786
  );


  not
  g1378
  (
    n1061,
    n724
  );


  buf
  g1379
  (
    n1006,
    n781
  );


  not
  g1380
  (
    n1362,
    n722
  );


  not
  g1381
  (
    n1572,
    n283
  );


  buf
  g1382
  (
    n1643,
    n579
  );


  buf
  g1383
  (
    n1152,
    n657
  );


  buf
  g1384
  (
    n1412,
    n782
  );


  not
  g1385
  (
    n1249,
    n284
  );


  not
  g1386
  (
    n872,
    n283
  );


  not
  g1387
  (
    n1379,
    n781
  );


  buf
  g1388
  (
    n1640,
    n777
  );


  not
  g1389
  (
    n1203,
    n733
  );


  buf
  g1390
  (
    n963,
    n635
  );


  not
  g1391
  (
    n1100,
    n628
  );


  not
  g1392
  (
    n804,
    n648
  );


  buf
  g1393
  (
    n1161,
    n584
  );


  not
  g1394
  (
    n1390,
    n722
  );


  not
  g1395
  (
    n987,
    n637
  );


  not
  g1396
  (
    n941,
    n586
  );


  buf
  g1397
  (
    n1045,
    n698
  );


  not
  g1398
  (
    n1086,
    n790
  );


  buf
  g1399
  (
    n1048,
    n709
  );


  not
  g1400
  (
    n840,
    n600
  );


  not
  g1401
  (
    n866,
    n333
  );


  not
  g1402
  (
    n1365,
    n697
  );


  not
  g1403
  (
    n850,
    n739
  );


  buf
  g1404
  (
    n1521,
    n609
  );


  buf
  g1405
  (
    n1532,
    n762
  );


  buf
  g1406
  (
    n1223,
    n636
  );


  not
  g1407
  (
    n868,
    n783
  );


  buf
  g1408
  (
    n1252,
    n779
  );


  buf
  g1409
  (
    n1596,
    n280
  );


  not
  g1410
  (
    n1673,
    n742
  );


  buf
  g1411
  (
    n1293,
    n765
  );


  buf
  g1412
  (
    n1214,
    n714
  );


  not
  g1413
  (
    n1120,
    n289
  );


  buf
  g1414
  (
    n1674,
    n601
  );


  buf
  g1415
  (
    n1247,
    n726
  );


  buf
  g1416
  (
    n1317,
    n281
  );


  buf
  g1417
  (
    n1097,
    n292
  );


  buf
  g1418
  (
    n1705,
    n574
  );


  not
  g1419
  (
    n1417,
    n687
  );


  buf
  g1420
  (
    n1101,
    n681
  );


  buf
  g1421
  (
    n1675,
    n719
  );


  buf
  g1422
  (
    n1718,
    n689
  );


  buf
  g1423
  (
    n1074,
    n749
  );


  buf
  g1424
  (
    n845,
    n610
  );


  buf
  g1425
  (
    n924,
    n743
  );


  buf
  g1426
  (
    n922,
    n755
  );


  not
  g1427
  (
    n1551,
    n787
  );


  not
  g1428
  (
    n1012,
    n712
  );


  buf
  g1429
  (
    n1720,
    n732
  );


  buf
  g1430
  (
    n908,
    n771
  );


  buf
  g1431
  (
    n1025,
    n677
  );


  not
  g1432
  (
    n836,
    n705
  );


  buf
  g1433
  (
    n1217,
    n332
  );


  not
  g1434
  (
    n1740,
    n661
  );


  buf
  g1435
  (
    n1309,
    n609
  );


  not
  g1436
  (
    n1105,
    n709
  );


  buf
  g1437
  (
    n1163,
    n443
  );


  not
  g1438
  (
    n1513,
    n731
  );


  not
  g1439
  (
    n997,
    n638
  );


  buf
  g1440
  (
    n1260,
    n625
  );


  not
  g1441
  (
    n1013,
    n760
  );


  buf
  g1442
  (
    n956,
    n722
  );


  buf
  g1443
  (
    n1690,
    n755
  );


  buf
  g1444
  (
    n1052,
    n595
  );


  buf
  g1445
  (
    n1331,
    n287
  );


  not
  g1446
  (
    n1140,
    n637
  );


  not
  g1447
  (
    n1509,
    n746
  );


  buf
  g1448
  (
    n1207,
    n694
  );


  buf
  g1449
  (
    n1537,
    n648
  );


  buf
  g1450
  (
    n1253,
    n591
  );


  buf
  g1451
  (
    KeyWire_0_21,
    n290
  );


  not
  g1452
  (
    n1516,
    n705
  );


  not
  g1453
  (
    n1539,
    n758
  );


  not
  g1454
  (
    n1475,
    n282
  );


  not
  g1455
  (
    n1471,
    n618
  );


  buf
  g1456
  (
    n1112,
    n748
  );


  not
  g1457
  (
    n1136,
    n697
  );


  not
  g1458
  (
    n1308,
    n769
  );


  buf
  g1459
  (
    n1683,
    n667
  );


  buf
  g1460
  (
    n1368,
    n635
  );


  not
  g1461
  (
    n1118,
    n645
  );


  not
  g1462
  (
    n1620,
    n638
  );


  not
  g1463
  (
    n1346,
    n441
  );


  buf
  g1464
  (
    n863,
    n599
  );


  not
  g1465
  (
    n1473,
    n707
  );


  buf
  g1466
  (
    n1035,
    n596
  );


  not
  g1467
  (
    n1479,
    n442
  );


  not
  g1468
  (
    n1111,
    n571
  );


  buf
  g1469
  (
    n1389,
    n745
  );


  not
  g1470
  (
    n1232,
    n704
  );


  buf
  g1471
  (
    n1167,
    n566
  );


  not
  g1472
  (
    n1477,
    n743
  );


  buf
  g1473
  (
    n822,
    n647
  );


  buf
  g1474
  (
    n1757,
    n790
  );


  buf
  g1475
  (
    n1124,
    n727
  );


  not
  g1476
  (
    n1028,
    n700
  );


  buf
  g1477
  (
    n1099,
    n663
  );


  not
  g1478
  (
    n1625,
    n736
  );


  not
  g1479
  (
    n1545,
    n770
  );


  not
  g1480
  (
    n891,
    n578
  );


  not
  g1481
  (
    n1261,
    n779
  );


  not
  g1482
  (
    n851,
    n730
  );


  buf
  g1483
  (
    n992,
    n752
  );


  not
  g1484
  (
    n1023,
    n666
  );


  not
  g1485
  (
    n1579,
    n570
  );


  not
  g1486
  (
    n1304,
    n608
  );


  not
  g1487
  (
    n1396,
    n711
  );


  not
  g1488
  (
    n910,
    n668
  );


  buf
  g1489
  (
    n1493,
    n583
  );


  buf
  g1490
  (
    n1455,
    n596
  );


  buf
  g1491
  (
    n1733,
    n763
  );


  not
  g1492
  (
    n1335,
    n643
  );


  not
  g1493
  (
    n878,
    n288
  );


  buf
  g1494
  (
    n985,
    n765
  );


  buf
  g1495
  (
    n1666,
    n589
  );


  not
  g1496
  (
    n1500,
    n639
  );


  buf
  g1497
  (
    n1450,
    n776
  );


  buf
  g1498
  (
    n1654,
    n657
  );


  buf
  g1499
  (
    n1386,
    n720
  );


  buf
  g1500
  (
    n988,
    n617
  );


  buf
  g1501
  (
    n1587,
    n673
  );


  not
  g1502
  (
    n1227,
    n706
  );


  not
  g1503
  (
    n1742,
    n569
  );


  buf
  g1504
  (
    n1256,
    n606
  );


  buf
  g1505
  (
    n961,
    n778
  );


  not
  g1506
  (
    n1612,
    n608
  );


  not
  g1507
  (
    n884,
    n445
  );


  buf
  g1508
  (
    n989,
    n712
  );


  not
  g1509
  (
    n1027,
    n757
  );


  buf
  g1510
  (
    n1538,
    n584
  );


  buf
  g1511
  (
    n1490,
    n704
  );


  buf
  g1512
  (
    n867,
    n772
  );


  buf
  g1513
  (
    n1324,
    n621
  );


  not
  g1514
  (
    n1729,
    n745
  );


  buf
  g1515
  (
    KeyWire_0_25,
    n800
  );


  buf
  g1516
  (
    n1480,
    n337
  );


  buf
  g1517
  (
    n984,
    n704
  );


  buf
  g1518
  (
    n1310,
    n731
  );


  buf
  g1519
  (
    n1029,
    n588
  );


  not
  g1520
  (
    n1282,
    n690
  );


  not
  g1521
  (
    n1146,
    n704
  );


  not
  g1522
  (
    n1103,
    n576
  );


  not
  g1523
  (
    n1129,
    n570
  );


  buf
  g1524
  (
    n805,
    n718
  );


  not
  g1525
  (
    n1508,
    n725
  );


  not
  g1526
  (
    n828,
    n337
  );


  buf
  g1527
  (
    n1682,
    n703
  );


  not
  g1528
  (
    n1108,
    n669
  );


  not
  g1529
  (
    n897,
    n706
  );


  not
  g1530
  (
    n1574,
    n290
  );


  buf
  g1531
  (
    n1603,
    n613
  );


  buf
  g1532
  (
    n1383,
    n711
  );


  not
  g1533
  (
    n1257,
    n685
  );


  not
  g1534
  (
    n1686,
    n638
  );


  buf
  g1535
  (
    n1759,
    n609
  );


  buf
  g1536
  (
    n1119,
    n610
  );


  not
  g1537
  (
    n1059,
    n683
  );


  buf
  g1538
  (
    n1726,
    n787
  );


  buf
  g1539
  (
    n1407,
    n622
  );


  buf
  g1540
  (
    n1714,
    n774
  );


  not
  g1541
  (
    n1218,
    n649
  );


  buf
  g1542
  (
    n1756,
    n588
  );


  buf
  g1543
  (
    n1213,
    n760
  );


  not
  g1544
  (
    n1337,
    n662
  );


  buf
  g1545
  (
    n1113,
    n703
  );


  buf
  g1546
  (
    n1410,
    n282
  );


  buf
  g1547
  (
    n1433,
    n749
  );


  not
  g1548
  (
    n1400,
    n292
  );


  not
  g1549
  (
    n1511,
    n799
  );


  not
  g1550
  (
    n843,
    n797
  );


  buf
  g1551
  (
    n978,
    n648
  );


  not
  g1552
  (
    n1098,
    n684
  );


  not
  g1553
  (
    n1716,
    n660
  );


  not
  g1554
  (
    n1699,
    n673
  );


  not
  g1555
  (
    n833,
    n642
  );


  buf
  g1556
  (
    n1088,
    n615
  );


  buf
  g1557
  (
    n1453,
    n288
  );


  not
  g1558
  (
    n900,
    n735
  );


  buf
  g1559
  (
    n1470,
    n766
  );


  buf
  g1560
  (
    n1648,
    n714
  );


  buf
  g1561
  (
    n869,
    n441
  );


  not
  g1562
  (
    n1436,
    n644
  );


  not
  g1563
  (
    n1032,
    n581
  );


  not
  g1564
  (
    n1463,
    n580
  );


  buf
  g1565
  (
    n1676,
    n701
  );


  buf
  g1566
  (
    n1353,
    n590
  );


  buf
  g1567
  (
    n1287,
    n759
  );


  buf
  g1568
  (
    n1527,
    n624
  );


  buf
  g1569
  (
    n1399,
    n622
  );


  buf
  g1570
  (
    n1440,
    n746
  );


  not
  g1571
  (
    n1435,
    n696
  );


  not
  g1572
  (
    n1325,
    n651
  );


  not
  g1573
  (
    n1592,
    n290
  );


  buf
  g1574
  (
    n1041,
    n777
  );


  buf
  g1575
  (
    n889,
    n803
  );


  buf
  g1576
  (
    n859,
    n701
  );


  not
  g1577
  (
    n1266,
    n676
  );


  not
  g1578
  (
    n1056,
    n647
  );


  buf
  g1579
  (
    n1754,
    n572
  );


  buf
  g1580
  (
    n1698,
    n802
  );


  not
  g1581
  (
    n1439,
    n796
  );


  buf
  g1582
  (
    n1242,
    n664
  );


  buf
  g1583
  (
    n1531,
    n792
  );


  buf
  g1584
  (
    n1244,
    n717
  );


  buf
  g1585
  (
    KeyWire_0_7,
    n280
  );


  not
  g1586
  (
    n1259,
    n595
  );


  buf
  g1587
  (
    n1498,
    n730
  );


  buf
  g1588
  (
    n1336,
    n779
  );


  buf
  g1589
  (
    n1418,
    n670
  );


  buf
  g1590
  (
    n1229,
    n714
  );


  not
  g1591
  (
    n1633,
    n612
  );


  not
  g1592
  (
    n1568,
    n574
  );


  buf
  g1593
  (
    n1660,
    n629
  );


  not
  g1594
  (
    n1197,
    n739
  );


  not
  g1595
  (
    n1566,
    n791
  );


  buf
  g1596
  (
    n830,
    n443
  );


  buf
  g1597
  (
    n1684,
    n711
  );


  buf
  g1598
  (
    n1018,
    n632
  );


  not
  g1599
  (
    n1619,
    n718
  );


  not
  g1600
  (
    n1409,
    n772
  );


  buf
  g1601
  (
    n1753,
    n624
  );


  buf
  g1602
  (
    n1668,
    n738
  );


  not
  g1603
  (
    n1078,
    n591
  );


  not
  g1604
  (
    n1131,
    n666
  );


  not
  g1605
  (
    n1665,
    n604
  );


  not
  g1606
  (
    n881,
    n616
  );


  not
  g1607
  (
    n1008,
    n754
  );


  not
  g1608
  (
    n1004,
    n445
  );


  not
  g1609
  (
    n967,
    n287
  );


  not
  g1610
  (
    n1697,
    n592
  );


  not
  g1611
  (
    n1528,
    n646
  );


  buf
  g1612
  (
    n1162,
    n572
  );


  buf
  g1613
  (
    n1461,
    n649
  );


  buf
  g1614
  (
    n1367,
    n573
  );


  not
  g1615
  (
    n942,
    n336
  );


  not
  g1616
  (
    n1606,
    n801
  );


  buf
  g1617
  (
    n1289,
    n621
  );


  not
  g1618
  (
    n1198,
    n739
  );


  not
  g1619
  (
    n1219,
    n334
  );


  not
  g1620
  (
    n954,
    n686
  );


  not
  g1621
  (
    n1014,
    n692
  );


  buf
  g1622
  (
    n1428,
    n633
  );


  buf
  g1623
  (
    n838,
    n785
  );


  not
  g1624
  (
    n856,
    n659
  );


  not
  g1625
  (
    n1563,
    n441
  );


  not
  g1626
  (
    n1374,
    n581
  );


  buf
  g1627
  (
    n849,
    n600
  );


  buf
  g1628
  (
    n1010,
    n602
  );


  buf
  g1629
  (
    n1444,
    n619
  );


  buf
  g1630
  (
    n1469,
    n766
  );


  buf
  g1631
  (
    n1468,
    n657
  );


  not
  g1632
  (
    n1066,
    n794
  );


  not
  g1633
  (
    n1694,
    n711
  );


  not
  g1634
  (
    n831,
    n632
  );


  not
  g1635
  (
    n1271,
    n578
  );


  not
  g1636
  (
    n1617,
    n669
  );


  buf
  g1637
  (
    n1188,
    n614
  );


  not
  g1638
  (
    n1080,
    n696
  );


  not
  g1639
  (
    n1651,
    n567
  );


  not
  g1640
  (
    n1327,
    n774
  );


  buf
  g1641
  (
    n1055,
    n693
  );


  not
  g1642
  (
    n911,
    n690
  );


  not
  g1643
  (
    n1314,
    n628
  );


  buf
  g1644
  (
    n1020,
    n595
  );


  buf
  g1645
  (
    n1489,
    n332
  );


  not
  g1646
  (
    n914,
    n566
  );


  buf
  g1647
  (
    n1505,
    n769
  );


  buf
  g1648
  (
    n1554,
    n729
  );


  buf
  g1649
  (
    n1267,
    n802
  );


  buf
  g1650
  (
    n1015,
    n651
  );


  buf
  g1651
  (
    n1494,
    n732
  );


  not
  g1652
  (
    n1077,
    n701
  );


  not
  g1653
  (
    n1212,
    n664
  );


  not
  g1654
  (
    n1484,
    n695
  );


  buf
  g1655
  (
    n1535,
    n698
  );


  buf
  g1656
  (
    n806,
    n635
  );


  not
  g1657
  (
    n1414,
    n795
  );


  buf
  g1658
  (
    n1749,
    n636
  );


  not
  g1659
  (
    n1356,
    n680
  );


  not
  g1660
  (
    n1174,
    n705
  );


  buf
  g1661
  (
    n1404,
    n652
  );


  buf
  g1662
  (
    n1091,
    n337
  );


  buf
  g1663
  (
    n1125,
    n620
  );


  not
  g1664
  (
    n1671,
    n747
  );


  buf
  g1665
  (
    n1382,
    n741
  );


  buf
  g1666
  (
    n1659,
    n735
  );


  not
  g1667
  (
    n879,
    n786
  );


  buf
  g1668
  (
    n1585,
    n642
  );


  buf
  g1669
  (
    n993,
    n291
  );


  not
  g1670
  (
    n1540,
    n283
  );


  buf
  g1671
  (
    n1597,
    n662
  );


  not
  g1672
  (
    n959,
    n708
  );


  not
  g1673
  (
    n1104,
    n749
  );


  buf
  g1674
  (
    n928,
    n639
  );


  buf
  g1675
  (
    n945,
    n696
  );


  buf
  g1676
  (
    n927,
    n567
  );


  not
  g1677
  (
    n1650,
    n713
  );


  not
  g1678
  (
    n1159,
    n336
  );


  not
  g1679
  (
    n1481,
    n441
  );


  buf
  g1680
  (
    n1237,
    n583
  );


  buf
  g1681
  (
    n1160,
    n587
  );


  not
  g1682
  (
    n1731,
    n574
  );


  buf
  g1683
  (
    n1333,
    n765
  );


  not
  g1684
  (
    n1114,
    n576
  );


  not
  g1685
  (
    n1366,
    n791
  );


  not
  g1686
  (
    n1276,
    n333
  );


  not
  g1687
  (
    n1037,
    n797
  );


  buf
  g1688
  (
    n1210,
    n335
  );


  buf
  g1689
  (
    n1076,
    n584
  );


  buf
  g1690
  (
    n1224,
    n652
  );


  not
  g1691
  (
    n1326,
    n641
  );


  buf
  g1692
  (
    n1413,
    n286
  );


  or
  g1693
  (
    n1627,
    n606,
    n687,
    n576,
    n585
  );


  xor
  g1694
  (
    n1533,
    n651,
    n603,
    n718,
    n655
  );


  and
  g1695
  (
    n1391,
    n742,
    n686,
    n582,
    n761
  );


  and
  g1696
  (
    n1719,
    n706,
    n700,
    n755,
    n674
  );


  nand
  g1697
  (
    n1728,
    n623,
    n757,
    n662,
    n708
  );


  and
  g1698
  (
    n1499,
    n784,
    n710,
    n646,
    n675
  );


  and
  g1699
  (
    n1349,
    n618,
    n726,
    n616,
    n282
  );


  or
  g1700
  (
    n882,
    n672,
    n793,
    n280,
    n637
  );


  and
  g1701
  (
    n1361,
    n627,
    n724,
    n725,
    n774
  );


  xor
  g1702
  (
    n813,
    n697,
    n790,
    n663,
    n590
  );


  nor
  g1703
  (
    n1737,
    n580,
    n565,
    n764,
    n691
  );


  xor
  g1704
  (
    n1347,
    n699,
    n588,
    n655,
    n279
  );


  or
  g1705
  (
    n1691,
    n743,
    n593,
    n587,
    n631
  );


  and
  g1706
  (
    n1703,
    n628,
    n650,
    n567,
    n742
  );


  xor
  g1707
  (
    n835,
    n699,
    n716,
    n574,
    n785
  );


  nand
  g1708
  (
    n1178,
    n733,
    n628,
    n289,
    n286
  );


  or
  g1709
  (
    n1663,
    n799,
    n746,
    n646,
    n292
  );


  or
  g1710
  (
    KeyWire_0_17,
    n695,
    n681,
    n334,
    n623
  );


  nand
  g1711
  (
    n1169,
    n785,
    n800,
    n647,
    n578
  );


  xor
  g1712
  (
    n844,
    n594,
    n658,
    n726,
    n613
  );


  nor
  g1713
  (
    n1000,
    n792,
    n715,
    n709,
    n640
  );


  nand
  g1714
  (
    n953,
    n792,
    n788,
    n757,
    n728
  );


  nor
  g1715
  (
    n1398,
    n586,
    n616,
    n693,
    n575
  );


  or
  g1716
  (
    n1529,
    n702,
    n658,
    n577,
    n334
  );


  xnor
  g1717
  (
    n1562,
    n801,
    n605,
    n281,
    n283
  );


  nand
  g1718
  (
    n936,
    n682,
    n641,
    n768,
    n796
  );


  or
  g1719
  (
    n1713,
    n645,
    n630,
    n634,
    n796
  );


  and
  g1720
  (
    n1329,
    n756,
    n728,
    n444,
    n658
  );


  or
  g1721
  (
    n1693,
    n629,
    n565,
    n671,
    n289
  );


  and
  g1722
  (
    n1565,
    n758,
    n572,
    n800,
    n613
  );


  and
  g1723
  (
    n1419,
    n738,
    n723,
    n709,
    n706
  );


  xnor
  g1724
  (
    n1132,
    n764,
    n568,
    n617,
    n336
  );


  xnor
  g1725
  (
    n1299,
    n677,
    n566,
    n280,
    n640
  );


  nor
  g1726
  (
    n1069,
    n639,
    n571,
    n611,
    n771
  );


  nand
  g1727
  (
    n2095,
    n1198,
    n985,
    n1042,
    n1354
  );


  nand
  g1728
  (
    n2170,
    n1257,
    n1148,
    n960,
    n1232
  );


  or
  g1729
  (
    n2534,
    n1176,
    n1034,
    n1119,
    n1009
  );


  nand
  g1730
  (
    n2194,
    n1376,
    n1585,
    n1108,
    n1078
  );


  xor
  g1731
  (
    n2114,
    n985,
    n1203,
    n1601,
    n1407
  );


  xor
  g1732
  (
    n2243,
    n1572,
    n1691,
    n1158,
    n1501
  );


  xnor
  g1733
  (
    n1921,
    n1361,
    n1235,
    n1589,
    n1552
  );


  xor
  g1734
  (
    n2350,
    n1563,
    n1135,
    n1064,
    n1485
  );


  nand
  g1735
  (
    n2592,
    n1448,
    n1727,
    n1699,
    n1705
  );


  nand
  g1736
  (
    n2079,
    n1672,
    n1313,
    n1495,
    n1542
  );


  xnor
  g1737
  (
    n2614,
    n1431,
    n1200,
    n1504,
    n1267
  );


  and
  g1738
  (
    n2311,
    n1291,
    n1501,
    n1410,
    n870
  );


  nor
  g1739
  (
    n2284,
    n1357,
    n1345,
    n1124,
    n1680
  );


  and
  g1740
  (
    n1865,
    n1583,
    n1721,
    n1252,
    n1708
  );


  nand
  g1741
  (
    n2389,
    n1553,
    n930,
    n1090,
    n1619
  );


  or
  g1742
  (
    n1771,
    n1500,
    n971,
    n1551,
    n823
  );


  nand
  g1743
  (
    n2601,
    n1604,
    n808,
    n1390,
    n1741
  );


  and
  g1744
  (
    n2027,
    n1477,
    n1233,
    n1058,
    n1344
  );


  or
  g1745
  (
    n2555,
    n1524,
    n1141,
    n1393,
    n1330
  );


  xor
  g1746
  (
    n1945,
    n1189,
    n994,
    n1732,
    n1401
  );


  and
  g1747
  (
    KeyWire_0_1,
    n1737,
    n813,
    n1075,
    n1565
  );


  nand
  g1748
  (
    n2251,
    n1745,
    n1431,
    n1643,
    n1531
  );


  and
  g1749
  (
    n2588,
    n1412,
    n1009,
    n1143,
    n1442
  );


  nor
  g1750
  (
    n2538,
    n1026,
    n1240,
    n1402,
    n1149
  );


  and
  g1751
  (
    n2238,
    n992,
    n1084,
    n1633,
    n929
  );


  and
  g1752
  (
    n2424,
    n1571,
    n1087,
    n1144,
    n1011
  );


  nand
  g1753
  (
    n2207,
    n965,
    n1617,
    n947,
    n1638
  );


  nand
  g1754
  (
    n2356,
    n1691,
    n926,
    n1512,
    n1528
  );


  or
  g1755
  (
    n2595,
    n1481,
    n1463,
    n881,
    n995
  );


  and
  g1756
  (
    n2625,
    n1527,
    n1499,
    n1505,
    n1215
  );


  xnor
  g1757
  (
    n2341,
    n1293,
    n1621,
    n1270,
    n1195
  );


  and
  g1758
  (
    n2075,
    n1533,
    n1451,
    n1385,
    n1511
  );


  xnor
  g1759
  (
    n1892,
    n1274,
    n1376,
    n828,
    n837
  );


  xor
  g1760
  (
    n2044,
    n1141,
    n1461,
    n1154,
    n1128
  );


  and
  g1761
  (
    n2411,
    n1125,
    n1241,
    n1269,
    n1174
  );


  nor
  g1762
  (
    n1998,
    n1231,
    n991,
    n1377,
    n1507
  );


  xor
  g1763
  (
    n2276,
    n1243,
    n958,
    n1364,
    n1699
  );


  nand
  g1764
  (
    n2458,
    n1104,
    n1467,
    n1499,
    n817
  );


  xnor
  g1765
  (
    n2107,
    n1716,
    n1040,
    n1414,
    n1239
  );


  xnor
  g1766
  (
    KeyWire_0_22,
    n1245,
    n1701,
    n1222,
    n1211
  );


  nand
  g1767
  (
    n2084,
    n1231,
    n1744,
    n1719,
    n865
  );


  and
  g1768
  (
    n2317,
    n1347,
    n807,
    n1653,
    n1673
  );


  xnor
  g1769
  (
    n2169,
    n1062,
    n1270,
    n1333,
    n1747
  );


  or
  g1770
  (
    n2320,
    n1383,
    n883,
    n1678,
    n1167
  );


  xnor
  g1771
  (
    n1935,
    n1063,
    n1690,
    n1204,
    n1550
  );


  nor
  g1772
  (
    n2496,
    n1486,
    n1714,
    n1565,
    n1057
  );


  or
  g1773
  (
    n2260,
    n1577,
    n1713,
    n1680,
    n1133
  );


  xor
  g1774
  (
    n2501,
    n1323,
    n1155,
    n943,
    n989
  );


  xnor
  g1775
  (
    n2149,
    n1720,
    n1527,
    n1309,
    n1459
  );


  nand
  g1776
  (
    n2228,
    n905,
    n1073,
    n1286,
    n1170
  );


  or
  g1777
  (
    n2670,
    n1328,
    n941,
    n1658,
    n932
  );


  and
  g1778
  (
    n2599,
    n1244,
    n1529,
    n920,
    n1088
  );


  or
  g1779
  (
    n2646,
    n1005,
    n1251,
    n1502,
    n1129
  );


  xor
  g1780
  (
    n2549,
    n994,
    n1490,
    n1465,
    n1181
  );


  nor
  g1781
  (
    n2286,
    n1658,
    n1495,
    n1202,
    n923
  );


  nand
  g1782
  (
    n2583,
    n1002,
    n1625,
    n1714,
    n1260
  );


  xor
  g1783
  (
    n2372,
    n1050,
    n1384,
    n1614,
    n1037
  );


  nor
  g1784
  (
    n2078,
    n1602,
    n1514,
    n1699,
    n963
  );


  nor
  g1785
  (
    n2427,
    n1238,
    n1679,
    n1288,
    n1505
  );


  or
  g1786
  (
    n2299,
    n1290,
    n1244,
    n954,
    n1589
  );


  xnor
  g1787
  (
    n1997,
    n1552,
    n1120,
    n1015,
    n896
  );


  nor
  g1788
  (
    n1859,
    n1361,
    n840,
    n1337,
    n1209
  );


  nand
  g1789
  (
    n2576,
    n1512,
    n1271,
    n1111,
    n1632
  );


  nand
  g1790
  (
    n2069,
    n1094,
    n1321,
    n1395,
    n1752
  );


  xor
  g1791
  (
    n2234,
    n1427,
    n1289,
    n1080,
    n1000
  );


  nor
  g1792
  (
    n2147,
    n1202,
    n1236,
    n1031,
    n1382
  );


  and
  g1793
  (
    n1894,
    n1555,
    n1063,
    n1077,
    n1656
  );


  or
  g1794
  (
    n1929,
    n1690,
    n1622,
    n1530,
    n1051
  );


  nand
  g1795
  (
    n2582,
    n1103,
    n1500,
    n1431,
    n1377
  );


  xor
  g1796
  (
    n1811,
    n1108,
    n1621,
    n1279,
    n1022
  );


  xor
  g1797
  (
    n2649,
    n1103,
    n1742,
    n1404,
    n1028
  );


  or
  g1798
  (
    n1959,
    n1021,
    n1357,
    n1374,
    n1249
  );


  xor
  g1799
  (
    n2213,
    n1435,
    n1483,
    n1688,
    n1468
  );


  nand
  g1800
  (
    n2021,
    n996,
    n1247,
    n1143,
    n1684
  );


  nor
  g1801
  (
    n2537,
    n1548,
    n1729,
    n1247,
    n1522
  );


  nor
  g1802
  (
    n2581,
    n1726,
    n892,
    n1015,
    n895
  );


  nor
  g1803
  (
    n2271,
    n1205,
    n1480,
    n1588,
    n1027
  );


  and
  g1804
  (
    n2418,
    n1542,
    n1744,
    n1295,
    n944
  );


  and
  g1805
  (
    n1854,
    n1238,
    n1560,
    n1703,
    n1325
  );


  nor
  g1806
  (
    n2435,
    n1285,
    n981,
    n1062,
    n1143
  );


  xor
  g1807
  (
    n2156,
    n1104,
    n1294,
    n1543,
    n1753
  );


  xor
  g1808
  (
    n2193,
    n1660,
    n1072,
    n1199,
    n894
  );


  nor
  g1809
  (
    n2010,
    n1460,
    n1184,
    n1046,
    n1749
  );


  xnor
  g1810
  (
    n2277,
    n1526,
    n1304,
    n890,
    n1468
  );


  xnor
  g1811
  (
    n2422,
    n1069,
    n1631,
    n1350,
    n1097
  );


  xnor
  g1812
  (
    n2065,
    n1325,
    n1461,
    n1064,
    n1430
  );


  nor
  g1813
  (
    n2158,
    n1162,
    n1189,
    n1242,
    n1260
  );


  and
  g1814
  (
    KeyWire_0_23,
    n1142,
    n1396,
    n1444,
    n1510
  );


  xor
  g1815
  (
    n2465,
    n1438,
    n1205,
    n1710,
    n1098
  );


  nor
  g1816
  (
    n1934,
    n1710,
    n1228,
    n1531,
    n1379
  );


  nor
  g1817
  (
    n1796,
    n1422,
    n1123,
    n810,
    n1302
  );


  and
  g1818
  (
    n2059,
    n1653,
    n1273,
    n1488,
    n1724
  );


  xnor
  g1819
  (
    n1938,
    n1635,
    n1746,
    n1596,
    n1509
  );


  nand
  g1820
  (
    n2070,
    n1492,
    n1263,
    n1597,
    n1529
  );


  and
  g1821
  (
    n2159,
    n1195,
    n1133,
    n1066,
    n1536
  );


  and
  g1822
  (
    n2133,
    n1040,
    n1454,
    n1379,
    n944
  );


  nor
  g1823
  (
    n2248,
    n1099,
    n1475,
    n921,
    n1442
  );


  nor
  g1824
  (
    n2641,
    n1548,
    n939,
    n1172,
    n1451
  );


  nor
  g1825
  (
    n1841,
    n1341,
    n1034,
    n1253,
    n1138
  );


  xor
  g1826
  (
    n1990,
    n1094,
    n1384,
    n1151,
    n1516
  );


  nand
  g1827
  (
    n2520,
    n1653,
    n1480,
    n1682,
    n1401
  );


  nor
  g1828
  (
    n2292,
    n1081,
    n1218,
    n1202,
    n1212
  );


  xnor
  g1829
  (
    n1888,
    n1264,
    n1070,
    n1465,
    n1664
  );


  xor
  g1830
  (
    n1821,
    n1023,
    n1022,
    n934,
    n1097
  );


  or
  g1831
  (
    n2314,
    n1131,
    n1389,
    n1022,
    n1315
  );


  xnor
  g1832
  (
    n2310,
    n1007,
    n1119,
    n1387,
    n1041
  );


  nor
  g1833
  (
    n2526,
    n1319,
    n967,
    n1602,
    n1376
  );


  or
  g1834
  (
    n2593,
    n1448,
    n1384,
    n1317,
    n1194
  );


  nor
  g1835
  (
    n2455,
    n1405,
    n965,
    n1313,
    n1215
  );


  nand
  g1836
  (
    n2144,
    n1438,
    n1749,
    n1071,
    n829
  );


  nor
  g1837
  (
    n2184,
    n1301,
    n1518,
    n979,
    n1382
  );


  and
  g1838
  (
    n2203,
    n1549,
    n1015,
    n1583,
    n1215
  );


  and
  g1839
  (
    n1770,
    n1733,
    n1652,
    n1604,
    n1126
  );


  xnor
  g1840
  (
    n2309,
    n1210,
    n1693,
    n1170,
    n1111
  );


  or
  g1841
  (
    n1874,
    n1210,
    n1231,
    n1473,
    n953
  );


  xnor
  g1842
  (
    n2060,
    n1295,
    n1639,
    n1204,
    n968
  );


  xor
  g1843
  (
    n2528,
    n968,
    n914,
    n1657,
    n1755
  );


  and
  g1844
  (
    n2420,
    n1372,
    n1371,
    n1287,
    n1465
  );


  xor
  g1845
  (
    n1940,
    n1363,
    n1013,
    n1177,
    n815
  );


  xnor
  g1846
  (
    n2196,
    n1360,
    n967,
    n1440,
    n1147
  );


  nand
  g1847
  (
    n2218,
    n1368,
    n1618,
    n1201,
    n1127
  );


  nand
  g1848
  (
    n2665,
    n975,
    n1254,
    n804,
    n1193
  );


  nand
  g1849
  (
    n2466,
    n1697,
    n1128,
    n1138,
    n1497
  );


  and
  g1850
  (
    n1810,
    n1751,
    n1183,
    n945,
    n1734
  );


  xor
  g1851
  (
    n2326,
    n1671,
    n1079,
    n882,
    n1286
  );


  and
  g1852
  (
    n1819,
    n876,
    n942,
    n1476,
    n1753
  );


  xor
  g1853
  (
    n2062,
    n1003,
    n1118,
    n1724,
    n1719
  );


  xor
  g1854
  (
    n1917,
    n903,
    n1326,
    n1048,
    n1107
  );


  and
  g1855
  (
    n2663,
    n1505,
    n1219,
    n965,
    n1030
  );


  or
  g1856
  (
    n2131,
    n887,
    n1607,
    n1216,
    n1440
  );


  xor
  g1857
  (
    n2616,
    n1675,
    n969,
    n1736,
    n1666
  );


  xor
  g1858
  (
    n2514,
    n1268,
    n1226,
    n1242,
    n1527
  );


  xnor
  g1859
  (
    n2383,
    n1713,
    n1100,
    n1346,
    n1332
  );


  nand
  g1860
  (
    n1769,
    n1222,
    n1535,
    n1088,
    n1105
  );


  or
  g1861
  (
    n1870,
    n1204,
    n1069,
    n1347,
    n1542
  );


  and
  g1862
  (
    n2072,
    n1187,
    n1398,
    n1660,
    n1433
  );


  xor
  g1863
  (
    n2227,
    n1700,
    n1104,
    n1105,
    n1337
  );


  nor
  g1864
  (
    n1999,
    n1284,
    n1071,
    n1504,
    n1018
  );


  or
  g1865
  (
    n2255,
    n1277,
    n1223,
    n915,
    n983
  );


  nand
  g1866
  (
    n2046,
    n1108,
    n1051,
    n810,
    n1079
  );


  nor
  g1867
  (
    n2483,
    n1130,
    n1299,
    n1119
  );


  nand
  g1868
  (
    n2369,
    n1559,
    n863,
    n1697,
    n1363
  );


  xor
  g1869
  (
    n2297,
    n1425,
    n1294,
    n1099,
    n1034
  );


  xnor
  g1870
  (
    n2175,
    n898,
    n1759,
    n1093,
    n1178
  );


  xnor
  g1871
  (
    n2305,
    n1526,
    n1064,
    n1714,
    n1221
  );


  nor
  g1872
  (
    n2385,
    n1489,
    n973,
    n1035,
    n822
  );


  xnor
  g1873
  (
    n2273,
    n927,
    n1516,
    n1512,
    n1691
  );


  or
  g1874
  (
    n2351,
    n1088,
    n1704,
    n917,
    n955
  );


  and
  g1875
  (
    n2198,
    n1059,
    n975,
    n1729,
    n1394
  );


  nor
  g1876
  (
    n2128,
    n1343,
    n1618,
    n1095,
    n1579
  );


  or
  g1877
  (
    n2524,
    n985,
    n1171,
    n1717,
    n1459
  );


  xor
  g1878
  (
    n1961,
    n1145,
    n1339,
    n1076,
    n1025
  );


  nor
  g1879
  (
    n2453,
    n1067,
    n1636,
    n1525,
    n1578
  );


  nand
  g1880
  (
    n2428,
    n1280,
    n1261,
    n1427,
    n1594
  );


  xnor
  g1881
  (
    n1979,
    n903,
    n1372,
    n1600,
    n959
  );


  nor
  g1882
  (
    n2347,
    n1266,
    n1433,
    n1434,
    n1073
  );


  and
  g1883
  (
    n2590,
    n1088,
    n1070,
    n1184,
    n1225
  );


  nand
  g1884
  (
    n2034,
    n1488,
    n934,
    n1319,
    n1403
  );


  or
  g1885
  (
    n1818,
    n1095,
    n1098,
    n1252,
    n923
  );


  xnor
  g1886
  (
    n1943,
    n1689,
    n1322,
    n1375,
    n1334
  );


  or
  g1887
  (
    n2470,
    n1311,
    n1662,
    n874,
    n1603
  );


  xor
  g1888
  (
    KeyWire_0_4,
    n1288,
    n1516,
    n1057,
    n1730
  );


  xor
  g1889
  (
    n2283,
    n1180,
    n1020,
    n1128,
    n1460
  );


  or
  g1890
  (
    n2058,
    n1554,
    n1568,
    n1380,
    n1258
  );


  or
  g1891
  (
    n2628,
    n1152,
    n899,
    n1753,
    n1348
  );


  or
  g1892
  (
    n1960,
    n1237,
    n1220,
    n1683,
    n1199
  );


  xnor
  g1893
  (
    n2000,
    n1067,
    n1567,
    n1687,
    n899
  );


  or
  g1894
  (
    n2637,
    n1744,
    n1144,
    n1596,
    n1226
  );


  and
  g1895
  (
    n1989,
    n808,
    n1142,
    n1182,
    n939
  );


  nand
  g1896
  (
    n2197,
    n993,
    n1424,
    n1641,
    n994
  );


  or
  g1897
  (
    n1987,
    n1733,
    n1120,
    n1174,
    n1350
  );


  nor
  g1898
  (
    n2190,
    n1212,
    n1023,
    n948,
    n1274
  );


  xor
  g1899
  (
    n1861,
    n1616,
    n981,
    n1227,
    n1193
  );


  or
  g1900
  (
    n2632,
    n1318,
    n1586,
    n1718,
    n1640
  );


  nand
  g1901
  (
    n2306,
    n977,
    n1711,
    n1736,
    n1012
  );


  xor
  g1902
  (
    n2368,
    n1369,
    n1292,
    n1419,
    n1055
  );


  xor
  g1903
  (
    n1918,
    n1432,
    n1635,
    n923,
    n1551
  );


  nor
  g1904
  (
    n2536,
    n1364,
    n1113,
    n1239,
    n1241
  );


  xor
  g1905
  (
    n1942,
    n997,
    n1682,
    n963,
    n1022
  );


  xor
  g1906
  (
    n2236,
    n1296,
    n1336,
    n841,
    n1084
  );


  nand
  g1907
  (
    n2244,
    n1399,
    n1094,
    n1453,
    n1253
  );


  nand
  g1908
  (
    n2071,
    n910,
    n1515,
    n867,
    n1236
  );


  nor
  g1909
  (
    n2199,
    n1715,
    n1334,
    n1701,
    n1219
  );


  and
  g1910
  (
    n2497,
    n1033,
    n915,
    n849,
    n1208
  );


  and
  g1911
  (
    n2030,
    n1214,
    n1128,
    n1217,
    n1340
  );


  xor
  g1912
  (
    n2519,
    n877,
    n1200,
    n1421,
    n1308
  );


  xnor
  g1913
  (
    n2357,
    n1485,
    n1113,
    n1314,
    n1165
  );


  xor
  g1914
  (
    n2460,
    n1010,
    n1208,
    n1260,
    n1230
  );


  and
  g1915
  (
    n2636,
    n1748,
    n948,
    n947,
    n1534
  );


  xnor
  g1916
  (
    n2507,
    n1031,
    n1716,
    n1437,
    n1710
  );


  xor
  g1917
  (
    n2316,
    n955,
    n958,
    n1259,
    n1148
  );


  and
  g1918
  (
    n2423,
    n1581,
    n1074,
    n1644,
    n816
  );


  xor
  g1919
  (
    n2250,
    n1046,
    n1693,
    n955,
    n1032
  );


  and
  g1920
  (
    n2402,
    n1149,
    n1624,
    n1075,
    n850
  );


  nor
  g1921
  (
    n2346,
    n869,
    n1036,
    n1517,
    n989
  );


  nor
  g1922
  (
    n2096,
    n1006,
    n945,
    n1266,
    n1649
  );


  xnor
  g1923
  (
    n1949,
    n1074,
    n896,
    n1607,
    n1121
  );


  nor
  g1924
  (
    n1970,
    n1052,
    n1634,
    n1584,
    n1126
  );


  xnor
  g1925
  (
    n2285,
    n1038,
    n1390,
    n869,
    n1117
  );


  nand
  g1926
  (
    n2480,
    n1165,
    n1304,
    n1352,
    n1391
  );


  xnor
  g1927
  (
    n1795,
    n1738,
    n1447,
    n1332,
    n1533
  );


  and
  g1928
  (
    n2038,
    n1367,
    n970,
    n996,
    n960
  );


  nor
  g1929
  (
    n2268,
    n1701,
    n1591,
    n1462,
    n1614
  );


  nand
  g1930
  (
    n2542,
    n1135,
    n1213,
    n1584,
    n906
  );


  nor
  g1931
  (
    n2404,
    n1615,
    n1756,
    n978,
    n1341
  );


  or
  g1932
  (
    n2444,
    n895,
    n1051,
    n1407,
    n1740
  );


  xnor
  g1933
  (
    n2565,
    n1562,
    n897,
    n838,
    n1711
  );


  xor
  g1934
  (
    n1972,
    n1090,
    n1670,
    n1188,
    n965
  );


  and
  g1935
  (
    n2490,
    n1585,
    n1494,
    n1720,
    n1555
  );


  or
  g1936
  (
    n2493,
    n1734,
    n946,
    n1195,
    n1349
  );


  xor
  g1937
  (
    n1909,
    n1453,
    n1151,
    n1628,
    n1208
  );


  nand
  g1938
  (
    n1830,
    n1584,
    n1122,
    n913,
    n1200
  );


  nand
  g1939
  (
    n2559,
    n843,
    n1505,
    n979,
    n817
  );


  and
  g1940
  (
    n2525,
    n1305,
    n1496,
    n1054,
    n1472
  );


  xnor
  g1941
  (
    n2267,
    n1702,
    n1074,
    n1025,
    n966
  );


  nand
  g1942
  (
    n1948,
    n973,
    n1648,
    n1398,
    n1667
  );


  nor
  g1943
  (
    n1893,
    n1026,
    n1147,
    n1157,
    n1131
  );


  and
  g1944
  (
    n2367,
    n1441,
    n1118,
    n1207,
    n907
  );


  nand
  g1945
  (
    n1809,
    n1180,
    n1739,
    n1209,
    n884
  );


  and
  g1946
  (
    n2382,
    n1506,
    n961,
    n1252,
    n977
  );


  or
  g1947
  (
    n1869,
    n1293,
    n1350,
    n1626,
    n1641
  );


  nand
  g1948
  (
    n2187,
    n1608,
    n1326,
    n1539,
    n1214
  );


  xor
  g1949
  (
    n2074,
    n951,
    n1068,
    n1371,
    n1577
  );


  nand
  g1950
  (
    n2415,
    n1671,
    n1083,
    n902,
    n1497
  );


  xor
  g1951
  (
    n2249,
    n1325,
    n1587,
    n1002,
    n821
  );


  nand
  g1952
  (
    n2613,
    n1165,
    n1048,
    n1392,
    n1706
  );


  xor
  g1953
  (
    n2660,
    n1050,
    n1117,
    n812,
    n1053
  );


  nor
  g1954
  (
    n1858,
    n907,
    n1737,
    n1188,
    n922
  );


  and
  g1955
  (
    n2139,
    n1297,
    n891,
    n940,
    n1625
  );


  xnor
  g1956
  (
    n1885,
    n1700,
    n1082,
    n1406,
    n1092
  );


  xor
  g1957
  (
    n1879,
    n1756,
    n1517,
    n1487,
    n835
  );


  xnor
  g1958
  (
    n2153,
    n952,
    n1445,
    n1308,
    n1614
  );


  xnor
  g1959
  (
    n1906,
    n1322,
    n1445,
    n1499,
    n1154
  );


  nor
  g1960
  (
    n2162,
    n1259,
    n1722,
    n1171,
    n1637
  );


  xor
  g1961
  (
    n2171,
    n1019,
    n1736,
    n1106,
    n1110
  );


  and
  g1962
  (
    n2028,
    n927,
    n1320,
    n1310,
    n1513
  );


  nand
  g1963
  (
    n2603,
    n1255,
    n1481,
    n1103,
    n1561
  );


  xnor
  g1964
  (
    n2242,
    n1595,
    n1087,
    n905,
    n1233
  );


  xor
  g1965
  (
    n1787,
    n1149,
    n1574,
    n1584,
    n1651
  );


  xnor
  g1966
  (
    n2093,
    n1272,
    n1471,
    n1757,
    n1311
  );


  xnor
  g1967
  (
    n2430,
    n824,
    n1126,
    n1390,
    n1254
  );


  or
  g1968
  (
    n2443,
    n1276,
    n1082,
    n1729,
    n1208
  );


  or
  g1969
  (
    n2361,
    n926,
    n987,
    n1443,
    n1158
  );


  nor
  g1970
  (
    n1848,
    n1409,
    n1257,
    n1236,
    n1151
  );


  nand
  g1971
  (
    n2553,
    n1753,
    n1039,
    n1168,
    n1725
  );


  xor
  g1972
  (
    n1814,
    n953,
    n1363,
    n1029,
    n1071
  );


  xor
  g1973
  (
    n2125,
    n1716,
    n1472,
    n1039,
    n1230
  );


  and
  g1974
  (
    n1844,
    n1364,
    n1581,
    n1689,
    n1115
  );


  and
  g1975
  (
    n2291,
    n1038,
    n1650,
    n1449,
    n903
  );


  xnor
  g1976
  (
    n2630,
    n1265,
    n901,
    n1634,
    n1030
  );


  xnor
  g1977
  (
    n2655,
    n1403,
    n1752,
    n1409,
    n1508
  );


  xnor
  g1978
  (
    n2598,
    n1550,
    n1036,
    n1549,
    n1597
  );


  nand
  g1979
  (
    n2226,
    n1494,
    n1739,
    n1454,
    n1712
  );


  nor
  g1980
  (
    n2138,
    n1562,
    n1476,
    n1295,
    n1719
  );


  xnor
  g1981
  (
    n2329,
    n835,
    n1667,
    n1652,
    n1636
  );


  nand
  g1982
  (
    n2323,
    n888,
    n1524,
    n1232,
    n933
  );


  xnor
  g1983
  (
    n2202,
    n911,
    n1058,
    n961,
    n1318
  );


  or
  g1984
  (
    n2106,
    n1355,
    n847,
    n1045,
    n806
  );


  and
  g1985
  (
    n2055,
    n921,
    n1401,
    n1648,
    n990
  );


  xor
  g1986
  (
    n1838,
    n1239,
    n1285,
    n1122,
    n1469
  );


  and
  g1987
  (
    n2080,
    n1598,
    n1037,
    n1268,
    n1705
  );


  and
  g1988
  (
    n1971,
    n1449,
    n1099,
    n1006,
    n1447
  );


  xnor
  g1989
  (
    n2403,
    n1055,
    n1333,
    n1487,
    n1166
  );


  xor
  g1990
  (
    n2011,
    n822,
    n1245,
    n1044,
    n1272
  );


  or
  g1991
  (
    n2573,
    n1535,
    n1600,
    n1435,
    n1035
  );


  xnor
  g1992
  (
    n1789,
    n1420,
    n1185,
    n976,
    n1706
  );


  or
  g1993
  (
    n2068,
    n1455,
    n904,
    n934,
    n957
  );


  nand
  g1994
  (
    n2451,
    n951,
    n1402,
    n1021,
    n966
  );


  and
  g1995
  (
    n2494,
    n1728,
    n1159,
    n1651,
    n1345
  );


  nand
  g1996
  (
    n2185,
    n1489,
    n1665,
    n1240,
    n1219
  );


  and
  g1997
  (
    n2315,
    n1353,
    n954,
    n1426,
    n1405
  );


  and
  g1998
  (
    n2167,
    n962,
    n956,
    n1659,
    n951
  );


  xor
  g1999
  (
    n2384,
    n1130,
    n1459,
    n901,
    n1219
  );


  nand
  g2000
  (
    n2041,
    n1595,
    n1380,
    n1407,
    n1046
  );


  xor
  g2001
  (
    n2391,
    n998,
    n1482,
    n898,
    n936
  );


  or
  g2002
  (
    n2166,
    n1386,
    n1538,
    n911,
    n1566
  );


  and
  g2003
  (
    n1820,
    n1000,
    n1383,
    n988,
    n1371
  );


  xnor
  g2004
  (
    n2092,
    n1747,
    n892,
    n1400,
    n1057
  );


  xor
  g2005
  (
    n1919,
    n956,
    n1513,
    n1551,
    n1339
  );


  xnor
  g2006
  (
    n2469,
    n1228,
    n1477,
    n1250
  );


  nor
  g2007
  (
    n1922,
    n1541,
    n1720,
    n1750,
    n1620
  );


  or
  g2008
  (
    n2364,
    n1489,
    n898,
    n904,
    n955
  );


  nand
  g2009
  (
    n2298,
    n1712,
    n952,
    n1115,
    n827
  );


  nand
  g2010
  (
    n2371,
    n1470,
    n1506,
    n1049,
    n951
  );


  or
  g2011
  (
    n2332,
    n1269,
    n1563,
    n1561,
    n1450
  );


  xnor
  g2012
  (
    n2529,
    n1133,
    n1606,
    n1012,
    n1406
  );


  and
  g2013
  (
    n2491,
    n1672,
    n1378,
    n1434,
    n1568
  );


  nand
  g2014
  (
    n2296,
    n1031,
    n1276,
    n1237,
    n1754
  );


  nor
  g2015
  (
    n2023,
    n1140,
    n1361,
    n1385,
    n1423
  );


  nand
  g2016
  (
    n1957,
    n936,
    n1443,
    n1642,
    n1065
  );


  xor
  g2017
  (
    n2447,
    n1263,
    n1682,
    n902,
    n1742
  );


  and
  g2018
  (
    n2132,
    n897,
    n1482,
    n932,
    n1127
  );


  xor
  g2019
  (
    n1864,
    n1743,
    n1717,
    n1675,
    n1469
  );


  nor
  g2020
  (
    KeyWire_0_16,
    n1606,
    n1435,
    n1247,
    n1016
  );


  nand
  g2021
  (
    n2508,
    n1042,
    n924,
    n1532,
    n1093
  );


  nand
  g2022
  (
    n2066,
    n1109,
    n1124,
    n1698,
    n1674
  );


  or
  g2023
  (
    n2280,
    n1077,
    n1633,
    n1117,
    n1721
  );


  nor
  g2024
  (
    n1825,
    n1144,
    n1522,
    n1602,
    n1159
  );


  nand
  g2025
  (
    n1761,
    n1515,
    n1506,
    n1462,
    n1498
  );


  nand
  g2026
  (
    n2449,
    n1479,
    n847,
    n1419,
    n1617
  );


  xor
  g2027
  (
    n2568,
    n1606,
    n1316,
    n1153,
    n1659
  );


  and
  g2028
  (
    n2115,
    n1113,
    n1374,
    n1120,
    n906
  );


  or
  g2029
  (
    n2281,
    n1604,
    n1598,
    n1541,
    n933
  );


  xnor
  g2030
  (
    n2584,
    n1093,
    n1650,
    n1586,
    n1500
  );


  nand
  g2031
  (
    n2394,
    n1688,
    n1667,
    n1093,
    n1048
  );


  xnor
  g2032
  (
    n2043,
    n928,
    n1280,
    n1518,
    n1395
  );


  nand
  g2033
  (
    n2634,
    n1601,
    n1061,
    n1418,
    n1007
  );


  and
  g2034
  (
    n1833,
    n1627,
    n1663,
    n1579,
    n1398
  );


  xor
  g2035
  (
    n2624,
    n1337,
    n830,
    n1281,
    n986
  );


  and
  g2036
  (
    n2275,
    n857,
    n1145,
    n1714,
    n1631
  );


  nand
  g2037
  (
    n2201,
    n1145,
    n970,
    n928,
    n1248
  );


  nand
  g2038
  (
    n2212,
    n1256,
    n1135,
    n1429,
    n1554
  );


  nand
  g2039
  (
    n2318,
    n1432,
    n1190,
    n1396,
    n1665
  );


  nor
  g2040
  (
    n1903,
    n971,
    n1746,
    n1365,
    n966
  );


  xnor
  g2041
  (
    n2256,
    n1556,
    n1545,
    n1752,
    n1635
  );


  nand
  g2042
  (
    n2589,
    n861,
    n967,
    n1415,
    n1409
  );


  or
  g2043
  (
    n2631,
    n1451,
    n1471,
    n1056,
    n816
  );


  xnor
  g2044
  (
    n2073,
    n1521,
    n1564,
    n959,
    n1687
  );


  and
  g2045
  (
    n2379,
    n1293,
    n1191,
    n1539,
    n1538
  );


  or
  g2046
  (
    n1932,
    n939,
    n1704,
    n1258,
    n919
  );


  or
  g2047
  (
    n1851,
    n1109,
    n1661,
    n1541,
    n837
  );


  xor
  g2048
  (
    n2473,
    n1046,
    n1284,
    n1129,
    n1383
  );


  nor
  g2049
  (
    n2586,
    n999,
    n1490,
    n860,
    n1167
  );


  xor
  g2050
  (
    n2206,
    n1646,
    n1052,
    n845,
    n1198
  );


  or
  g2051
  (
    n2219,
    n1227,
    n885,
    n891,
    n1256
  );


  xor
  g2052
  (
    n2407,
    n1250,
    n1224,
    n1671,
    n1492
  );


  xnor
  g2053
  (
    n2548,
    n1643,
    n1367,
    n1445,
    n1453
  );


  nor
  g2054
  (
    n2173,
    n1053,
    n1452,
    n1543,
    n1256
  );


  and
  g2055
  (
    n1797,
    n1060,
    n1316,
    n1418,
    n1399
  );


  and
  g2056
  (
    n2145,
    n1187,
    n1595,
    n1739,
    n1014
  );


  and
  g2057
  (
    n2122,
    n1356,
    n1608,
    n1230,
    n1073
  );


  nor
  g2058
  (
    n2342,
    n1664,
    n1388,
    n1583,
    n1318
  );


  xnor
  g2059
  (
    n2554,
    n885,
    n1243,
    n1054,
    n964
  );


  nand
  g2060
  (
    n2014,
    n1050,
    n1204,
    n1197,
    n1098
  );


  nand
  g2061
  (
    n2179,
    n1060,
    n1127,
    n1577,
    n1169
  );


  or
  g2062
  (
    n2373,
    n1125,
    n852,
    n1024,
    n1084
  );


  nand
  g2063
  (
    n2178,
    n1678,
    n1602,
    n1586,
    n875
  );


  xnor
  g2064
  (
    n2091,
    n990,
    n1578,
    n1638,
    n1545
  );


  and
  g2065
  (
    n2333,
    n1506,
    n1134,
    n1443,
    n1291
  );


  and
  g2066
  (
    n1780,
    n1101,
    n1274,
    n934,
    n1347
  );


  nor
  g2067
  (
    n2456,
    n1538,
    n1020,
    n1192,
    n1064
  );


  xor
  g2068
  (
    n2002,
    n1428,
    n1317,
    n1166,
    n1757
  );


  xnor
  g2069
  (
    n2359,
    n1493,
    n1303,
    n966,
    n851
  );


  xor
  g2070
  (
    n2355,
    n1331,
    n1684,
    n1726,
    n1145
  );


  nor
  g2071
  (
    n2262,
    n969,
    n1202,
    n963,
    n1537
  );


  xnor
  g2072
  (
    n2653,
    n1228,
    n1568,
    n1588
  );


  nand
  g2073
  (
    n1835,
    n1289,
    n1619,
    n882,
    n1156
  );


  and
  g2074
  (
    n2432,
    n1603,
    n1455,
    n1470,
    n1373
  );


  nor
  g2075
  (
    n2121,
    n989,
    n900,
    n894,
    n1600
  );


  and
  g2076
  (
    n2076,
    n1178,
    n1641,
    n1435,
    n1055
  );


  or
  g2077
  (
    n2245,
    n1326,
    n1338,
    n1221,
    n1375
  );


  and
  g2078
  (
    n2378,
    n1094,
    n1229,
    n1283,
    n1080
  );


  or
  g2079
  (
    n2104,
    n1630,
    n1296,
    n1456,
    n1137
  );


  or
  g2080
  (
    n2547,
    n930,
    n1529,
    n1538,
    n1182
  );


  xnor
  g2081
  (
    n1950,
    n1251,
    n1130,
    n983,
    n1436
  );


  xnor
  g2082
  (
    n2142,
    n1029,
    n1319,
    n805,
    n1641
  );


  xnor
  g2083
  (
    n2054,
    n1514,
    n1751,
    n859,
    n899
  );


  or
  g2084
  (
    n2552,
    n993,
    n1425,
    n1302,
    n1599
  );


  or
  g2085
  (
    n2664,
    n1629,
    n1482,
    n1514,
    n1214
  );


  or
  g2086
  (
    n2087,
    n1648,
    n1284,
    n878,
    n863
  );


  and
  g2087
  (
    n1983,
    n1689,
    n1225,
    n1735,
    n1249
  );


  nand
  g2088
  (
    n2141,
    n1759,
    n1652,
    n1431,
    n1342
  );


  xor
  g2089
  (
    n2176,
    n1366,
    n1032,
    n1155,
    n1398
  );


  xnor
  g2090
  (
    n1930,
    n1091,
    n1003,
    n1617,
    n917
  );


  nor
  g2091
  (
    n2408,
    n1464,
    n1434,
    n1354,
    n1112
  );


  or
  g2092
  (
    n2241,
    n1501,
    n1702,
    n858,
    n1158
  );


  xor
  g2093
  (
    n1955,
    n1016,
    n1312,
    n1687,
    n1637
  );


  nand
  g2094
  (
    n2116,
    n1310,
    n1152,
    n1302,
    n1484
  );


  xnor
  g2095
  (
    n2258,
    n1731,
    n1560,
    n1646,
    n1420
  );


  or
  g2096
  (
    n1828,
    n1152,
    n1073,
    n1675,
    n1299
  );


  or
  g2097
  (
    n1975,
    n1654,
    n1297,
    n1610,
    n1475
  );


  xor
  g2098
  (
    n2414,
    n838,
    n1452,
    n1203,
    n1374
  );


  xnor
  g2099
  (
    n2410,
    n1352,
    n1676,
    n1294,
    n1188
  );


  xnor
  g2100
  (
    n2531,
    n1044,
    n1484,
    n1120,
    n940
  );


  xnor
  g2101
  (
    n2024,
    n1471,
    n1335,
    n1690,
    n1019
  );


  and
  g2102
  (
    n2182,
    n1213,
    n1156,
    n1637,
    n1715
  );


  or
  g2103
  (
    n2591,
    n1531,
    n1650,
    n1748,
    n937
  );


  or
  g2104
  (
    n2401,
    n1237,
    n1518,
    n1179,
    n1091
  );


  xnor
  g2105
  (
    n2381,
    n1672,
    n1116,
    n1596,
    n1028
  );


  or
  g2106
  (
    n1782,
    n1351,
    n1595,
    n1599,
    n1061
  );


  xnor
  g2107
  (
    n2604,
    n1456,
    n1446,
    n887,
    n903
  );


  or
  g2108
  (
    n2579,
    n1674,
    n1010,
    n1265,
    n932
  );


  nand
  g2109
  (
    n1877,
    n1511,
    n998,
    n1751,
    n1330
  );


  xor
  g2110
  (
    n2152,
    n958,
    n906,
    n1163,
    n1152
  );


  nor
  g2111
  (
    n2438,
    n898,
    n1263,
    n1483,
    n1660
  );


  nand
  g2112
  (
    n1964,
    n1743,
    n1560,
    n1021,
    n1751
  );


  nor
  g2113
  (
    n2446,
    n1486,
    n818,
    n871,
    n1279
  );


  nand
  g2114
  (
    n2056,
    n1418,
    n1478,
    n1518,
    n896
  );


  or
  g2115
  (
    n1778,
    n1182,
    n1390,
    n1509,
    n1192
  );


  xnor
  g2116
  (
    n2392,
    n1519,
    n1270,
    n998,
    n1610
  );


  xor
  g2117
  (
    n2431,
    n1138,
    n1743,
    n1075,
    n879
  );


  xor
  g2118
  (
    n2609,
    n916,
    n889,
    n1282,
    n1056
  );


  or
  g2119
  (
    n2192,
    n1429,
    n1328,
    n1297,
    n1023
  );


  and
  g2120
  (
    n2409,
    n1715,
    n1154,
    n1158,
    n1345
  );


  nor
  g2121
  (
    n2658,
    n1496,
    n1127,
    n1207,
    n1351
  );


  xor
  g2122
  (
    n1981,
    n1209,
    n1227,
    n1525,
    n1363
  );


  nor
  g2123
  (
    n2475,
    n1097,
    n1639,
    n856,
    n1694
  );


  and
  g2124
  (
    n1899,
    n1360,
    n988,
    n1649,
    n948
  );


  xnor
  g2125
  (
    n2077,
    n1436,
    n1063,
    n1579,
    n1669
  );


  nand
  g2126
  (
    n2083,
    n930,
    n937,
    n1077,
    n1216
  );


  or
  g2127
  (
    n2160,
    n942,
    n1399,
    n909,
    n1524
  );


  xnor
  g2128
  (
    n1766,
    n1026,
    n1659,
    n1102,
    n1597
  );


  xnor
  g2129
  (
    n1785,
    n1400,
    n947,
    n1340,
    n982
  );


  xor
  g2130
  (
    n2331,
    n825,
    n1083,
    n1058,
    n1442
  );


  and
  g2131
  (
    n2596,
    n984,
    n1662,
    n1175,
    n1282
  );


  and
  g2132
  (
    n2619,
    n1482,
    n1534,
    n1335,
    n1582
  );


  or
  g2133
  (
    n1976,
    n1650,
    n979,
    n1723,
    n1330
  );


  and
  g2134
  (
    n2231,
    n957,
    n1636,
    n1086,
    n1067
  );


  and
  g2135
  (
    n2278,
    n1169,
    n935,
    n1018,
    n910
  );


  nor
  g2136
  (
    n2161,
    n1380,
    n1510,
    n1036,
    n1161
  );


  and
  g2137
  (
    n2585,
    n1523,
    n1065,
    n1569,
    n1253
  );


  or
  g2138
  (
    n2050,
    n1524,
    n849,
    n1110,
    n950
  );


  xnor
  g2139
  (
    n2398,
    n1623,
    n1622,
    n1703,
    n1273
  );


  and
  g2140
  (
    n2421,
    n952,
    n954,
    n1489,
    n978
  );


  and
  g2141
  (
    n1973,
    n1015,
    n1354,
    n1222,
    n1373
  );


  nor
  g2142
  (
    n2594,
    n911,
    n1150,
    n964,
    n1708
  );


  or
  g2143
  (
    n1985,
    n1163,
    n1405,
    n1741,
    n1071
  );


  nand
  g2144
  (
    n2321,
    n1528,
    n1042,
    n1039,
    n1685
  );


  and
  g2145
  (
    n1837,
    n1362,
    n1626,
    n941,
    n1529
  );


  xnor
  g2146
  (
    n2433,
    n1169,
    n905,
    n1141,
    n990
  );


  nand
  g2147
  (
    n2123,
    n1522,
    n1609,
    n917,
    n912
  );


  nand
  g2148
  (
    n1896,
    n1000,
    n1646,
    n1043,
    n1267
  );


  nand
  g2149
  (
    n2354,
    n1159,
    n1680,
    n920,
    n1623
  );


  and
  g2150
  (
    n2163,
    n1573,
    n1570,
    n1733,
    n1004
  );


  xor
  g2151
  (
    n1897,
    n1422,
    n1553,
    n867,
    n1558
  );


  xnor
  g2152
  (
    n1808,
    n1439,
    n1369,
    n1308,
    n909
  );


  xor
  g2153
  (
    n2288,
    n1192,
    n18,
    n1201,
    n1357
  );


  and
  g2154
  (
    n2180,
    n1661,
    n1106,
    n899,
    n1686
  );


  nand
  g2155
  (
    n1857,
    n870,
    n922,
    n807,
    n1336
  );


  nand
  g2156
  (
    n2643,
    n1345,
    n1704,
    n1503,
    n1245
  );


  and
  g2157
  (
    n2602,
    n994,
    n1176,
    n1191,
    n992
  );


  xnor
  g2158
  (
    n2265,
    n1140,
    n1087,
    n1619,
    n1024
  );


  nor
  g2159
  (
    n1846,
    n1739,
    n1580,
    n1433,
    n1157
  );


  and
  g2160
  (
    n2308,
    n1197,
    n1624,
    n1006,
    n1634
  );


  xnor
  g2161
  (
    n2541,
    n1459,
    n1686,
    n1559,
    n1018
  );


  xor
  g2162
  (
    n2452,
    n1580,
    n1681,
    n881,
    n1067
  );


  xnor
  g2163
  (
    n2137,
    n1375,
    n992,
    n1327,
    n1655
  );


  and
  g2164
  (
    n1760,
    n1298,
    n868,
    n1685,
    n1658
  );


  nand
  g2165
  (
    n2340,
    n1254,
    n1040,
    n1329,
    n1241
  );


  nand
  g2166
  (
    n1876,
    n1261,
    n1044,
    n1220,
    n1246
  );


  nand
  g2167
  (
    n2090,
    n1386,
    n1365,
    n1395,
    n1164
  );


  nand
  g2168
  (
    n2345,
    n1162,
    n1096,
    n949,
    n1414
  );


  xnor
  g2169
  (
    n2022,
    n1255,
    n824,
    n921,
    n1394
  );


  nor
  g2170
  (
    n2289,
    n1214,
    n1083,
    n962,
    n901
  );


  or
  g2171
  (
    n1882,
    n1301,
    n912,
    n1394,
    n989
  );


  xor
  g2172
  (
    n2257,
    n1217,
    n1356,
    n1519,
    n1134
  );


  nand
  g2173
  (
    n2484,
    n1629,
    n806,
    n969,
    n1402
  );


  nand
  g2174
  (
    n2437,
    n1508,
    n1053,
    n1608,
    n1456
  );


  xnor
  g2175
  (
    n2532,
    n938,
    n1242,
    n1147,
    n1140
  );


  nor
  g2176
  (
    n2642,
    n1517,
    n1629,
    n1382,
    n1620
  );


  xnor
  g2177
  (
    n2029,
    n812,
    n1644,
    n1582,
    n982
  );


  or
  g2178
  (
    n2031,
    n1199,
    n1077,
    n1102,
    n873
  );


  or
  g2179
  (
    n1798,
    n1221,
    n900,
    n1523,
    n1181
  );


  nor
  g2180
  (
    n1840,
    n894,
    n1337,
    n1464,
    n984
  );


  nand
  g2181
  (
    n2300,
    n1381,
    n1292,
    n893,
    n1255
  );


  and
  g2182
  (
    n2304,
    n1150,
    n1049,
    n1467,
    n997
  );


  or
  g2183
  (
    n1832,
    n1481,
    n1293,
    n1723,
    n1207
  );


  and
  g2184
  (
    n2560,
    n1750,
    n1654,
    n1278,
    n820
  );


  nor
  g2185
  (
    n1777,
    n1748,
    n1136,
    n935,
    n943
  );


  nand
  g2186
  (
    n2210,
    n1469,
    n949,
    n1321,
    n1035
  );


  and
  g2187
  (
    n1947,
    n962,
    n1175,
    n1255,
    n1652
  );


  and
  g2188
  (
    n1920,
    n895,
    n914,
    n1515,
    n1137
  );


  and
  g2189
  (
    n1915,
    n1024,
    n1692,
    n1589,
    n1461
  );


  nor
  g2190
  (
    n2419,
    n1180,
    n1050,
    n1310,
    n1331
  );


  and
  g2191
  (
    n1826,
    n1615,
    n1347,
    n1223,
    n995
  );


  or
  g2192
  (
    n1891,
    n1467,
    n1552,
    n1724,
    n1167
  );


  xor
  g2193
  (
    n2264,
    n1732,
    n1049,
    n1382,
    n1146
  );


  nor
  g2194
  (
    n1816,
    n1373,
    n1017,
    n1007,
    n1218
  );


  nand
  g2195
  (
    n2270,
    n1608,
    n1185,
    n1264,
    n1121
  );


  xnor
  g2196
  (
    n1856,
    n1532,
    n811,
    n1540,
    n1700
  );


  xnor
  g2197
  (
    n2165,
    n1057,
    n1626,
    n1417,
    n1715
  );


  nor
  g2198
  (
    n2656,
    n1121,
    n1406,
    n1525,
    n805
  );


  xor
  g2199
  (
    KeyWire_0_20,
    n1346,
    n1703,
    n1737,
    n1724
  );


  or
  g2200
  (
    n2638,
    n1176,
    n1386,
    n1273,
    n1271
  );


  nand
  g2201
  (
    KeyWire_0_6,
    n1348,
    n1258,
    n1261,
    n1157
  );


  xor
  g2202
  (
    n2110,
    n1668,
    n1333,
    n1223,
    n1311
  );


  xor
  g2203
  (
    n2518,
    n1177,
    n1341,
    n1251,
    n1497
  );


  nand
  g2204
  (
    n2259,
    n1307,
    n1493,
    n1166,
    n1285
  );


  and
  g2205
  (
    n1872,
    n1552,
    n907,
    n1212,
    n1327
  );


  and
  g2206
  (
    n1887,
    n998,
    n1670,
    n1533,
    n931
  );


  xor
  g2207
  (
    n2088,
    n1495,
    n1663,
    n1574,
    n1013
  );


  and
  g2208
  (
    n2319,
    n1365,
    n1721,
    n1475,
    n916
  );


  and
  g2209
  (
    n2416,
    n1436,
    n1286,
    n1098,
    n916
  );


  xnor
  g2210
  (
    n2287,
    n1666,
    n1139,
    n1096,
    n1615
  );


  xnor
  g2211
  (
    n1916,
    n1679,
    n1683,
    n1036,
    n859
  );


  nand
  g2212
  (
    n2558,
    n843,
    n1246,
    n1361,
    n1351
  );


  xnor
  g2213
  (
    n2148,
    n1536,
    n1298,
    n1379,
    n809
  );


  xor
  g2214
  (
    n2672,
    n1461,
    n1061,
    n984,
    n1181
  );


  xor
  g2215
  (
    n2500,
    n1099,
    n1187,
    n1368,
    n935
  );


  or
  g2216
  (
    n2654,
    n963,
    n1655,
    n1480,
    n1226
  );


  nor
  g2217
  (
    n2650,
    n1232,
    n1557,
    n1683,
    n1727
  );


  or
  g2218
  (
    n2506,
    n1228,
    n1085,
    n1483,
    n1173
  );


  xor
  g2219
  (
    n1866,
    n1416,
    n1423,
    n826,
    n1437
  );


  xor
  g2220
  (
    n2151,
    n1557,
    n1566,
    n1612,
    n1112
  );


  nand
  g2221
  (
    n2540,
    n1193,
    n1362,
    n1315,
    n1654
  );


  xor
  g2222
  (
    n2617,
    n990,
    n1373,
    n872,
    n1530
  );


  xnor
  g2223
  (
    n1823,
    n1244,
    n1758,
    n1132,
    n1618
  );


  or
  g2224
  (
    n2105,
    n1598,
    n1655,
    n1679
  );


  xnor
  g2225
  (
    n2223,
    n942,
    n1114,
    n918,
    n840
  );


  or
  g2226
  (
    n1883,
    n1415,
    n1729,
    n1442,
    n1017
  );


  xnor
  g2227
  (
    n2468,
    n938,
    n1291,
    n1338,
    n1580
  );


  and
  g2228
  (
    n1875,
    n1272,
    n1559,
    n1366,
    n1478
  );


  or
  g2229
  (
    n2505,
    n1668,
    n1605,
    n1562,
    n1162
  );


  nor
  g2230
  (
    n2400,
    n1175,
    n988,
    n1409,
    n972
  );


  xor
  g2231
  (
    n1822,
    n1306,
    n1001,
    n1509,
    n1324
  );


  nor
  g2232
  (
    n1827,
    n1596,
    n1043,
    n1590,
    n1234
  );


  xor
  g2233
  (
    n1790,
    n1694,
    n1629,
    n1601,
    n1072
  );


  and
  g2234
  (
    n2035,
    n1424,
    n1111,
    n1593,
    n1656
  );


  xnor
  g2235
  (
    n2562,
    n1192,
    n980,
    n1447,
    n1001
  );


  nand
  g2236
  (
    n2543,
    n1146,
    n1339,
    n1400,
    n919
  );


  xnor
  g2237
  (
    n2215,
    n1573,
    n1183,
    n1252,
    n1496
  );


  or
  g2238
  (
    n2395,
    n1179,
    n985,
    n1486,
    n1662
  );


  xor
  g2239
  (
    n2052,
    n1654,
    n1052,
    n862,
    n991
  );


  nand
  g2240
  (
    n2150,
    n1755,
    n1639,
    n1276,
    n1223
  );


  xor
  g2241
  (
    n2282,
    n1100,
    n1290,
    n1359,
    n1287
  );


  and
  g2242
  (
    n2486,
    n1296,
    n1182,
    n1235,
    n1701
  );


  and
  g2243
  (
    n2515,
    n1323,
    n922,
    n1427,
    n883
  );


  or
  g2244
  (
    n2523,
    n1757,
    n984,
    n931,
    n1452
  );


  nand
  g2245
  (
    n2334,
    n968,
    n1090,
    n980,
    n1217
  );


  xor
  g2246
  (
    n1954,
    n1520,
    n919,
    n1404,
    n1300
  );


  xnor
  g2247
  (
    n2086,
    n897,
    n1583,
    n909,
    n1327
  );


  xnor
  g2248
  (
    n2426,
    n1368,
    n902,
    n1649,
    n967
  );


  or
  g2249
  (
    n1910,
    n1068,
    n1316,
    n908,
    n1593
  );


  and
  g2250
  (
    n1901,
    n1507,
    n1195,
    n1199,
    n1481
  );


  nor
  g2251
  (
    n2017,
    n1640,
    n1020,
    n1079,
    n1559
  );


  and
  g2252
  (
    n2511,
    n1150,
    n1663,
    n974,
    n1218
  );


  or
  g2253
  (
    n2154,
    n1645,
    n957,
    n1496,
    n1479
  );


  xnor
  g2254
  (
    n1803,
    n1422,
    n818,
    n1685,
    n1189
  );


  xnor
  g2255
  (
    n1927,
    n1184,
    n1569,
    n1320,
    n1609
  );


  or
  g2256
  (
    n2472,
    n1735,
    n1643,
    n1452,
    n1631
  );


  nor
  g2257
  (
    n2374,
    n1300,
    n1313,
    n1484,
    n1302
  );


  and
  g2258
  (
    n2313,
    n1375,
    n1623,
    n1575,
    n1427
  );


  xor
  g2259
  (
    n2633,
    n1211,
    n1091,
    n1178,
    n1451
  );


  xor
  g2260
  (
    n2615,
    n1001,
    n1110,
    n1679,
    n1620
  );


  nand
  g2261
  (
    n2434,
    n1254,
    n839,
    n1324,
    n1681
  );


  nor
  g2262
  (
    n1781,
    n1194,
    n1354,
    n1420,
    n950
  );


  nor
  g2263
  (
    n2572,
    n1745,
    n1187,
    n1520,
    n1630
  );


  xnor
  g2264
  (
    n2232,
    n926,
    n1532,
    n1755,
    n1271
  );


  nor
  g2265
  (
    n2387,
    n1696,
    n1560,
    n900,
    n1137
  );


  and
  g2266
  (
    n2183,
    n1262,
    n1466,
    n952,
    n1612
  );


  xor
  g2267
  (
    n1773,
    n1013,
    n1247,
    n1448,
    n1225
  );


  xnor
  g2268
  (
    n2204,
    n1700,
    n1059,
    n1135,
    n1378
  );


  xor
  g2269
  (
    n2295,
    n1042,
    n1172,
    n1256,
    n1196
  );


  xnor
  g2270
  (
    n2393,
    n1186,
    n1008,
    n1179,
    n938
  );


  or
  g2271
  (
    n2360,
    n1215,
    n1160,
    n1358,
    n1136
  );


  nand
  g2272
  (
    n2127,
    n1689,
    n1549,
    n1513,
    n1727
  );


  xor
  g2273
  (
    n2003,
    n1737,
    n1497,
    n1546,
    n1116
  );


  xnor
  g2274
  (
    n1817,
    n846,
    n1511,
    n1667,
    n1712
  );


  nor
  g2275
  (
    n2126,
    n924,
    n982,
    n943,
    n1632
  );


  or
  g2276
  (
    n1812,
    n1001,
    n1168,
    n935,
    n1468
  );


  xor
  g2277
  (
    n1852,
    n1123,
    n853,
    n909,
    n896
  );


  nor
  g2278
  (
    n1993,
    n1234,
    n1633,
    n1416,
    n1684
  );


  xor
  g2279
  (
    n2339,
    n1669,
    n1616,
    n1603,
    n1320
  );


  or
  g2280
  (
    n2377,
    n1438,
    n1387,
    n918,
    n1249
  );


  or
  g2281
  (
    n1868,
    n1526,
    n1264,
    n815,
    n1327
  );


  nand
  g2282
  (
    n2363,
    n1613,
    n1024,
    n917,
    n1095
  );


  nand
  g2283
  (
    n1793,
    n1397,
    n1342,
    n980,
    n1379
  );


  nor
  g2284
  (
    n2477,
    n1151,
    n1186,
    n1474,
    n1030
  );


  nor
  g2285
  (
    n2188,
    n972,
    n866,
    n1441,
    n1300
  );


  or
  g2286
  (
    n2669,
    n1147,
    n832,
    n848,
    n1546
  );


  nand
  g2287
  (
    n1804,
    n833,
    n1322,
    n1600,
    n1611
  );


  xnor
  g2288
  (
    n1839,
    n923,
    n1384,
    n1282,
    n1423
  );


  xor
  g2289
  (
    n2485,
    n1305,
    n1486,
    n1362,
    n925
  );


  nand
  g2290
  (
    n1863,
    n1713,
    n1038,
    n831,
    n1587
  );


  or
  g2291
  (
    n2099,
    n1216,
    n1245,
    n1585,
    n1338
  );


  nand
  g2292
  (
    n2181,
    n1455,
    n1519,
    n1149,
    n1160
  );


  nor
  g2293
  (
    n2425,
    n1579,
    n1249,
    n1565,
    n1735
  );


  or
  g2294
  (
    n2246,
    n1612,
    n1492,
    n1027,
    n1106
  );


  nor
  g2295
  (
    n2009,
    n1349,
    n1387,
    n930,
    n1591
  );


  or
  g2296
  (
    n2545,
    n1507,
    n983,
    n866,
    n1458
  );


  nand
  g2297
  (
    n1924,
    n1588,
    n1321,
    n1011,
    n900
  );


  or
  g2298
  (
    n2303,
    n1547,
    n1371,
    n1264,
    n1325
  );


  xor
  g2299
  (
    n2612,
    n1123,
    n1016,
    n1620,
    n1184
  );


  and
  g2300
  (
    n1992,
    n1599,
    n1197,
    n1695,
    n1297
  );


  xnor
  g2301
  (
    n1849,
    n936,
    n1395,
    n927,
    n1745
  );


  and
  g2302
  (
    n1831,
    n890,
    n1498,
    n1109,
    n960
  );


  xor
  g2303
  (
    n1842,
    n1368,
    n1722,
    n1008,
    n948
  );


  nor
  g2304
  (
    n2330,
    n1003,
    n1279,
    n1089,
    n1105
  );


  and
  g2305
  (
    n2097,
    n1677,
    n1404,
    n1759,
    n1696
  );


  nand
  g2306
  (
    n2492,
    n1229,
    n1580,
    n1721,
    n1575
  );


  xnor
  g2307
  (
    n2623,
    n1447,
    n1011,
    n978,
    n1527
  );


  xnor
  g2308
  (
    n2610,
    n1349,
    n1673,
    n1178,
    n1719
  );


  nor
  g2309
  (
    n2412,
    n1709,
    n1340,
    n1047,
    n1072
  );


  or
  g2310
  (
    n1762,
    n1665,
    n1381,
    n1709,
    n1326
  );


  or
  g2311
  (
    n2495,
    n1317,
    n1642,
    n1491,
    n1171
  );


  and
  g2312
  (
    n1881,
    n1275,
    n1750,
    n1086,
    n1033
  );


  and
  g2313
  (
    n1968,
    n1270,
    n1564,
    n1417,
    n1021
  );


  and
  g2314
  (
    n2109,
    n1338,
    n1712,
    n1569,
    n1677
  );


  xor
  g2315
  (
    n2516,
    n1416,
    n1025,
    n1625,
    n929
  );


  or
  g2316
  (
    n1768,
    n860,
    n1004,
    n1312,
    n1676
  );


  nor
  g2317
  (
    n2279,
    n1420,
    n995,
    n1118,
    n949
  );


  and
  g2318
  (
    n1889,
    n1170,
    n1008,
    n1314,
    n1647
  );


  nor
  g2319
  (
    n2439,
    n1622,
    n1290,
    n1173,
    n921
  );


  or
  g2320
  (
    n2253,
    n834,
    n1265,
    n924,
    n913
  );


  or
  g2321
  (
    n1900,
    n1543,
    n956,
    n1206,
    n960
  );


  or
  g2322
  (
    n1926,
    n873,
    n821,
    n1109,
    n1696
  );


  xor
  g2323
  (
    n2563,
    n1446,
    n1037,
    n1321,
    n839
  );


  nand
  g2324
  (
    n2235,
    n1060,
    n1367,
    n1520,
    n1087
  );


  or
  g2325
  (
    n2557,
    n1726,
    n1426,
    n1540,
    n1463
  );


  nor
  g2326
  (
    n2327,
    n878,
    n1224,
    n1501,
    n940
  );


  xor
  g2327
  (
    KeyWire_0_30,
    n1642,
    n836,
    n1171,
    n1687
  );


  nand
  g2328
  (
    n2608,
    n1068,
    n1259,
    n886,
    n1474
  );


  and
  g2329
  (
    n1772,
    n1546,
    n908,
    n1603,
    n1556
  );


  and
  g2330
  (
    n1878,
    n1191,
    n1502,
    n1193,
    n983
  );


  xor
  g2331
  (
    n2644,
    n1262,
    n1587,
    n1640,
    n1211
  );


  xnor
  g2332
  (
    n2429,
    n1276,
    n1013,
    n1449,
    n1592
  );


  and
  g2333
  (
    n2209,
    n1359,
    n901,
    n1717,
    n1027
  );


  xor
  g2334
  (
    n1953,
    n946,
    n1632,
    n937,
    n1034
  );


  or
  g2335
  (
    n2667,
    n1153,
    n1210,
    n1349,
    n1411
  );


  or
  g2336
  (
    n2301,
    n986,
    n1717,
    n1438,
    n997
  );


  xor
  g2337
  (
    n2200,
    n830,
    n1277,
    n1510,
    n1446
  );


  and
  g2338
  (
    n2567,
    n907,
    n1740,
    n1203,
    n1259
  );


  or
  g2339
  (
    n2611,
    n1613,
    n1408,
    n941,
    n1521
  );


  and
  g2340
  (
    n2580,
    n1638,
    n1059,
    n1388,
    n906
  );


  and
  g2341
  (
    n2049,
    n1353,
    n1702,
    n1703,
    n1578
  );


  nand
  g2342
  (
    n2189,
    n1628,
    n1393,
    n1343,
    n1611
  );


  or
  g2343
  (
    KeyWire_0_3,
    n1190,
    n1020,
    n1335,
    n1756
  );


  nor
  g2344
  (
    n1996,
    n1532,
    n1116,
    n1043,
    n1307
  );


  nor
  g2345
  (
    n1925,
    n1517,
    n1285,
    n1617,
    n1408
  );


  and
  g2346
  (
    n2117,
    n1309,
    n1183,
    n1671,
    n1023
  );


  xnor
  g2347
  (
    n2647,
    n1101,
    n1597,
    n1576,
    n1439
  );


  xor
  g2348
  (
    n2328,
    n1630,
    n1359,
    n1470,
    n1358
  );


  nand
  g2349
  (
    n2335,
    n1418,
    n1440,
    n1494,
    n1316
  );


  xnor
  g2350
  (
    n2622,
    n1392,
    n1466,
    n1472,
    n1244
  );


  xnor
  g2351
  (
    n2551,
    n1439,
    n1656,
    n1177,
    n1179
  );


  and
  g2352
  (
    n2380,
    n1172,
    n857,
    n894,
    n1657
  );


  nor
  g2353
  (
    n2606,
    n1515,
    n1164,
    n1113,
    n1030
  );


  xor
  g2354
  (
    n2499,
    n1504,
    n1200,
    n1750,
    n918
  );


  nand
  g2355
  (
    n2100,
    n1740,
    n1429,
    n1713,
    n1741
  );


  xnor
  g2356
  (
    n2569,
    n1268,
    n1445,
    n1229,
    n1742
  );


  xor
  g2357
  (
    n2146,
    n1407,
    n1010,
    n804,
    n1216
  );


  nand
  g2358
  (
    n2348,
    n1331,
    n1539,
    n1082,
    n1606
  );


  xnor
  g2359
  (
    n1951,
    n1491,
    n905,
    n1664,
    n1444
  );


  or
  g2360
  (
    n2120,
    n1499,
    n1718,
    n1085,
    n959
  );


  nor
  g2361
  (
    n1884,
    n1315,
    n1503,
    n1190,
    n1066
  );


  nor
  g2362
  (
    n2119,
    n1045,
    n1455,
    n1674,
    n1450
  );


  or
  g2363
  (
    n2186,
    n1222,
    n1456,
    n1060,
    n1690
  );


  or
  g2364
  (
    n1767,
    n1180,
    n1734,
    n855,
    n1198
  );


  xor
  g2365
  (
    n2108,
    n931,
    n1234,
    n1399,
    n1466
  );


  xnor
  g2366
  (
    n2645,
    n1312,
    n1005,
    n1271,
    n845
  );


  nand
  g2367
  (
    n1800,
    n897,
    n1194,
    n1212,
    n954
  );


  nor
  g2368
  (
    n1791,
    n1426,
    n1032,
    n1537,
    n1722
  );


  xor
  g2369
  (
    n2388,
    n1066,
    n1133,
    n1747,
    n1386
  );


  nand
  g2370
  (
    n1995,
    n1364,
    n925,
    n1410,
    n1670
  );


  xnor
  g2371
  (
    n2124,
    n1313,
    n1443,
    n1237,
    n1017
  );


  nor
  g2372
  (
    n1765,
    n970,
    n1381,
    n975,
    n1709
  );


  nand
  g2373
  (
    n2103,
    n1161,
    n950,
    n1605,
    n1471
  );


  xor
  g2374
  (
    n2512,
    n1647,
    n1485,
    n1642,
    n1535
  );


  or
  g2375
  (
    n1958,
    n956,
    n1526,
    n1211,
    n1069
  );


  xor
  g2376
  (
    n2503,
    n1709,
    n1230,
    n892,
    n912
  );


  xnor
  g2377
  (
    n2016,
    n1740,
    n1136,
    n1142,
    n1479
  );


  nor
  g2378
  (
    n2261,
    n1546,
    n1604,
    n1454,
    n913
  );


  and
  g2379
  (
    n2436,
    n1365,
    n1055,
    n1003,
    n1591
  );


  nand
  g2380
  (
    n2652,
    n1218,
    n1065,
    n1693,
    n1353
  );


  or
  g2381
  (
    n1862,
    n928,
    n1201,
    n1490,
    n1140
  );


  nor
  g2382
  (
    n2578,
    n1176,
    n1035,
    n1051,
    n1569
  );


  and
  g2383
  (
    n2111,
    n1078,
    n1521,
    n1474,
    n1360
  );


  nand
  g2384
  (
    n1941,
    n1332,
    n1330,
    n846,
    n1311
  );


  xor
  g2385
  (
    n2012,
    n1537,
    n1630,
    n1124,
    n1241
  );


  or
  g2386
  (
    n2048,
    n938,
    n1108,
    n1706,
    n1101
  );


  xor
  g2387
  (
    n2461,
    n1027,
    n1262,
    n1167,
    n1372
  );


  nand
  g2388
  (
    n1786,
    n1076,
    n1647,
    n886,
    n1391
  );


  or
  g2389
  (
    n1911,
    n1132,
    n1002,
    n908,
    n1343
  );


  xnor
  g2390
  (
    n2550,
    n1303,
    n819,
    n1047,
    n1260
  );


  or
  g2391
  (
    n2013,
    n1389,
    n1335,
    n1170,
    n1678
  );


  xor
  g2392
  (
    n2047,
    n1239,
    n1711,
    n1484,
    n1106
  );


  xor
  g2393
  (
    n2094,
    n996,
    n1114,
    n988,
    n1378
  );


  or
  g2394
  (
    n2353,
    n1544,
    n852,
    n841,
    n1004
  );


  xnor
  g2395
  (
    n2448,
    n929,
    n1707,
    n1428,
    n1173
  );


  and
  g2396
  (
    n2129,
    n1657,
    n1010,
    n893,
    n1009
  );


  xnor
  g2397
  (
    n1969,
    n1262,
    n1033,
    n1733,
    n1310
  );


  and
  g2398
  (
    n1873,
    n1540,
    n1473,
    n1033,
    n1553
  );


  nor
  g2399
  (
    n2263,
    n1388,
    n1353,
    n1555,
    n1516
  );


  nand
  g2400
  (
    n2057,
    n1646,
    n1745,
    n1299,
    n925
  );


  nand
  g2401
  (
    n2441,
    n819,
    n1680,
    n1494,
    n1571
  );


  nand
  g2402
  (
    n2370,
    n1631,
    n1696,
    n1350,
    n1677
  );


  nand
  g2403
  (
    n2174,
    n1697,
    n1226,
    n1236,
    n1570
  );


  and
  g2404
  (
    n2564,
    n1257,
    n1695,
    n1081,
    n1628
  );


  nand
  g2405
  (
    n1914,
    n1336,
    n1746,
    n1148,
    n1585
  );


  nor
  g2406
  (
    n2509,
    n1722,
    n1261,
    n1542,
    n912
  );


  xnor
  g2407
  (
    n2214,
    n1061,
    n1288,
    n1488,
    n879
  );


  nand
  g2408
  (
    n2221,
    n889,
    n1275,
    n1188,
    n1758
  );


  xnor
  g2409
  (
    n2312,
    n920,
    n1082,
    n933,
    n1392
  );


  nand
  g2410
  (
    n1855,
    n1070,
    n1421,
    n1669,
    n902
  );


  nand
  g2411
  (
    n2208,
    n968,
    n1277,
    n987,
    n1165
  );


  xnor
  g2412
  (
    n2489,
    n1705,
    n1079,
    n1692,
    n1000
  );


  xor
  g2413
  (
    n1988,
    n1008,
    n1547,
    n1716,
    n1410
  );


  xnor
  g2414
  (
    n1788,
    n1425,
    n1104,
    n1639,
    n1231
  );


  nor
  g2415
  (
    n2533,
    n1571,
    n1725,
    n976,
    n1062
  );


  and
  g2416
  (
    n1886,
    n1662,
    n829,
    n1581,
    n1736
  );


  or
  g2417
  (
    n2004,
    n915,
    n1045,
    n1593,
    n1428
  );


  nor
  g2418
  (
    n1967,
    n1394,
    n1014,
    n1591,
    n858
  );


  and
  g2419
  (
    n2118,
    n1732,
    n1075,
    n1388,
    n925
  );


  nand
  g2420
  (
    n2040,
    n1628,
    n1117,
    n1250,
    n1572
  );


  nor
  g2421
  (
    n2195,
    n957,
    n1519,
    n973,
    n1402
  );


  or
  g2422
  (
    n2535,
    n1153,
    n911,
    n1575,
    n975
  );


  nor
  g2423
  (
    n2413,
    n1493,
    n1444,
    n1056,
    n836
  );


  nand
  g2424
  (
    n2033,
    n1198,
    n1009,
    n1582,
    n1508
  );


  nand
  g2425
  (
    n2626,
    n1448,
    n1430,
    n1243,
    n1758
  );


  xnor
  g2426
  (
    n2390,
    n1348,
    n1674,
    n1111,
    n1632
  );


  or
  g2427
  (
    n2102,
    n1346,
    n853,
    n1754,
    n1570
  );


  and
  g2428
  (
    n2290,
    n1385,
    n1677,
    n1465,
    n1078
  );


  xnor
  g2429
  (
    n1908,
    n958,
    n1168,
    n1403,
    n1275
  );


  or
  g2430
  (
    n2478,
    n1473,
    n1458,
    n1566,
    n1498
  );


  nand
  g2431
  (
    n1775,
    n904,
    n1377,
    n1155,
    n1213
  );


  and
  g2432
  (
    n2026,
    n1664,
    n1105,
    n1411,
    n1318
  );


  nand
  g2433
  (
    n2135,
    n851,
    n1668,
    n1299,
    n1699
  );


  xnor
  g2434
  (
    n1860,
    n1161,
    n1633,
    n1581,
    n946
  );


  or
  g2435
  (
    n2659,
    n1143,
    n1160,
    n1154,
    n1303
  );


  and
  g2436
  (
    n2440,
    n864,
    n1665,
    n1522,
    n1556
  );


  xnor
  g2437
  (
    n2561,
    n1609,
    n1688,
    n1242,
    n1097
  );


  nand
  g2438
  (
    n1928,
    n1457,
    n1369,
    n1206,
    n1037
  );


  xor
  g2439
  (
    n1853,
    n1044,
    n1563,
    n981,
    n1413
  );


  xor
  g2440
  (
    n2464,
    n1054,
    n1062,
    n953,
    n1186
  );


  xnor
  g2441
  (
    n1978,
    n1383,
    n1328,
    n1329,
    n1487
  );


  or
  g2442
  (
    n2293,
    n820,
    n1728,
    n1684,
    n1362
  );


  or
  g2443
  (
    n2063,
    n1412,
    n1693,
    n1355,
    n1458
  );


  and
  g2444
  (
    n2136,
    n1309,
    n949,
    n993,
    n1728
  );


  and
  g2445
  (
    n1952,
    n1511,
    n1645,
    n1479,
    n1657
  );


  xnor
  g2446
  (
    n2269,
    n1041,
    n918,
    n1450,
    n1392
  );


  nor
  g2447
  (
    n2544,
    n1738,
    n1137,
    n1698,
    n910
  );


  nand
  g2448
  (
    n2527,
    n1528,
    n1351,
    n1139,
    n1478
  );


  nor
  g2449
  (
    n2140,
    n1592,
    n1391,
    n1573,
    n1305
  );


  xor
  g2450
  (
    n2454,
    n1433,
    n1536,
    n1676,
    n924
  );


  xnor
  g2451
  (
    n1783,
    n1681,
    n1567,
    n1400,
    n856
  );


  nand
  g2452
  (
    n2459,
    n1348,
    n875,
    n1181,
    n1019
  );


  xnor
  g2453
  (
    n1871,
    n1343,
    n926,
    n1510,
    n1303
  );


  xnor
  g2454
  (
    n1824,
    n1059,
    n1446,
    n1107,
    n880
  );


  and
  g2455
  (
    n2386,
    n1412,
    n1076,
    n1144,
    n1287
  );


  nand
  g2456
  (
    n2164,
    n1539,
    n1749,
    n809,
    n1698
  );


  or
  g2457
  (
    n2620,
    n1185,
    n929,
    n1139,
    n915
  );


  xor
  g2458
  (
    n2272,
    n1460,
    n1678,
    n1458,
    n1278
  );


  xor
  g2459
  (
    n2479,
    n1423,
    n1421,
    n1014,
    n1118
  );


  nor
  g2460
  (
    n2600,
    n1473,
    n1283,
    n1056,
    n1415
  );


  or
  g2461
  (
    n2101,
    n1040,
    n1411,
    n1248,
    n1621
  );


  or
  g2462
  (
    n2025,
    n914,
    n1644,
    n1092,
    n1422
  );


  xor
  g2463
  (
    n2061,
    n1269,
    n1206,
    n991,
    n1238
  );


  and
  g2464
  (
    n2662,
    n1146,
    n1547,
    n1346,
    n1301
  );


  or
  g2465
  (
    n2157,
    n1012,
    n1168,
    n973,
    n913
  );


  and
  g2466
  (
    n2639,
    n1359,
    n1052,
    n1134,
    n1405
  );


  nand
  g2467
  (
    n2463,
    n1554,
    n1624,
    n1698,
    n1416
  );


  and
  g2468
  (
    n1905,
    n1523,
    n877,
    n1437,
    n834
  );


  xnor
  g2469
  (
    n2629,
    n1072,
    n1564,
    n1413
  );


  xnor
  g2470
  (
    n2481,
    n1138,
    n1415,
    n1562,
    n980
  );


  xnor
  g2471
  (
    n2556,
    n1492,
    n1086,
    n1191,
    n1561
  );


  nand
  g2472
  (
    n1834,
    n1265,
    n1070,
    n1174,
    n1322
  );


  and
  g2473
  (
    n2358,
    n1682,
    n1012,
    n1660,
    n1570
  );


  xnor
  g2474
  (
    n2130,
    n1686,
    n1122,
    n1470,
    n987
  );


  nand
  g2475
  (
    n2112,
    n1277,
    n1550,
    n1457,
    n1306
  );


  xnor
  g2476
  (
    n1956,
    n1085,
    n1248,
    n1555,
    n1100
  );


  xor
  g2477
  (
    n2574,
    n1130,
    n1428,
    n1319,
    n974
  );


  nand
  g2478
  (
    n2211,
    n1295,
    n1582,
    n1417,
    n1028
  );


  and
  g2479
  (
    n2081,
    n1417,
    n1616,
    n1196,
    n1533
  );


  xor
  g2480
  (
    n2325,
    n1710,
    n1107,
    n1462,
    n1523
  );


  xnor
  g2481
  (
    n2085,
    n1280,
    n1566,
    n1454,
    n1089
  );


  nor
  g2482
  (
    n1850,
    n1707,
    n1637,
    n1759,
    n871
  );


  nand
  g2483
  (
    n1974,
    n1246,
    n914,
    n884,
    n1086
  );


  nand
  g2484
  (
    n2007,
    n1502,
    n1520,
    n1089,
    n1613
  );


  xor
  g2485
  (
    n2089,
    n1220,
    n1201,
    n1115,
    n1096
  );


  or
  g2486
  (
    n2230,
    n1613,
    n1280,
    n982,
    n1129
  );


  nand
  g2487
  (
    n2240,
    n1389,
    n1314,
    n1692,
    n1488
  );


  nor
  g2488
  (
    n2222,
    n1704,
    n1232,
    n1476,
    n1508
  );


  and
  g2489
  (
    n1843,
    n1571,
    n1317,
    n1278,
    n1263
  );


  or
  g2490
  (
    n1931,
    n862,
    n1594,
    n1661,
    n1401
  );


  or
  g2491
  (
    n2217,
    n1742,
    n971,
    n1253,
    n1220
  );


  or
  g2492
  (
    n2191,
    n1588,
    n999,
    n1019,
    n1673
  );


  or
  g2493
  (
    n2233,
    n1085,
    n1643,
    n1467,
    n1136
  );


  xnor
  g2494
  (
    n1836,
    n1289,
    n1592,
    n1624,
    n1556
  );


  nor
  g2495
  (
    n2488,
    n1702,
    n1334,
    n827,
    n1123
  );


  or
  g2496
  (
    n2376,
    n1509,
    n919,
    n1626,
    n1574
  );


  nor
  g2497
  (
    n1794,
    n868,
    n916,
    n1513,
    n1197
  );


  nor
  g2498
  (
    n2570,
    n1707,
    n1463,
    n1053,
    n1069
  );


  nor
  g2499
  (
    n1904,
    n1688,
    n971,
    n1578,
    n1567
  );


  xor
  g2500
  (
    n2375,
    n1017,
    n1298,
    n1344,
    n1610
  );


  xnor
  g2501
  (
    n2302,
    n981,
    n1288,
    n1457,
    n1250
  );


  and
  g2502
  (
    n2504,
    n1332,
    n1487,
    n1233,
    n1673
  );


  or
  g2503
  (
    n2571,
    n1705,
    n1173,
    n1413,
    n872
  );


  or
  g2504
  (
    n2666,
    n964,
    n1598,
    n1670,
    n1142
  );


  xnor
  g2505
  (
    n2064,
    n1412,
    n1480,
    n1658,
    n1615
  );


  or
  g2506
  (
    n2018,
    n1352,
    n1651,
    n1393,
    n1404
  );


  and
  g2507
  (
    n1965,
    n1692,
    n937,
    n1369,
    n893
  );


  nand
  g2508
  (
    n2482,
    n943,
    n1278,
    n1414,
    n1209
  );


  xor
  g2509
  (
    n2134,
    n1132,
    n1312,
    n1732,
    n1221
  );


  nor
  g2510
  (
    n1946,
    n977,
    n1468,
    n1491,
    n946
  );


  nor
  g2511
  (
    n2039,
    n1576,
    n1287,
    n842,
    n1430
  );


  or
  g2512
  (
    n1984,
    n1032,
    n1625,
    n1091,
    n1490
  );


  nor
  g2513
  (
    n2168,
    n1411,
    n1530,
    n1396,
    n1112
  );


  nand
  g2514
  (
    n1962,
    n1695,
    n1525,
    n1163,
    n1449
  );


  and
  g2515
  (
    n1902,
    n953,
    n1305,
    n1574,
    n1356
  );


  xnor
  g2516
  (
    n1779,
    n1315,
    n970,
    n920,
    n1528
  );


  nand
  g2517
  (
    n2036,
    n1396,
    n1283,
    n1125,
    n1102
  );


  and
  g2518
  (
    n2668,
    n1711,
    n1612,
    n1367,
    n1541
  );


  and
  g2519
  (
    n2307,
    n1649,
    n1029,
    n1676,
    n813
  );


  xor
  g2520
  (
    n1936,
    n1535,
    n1286,
    n1029,
    n1333
  );


  nand
  g2521
  (
    n2001,
    n1672,
    n1114,
    n1007,
    n1329
  );


  and
  g2522
  (
    n2155,
    n999,
    n1472,
    n1450,
    n1586
  );


  nor
  g2523
  (
    n2220,
    n888,
    n1358,
    n1092,
    n1685
  );


  and
  g2524
  (
    n2487,
    n1594,
    n1357,
    n940,
    n1132
  );


  nor
  g2525
  (
    n2618,
    n961,
    n1041,
    n1618,
    n1476
  );


  xnor
  g2526
  (
    n2343,
    n1477,
    n1419,
    n1627,
    n1741
  );


  xnor
  g2527
  (
    n2020,
    n1006,
    n1092,
    n1342,
    n1356
  );


  nand
  g2528
  (
    n2336,
    n855,
    n1756,
    n842,
    n1592
  );


  nand
  g2529
  (
    n2566,
    n1545,
    n850,
    n1126,
    n1441
  );


  xnor
  g2530
  (
    n2457,
    n1370,
    n1122,
    n844,
    n1635
  );


  xor
  g2531
  (
    n2657,
    n1668,
    n1440,
    n861,
    n1474
  );


  nor
  g2532
  (
    n1763,
    n1240,
    n1547,
    n823,
    n1536
  );


  nand
  g2533
  (
    n1994,
    n1754,
    n864,
    n1058,
    n1229
  );


  and
  g2534
  (
    n2082,
    n997,
    n1614,
    n1300,
    n1103
  );


  xor
  g2535
  (
    n2053,
    n1393,
    n1385,
    n1227,
    n1557
  );


  xor
  g2536
  (
    n1764,
    n865,
    n1304,
    n1397,
    n1156
  );


  and
  g2537
  (
    n2546,
    n1590,
    n1387,
    n1558,
    n1647
  );


  or
  g2538
  (
    n2051,
    n1174,
    n1534,
    n1078,
    n1551
  );


  nand
  g2539
  (
    n2224,
    n814,
    n1609,
    n1308,
    n1074
  );


  xor
  g2540
  (
    n1806,
    n1410,
    n978,
    n1413,
    n1485
  );


  and
  g2541
  (
    n2521,
    n1694,
    n1755,
    n1557,
    n1718
  );


  nor
  g2542
  (
    n1829,
    n1548,
    n1397,
    n974,
    n1089
  );


  xnor
  g2543
  (
    n2294,
    n1530,
    n1283,
    n1550,
    n995
  );


  xor
  g2544
  (
    n2362,
    n1355,
    n1500,
    n1102,
    n1190
  );


  nand
  g2545
  (
    n2605,
    n1049,
    n1134,
    n1028,
    n1274
  );


  xnor
  g2546
  (
    n2648,
    n1161,
    n1240,
    n1601,
    n959
  );


  xor
  g2547
  (
    n2037,
    n1309,
    n1744,
    n1169,
    n1320
  );


  and
  g2548
  (
    n1939,
    n1157,
    n1735,
    n1186,
    n1548
  );


  xor
  g2549
  (
    n2352,
    n1306,
    n848,
    n1323,
    n1619
  );


  nor
  g2550
  (
    n1784,
    n1121,
    n1043,
    n976,
    n1115
  );


  nor
  g2551
  (
    n2042,
    n1246,
    n950,
    n1081,
    n1503
  );


  or
  g2552
  (
    n1982,
    n1757,
    n1544,
    n1607,
    n999
  );


  xor
  g2553
  (
    n1923,
    n979,
    n1066,
    n944,
    n931
  );


  xor
  g2554
  (
    n2445,
    n941,
    n1634,
    n1424,
    n1734
  );


  and
  g2555
  (
    n1933,
    n1743,
    n1421,
    n1656,
    n928
  );


  nand
  g2556
  (
    n2539,
    n1437,
    n1164,
    n1342,
    n1076
  );


  or
  g2557
  (
    n2442,
    n1039,
    n942,
    n1380,
    n1281
  );


  and
  g2558
  (
    n2522,
    n833,
    n1669,
    n1328,
    n831
  );


  xnor
  g2559
  (
    n1966,
    n1432,
    n1408,
    n1065,
    n1334
  );


  and
  g2560
  (
    n2032,
    n814,
    n1336,
    n1081,
    n1298
  );


  or
  g2561
  (
    n2396,
    n1746,
    n1352,
    n1114,
    n1436
  );


  xor
  g2562
  (
    n2205,
    n1162,
    n1638,
    n1172,
    n1005
  );


  and
  g2563
  (
    n2015,
    n1754,
    n1540,
    n1607,
    n1686
  );


  or
  g2564
  (
    n2113,
    n1498,
    n1483,
    n1605,
    n1512
  );


  xor
  g2565
  (
    n2344,
    n1243,
    n1014,
    n874,
    n1358
  );


  nor
  g2566
  (
    n1937,
    n1026,
    n932,
    n1695,
    n1434
  );


  nor
  g2567
  (
    n1880,
    n1002,
    n1659,
    n1648,
    n854
  );


  nand
  g2568
  (
    n2177,
    n880,
    n1636,
    n993,
    n1360
  );


  xor
  g2569
  (
    n1907,
    n1537,
    n1159,
    n1425,
    n1129
  );


  nand
  g2570
  (
    n2450,
    n977,
    n1464,
    n1378,
    n1124
  );


  or
  g2571
  (
    n1890,
    n1534,
    n1565,
    n1503,
    n1466
  );


  or
  g2572
  (
    n2172,
    n1101,
    n1587,
    n1080,
    n1238
  );


  and
  g2573
  (
    n2252,
    n1738,
    n1339,
    n1572,
    n1141
  );


  nor
  g2574
  (
    n2467,
    n1160,
    n1543,
    n1554,
    n1054
  );


  nor
  g2575
  (
    n2651,
    n1217,
    n1419,
    n1292,
    n1430
  );


  xor
  g2576
  (
    n2019,
    n1068,
    n1205,
    n1610,
    n1645
  );


  nor
  g2577
  (
    n2008,
    n1282,
    n1651,
    n1372,
    n1730
  );


  nand
  g2578
  (
    n2266,
    n1366,
    n1730,
    n1457,
    n1558
  );


  nand
  g2579
  (
    n2597,
    n1575,
    n1025,
    n1545,
    n1747
  );


  or
  g2580
  (
    n1977,
    n1683,
    n1266,
    n1408,
    n1150
  );


  xnor
  g2581
  (
    n1895,
    n828,
    n1110,
    n1752,
    n1206
  );


  xnor
  g2582
  (
    n2417,
    n1475,
    n974,
    n1331,
    n1561
  );


  xnor
  g2583
  (
    n2366,
    n1183,
    n1622,
    n1116,
    n1605
  );


  or
  g2584
  (
    n2405,
    n1691,
    n1563,
    n1706,
    n1391
  );


  xnor
  g2585
  (
    n2337,
    n1257,
    n1268,
    n1011,
    n1491
  );


  xor
  g2586
  (
    n2513,
    n1726,
    n1196,
    n1258,
    n936
  );


  or
  g2587
  (
    n1845,
    n1344,
    n1289,
    n972,
    n1611
  );


  nor
  g2588
  (
    n1802,
    n1572,
    n1341,
    n1275,
    n1429
  );


  or
  g2589
  (
    n1774,
    n1728,
    n1621,
    n1748,
    n1290
  );


  nor
  g2590
  (
    n2045,
    n1063,
    n1148,
    n1131,
    n1661
  );


  or
  g2591
  (
    n1980,
    n1544,
    n1381,
    n1640,
    n1284
  );


  or
  g2592
  (
    n2239,
    n1507,
    n992,
    n1460,
    n1084
  );


  xor
  g2593
  (
    n2502,
    n1426,
    n1031,
    n1273,
    n1041
  );


  xor
  g2594
  (
    n2349,
    n996,
    n1047,
    n1567,
    n1720
  );


  and
  g2595
  (
    n1807,
    n904,
    n1731,
    n1185,
    n962
  );


  nand
  g2596
  (
    n2247,
    n1307,
    n1495,
    n811,
    n1090
  );


  and
  g2597
  (
    n1801,
    n1627,
    n1694,
    n1389,
    n1131
  );


  xnor
  g2598
  (
    n2474,
    n961,
    n1366,
    n1644,
    n1203
  );


  nor
  g2599
  (
    n2397,
    n1653,
    n1727,
    n1627,
    n1235
  );


  nor
  g2600
  (
    n2225,
    n1469,
    n1441,
    n1323,
    n1196
  );


  and
  g2601
  (
    n1913,
    n1444,
    n1576,
    n892,
    n1675
  );


  nor
  g2602
  (
    n1867,
    n1544,
    n1304,
    n1453,
    n1504
  );


  xnor
  g2603
  (
    n2274,
    n1553,
    n1146,
    n986,
    n1296
  );


  nor
  g2604
  (
    n1912,
    n1463,
    n1666,
    n1314,
    n1324
  );


  xor
  g2605
  (
    n2338,
    n1376,
    n1725,
    n1749,
    n1397
  );


  or
  g2606
  (
    n1813,
    n1281,
    n1175,
    n1018,
    n1272
  );


  and
  g2607
  (
    n2399,
    n944,
    n1697,
    n922,
    n1166
  );


  and
  g2608
  (
    n2406,
    n987,
    n1266,
    n1623,
    n1758
  );


  and
  g2609
  (
    n2254,
    n1153,
    n1100,
    n1549,
    n1294
  );


  nand
  g2610
  (
    n2143,
    n1558,
    n1139,
    n1163,
    n1514
  );


  xnor
  g2611
  (
    n2067,
    n825,
    n1521,
    n1370,
    n1531
  );


  xnor
  g2612
  (
    n2661,
    n469,
    n1224,
    n1723,
    n945
  );


  and
  g2613
  (
    n1815,
    n1107,
    n947,
    n1205,
    n1589
  );


  nor
  g2614
  (
    n2587,
    n933,
    n1048,
    n1233,
    n1096
  );


  xnor
  g2615
  (
    n1805,
    n1083,
    n1573,
    n1210,
    n1251
  );


  xnor
  g2616
  (
    n2627,
    n1125,
    n1189,
    n844,
    n1590
  );


  xnor
  g2617
  (
    n2577,
    n1095,
    n1194,
    n1462,
    n1666
  );


  and
  g2618
  (
    n1991,
    n1340,
    n1155,
    n945,
    n910
  );


  or
  g2619
  (
    n2498,
    n1301,
    n1005,
    n1306,
    n964
  );


  xor
  g2620
  (
    n2575,
    n1355,
    n1377,
    n1593,
    n1403
  );


  xnor
  g2621
  (
    n2517,
    n1576,
    n1681,
    n969,
    n976
  );


  nand
  g2622
  (
    n1986,
    n1213,
    n1281,
    n1406,
    n1611
  );


  nor
  g2623
  (
    KeyWire_0_8,
    n1478,
    n1307,
    n1731,
    n1708
  );


  nand
  g2624
  (
    n2229,
    n1344,
    n1502,
    n1248,
    n1112
  );


  or
  g2625
  (
    n2005,
    n1374,
    n1225,
    n1599,
    n854
  );


  xnor
  g2626
  (
    n1963,
    n908,
    n1045,
    n1663,
    n1594
  );


  nand
  g2627
  (
    n1898,
    n1177,
    n1370,
    n1080,
    n1004
  );


  and
  g2628
  (
    n2640,
    n1731,
    n1329,
    n927,
    n891
  );


  xnor
  g2629
  (
    n1776,
    n1235,
    n991,
    n1207,
    n1738
  );


  xor
  g2630
  (
    n2635,
    n1730,
    n1156,
    n1414,
    n876
  );


  nor
  g2631
  (
    n2530,
    n1645,
    n832,
    n1616,
    n1577
  );


  and
  g2632
  (
    n2621,
    n1370,
    n1432,
    n972,
    n1224
  );


  or
  g2633
  (
    n2471,
    n1279,
    n891,
    n1718,
    n1723
  );


  nor
  g2634
  (
    n2365,
    n1291,
    n1164,
    n1439,
    n1267
  );


  or
  g2635
  (
    n2476,
    n1324,
    n1038,
    n1292,
    n1708
  );


  nand
  g2636
  (
    n2324,
    n1493,
    n1464,
    n1234,
    n895
  );


  and
  g2637
  (
    n2510,
    n826,
    n986,
    n1424,
    n1267
  );


  xor
  g2638
  (
    n2006,
    n1016,
    n1707,
    n1269,
    n893
  );


  nand
  g2639
  (
    n2237,
    n1725,
    n1047,
    n939,
    n1590
  );


  nand
  g2640
  (
    n2899,
    n1998,
    n2265,
    n2148,
    n1823
  );


  nor
  g2641
  (
    n2687,
    n2055,
    n1973,
    n1883,
    n2091
  );


  and
  g2642
  (
    n2681,
    n2203,
    n2134,
    n556,
    n2612
  );


  and
  g2643
  (
    n2805,
    n2369,
    n2393,
    n2464,
    n2586
  );


  nor
  g2644
  (
    n2748,
    n1980,
    n1984,
    n536,
    n2138
  );


  or
  g2645
  (
    n2695,
    n1793,
    n2497,
    n2085,
    n2040
  );


  nor
  g2646
  (
    n2816,
    n2246,
    n2582,
    n1783,
    n1847
  );


  xor
  g2647
  (
    n2901,
    n2263,
    n2509,
    n547,
    n1787
  );


  nand
  g2648
  (
    n2785,
    n1913,
    n1842,
    n2074,
    n2037
  );


  nor
  g2649
  (
    n2743,
    n2108,
    n1767,
    n2628,
    n2014
  );


  or
  g2650
  (
    n2903,
    n1914,
    n2450,
    n2529,
    n2648
  );


  nand
  g2651
  (
    n2843,
    n1854,
    n2064,
    n554,
    n2607
  );


  or
  g2652
  (
    n2845,
    n2201,
    n2240,
    n543,
    n2153
  );


  xor
  g2653
  (
    n2931,
    n1948,
    n1778,
    n559,
    n2069
  );


  nand
  g2654
  (
    n2862,
    n1877,
    n1918,
    n2645,
    n2062
  );


  nor
  g2655
  (
    n2918,
    n2462,
    n1929,
    n2295,
    n2411
  );


  and
  g2656
  (
    n2930,
    n2653,
    n547,
    n1795,
    n2538
  );


  or
  g2657
  (
    n2747,
    n2379,
    n1788,
    n544,
    n2116
  );


  xnor
  g2658
  (
    n2764,
    n2207,
    n2121,
    n2358,
    n2542
  );


  xnor
  g2659
  (
    n2821,
    n2096,
    n2182,
    n1760,
    n2010
  );


  and
  g2660
  (
    n2834,
    n2565,
    n2485,
    n2404,
    n2094
  );


  xnor
  g2661
  (
    n2803,
    n1899,
    n1863,
    n2083,
    n551
  );


  xor
  g2662
  (
    n2894,
    n2401,
    n2098,
    n1908,
    n2616
  );


  nand
  g2663
  (
    n2877,
    n2600,
    n537,
    n1840,
    n2343
  );


  nand
  g2664
  (
    n2674,
    n548,
    n534,
    n2657,
    n2321
  );


  nand
  g2665
  (
    n2910,
    n1828,
    n2534,
    n2076,
    n2079
  );


  or
  g2666
  (
    n2818,
    n541,
    n2298,
    n1796,
    n2031
  );


  nand
  g2667
  (
    n2879,
    n2621,
    n1844,
    n545,
    n560
  );


  and
  g2668
  (
    n2864,
    n2054,
    n2104,
    n2171,
    n1798
  );


  xnor
  g2669
  (
    n2753,
    n553,
    n2111,
    n1949,
    n2239
  );


  nor
  g2670
  (
    n2745,
    n551,
    n2555,
    n547,
    n2232
  );


  xor
  g2671
  (
    n2817,
    n1774,
    n540,
    n2258,
    n2328
  );


  or
  g2672
  (
    n2915,
    n2608,
    n1845,
    n2429,
    n2603
  );


  nor
  g2673
  (
    n2740,
    n2067,
    n2662,
    n1993,
    n2589
  );


  xnor
  g2674
  (
    n2923,
    n559,
    n1821,
    n544,
    n2424
  );


  nor
  g2675
  (
    n2788,
    n1763,
    n2660,
    n2101,
    n2456
  );


  xor
  g2676
  (
    n2784,
    n2403,
    n1806,
    n1925,
    n560
  );


  or
  g2677
  (
    n2715,
    n1895,
    n552,
    n2472,
    n2453
  );


  nor
  g2678
  (
    n2851,
    n2493,
    n1762,
    n2309,
    n542
  );


  xnor
  g2679
  (
    n2934,
    n2044,
    n2592,
    n2306,
    n2194
  );


  and
  g2680
  (
    n2812,
    n2564,
    n2231,
    n1898,
    n2090
  );


  nand
  g2681
  (
    n2770,
    n1979,
    n1983,
    n2406,
    n2544
  );


  nand
  g2682
  (
    n2850,
    n2305,
    n2155,
    n541,
    n559
  );


  or
  g2683
  (
    n2854,
    n2417,
    n2444,
    n551,
    n2262
  );


  or
  g2684
  (
    n2893,
    n1901,
    n2385,
    n2507,
    n2519
  );


  or
  g2685
  (
    n2677,
    n2303,
    n541,
    n554,
    n2034
  );


  and
  g2686
  (
    n2880,
    n2291,
    n2282,
    n539,
    n1961
  );


  or
  g2687
  (
    n2928,
    n1982,
    n1967,
    n1900,
    n540
  );


  or
  g2688
  (
    n2792,
    n2526,
    n2293,
    n2151,
    n2132
  );


  nor
  g2689
  (
    n2723,
    n2212,
    n2118,
    n2089,
    n2073
  );


  nand
  g2690
  (
    n2756,
    n1791,
    n2256,
    n533,
    n2136
  );


  and
  g2691
  (
    n2712,
    n2123,
    n2187,
    n2436,
    n2566
  );


  nor
  g2692
  (
    n2720,
    n1825,
    n2276,
    n2413,
    n553
  );


  xnor
  g2693
  (
    n2701,
    n2528,
    n2122,
    n1764,
    n2313
  );


  xor
  g2694
  (
    n2824,
    n1897,
    n2179,
    n2405,
    n2665
  );


  and
  g2695
  (
    n2733,
    n531,
    n544,
    n2659,
    n553
  );


  or
  g2696
  (
    n2833,
    n2381,
    n2340,
    n2466,
    n2552
  );


  nor
  g2697
  (
    n2693,
    n2113,
    n1880,
    n2125,
    n2220
  );


  or
  g2698
  (
    n2800,
    n1959,
    n2556,
    n2103,
    n2460
  );


  xor
  g2699
  (
    n2813,
    n2052,
    n549,
    n2557,
    n2081
  );


  and
  g2700
  (
    n2705,
    n2004,
    n559,
    n558,
    n538
  );


  nor
  g2701
  (
    n2684,
    n1892,
    n2175,
    n2233,
    n2003
  );


  xor
  g2702
  (
    n2755,
    n532,
    n2334,
    n542,
    n2513
  );


  nor
  g2703
  (
    n2832,
    n563,
    n2189,
    n2409,
    n1893
  );


  xor
  g2704
  (
    n2709,
    n2229,
    n550,
    n2013,
    n2654
  );


  and
  g2705
  (
    n2922,
    n1938,
    n2541,
    n2366,
    n2459
  );


  and
  g2706
  (
    n2891,
    n539,
    n2102,
    n1891,
    n548
  );


  xnor
  g2707
  (
    n2916,
    n1920,
    n2290,
    n2152,
    n535
  );


  nor
  g2708
  (
    n2781,
    n2162,
    n1860,
    n536,
    n1830
  );


  nor
  g2709
  (
    n2819,
    n1906,
    n2144,
    n1775,
    n2188
  );


  xnor
  g2710
  (
    n2920,
    n1894,
    n2433,
    n2086,
    n2224
  );


  xnor
  g2711
  (
    n2734,
    n1997,
    n552,
    n2249,
    n2389
  );


  nand
  g2712
  (
    n2777,
    n1857,
    n2065,
    n2667,
    n1810
  );


  or
  g2713
  (
    n2768,
    n534,
    n2584,
    n2384,
    n550
  );


  xor
  g2714
  (
    n2758,
    n555,
    n2025,
    n2341,
    n2095
  );


  or
  g2715
  (
    n2914,
    n2351,
    n2668,
    n543,
    n2169
  );


  xnor
  g2716
  (
    n2908,
    n1808,
    n2011,
    n2627,
    n2092
  );


  nand
  g2717
  (
    n2856,
    n557,
    n1786,
    n2312,
    n2451
  );


  or
  g2718
  (
    n2921,
    n562,
    n2088,
    n2043,
    n2082
  );


  and
  g2719
  (
    n2749,
    n2183,
    n2614,
    n2364,
    n2039
  );


  xor
  g2720
  (
    n2895,
    n1849,
    n2075,
    n2651,
    n550
  );


  nor
  g2721
  (
    n2700,
    n2524,
    n532,
    n2310,
    n1996
  );


  nor
  g2722
  (
    n2759,
    n2007,
    n2506,
    n1820,
    n2247
  );


  nand
  g2723
  (
    n2860,
    n1989,
    n1861,
    n2147,
    n2511
  );


  and
  g2724
  (
    n2760,
    n533,
    n2211,
    n1813,
    n535
  );


  xor
  g2725
  (
    n2841,
    n2269,
    n2235,
    n2480,
    n1922
  );


  and
  g2726
  (
    n2796,
    n2346,
    n2471,
    n2015,
    n2397
  );


  nand
  g2727
  (
    n2898,
    n1812,
    n2489,
    n1896,
    n2392
  );


  or
  g2728
  (
    n2885,
    n1927,
    n2241,
    n1807,
    n2546
  );


  xnor
  g2729
  (
    n2874,
    n2289,
    n2613,
    n1839,
    n546
  );


  nand
  g2730
  (
    KeyWire_0_0,
    n563,
    n1819,
    n2170,
    n2443
  );


  nand
  g2731
  (
    n2842,
    n2629,
    n2331,
    n1995,
    n535
  );


  and
  g2732
  (
    n2829,
    n1785,
    n2448,
    n1831,
    n1972
  );


  nor
  g2733
  (
    n2929,
    n2315,
    n2377,
    n2537,
    n2056
  );


  nand
  g2734
  (
    n2838,
    n2597,
    n2322,
    n538,
    n2483
  );


  xor
  g2735
  (
    n2791,
    n1962,
    n2458,
    n2033,
    n2338
  );


  xor
  g2736
  (
    n2811,
    n2661,
    n2349,
    n2260,
    n540
  );


  nand
  g2737
  (
    n2673,
    n1781,
    n544,
    n2540,
    n1815
  );


  or
  g2738
  (
    n2896,
    n1941,
    n2640,
    n2484,
    n2469
  );


  nor
  g2739
  (
    n2825,
    n564,
    n2470,
    n2045,
    n1957
  );


  and
  g2740
  (
    n2773,
    n2286,
    n2160,
    n1772,
    n2317
  );


  xnor
  g2741
  (
    n2775,
    n2307,
    n1951,
    n2219,
    n1946
  );


  nand
  g2742
  (
    n2927,
    n1974,
    n2359,
    n1924,
    n2165
  );


  nand
  g2743
  (
    n2859,
    n2617,
    n2588,
    n2655,
    n1987
  );


  xnor
  g2744
  (
    n2807,
    n1872,
    n2129,
    n2029,
    n1867
  );


  or
  g2745
  (
    n2762,
    n539,
    n2656,
    n2311,
    n1960
  );


  nand
  g2746
  (
    n2878,
    n1994,
    n2163,
    n2634,
    n2422
  );


  xor
  g2747
  (
    n2875,
    n2070,
    n1888,
    n2105,
    n537
  );


  nor
  g2748
  (
    n2872,
    n529,
    n2242,
    n555,
    n1809
  );


  xor
  g2749
  (
    n2865,
    n2330,
    n1838,
    n1910,
    n1869
  );


  and
  g2750
  (
    n2804,
    n1818,
    n1865,
    n2498,
    n1904
  );


  xor
  g2751
  (
    n2909,
    n2535,
    n2314,
    n2585,
    n2058
  );


  and
  g2752
  (
    n2766,
    n2402,
    n2461,
    n2439,
    n2467
  );


  nand
  g2753
  (
    n2884,
    n1968,
    n1976,
    n2142,
    n2623
  );


  xnor
  g2754
  (
    n2849,
    n2371,
    n2124,
    n556,
    n2005
  );


  nor
  g2755
  (
    n2754,
    n2195,
    n2042,
    n533,
    n2490
  );


  nand
  g2756
  (
    n2913,
    n2287,
    n2583,
    n1803,
    n1955
  );


  xnor
  g2757
  (
    n2774,
    n2624,
    n2531,
    n1903,
    n19
  );


  xor
  g2758
  (
    n2806,
    n2375,
    n2325,
    n2333,
    n1804
  );


  or
  g2759
  (
    n2726,
    n1766,
    n2173,
    n2492,
    n2591
  );


  or
  g2760
  (
    n2765,
    n1848,
    n2022,
    n2202,
    n2077
  );


  or
  g2761
  (
    n2683,
    n2251,
    n1969,
    n1928,
    n2057
  );


  or
  g2762
  (
    n2732,
    n1921,
    n2133,
    n2590,
    n555
  );


  xnor
  g2763
  (
    n2675,
    n531,
    n2639,
    n2353,
    n2598
  );


  and
  g2764
  (
    n2696,
    n2185,
    n2264,
    n2087,
    n2271
  );


  and
  g2765
  (
    n2706,
    n2178,
    n2255,
    n1912,
    n2294
  );


  nand
  g2766
  (
    n2846,
    n2354,
    n2652,
    n19,
    n2465
  );


  nand
  g2767
  (
    n2897,
    n2177,
    n2299,
    n2633,
    n2391
  );


  nor
  g2768
  (
    n2847,
    n1931,
    n534,
    n2505,
    n2669
  );


  xor
  g2769
  (
    n2855,
    n2197,
    n560,
    n2259,
    n1858
  );


  xnor
  g2770
  (
    n2721,
    n2140,
    n1871,
    n1970,
    n1799
  );


  nand
  g2771
  (
    n2757,
    n1874,
    n2644,
    n1954,
    n1887
  );


  nand
  g2772
  (
    n2799,
    n2109,
    n1800,
    n1769,
    n2428
  );


  nand
  g2773
  (
    n2868,
    n2018,
    n1965,
    n2559,
    n2440
  );


  nand
  g2774
  (
    n2702,
    n2622,
    n1878,
    n2410,
    n1963
  );


  or
  g2775
  (
    n2797,
    n2210,
    n2571,
    n2320,
    n1966
  );


  xnor
  g2776
  (
    n2685,
    n2107,
    n540,
    n2352,
    n1853
  );


  and
  g2777
  (
    n2907,
    n2049,
    n2512,
    n2006,
    n2337
  );


  nand
  g2778
  (
    n2704,
    n2072,
    n1761,
    n2008,
    n2510
  );


  or
  g2779
  (
    n2919,
    n2275,
    n2390,
    n2036,
    n2431
  );


  xor
  g2780
  (
    n2926,
    n2180,
    n546,
    n2416,
    n1881
  );


  nand
  g2781
  (
    n2873,
    n2002,
    n1864,
    n2604,
    n1905
  );


  xnor
  g2782
  (
    n2912,
    n2618,
    n2615,
    n545,
    n2161
  );


  nor
  g2783
  (
    n2776,
    n2174,
    n1919,
    n2475,
    n1992
  );


  nand
  g2784
  (
    n2814,
    n2281,
    n2131,
    n533,
    n2327
  );


  xnor
  g2785
  (
    n2778,
    n2396,
    n2488,
    n536,
    n1953
  );


  and
  g2786
  (
    n2790,
    n2380,
    n2270,
    n530,
    n2225
  );


  xor
  g2787
  (
    n2871,
    n2209,
    n1822,
    n2503,
    n532
  );


  xor
  g2788
  (
    n2857,
    n2019,
    n2670,
    n2620,
    n547
  );


  or
  g2789
  (
    n2780,
    n2273,
    n1936,
    n534,
    n2370
  );


  or
  g2790
  (
    n2870,
    n1986,
    n564,
    n1876,
    n2110
  );


  or
  g2791
  (
    n2828,
    n2355,
    n535,
    n1836,
    n2135
  );


  xnor
  g2792
  (
    n2782,
    n2230,
    n2601,
    n2030,
    n1833
  );


  xnor
  g2793
  (
    n2911,
    n543,
    n1846,
    n2218,
    n2248
  );


  or
  g2794
  (
    n2787,
    n2227,
    n2641,
    n2205,
    n2336
  );


  xor
  g2795
  (
    n2746,
    n2176,
    n2452,
    n2097,
    n2572
  );


  nor
  g2796
  (
    n2917,
    n2494,
    n1829,
    n2468,
    n2017
  );


  nand
  g2797
  (
    n2802,
    n541,
    n548,
    n2560,
    n1868
  );


  or
  g2798
  (
    n2730,
    n2252,
    n552,
    n2001,
    n2344
  );


  nor
  g2799
  (
    n2707,
    n2549,
    n2570,
    n2166,
    n530
  );


  nand
  g2800
  (
    n2826,
    n1837,
    n2296,
    n2243,
    n1777
  );


  nor
  g2801
  (
    n2761,
    n2398,
    n2184,
    n2671,
    n2474
  );


  nor
  g2802
  (
    n2703,
    n2548,
    n1834,
    n2143,
    n1958
  );


  and
  g2803
  (
    n2682,
    n2345,
    n2527,
    n1942,
    n2332
  );


  nand
  g2804
  (
    n2881,
    n2316,
    n2525,
    n557,
    n2536
  );


  or
  g2805
  (
    n2801,
    n2035,
    n1889,
    n2139,
    n2159
  );


  nand
  g2806
  (
    n2837,
    n1981,
    n536,
    n2362,
    n1835
  );


  nor
  g2807
  (
    n2738,
    n2360,
    n2192,
    n2575,
    n2223
  );


  xnor
  g2808
  (
    n2751,
    n2181,
    n551,
    n1907,
    n1862
  );


  and
  g2809
  (
    n2925,
    n1930,
    n2473,
    n2630,
    n550
  );


  or
  g2810
  (
    n2727,
    n554,
    n2574,
    n2532,
    n2382
  );


  nand
  g2811
  (
    n2853,
    n561,
    n1790,
    n1826,
    n2164
  );


  nor
  g2812
  (
    n2716,
    n2288,
    n2020,
    n2516,
    n2193
  );


  or
  g2813
  (
    n2713,
    n2567,
    n1870,
    n2078,
    n2114
  );


  xnor
  g2814
  (
    n2731,
    n2491,
    n1816,
    n558,
    n2602
  );


  nand
  g2815
  (
    n2699,
    n2539,
    n2388,
    n2228,
    n1977
  );


  xor
  g2816
  (
    n2767,
    n2646,
    n561,
    n2420,
    n1882
  );


  nor
  g2817
  (
    n2886,
    n2477,
    n1917,
    n2245,
    n2547
  );


  xnor
  g2818
  (
    n2839,
    n2569,
    n1952,
    n1782,
    n1950
  );


  xor
  g2819
  (
    n2711,
    n2579,
    n2666,
    n2244,
    n2186
  );


  and
  g2820
  (
    n2831,
    n2284,
    n2515,
    n1776,
    n2545
  );


  and
  g2821
  (
    n2904,
    n2323,
    n546,
    n2376,
    n2374
  );


  or
  g2822
  (
    n2694,
    n2635,
    n1909,
    n2204,
    n2280
  );


  nor
  g2823
  (
    n2889,
    n2348,
    n2261,
    n545,
    n1944
  );


  or
  g2824
  (
    n2680,
    n2606,
    n2300,
    n2449,
    n2658
  );


  nand
  g2825
  (
    n2809,
    n542,
    n2196,
    n2217,
    n562
  );


  or
  g2826
  (
    n2836,
    n2533,
    n562,
    n2550,
    n556
  );


  nand
  g2827
  (
    n2793,
    n2499,
    n1780,
    n2080,
    n561
  );


  xnor
  g2828
  (
    n2810,
    n2430,
    n2191,
    n2495,
    n2266
  );


  nand
  g2829
  (
    n2724,
    n2253,
    n2500,
    n2415,
    n558
  );


  nand
  g2830
  (
    n2905,
    n1765,
    n2558,
    n538,
    n1886
  );


  and
  g2831
  (
    n2725,
    n538,
    n2368,
    n1794,
    n2543
  );


  nand
  g2832
  (
    n2840,
    n2339,
    n2383,
    n564,
    n1943
  );


  and
  g2833
  (
    n2867,
    n2577,
    n2117,
    n1975,
    n1814
  );


  or
  g2834
  (
    n2735,
    n1805,
    n2100,
    n1792,
    n530
  );


  xor
  g2835
  (
    n2932,
    n2326,
    n562,
    n2518,
    n563
  );


  nand
  g2836
  (
    n2718,
    n2206,
    n2372,
    n556,
    n561
  );


  or
  g2837
  (
    n2692,
    n2664,
    n548,
    n537,
    n1859
  );


  xor
  g2838
  (
    n2858,
    n2038,
    n2016,
    n2084,
    n1784
  );


  nor
  g2839
  (
    n2887,
    n2427,
    n2520,
    n1850,
    n2277
  );


  and
  g2840
  (
    n2906,
    n2580,
    n2576,
    n2400,
    n2168
  );


  nand
  g2841
  (
    n2900,
    n537,
    n2154,
    n2551,
    n2254
  );


  nand
  g2842
  (
    n2795,
    n555,
    n2208,
    n2446,
    n1971
  );


  nor
  g2843
  (
    n2736,
    n1856,
    n2093,
    n2009,
    n2128
  );


  xnor
  g2844
  (
    n2714,
    n2611,
    n1852,
    n532,
    n2071
  );


  xor
  g2845
  (
    n2902,
    n2553,
    n2454,
    n557,
    n2050
  );


  or
  g2846
  (
    n2690,
    n2496,
    n1999,
    n2365,
    n552
  );


  or
  g2847
  (
    n2892,
    n2399,
    n2599,
    n2441,
    n1947
  );


  xnor
  g2848
  (
    n2686,
    n531,
    n2407,
    n2221,
    n1770
  );


  xor
  g2849
  (
    n2861,
    n1939,
    n2156,
    n2149,
    n2373
  );


  xnor
  g2850
  (
    n2883,
    n2663,
    n2274,
    n2357,
    n1811
  );


  xnor
  g2851
  (
    n2936,
    n2000,
    n2061,
    n1964,
    n1801
  );


  and
  g2852
  (
    n2789,
    n1851,
    n2502,
    n1843,
    n2047
  );


  xnor
  g2853
  (
    n2844,
    n2363,
    n1885,
    n2554,
    n1956
  );


  nand
  g2854
  (
    n2741,
    n549,
    n2051,
    n2463,
    n2412
  );


  xor
  g2855
  (
    n2798,
    n1873,
    n2200,
    n1935,
    n2522
  );


  xor
  g2856
  (
    n2697,
    n2234,
    n1841,
    n2115,
    n549
  );


  or
  g2857
  (
    n2786,
    n530,
    n1802,
    n2435,
    n545
  );


  or
  g2858
  (
    n2830,
    n2053,
    n2041,
    n2395,
    n2158
  );


  xnor
  g2859
  (
    n2933,
    n2632,
    n2021,
    n1934,
    n1916
  );


  xor
  g2860
  (
    n2698,
    n2426,
    n2610,
    n2425,
    n2442
  );


  nor
  g2861
  (
    n2808,
    n2026,
    n2347,
    n2157,
    n2238
  );


  xnor
  g2862
  (
    n2689,
    n2573,
    n2350,
    n539,
    n2578
  );


  and
  g2863
  (
    n2848,
    n2012,
    n531,
    n2650,
    n2479
  );


  xnor
  g2864
  (
    n2769,
    n2285,
    n2215,
    n2421,
    n2478
  );


  xor
  g2865
  (
    n2679,
    n558,
    n2605,
    n2387,
    n2126
  );


  xor
  g2866
  (
    n2827,
    n1817,
    n2563,
    n2408,
    n2523
  );


  nor
  g2867
  (
    n2691,
    n1978,
    n2146,
    n2267,
    n2561
  );


  xnor
  g2868
  (
    n2783,
    n543,
    n2023,
    n1773,
    n2481
  );


  nor
  g2869
  (
    n2882,
    n2447,
    n2642,
    n2587,
    n1991
  );


  or
  g2870
  (
    n2876,
    n2130,
    n2595,
    n1866,
    n2272
  );


  nor
  g2871
  (
    n2737,
    n2637,
    n1789,
    n2568,
    n2626
  );


  or
  g2872
  (
    n2719,
    n2418,
    n2419,
    n2342,
    n2127
  );


  xor
  g2873
  (
    n2869,
    n2521,
    n2643,
    n2060,
    n2236
  );


  or
  g2874
  (
    n2924,
    n2268,
    n1940,
    n1933,
    n557
  );


  and
  g2875
  (
    n2835,
    n2226,
    n2190,
    n1768,
    n2432
  );


  xor
  g2876
  (
    KeyWire_0_15,
    n549,
    n2137,
    n2455,
    n554
  );


  or
  g2877
  (
    n2820,
    n1990,
    n1988,
    n563,
    n2517
  );


  nor
  g2878
  (
    n2722,
    n2501,
    n1915,
    n2476,
    n2356
  );


  and
  g2879
  (
    n2863,
    n2625,
    n2257,
    n2048,
    n2059
  );


  xor
  g2880
  (
    n2739,
    n2672,
    n1945,
    n2214,
    n553
  );


  xnor
  g2881
  (
    n2742,
    n2562,
    n2027,
    n2024,
    n2457
  );


  nor
  g2882
  (
    n2794,
    n2237,
    n2106,
    n2308,
    n2394
  );


  xor
  g2883
  (
    n2890,
    n2647,
    n2486,
    n1879,
    n2046
  );


  or
  g2884
  (
    n2676,
    n2066,
    n2292,
    n2150,
    n1855
  );


  xnor
  g2885
  (
    n2822,
    n2361,
    n2145,
    n1911,
    n1827
  );


  and
  g2886
  (
    n2771,
    n2028,
    n2386,
    n2631,
    n2504
  );


  xnor
  g2887
  (
    n2728,
    n2530,
    n546,
    n2636,
    n2581
  );


  nor
  g2888
  (
    n2815,
    n2319,
    n2508,
    n1890,
    n1824
  );


  xnor
  g2889
  (
    n2823,
    n2198,
    n2619,
    n1884,
    n2283
  );


  xnor
  g2890
  (
    n2710,
    n2172,
    n2434,
    n1985,
    n2120
  );


  and
  g2891
  (
    n2772,
    n1937,
    n2638,
    n2063,
    n2594
  );


  or
  g2892
  (
    n2888,
    n2216,
    n2593,
    n2318,
    n2199
  );


  xnor
  g2893
  (
    n2688,
    n2487,
    n2423,
    n2514,
    n1771
  );


  xnor
  g2894
  (
    n2935,
    n2367,
    n2302,
    n2304,
    n2068
  );


  xnor
  g2895
  (
    n2708,
    n560,
    n2119,
    n2649,
    n2335
  );


  or
  g2896
  (
    n2717,
    n2301,
    n2279,
    n542,
    n1926
  );


  xor
  g2897
  (
    n2752,
    n2167,
    n2222,
    n2250,
    n2445
  );


  or
  g2898
  (
    n2729,
    n2378,
    n1923,
    n2213,
    n2482
  );


  nand
  g2899
  (
    n2678,
    n2609,
    n2141,
    n2112,
    n1875
  );


  xor
  g2900
  (
    n2763,
    n2278,
    n1932,
    n1832,
    n1779
  );


  xnor
  g2901
  (
    n2852,
    n564,
    n2596,
    n2324,
    n1902
  );


  xor
  g2902
  (
    n2750,
    n2437,
    n2414,
    n1797,
    n2329
  );


  and
  g2903
  (
    n2779,
    n2438,
    n2099,
    n2032,
    n2297
  );


  xnor
  g2904
  (
    n2988,
    n2861,
    n2873,
    n2924,
    n2682
  );


  nor
  g2905
  (
    n2986,
    n2911,
    n2746,
    n2830,
    n2725
  );


  or
  g2906
  (
    n2947,
    n2838,
    n2818,
    n2887,
    n2875
  );


  xnor
  g2907
  (
    n2957,
    n2835,
    n2878,
    n2865,
    n2817
  );


  xnor
  g2908
  (
    n2970,
    n2919,
    n2900,
    n2772,
    n2715
  );


  and
  g2909
  (
    n2981,
    n2708,
    n2859,
    n2773,
    n2793
  );


  xor
  g2910
  (
    n2991,
    n2781,
    n2896,
    n2931,
    n2706
  );


  nor
  g2911
  (
    n3002,
    n2871,
    n2720,
    n2744,
    n2893
  );


  nand
  g2912
  (
    n2990,
    n2918,
    n2680,
    n2740,
    n2685
  );


  nor
  g2913
  (
    n3000,
    n2925,
    n2770,
    n2674,
    n2867
  );


  nor
  g2914
  (
    n2976,
    n2749,
    n2774,
    n2805,
    n2762
  );


  nand
  g2915
  (
    n2952,
    n2910,
    n2935,
    n2872,
    n2771
  );


  or
  g2916
  (
    n2940,
    n2903,
    n2876,
    n2687,
    n2756
  );


  or
  g2917
  (
    n2984,
    n2791,
    n2747,
    n2798,
    n2923
  );


  xnor
  g2918
  (
    n2972,
    n2928,
    n2738,
    n2832,
    n2842
  );


  or
  g2919
  (
    n2966,
    n2857,
    n2922,
    n2902,
    n2884
  );


  or
  g2920
  (
    n2983,
    n2863,
    n2727,
    n2702,
    n2881
  );


  nand
  g2921
  (
    n2998,
    n2840,
    n2719,
    n2778,
    n2731
  );


  xor
  g2922
  (
    n2955,
    n2752,
    n2811,
    n2797,
    n2689
  );


  nand
  g2923
  (
    n2968,
    n2834,
    n2792,
    n2823,
    n2898
  );


  or
  g2924
  (
    n2941,
    n2717,
    n2850,
    n2849,
    n2809
  );


  xnor
  g2925
  (
    n2948,
    n2906,
    n2782,
    n2754,
    n2750
  );


  nor
  g2926
  (
    n2975,
    n2803,
    n2844,
    n2882,
    n2721
  );


  xor
  g2927
  (
    KeyWire_0_24,
    n2733,
    n2712,
    n2877,
    n2810
  );


  nand
  g2928
  (
    n2946,
    n2814,
    n2710,
    n2776,
    n2693
  );


  nand
  g2929
  (
    n2959,
    n2930,
    n2933,
    n2934,
    n2794
  );


  nor
  g2930
  (
    n2994,
    n2913,
    n2815,
    n2723,
    n2788
  );


  and
  g2931
  (
    n2939,
    n2886,
    n2899,
    n2713,
    n2914
  );


  and
  g2932
  (
    n2963,
    n2711,
    n2737,
    n2856,
    n2845
  );


  nand
  g2933
  (
    n2956,
    n2885,
    n2764,
    n2783,
    n2890
  );


  xor
  g2934
  (
    n2942,
    n2769,
    n2826,
    n2676,
    n2912
  );


  or
  g2935
  (
    n2973,
    n2908,
    n2880,
    n2801,
    n2833
  );


  xnor
  g2936
  (
    n2945,
    n2780,
    n2707,
    n2868,
    n2795
  );


  or
  g2937
  (
    n2954,
    n2714,
    n2690,
    n2800,
    n2821
  );


  nor
  g2938
  (
    n2951,
    n2837,
    n2929,
    n2848,
    n2820
  );


  and
  g2939
  (
    n2969,
    n2894,
    n2813,
    n2681,
    n2870
  );


  or
  g2940
  (
    n2965,
    n2785,
    n2866,
    n2812,
    n2828
  );


  nor
  g2941
  (
    n2996,
    n2879,
    n2757,
    n2745,
    n2921
  );


  xor
  g2942
  (
    n3001,
    n2704,
    n2694,
    n2824,
    n2915
  );


  nand
  g2943
  (
    n2985,
    n2829,
    n2728,
    n2718,
    n2730
  );


  xor
  g2944
  (
    n2958,
    n2796,
    n2843,
    n2678,
    n2790
  );


  xor
  g2945
  (
    n2977,
    n2751,
    n2724,
    n2787,
    n2777
  );


  and
  g2946
  (
    n2961,
    n2860,
    n2729,
    n2864,
    n2767
  );


  and
  g2947
  (
    n2980,
    n2858,
    n2853,
    n2831,
    n2722
  );


  xnor
  g2948
  (
    n2964,
    n2869,
    n2716,
    n2734,
    n2804
  );


  nand
  g2949
  (
    n2989,
    n2761,
    n2735,
    n2802,
    n2698
  );


  xor
  g2950
  (
    n2950,
    n2688,
    n2695,
    n2736,
    n2768
  );


  nand
  g2951
  (
    n2987,
    n2841,
    n2808,
    n2763,
    n2679
  );


  xnor
  g2952
  (
    n2960,
    n2700,
    n2836,
    n2748,
    n2799
  );


  or
  g2953
  (
    n2997,
    n2839,
    n2904,
    n2901,
    n2909
  );


  nand
  g2954
  (
    n2962,
    n2701,
    n2692,
    n2784,
    n2917
  );


  nand
  g2955
  (
    n2953,
    n2789,
    n2807,
    n2726,
    n2753
  );


  and
  g2956
  (
    n2943,
    n2932,
    n2743,
    n2892,
    n2779
  );


  xor
  g2957
  (
    n2999,
    n2907,
    n2883,
    n2677,
    n2895
  );


  or
  g2958
  (
    n2979,
    n2897,
    n2755,
    n2675,
    n2739
  );


  nand
  g2959
  (
    n2995,
    n2825,
    n2742,
    n2891,
    n2775
  );


  nor
  g2960
  (
    n2944,
    n2816,
    n2936,
    n2889,
    n2847
  );


  and
  g2961
  (
    n2992,
    n2697,
    n2926,
    n2827,
    n2905
  );


  xnor
  g2962
  (
    n2982,
    n2691,
    n2684,
    n2683,
    n2732
  );


  or
  g2963
  (
    n2949,
    n2741,
    n2699,
    n2854,
    n2822
  );


  nand
  g2964
  (
    n2974,
    n2862,
    n2874,
    n2806,
    n2765
  );


  or
  g2965
  (
    n2971,
    n2920,
    n2851,
    n2927,
    n2673
  );


  xor
  g2966
  (
    n2967,
    n2758,
    n2916,
    n2759,
    n2696
  );


  nand
  g2967
  (
    n2937,
    n2888,
    n2760,
    n2855,
    n2686
  );


  nor
  g2968
  (
    n2938,
    n2705,
    n2819,
    n2786,
    n2709
  );


  nand
  g2969
  (
    n2978,
    n2846,
    n2703,
    n2766,
    n2852
  );


  nand
  g2970
  (
    n3011,
    n2979,
    n2966,
    n2940,
    n2975
  );


  and
  g2971
  (
    n3015,
    n2959,
    n2954,
    n21,
    n2978
  );


  xor
  g2972
  (
    n3023,
    n26,
    n2984,
    n2938,
    n23
  );


  xnor
  g2973
  (
    n3018,
    n3000,
    n2955,
    n2945,
    n27
  );


  xnor
  g2974
  (
    n3030,
    n25,
    n2951,
    n31,
    n27
  );


  and
  g2975
  (
    n3019,
    n2976,
    n19,
    n2977,
    n24
  );


  nand
  g2976
  (
    n3025,
    n2953,
    n23,
    n2937,
    n22
  );


  xnor
  g2977
  (
    n3022,
    n2999,
    n2967,
    n2972,
    n27
  );


  nor
  g2978
  (
    n3012,
    n20,
    n2949,
    n2985,
    n32
  );


  or
  g2979
  (
    n3020,
    n29,
    n21,
    n27,
    n24
  );


  or
  g2980
  (
    n3006,
    n29,
    n2941,
    n24,
    n25
  );


  nand
  g2981
  (
    n3008,
    n26,
    n21,
    n2965,
    n2939
  );


  nor
  g2982
  (
    n3007,
    n19,
    n2944,
    n30,
    n2943
  );


  nand
  g2983
  (
    n3004,
    n2980,
    n20,
    n2986,
    n29
  );


  and
  g2984
  (
    n3028,
    n23,
    n28,
    n2987
  );


  nor
  g2985
  (
    n3016,
    n32,
    n2990,
    n2970,
    n2969
  );


  or
  g2986
  (
    n3003,
    n2994,
    n2961,
    n26,
    n30
  );


  and
  g2987
  (
    n3026,
    n26,
    n2981,
    n2974,
    n2950
  );


  nor
  g2988
  (
    n3009,
    n2991,
    n2963,
    n21,
    n2962
  );


  nor
  g2989
  (
    n3017,
    n2996,
    n31,
    n22
  );


  xor
  g2990
  (
    n3021,
    n2958,
    n2971,
    n2960,
    n2993
  );


  xnor
  g2991
  (
    n3032,
    n2948,
    n3001,
    n2995,
    n23
  );


  xnor
  g2992
  (
    n3027,
    n2989,
    n29,
    n2973,
    n2968
  );


  xor
  g2993
  (
    n3013,
    n28,
    n3002,
    n2947,
    n2983
  );


  xnor
  g2994
  (
    n3029,
    n2946,
    n22,
    n30,
    n32
  );


  xor
  g2995
  (
    n3010,
    n2997,
    n2942,
    n24,
    n2964
  );


  xor
  g2996
  (
    n3005,
    n2998,
    n2992,
    n30,
    n20
  );


  nand
  g2997
  (
    n3024,
    n25,
    n2957,
    n31,
    n2956
  );


  and
  g2998
  (
    n3014,
    n32,
    n20,
    n31,
    n25
  );


  or
  g2999
  (
    n3031,
    n2952,
    n2988,
    n2982,
    n28
  );


  xor
  KeyGate_0_0
  (
    n2744,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n2671,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n1092,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n2216,
    keyIn_0_3,
    KeyWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n2462,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n725,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1847,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n1283,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1792,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n737,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n1429,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n312,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n433,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n1144,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n185,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n2866,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1799,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n1323,
    keyIn_0_17,
    KeyWire_0_17
  );


  xnor
  KeyGate_0_18
  (
    n697,
    keyIn_0_18,
    KeyWire_0_18
  );


  xnor
  KeyGate_0_19
  (
    n1081,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1944,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    n1005,
    keyIn_0_21,
    KeyWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n2098,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n2607,
    keyIn_0_23,
    KeyWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n2993,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n1183,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1151,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n983,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1300,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n904,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n2322,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n779,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


