

module Stat_2749_29_1
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n2466,
  n2459,
  n2515,
  n2748,
  n2757,
  n2770,
  n2755,
  n2774,
  n2759,
  n2742,
  n2766,
  n2747,
  n2773,
  n2743,
  n2772,
  n2761,
  n2749,
  n2752,
  n2763,
  n2746,
  n2762,
  n2768,
  n2758,
  n2741,
  n2753,
  n2764,
  n2751,
  n2767,
  n2750,
  n2756,
  n2745,
  n2769,
  n2760,
  n2765,
  n2744,
  n2754,
  n2771
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n2466;output n2459;output n2515;output n2748;output n2757;output n2770;output n2755;output n2774;output n2759;output n2742;output n2766;output n2747;output n2773;output n2743;output n2772;output n2761;output n2749;output n2752;output n2763;output n2746;output n2762;output n2768;output n2758;output n2741;output n2753;output n2764;output n2751;output n2767;output n2750;output n2756;output n2745;output n2769;output n2760;output n2765;output n2744;output n2754;output n2771;
  wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  buf
  g0
  (
    n88,
    n12
  );


  buf
  g1
  (
    n105,
    n9
  );


  not
  g2
  (
    n90,
    n13
  );


  buf
  g3
  (
    n106,
    n9
  );


  buf
  g4
  (
    n92,
    n19
  );


  buf
  g5
  (
    n63,
    n7
  );


  not
  g6
  (
    n57,
    n13
  );


  buf
  g7
  (
    n77,
    n5
  );


  not
  g8
  (
    n66,
    n2
  );


  not
  g9
  (
    n85,
    n6
  );


  buf
  g10
  (
    n50,
    n16
  );


  not
  g11
  (
    n47,
    n4
  );


  buf
  g12
  (
    n40,
    n19
  );


  not
  g13
  (
    n51,
    n4
  );


  buf
  g14
  (
    n84,
    n15
  );


  not
  g15
  (
    n37,
    n4
  );


  not
  g16
  (
    n30,
    n5
  );


  not
  g17
  (
    n73,
    n21
  );


  not
  g18
  (
    n75,
    n19
  );


  not
  g19
  (
    n97,
    n18
  );


  buf
  g20
  (
    n98,
    n3
  );


  buf
  g21
  (
    n76,
    n8
  );


  buf
  g22
  (
    n48,
    n8
  );


  buf
  g23
  (
    n46,
    n6
  );


  buf
  g24
  (
    n29,
    n3
  );


  buf
  g25
  (
    n100,
    n20
  );


  not
  g26
  (
    n86,
    n13
  );


  not
  g27
  (
    n42,
    n2
  );


  buf
  g28
  (
    n59,
    n12
  );


  not
  g29
  (
    n81,
    n17
  );


  not
  g30
  (
    n104,
    n18
  );


  buf
  g31
  (
    n55,
    n14
  );


  buf
  g32
  (
    n53,
    n6
  );


  buf
  g33
  (
    n83,
    n14
  );


  not
  g34
  (
    n28,
    n20
  );


  buf
  g35
  (
    n54,
    n14
  );


  not
  g36
  (
    n101,
    n3
  );


  buf
  g37
  (
    n33,
    n9
  );


  not
  g38
  (
    n45,
    n7
  );


  buf
  g39
  (
    n64,
    n5
  );


  not
  g40
  (
    n102,
    n17
  );


  not
  g41
  (
    n89,
    n2
  );


  not
  g42
  (
    n44,
    n9
  );


  not
  g43
  (
    KeyWire_0_31,
    n15
  );


  not
  g44
  (
    n68,
    n1
  );


  not
  g45
  (
    n43,
    n10
  );


  not
  g46
  (
    n74,
    n1
  );


  not
  g47
  (
    n65,
    n18
  );


  buf
  g48
  (
    n60,
    n16
  );


  not
  g49
  (
    n26,
    n12
  );


  buf
  g50
  (
    n34,
    n5
  );


  buf
  g51
  (
    n35,
    n19
  );


  buf
  g52
  (
    n52,
    n15
  );


  buf
  g53
  (
    n78,
    n17
  );


  buf
  g54
  (
    n71,
    n7
  );


  buf
  g55
  (
    n31,
    n1
  );


  not
  g56
  (
    n61,
    n17
  );


  not
  g57
  (
    n36,
    n14
  );


  buf
  g58
  (
    n38,
    n1
  );


  buf
  g59
  (
    n87,
    n11
  );


  not
  g60
  (
    n41,
    n12
  );


  buf
  g61
  (
    n67,
    n11
  );


  not
  g62
  (
    n70,
    n3
  );


  not
  g63
  (
    n94,
    n10
  );


  buf
  g64
  (
    n96,
    n4
  );


  buf
  g65
  (
    n103,
    n18
  );


  buf
  g66
  (
    n39,
    n16
  );


  buf
  g67
  (
    n49,
    n11
  );


  not
  g68
  (
    n32,
    n10
  );


  not
  g69
  (
    n91,
    n16
  );


  not
  g70
  (
    n93,
    n20
  );


  not
  g71
  (
    n95,
    n13
  );


  not
  g72
  (
    n99,
    n2
  );


  not
  g73
  (
    n62,
    n7
  );


  buf
  g74
  (
    n58,
    n11
  );


  buf
  g75
  (
    n82,
    n20
  );


  buf
  g76
  (
    n80,
    n8
  );


  not
  g77
  (
    n69,
    n15
  );


  buf
  g78
  (
    n72,
    n10
  );


  buf
  g79
  (
    n56,
    n8
  );


  buf
  g80
  (
    n27,
    n6
  );


  buf
  g81
  (
    n330,
    n60
  );


  not
  g82
  (
    n410,
    n32
  );


  not
  g83
  (
    n411,
    n30
  );


  buf
  g84
  (
    n159,
    n36
  );


  not
  g85
  (
    n109,
    n81
  );


  buf
  g86
  (
    n336,
    n92
  );


  buf
  g87
  (
    n230,
    n36
  );


  not
  g88
  (
    n279,
    n45
  );


  buf
  g89
  (
    n254,
    n46
  );


  buf
  g90
  (
    n396,
    n43
  );


  buf
  g91
  (
    n133,
    n44
  );


  not
  g92
  (
    n340,
    n96
  );


  buf
  g93
  (
    n256,
    n90
  );


  buf
  g94
  (
    n343,
    n102
  );


  not
  g95
  (
    n223,
    n39
  );


  not
  g96
  (
    n124,
    n101
  );


  not
  g97
  (
    n320,
    n95
  );


  buf
  g98
  (
    n354,
    n49
  );


  buf
  g99
  (
    n355,
    n104
  );


  not
  g100
  (
    n307,
    n37
  );


  not
  g101
  (
    n260,
    n85
  );


  not
  g102
  (
    n383,
    n80
  );


  buf
  g103
  (
    n392,
    n104
  );


  buf
  g104
  (
    n333,
    n46
  );


  buf
  g105
  (
    n132,
    n94
  );


  not
  g106
  (
    n121,
    n95
  );


  buf
  g107
  (
    n128,
    n47
  );


  buf
  g108
  (
    n202,
    n50
  );


  buf
  g109
  (
    n306,
    n74
  );


  buf
  g110
  (
    n193,
    n90
  );


  not
  g111
  (
    n118,
    n47
  );


  buf
  g112
  (
    n135,
    n44
  );


  buf
  g113
  (
    n196,
    n99
  );


  buf
  g114
  (
    n273,
    n46
  );


  not
  g115
  (
    n235,
    n104
  );


  not
  g116
  (
    n155,
    n76
  );


  not
  g117
  (
    n368,
    n30
  );


  buf
  g118
  (
    n374,
    n66
  );


  not
  g119
  (
    n208,
    n40
  );


  not
  g120
  (
    n263,
    n81
  );


  not
  g121
  (
    n236,
    n86
  );


  not
  g122
  (
    n324,
    n71
  );


  buf
  g123
  (
    n421,
    n89
  );


  buf
  g124
  (
    n394,
    n44
  );


  not
  g125
  (
    n364,
    n43
  );


  not
  g126
  (
    n420,
    n82
  );


  buf
  g127
  (
    n348,
    n27
  );


  buf
  g128
  (
    n220,
    n63
  );


  buf
  g129
  (
    n422,
    n70
  );


  not
  g130
  (
    n325,
    n52
  );


  buf
  g131
  (
    n402,
    n77
  );


  not
  g132
  (
    n321,
    n50
  );


  buf
  g133
  (
    n184,
    n103
  );


  buf
  g134
  (
    n219,
    n54
  );


  not
  g135
  (
    n244,
    n56
  );


  not
  g136
  (
    n268,
    n88
  );


  buf
  g137
  (
    n391,
    n41
  );


  not
  g138
  (
    n186,
    n99
  );


  buf
  g139
  (
    n185,
    n35
  );


  buf
  g140
  (
    n406,
    n79
  );


  buf
  g141
  (
    n258,
    n58
  );


  buf
  g142
  (
    n141,
    n99
  );


  buf
  g143
  (
    n337,
    n78
  );


  buf
  g144
  (
    n351,
    n52
  );


  buf
  g145
  (
    n115,
    n64
  );


  buf
  g146
  (
    n416,
    n42
  );


  not
  g147
  (
    n366,
    n29
  );


  buf
  g148
  (
    n281,
    n75
  );


  buf
  g149
  (
    n180,
    n82
  );


  buf
  g150
  (
    n187,
    n77
  );


  not
  g151
  (
    n171,
    n89
  );


  buf
  g152
  (
    n267,
    n101
  );


  buf
  g153
  (
    n117,
    n70
  );


  not
  g154
  (
    n203,
    n77
  );


  not
  g155
  (
    n216,
    n80
  );


  buf
  g156
  (
    n127,
    n75
  );


  buf
  g157
  (
    n301,
    n49
  );


  not
  g158
  (
    n151,
    n61
  );


  buf
  g159
  (
    n309,
    n92
  );


  buf
  g160
  (
    KeyWire_0_4,
    n102
  );


  buf
  g161
  (
    n249,
    n97
  );


  not
  g162
  (
    n169,
    n96
  );


  buf
  g163
  (
    n362,
    n86
  );


  not
  g164
  (
    n125,
    n27
  );


  not
  g165
  (
    n298,
    n72
  );


  buf
  g166
  (
    n276,
    n67
  );


  not
  g167
  (
    n190,
    n96
  );


  not
  g168
  (
    n363,
    n66
  );


  buf
  g169
  (
    n404,
    n62
  );


  buf
  g170
  (
    n111,
    n63
  );


  buf
  g171
  (
    n382,
    n63
  );


  buf
  g172
  (
    n405,
    n92
  );


  buf
  g173
  (
    n138,
    n26
  );


  buf
  g174
  (
    n367,
    n53
  );


  not
  g175
  (
    n308,
    n42
  );


  not
  g176
  (
    n409,
    n87
  );


  not
  g177
  (
    n142,
    n28
  );


  buf
  g178
  (
    n126,
    n34
  );


  buf
  g179
  (
    n418,
    n44
  );


  buf
  g180
  (
    n311,
    n78
  );


  not
  g181
  (
    n250,
    n67
  );


  buf
  g182
  (
    n211,
    n47
  );


  buf
  g183
  (
    n120,
    n59
  );


  buf
  g184
  (
    n173,
    n104
  );


  not
  g185
  (
    n417,
    n33
  );


  buf
  g186
  (
    n357,
    n89
  );


  not
  g187
  (
    n174,
    n42
  );


  buf
  g188
  (
    n144,
    n31
  );


  buf
  g189
  (
    n261,
    n51
  );


  not
  g190
  (
    n122,
    n66
  );


  buf
  g191
  (
    n361,
    n77
  );


  buf
  g192
  (
    n365,
    n29
  );


  buf
  g193
  (
    n304,
    n31
  );


  not
  g194
  (
    n168,
    n48
  );


  not
  g195
  (
    n302,
    n59
  );


  not
  g196
  (
    n401,
    n76
  );


  buf
  g197
  (
    n188,
    n49
  );


  buf
  g198
  (
    n242,
    n37
  );


  not
  g199
  (
    n269,
    n60
  );


  buf
  g200
  (
    n257,
    n30
  );


  buf
  g201
  (
    n136,
    n37
  );


  not
  g202
  (
    n339,
    n38
  );


  buf
  g203
  (
    n240,
    n50
  );


  not
  g204
  (
    n214,
    n38
  );


  buf
  g205
  (
    n295,
    n55
  );


  buf
  g206
  (
    n114,
    n97
  );


  not
  g207
  (
    n403,
    n55
  );


  buf
  g208
  (
    n108,
    n64
  );


  not
  g209
  (
    n386,
    n79
  );


  not
  g210
  (
    n356,
    n86
  );


  not
  g211
  (
    n318,
    n81
  );


  buf
  g212
  (
    n177,
    n47
  );


  not
  g213
  (
    n119,
    n65
  );


  not
  g214
  (
    n413,
    n85
  );


  not
  g215
  (
    n226,
    n88
  );


  not
  g216
  (
    n253,
    n33
  );


  buf
  g217
  (
    n369,
    n73
  );


  buf
  g218
  (
    n234,
    n34
  );


  buf
  g219
  (
    n229,
    n33
  );


  buf
  g220
  (
    n389,
    n58
  );


  buf
  g221
  (
    n313,
    n84
  );


  not
  g222
  (
    n178,
    n90
  );


  not
  g223
  (
    n210,
    n70
  );


  buf
  g224
  (
    n205,
    n60
  );


  buf
  g225
  (
    n310,
    n60
  );


  buf
  g226
  (
    n189,
    n28
  );


  buf
  g227
  (
    n238,
    n83
  );


  not
  g228
  (
    n140,
    n76
  );


  buf
  g229
  (
    n329,
    n98
  );


  not
  g230
  (
    n378,
    n65
  );


  buf
  g231
  (
    n291,
    n102
  );


  buf
  g232
  (
    n283,
    n101
  );


  buf
  g233
  (
    n160,
    n45
  );


  not
  g234
  (
    n282,
    n29
  );


  buf
  g235
  (
    n312,
    n49
  );


  buf
  g236
  (
    n350,
    n32
  );


  buf
  g237
  (
    n342,
    n91
  );


  not
  g238
  (
    n262,
    n61
  );


  buf
  g239
  (
    n370,
    n88
  );


  buf
  g240
  (
    n259,
    n93
  );


  buf
  g241
  (
    n194,
    n29
  );


  not
  g242
  (
    n130,
    n62
  );


  buf
  g243
  (
    n204,
    n68
  );


  not
  g244
  (
    n266,
    n71
  );


  not
  g245
  (
    n233,
    n41
  );


  buf
  g246
  (
    n395,
    n68
  );


  buf
  g247
  (
    n264,
    n69
  );


  not
  g248
  (
    n148,
    n56
  );


  not
  g249
  (
    n349,
    n69
  );


  not
  g250
  (
    n317,
    n83
  );


  buf
  g251
  (
    n110,
    n53
  );


  not
  g252
  (
    n407,
    n74
  );


  buf
  g253
  (
    n289,
    n69
  );


  buf
  g254
  (
    n344,
    n64
  );


  buf
  g255
  (
    n326,
    n80
  );


  not
  g256
  (
    n284,
    n78
  );


  buf
  g257
  (
    n373,
    n28
  );


  not
  g258
  (
    n166,
    n32
  );


  buf
  g259
  (
    n172,
    n35
  );


  buf
  g260
  (
    n359,
    n68
  );


  not
  g261
  (
    n247,
    n96
  );


  not
  g262
  (
    n241,
    n57
  );


  buf
  g263
  (
    n332,
    n83
  );


  buf
  g264
  (
    n319,
    n64
  );


  buf
  g265
  (
    n143,
    n55
  );


  not
  g266
  (
    n314,
    n51
  );


  buf
  g267
  (
    n360,
    n85
  );


  buf
  g268
  (
    n248,
    n45
  );


  buf
  g269
  (
    n182,
    n56
  );


  buf
  g270
  (
    n290,
    n78
  );


  buf
  g271
  (
    n346,
    n35
  );


  not
  g272
  (
    n154,
    n54
  );


  buf
  g273
  (
    n408,
    n94
  );


  not
  g274
  (
    n165,
    n51
  );


  not
  g275
  (
    n293,
    n65
  );


  buf
  g276
  (
    n162,
    n98
  );


  buf
  g277
  (
    n251,
    n98
  );


  not
  g278
  (
    n224,
    n74
  );


  buf
  g279
  (
    n137,
    n54
  );


  not
  g280
  (
    n399,
    n100
  );


  buf
  g281
  (
    n227,
    n84
  );


  not
  g282
  (
    n419,
    n83
  );


  buf
  g283
  (
    n222,
    n61
  );


  not
  g284
  (
    n385,
    n70
  );


  not
  g285
  (
    n153,
    n102
  );


  not
  g286
  (
    n278,
    n100
  );


  not
  g287
  (
    n334,
    n73
  );


  buf
  g288
  (
    n287,
    n69
  );


  buf
  g289
  (
    n305,
    n46
  );


  not
  g290
  (
    n272,
    n36
  );


  not
  g291
  (
    n371,
    n95
  );


  buf
  g292
  (
    n175,
    n58
  );


  not
  g293
  (
    n200,
    n90
  );


  not
  g294
  (
    n397,
    n97
  );


  buf
  g295
  (
    n294,
    n52
  );


  buf
  g296
  (
    n280,
    n100
  );


  not
  g297
  (
    n335,
    n45
  );


  buf
  g298
  (
    n237,
    n42
  );


  not
  g299
  (
    n163,
    n84
  );


  buf
  g300
  (
    n331,
    n74
  );


  not
  g301
  (
    n167,
    n99
  );


  buf
  g302
  (
    n255,
    n38
  );


  buf
  g303
  (
    n415,
    n39
  );


  not
  g304
  (
    n164,
    n26
  );


  buf
  g305
  (
    n183,
    n73
  );


  not
  g306
  (
    n303,
    n27
  );


  not
  g307
  (
    n381,
    n57
  );


  not
  g308
  (
    n323,
    n65
  );


  not
  g309
  (
    n379,
    n91
  );


  buf
  g310
  (
    n412,
    n87
  );


  buf
  g311
  (
    n400,
    n56
  );


  buf
  g312
  (
    n372,
    n71
  );


  buf
  g313
  (
    n129,
    n89
  );


  not
  g314
  (
    n384,
    n75
  );


  buf
  g315
  (
    n112,
    n35
  );


  buf
  g316
  (
    n245,
    n75
  );


  buf
  g317
  (
    KeyWire_0_30,
    n63
  );


  not
  g318
  (
    n116,
    n43
  );


  buf
  g319
  (
    n288,
    n72
  );


  not
  g320
  (
    n286,
    n91
  );


  not
  g321
  (
    n158,
    n97
  );


  buf
  g322
  (
    n156,
    n54
  );


  buf
  g323
  (
    n265,
    n50
  );


  not
  g324
  (
    n231,
    n36
  );


  not
  g325
  (
    n145,
    n95
  );


  buf
  g326
  (
    n358,
    n68
  );


  not
  g327
  (
    n375,
    n103
  );


  buf
  g328
  (
    n297,
    n28
  );


  buf
  g329
  (
    n315,
    n48
  );


  not
  g330
  (
    n414,
    n66
  );


  buf
  g331
  (
    n218,
    n34
  );


  not
  g332
  (
    n192,
    n85
  );


  not
  g333
  (
    n191,
    n62
  );


  not
  g334
  (
    n274,
    n93
  );


  buf
  g335
  (
    n341,
    n87
  );


  buf
  g336
  (
    n207,
    n94
  );


  buf
  g337
  (
    n398,
    n61
  );


  not
  g338
  (
    n387,
    n55
  );


  not
  g339
  (
    n376,
    n38
  );


  not
  g340
  (
    n328,
    n58
  );


  buf
  g341
  (
    n139,
    n30
  );


  not
  g342
  (
    n179,
    n48
  );


  not
  g343
  (
    n345,
    n73
  );


  buf
  g344
  (
    n292,
    n67
  );


  not
  g345
  (
    n327,
    n98
  );


  buf
  g346
  (
    n149,
    n81
  );


  buf
  g347
  (
    n201,
    n59
  );


  not
  g348
  (
    n161,
    n41
  );


  not
  g349
  (
    n390,
    n51
  );


  buf
  g350
  (
    n146,
    n82
  );


  not
  g351
  (
    n107,
    n27
  );


  buf
  g352
  (
    n195,
    n62
  );


  not
  g353
  (
    n170,
    n79
  );


  not
  g354
  (
    n181,
    n52
  );


  not
  g355
  (
    n299,
    n37
  );


  not
  g356
  (
    n388,
    n72
  );


  buf
  g357
  (
    n232,
    n101
  );


  buf
  g358
  (
    n296,
    n67
  );


  buf
  g359
  (
    n217,
    n39
  );


  buf
  g360
  (
    n277,
    n79
  );


  buf
  g361
  (
    n197,
    n93
  );


  buf
  g362
  (
    n199,
    n86
  );


  not
  g363
  (
    n221,
    n41
  );


  not
  g364
  (
    n252,
    n40
  );


  not
  g365
  (
    n209,
    n92
  );


  not
  g366
  (
    n338,
    n34
  );


  not
  g367
  (
    n380,
    n57
  );


  not
  g368
  (
    n131,
    n59
  );


  buf
  g369
  (
    n134,
    n80
  );


  not
  g370
  (
    n150,
    n103
  );


  not
  g371
  (
    n215,
    n91
  );


  not
  g372
  (
    n157,
    n31
  );


  not
  g373
  (
    n147,
    n87
  );


  not
  g374
  (
    n347,
    n53
  );


  not
  g375
  (
    n352,
    n31
  );


  not
  g376
  (
    n228,
    n100
  );


  buf
  g377
  (
    n212,
    n43
  );


  buf
  g378
  (
    n316,
    n40
  );


  not
  g379
  (
    n243,
    n53
  );


  not
  g380
  (
    n152,
    n76
  );


  not
  g381
  (
    n246,
    n33
  );


  not
  g382
  (
    n271,
    n88
  );


  not
  g383
  (
    n300,
    n40
  );


  not
  g384
  (
    n322,
    n82
  );


  buf
  g385
  (
    n377,
    n94
  );


  not
  g386
  (
    n225,
    n32
  );


  buf
  g387
  (
    n113,
    n26
  );


  not
  g388
  (
    n176,
    n93
  );


  not
  g389
  (
    n353,
    n39
  );


  buf
  g390
  (
    n239,
    n71
  );


  not
  g391
  (
    n206,
    n72
  );


  not
  g392
  (
    n275,
    n26
  );


  not
  g393
  (
    n198,
    n84
  );


  not
  g394
  (
    n270,
    n48
  );


  not
  g395
  (
    n213,
    n57
  );


  not
  g396
  (
    n285,
    n103
  );


  not
  g397
  (
    n651,
    n303
  );


  not
  g398
  (
    n1268,
    n407
  );


  not
  g399
  (
    n1030,
    n240
  );


  not
  g400
  (
    n886,
    n151
  );


  not
  g401
  (
    n1204,
    n239
  );


  buf
  g402
  (
    n1128,
    n374
  );


  not
  g403
  (
    n1091,
    n174
  );


  buf
  g404
  (
    n1545,
    n392
  );


  buf
  g405
  (
    n798,
    n313
  );


  not
  g406
  (
    n1044,
    n252
  );


  not
  g407
  (
    n1616,
    n265
  );


  buf
  g408
  (
    n1640,
    n362
  );


  not
  g409
  (
    n1067,
    n404
  );


  not
  g410
  (
    n496,
    n202
  );


  not
  g411
  (
    n1312,
    n171
  );


  not
  g412
  (
    n1353,
    n421
  );


  not
  g413
  (
    n1038,
    n107
  );


  buf
  g414
  (
    n581,
    n142
  );


  not
  g415
  (
    n826,
    n238
  );


  not
  g416
  (
    n1025,
    n331
  );


  buf
  g417
  (
    n1114,
    n335
  );


  not
  g418
  (
    n1408,
    n419
  );


  not
  g419
  (
    n836,
    n383
  );


  not
  g420
  (
    n915,
    n397
  );


  buf
  g421
  (
    n674,
    n166
  );


  not
  g422
  (
    n440,
    n414
  );


  not
  g423
  (
    n1051,
    n218
  );


  buf
  g424
  (
    n1306,
    n171
  );


  not
  g425
  (
    n1130,
    n140
  );


  not
  g426
  (
    n1646,
    n217
  );


  buf
  g427
  (
    n1533,
    n321
  );


  buf
  g428
  (
    n1496,
    n163
  );


  buf
  g429
  (
    n788,
    n196
  );


  buf
  g430
  (
    n525,
    n177
  );


  not
  g431
  (
    n743,
    n253
  );


  buf
  g432
  (
    n438,
    n346
  );


  buf
  g433
  (
    n458,
    n333
  );


  not
  g434
  (
    n775,
    n379
  );


  not
  g435
  (
    n617,
    n294
  );


  buf
  g436
  (
    n1278,
    n185
  );


  not
  g437
  (
    n1056,
    n390
  );


  not
  g438
  (
    n938,
    n337
  );


  buf
  g439
  (
    n1052,
    n359
  );


  buf
  g440
  (
    n570,
    n404
  );


  not
  g441
  (
    n1347,
    n367
  );


  not
  g442
  (
    n907,
    n348
  );


  not
  g443
  (
    n1265,
    n161
  );


  buf
  g444
  (
    n1614,
    n223
  );


  buf
  g445
  (
    n999,
    n187
  );


  buf
  g446
  (
    n1293,
    n157
  );


  not
  g447
  (
    n1491,
    n220
  );


  buf
  g448
  (
    n538,
    n211
  );


  not
  g449
  (
    n585,
    n322
  );


  buf
  g450
  (
    n903,
    n145
  );


  buf
  g451
  (
    n1003,
    n351
  );


  not
  g452
  (
    n1463,
    n277
  );


  buf
  g453
  (
    n1097,
    n347
  );


  buf
  g454
  (
    n856,
    n299
  );


  not
  g455
  (
    n1156,
    n193
  );


  buf
  g456
  (
    n1064,
    n410
  );


  buf
  g457
  (
    n771,
    n184
  );


  buf
  g458
  (
    n567,
    n228
  );


  buf
  g459
  (
    n919,
    n395
  );


  buf
  g460
  (
    n709,
    n255
  );


  not
  g461
  (
    n1193,
    n280
  );


  not
  g462
  (
    n1512,
    n284
  );


  buf
  g463
  (
    n1477,
    n250
  );


  not
  g464
  (
    n1604,
    n351
  );


  not
  g465
  (
    n1664,
    n301
  );


  not
  g466
  (
    n618,
    n355
  );


  buf
  g467
  (
    n573,
    n170
  );


  buf
  g468
  (
    n1569,
    n134
  );


  buf
  g469
  (
    n1652,
    n310
  );


  buf
  g470
  (
    n610,
    n170
  );


  buf
  g471
  (
    n1279,
    n198
  );


  buf
  g472
  (
    n1162,
    n197
  );


  not
  g473
  (
    n1473,
    n316
  );


  buf
  g474
  (
    n1682,
    n247
  );


  buf
  g475
  (
    n833,
    n131
  );


  not
  g476
  (
    n1553,
    n416
  );


  buf
  g477
  (
    n1529,
    n225
  );


  not
  g478
  (
    n435,
    n300
  );


  buf
  g479
  (
    n1430,
    n380
  );


  buf
  g480
  (
    n888,
    n384
  );


  not
  g481
  (
    n948,
    n162
  );


  buf
  g482
  (
    n757,
    n116
  );


  buf
  g483
  (
    n582,
    n288
  );


  buf
  g484
  (
    n1208,
    n386
  );


  not
  g485
  (
    n443,
    n270
  );


  not
  g486
  (
    n1191,
    n293
  );


  buf
  g487
  (
    n656,
    n365
  );


  not
  g488
  (
    n866,
    n173
  );


  buf
  g489
  (
    n859,
    n267
  );


  buf
  g490
  (
    n428,
    n123
  );


  not
  g491
  (
    n1339,
    n360
  );


  buf
  g492
  (
    n1543,
    n222
  );


  not
  g493
  (
    n1550,
    n401
  );


  not
  g494
  (
    n1078,
    n189
  );


  buf
  g495
  (
    n1443,
    n261
  );


  buf
  g496
  (
    n1133,
    n114
  );


  buf
  g497
  (
    n801,
    n379
  );


  buf
  g498
  (
    n532,
    n307
  );


  not
  g499
  (
    n621,
    n376
  );


  not
  g500
  (
    n1547,
    n185
  );


  buf
  g501
  (
    n1615,
    n265
  );


  not
  g502
  (
    n1027,
    n301
  );


  buf
  g503
  (
    n1618,
    n282
  );


  buf
  g504
  (
    n764,
    n143
  );


  buf
  g505
  (
    n1358,
    n200
  );


  not
  g506
  (
    n1561,
    n395
  );


  buf
  g507
  (
    n624,
    n224
  );


  not
  g508
  (
    n756,
    n241
  );


  not
  g509
  (
    n1313,
    n378
  );


  not
  g510
  (
    n1062,
    n124
  );


  buf
  g511
  (
    n975,
    n164
  );


  not
  g512
  (
    n639,
    n107
  );


  not
  g513
  (
    n664,
    n279
  );


  not
  g514
  (
    n1511,
    n258
  );


  buf
  g515
  (
    n1404,
    n357
  );


  buf
  g516
  (
    n1612,
    n160
  );


  buf
  g517
  (
    n1518,
    n264
  );


  not
  g518
  (
    n831,
    n209
  );


  not
  g519
  (
    n569,
    n385
  );


  not
  g520
  (
    n1623,
    n392
  );


  buf
  g521
  (
    n1455,
    n325
  );


  buf
  g522
  (
    n1231,
    n205
  );


  not
  g523
  (
    n998,
    n268
  );


  buf
  g524
  (
    n1548,
    n175
  );


  not
  g525
  (
    n464,
    n314
  );


  buf
  g526
  (
    n1377,
    n274
  );


  not
  g527
  (
    n712,
    n371
  );


  buf
  g528
  (
    n1402,
    n192
  );


  buf
  g529
  (
    n1409,
    n252
  );


  buf
  g530
  (
    n970,
    n307
  );


  not
  g531
  (
    n901,
    n165
  );


  buf
  g532
  (
    n1461,
    n202
  );


  buf
  g533
  (
    n657,
    n308
  );


  not
  g534
  (
    n462,
    n197
  );


  buf
  g535
  (
    n916,
    n236
  );


  not
  g536
  (
    n855,
    n286
  );


  not
  g537
  (
    n439,
    n312
  );


  not
  g538
  (
    n746,
    n248
  );


  buf
  g539
  (
    n1144,
    n261
  );


  buf
  g540
  (
    n1571,
    n333
  );


  not
  g541
  (
    KeyWire_0_28,
    n299
  );


  not
  g542
  (
    n1656,
    n268
  );


  buf
  g543
  (
    n549,
    n133
  );


  not
  g544
  (
    n1609,
    n109
  );


  buf
  g545
  (
    n1648,
    n229
  );


  not
  g546
  (
    n1601,
    n239
  );


  buf
  g547
  (
    n1307,
    n361
  );


  not
  g548
  (
    n1223,
    n335
  );


  not
  g549
  (
    n542,
    n269
  );


  not
  g550
  (
    n1387,
    n288
  );


  not
  g551
  (
    n739,
    n326
  );


  buf
  g552
  (
    n981,
    n359
  );


  buf
  g553
  (
    n1102,
    n317
  );


  buf
  g554
  (
    n1633,
    n340
  );


  not
  g555
  (
    n1600,
    n410
  );


  buf
  g556
  (
    n1281,
    n416
  );


  buf
  g557
  (
    n780,
    n224
  );


  buf
  g558
  (
    n620,
    n417
  );


  buf
  g559
  (
    n1292,
    n321
  );


  not
  g560
  (
    n654,
    n421
  );


  not
  g561
  (
    n1254,
    n374
  );


  buf
  g562
  (
    n1126,
    n366
  );


  buf
  g563
  (
    n1369,
    n117
  );


  buf
  g564
  (
    n425,
    n283
  );


  not
  g565
  (
    n1450,
    n181
  );


  not
  g566
  (
    n1579,
    n374
  );


  buf
  g567
  (
    n1636,
    n233
  );


  not
  g568
  (
    n518,
    n405
  );


  buf
  g569
  (
    n1673,
    n385
  );


  buf
  g570
  (
    n666,
    n406
  );


  buf
  g571
  (
    n744,
    n270
  );


  not
  g572
  (
    n619,
    n125
  );


  not
  g573
  (
    n544,
    n177
  );


  not
  g574
  (
    n734,
    n248
  );


  buf
  g575
  (
    n1232,
    n419
  );


  not
  g576
  (
    n885,
    n227
  );


  not
  g577
  (
    n1419,
    n164
  );


  not
  g578
  (
    n467,
    n375
  );


  not
  g579
  (
    n1457,
    n259
  );


  not
  g580
  (
    n471,
    n114
  );


  not
  g581
  (
    n973,
    n195
  );


  buf
  g582
  (
    n1053,
    n128
  );


  not
  g583
  (
    n1414,
    n300
  );


  not
  g584
  (
    n1163,
    n378
  );


  not
  g585
  (
    n1176,
    n293
  );


  buf
  g586
  (
    n936,
    n348
  );


  not
  g587
  (
    n1017,
    n208
  );


  buf
  g588
  (
    n1494,
    n236
  );


  buf
  g589
  (
    n1077,
    n240
  );


  buf
  g590
  (
    n926,
    n108
  );


  buf
  g591
  (
    n1207,
    n417
  );


  buf
  g592
  (
    n632,
    n378
  );


  buf
  g593
  (
    n784,
    n405
  );


  buf
  g594
  (
    n1337,
    n210
  );


  buf
  g595
  (
    n1345,
    n169
  );


  buf
  g596
  (
    n1079,
    n201
  );


  buf
  g597
  (
    n898,
    n275
  );


  buf
  g598
  (
    n884,
    n207
  );


  buf
  g599
  (
    n1523,
    n377
  );


  buf
  g600
  (
    n495,
    n253
  );


  buf
  g601
  (
    n956,
    n337
  );


  buf
  g602
  (
    n1197,
    n176
  );


  not
  g603
  (
    n1563,
    n339
  );


  buf
  g604
  (
    n929,
    n163
  );


  buf
  g605
  (
    n1214,
    n120
  );


  not
  g606
  (
    n1624,
    n388
  );


  buf
  g607
  (
    n1593,
    n365
  );


  buf
  g608
  (
    n1532,
    n206
  );


  buf
  g609
  (
    n676,
    n358
  );


  not
  g610
  (
    n1297,
    n314
  );


  not
  g611
  (
    n1684,
    n213
  );


  buf
  g612
  (
    n672,
    n243
  );


  buf
  g613
  (
    n1479,
    n308
  );


  buf
  g614
  (
    n670,
    n344
  );


  not
  g615
  (
    n1177,
    n377
  );


  not
  g616
  (
    n1088,
    n246
  );


  buf
  g617
  (
    n1249,
    n241
  );


  not
  g618
  (
    n700,
    n133
  );


  buf
  g619
  (
    n953,
    n389
  );


  not
  g620
  (
    n993,
    n195
  );


  not
  g621
  (
    n842,
    n277
  );


  not
  g622
  (
    n485,
    n236
  );


  buf
  g623
  (
    n810,
    n269
  );


  not
  g624
  (
    n1354,
    n115
  );


  not
  g625
  (
    n1334,
    n269
  );


  not
  g626
  (
    n447,
    n258
  );


  not
  g627
  (
    n1273,
    n282
  );


  not
  g628
  (
    n1438,
    n232
  );


  buf
  g629
  (
    n730,
    n136
  );


  buf
  g630
  (
    n942,
    n110
  );


  buf
  g631
  (
    n1662,
    n216
  );


  buf
  g632
  (
    n694,
    n415
  );


  not
  g633
  (
    n701,
    n310
  );


  buf
  g634
  (
    n1350,
    n411
  );


  buf
  g635
  (
    n851,
    n236
  );


  not
  g636
  (
    n850,
    n247
  );


  buf
  g637
  (
    n1597,
    n139
  );


  not
  g638
  (
    n590,
    n365
  );


  buf
  g639
  (
    n1186,
    n346
  );


  buf
  g640
  (
    n649,
    n120
  );


  buf
  g641
  (
    n1531,
    n407
  );


  buf
  g642
  (
    n1021,
    n323
  );


  not
  g643
  (
    n1008,
    n414
  );


  not
  g644
  (
    n1653,
    n400
  );


  buf
  g645
  (
    n655,
    n394
  );


  buf
  g646
  (
    n1175,
    n353
  );


  buf
  g647
  (
    n1514,
    n413
  );


  not
  g648
  (
    n1014,
    n110
  );


  not
  g649
  (
    n691,
    n112
  );


  not
  g650
  (
    n605,
    n203
  );


  not
  g651
  (
    n935,
    n204
  );


  not
  g652
  (
    n1433,
    n118
  );


  not
  g653
  (
    n738,
    n363
  );


  not
  g654
  (
    n1449,
    n279
  );


  not
  g655
  (
    n545,
    n180
  );


  buf
  g656
  (
    n586,
    n353
  );


  not
  g657
  (
    n1559,
    n158
  );


  buf
  g658
  (
    n943,
    n284
  );


  not
  g659
  (
    n1210,
    n146
  );


  buf
  g660
  (
    n1356,
    n233
  );


  buf
  g661
  (
    n1309,
    n320
  );


  buf
  g662
  (
    n1539,
    n206
  );


  buf
  g663
  (
    n1493,
    n372
  );


  not
  g664
  (
    n494,
    n209
  );


  buf
  g665
  (
    n1229,
    n364
  );


  buf
  g666
  (
    n722,
    n131
  );


  buf
  g667
  (
    n1431,
    n297
  );


  not
  g668
  (
    n524,
    n110
  );


  not
  g669
  (
    n1454,
    n317
  );


  not
  g670
  (
    n949,
    n353
  );


  buf
  g671
  (
    n865,
    n227
  );


  not
  g672
  (
    n977,
    n276
  );


  buf
  g673
  (
    n1280,
    n276
  );


  not
  g674
  (
    n768,
    n179
  );


  not
  g675
  (
    n1425,
    n201
  );


  not
  g676
  (
    n1002,
    n134
  );


  buf
  g677
  (
    n776,
    n235
  );


  buf
  g678
  (
    n578,
    n221
  );


  not
  g679
  (
    n1150,
    n237
  );


  not
  g680
  (
    n1073,
    n378
  );


  buf
  g681
  (
    n1226,
    n167
  );


  not
  g682
  (
    n1271,
    n128
  );


  not
  g683
  (
    n1023,
    n418
  );


  buf
  g684
  (
    n767,
    n168
  );


  not
  g685
  (
    n719,
    n156
  );


  not
  g686
  (
    n832,
    n109
  );


  buf
  g687
  (
    n520,
    n108
  );


  not
  g688
  (
    n1360,
    n198
  );


  not
  g689
  (
    n910,
    n335
  );


  not
  g690
  (
    n614,
    n161
  );


  not
  g691
  (
    n733,
    n362
  );


  not
  g692
  (
    n1185,
    n286
  );


  not
  g693
  (
    n1215,
    n111
  );


  buf
  g694
  (
    n1372,
    n209
  );


  not
  g695
  (
    n822,
    n237
  );


  buf
  g696
  (
    n1534,
    n380
  );


  buf
  g697
  (
    n1109,
    n406
  );


  buf
  g698
  (
    n1098,
    n350
  );


  buf
  g699
  (
    n1211,
    n290
  );


  buf
  g700
  (
    n952,
    n366
  );


  buf
  g701
  (
    n976,
    n370
  );


  not
  g702
  (
    n1535,
    n259
  );


  buf
  g703
  (
    n627,
    n143
  );


  not
  g704
  (
    n1467,
    n319
  );


  buf
  g705
  (
    n1040,
    n313
  );


  buf
  g706
  (
    n1359,
    n112
  );


  buf
  g707
  (
    n747,
    n387
  );


  not
  g708
  (
    n1606,
    n163
  );


  buf
  g709
  (
    n1300,
    n326
  );


  buf
  g710
  (
    n1287,
    n258
  );


  buf
  g711
  (
    n1391,
    n413
  );


  not
  g712
  (
    n1244,
    n206
  );


  not
  g713
  (
    n1024,
    n303
  );


  not
  g714
  (
    n1448,
    n403
  );


  buf
  g715
  (
    n1240,
    n251
  );


  not
  g716
  (
    n1367,
    n205
  );


  not
  g717
  (
    n553,
    n222
  );


  buf
  g718
  (
    n516,
    n256
  );


  buf
  g719
  (
    n1153,
    n252
  );


  buf
  g720
  (
    n1355,
    n247
  );


  not
  g721
  (
    n1295,
    n173
  );


  buf
  g722
  (
    n482,
    n207
  );


  buf
  g723
  (
    n1198,
    n373
  );


  buf
  g724
  (
    n1217,
    n125
  );


  not
  g725
  (
    n896,
    n308
  );


  not
  g726
  (
    n491,
    n157
  );


  not
  g727
  (
    n797,
    n255
  );


  buf
  g728
  (
    n1299,
    n284
  );


  buf
  g729
  (
    n772,
    n191
  );


  buf
  g730
  (
    n1241,
    n249
  );


  buf
  g731
  (
    n1131,
    n395
  );


  not
  g732
  (
    n1421,
    n194
  );


  not
  g733
  (
    n1000,
    n393
  );


  buf
  g734
  (
    n880,
    n152
  );


  not
  g735
  (
    n1283,
    n259
  );


  buf
  g736
  (
    n1630,
    n382
  );


  buf
  g737
  (
    n720,
    n330
  );


  not
  g738
  (
    n668,
    n200
  );


  buf
  g739
  (
    n1272,
    n415
  );


  not
  g740
  (
    n870,
    n355
  );


  not
  g741
  (
    n1092,
    n324
  );


  buf
  g742
  (
    n1143,
    n389
  );


  not
  g743
  (
    n1351,
    n204
  );


  not
  g744
  (
    n450,
    n167
  );


  not
  g745
  (
    n812,
    n172
  );


  not
  g746
  (
    n761,
    n158
  );


  buf
  g747
  (
    n459,
    n134
  );


  not
  g748
  (
    n890,
    n145
  );


  buf
  g749
  (
    n1440,
    n292
  );


  not
  g750
  (
    n827,
    n272
  );


  not
  g751
  (
    n1558,
    n213
  );


  buf
  g752
  (
    n1298,
    n399
  );


  not
  g753
  (
    n1034,
    n245
  );


  not
  g754
  (
    n522,
    n114
  );


  not
  g755
  (
    n579,
    n336
  );


  not
  g756
  (
    n873,
    n262
  );


  buf
  g757
  (
    n1598,
    n295
  );


  not
  g758
  (
    n1196,
    n342
  );


  not
  g759
  (
    n1517,
    n294
  );


  buf
  g760
  (
    n1560,
    n261
  );


  not
  g761
  (
    n457,
    n395
  );


  buf
  g762
  (
    n882,
    n307
  );


  not
  g763
  (
    n592,
    n317
  );


  buf
  g764
  (
    n1666,
    n295
  );


  not
  g765
  (
    n1058,
    n363
  );


  not
  g766
  (
    n714,
    n380
  );


  buf
  g767
  (
    n1480,
    n242
  );


  buf
  g768
  (
    n741,
    n108
  );


  buf
  g769
  (
    n1031,
    n140
  );


  not
  g770
  (
    n1575,
    n192
  );


  not
  g771
  (
    n692,
    n152
  );


  buf
  g772
  (
    n1263,
    n408
  );


  not
  g773
  (
    n785,
    n371
  );


  buf
  g774
  (
    n1610,
    n256
  );


  buf
  g775
  (
    n753,
    n413
  );


  buf
  g776
  (
    n1371,
    n366
  );


  buf
  g777
  (
    n779,
    n150
  );


  not
  g778
  (
    n623,
    n285
  );


  not
  g779
  (
    n951,
    n214
  );


  not
  g780
  (
    n1202,
    n229
  );


  not
  g781
  (
    n1234,
    n265
  );


  buf
  g782
  (
    n1066,
    n142
  );


  not
  g783
  (
    n642,
    n190
  );


  buf
  g784
  (
    n1582,
    n153
  );


  not
  g785
  (
    n807,
    n183
  );


  not
  g786
  (
    n823,
    n198
  );


  buf
  g787
  (
    n960,
    n119
  );


  not
  g788
  (
    n511,
    n183
  );


  not
  g789
  (
    n726,
    n352
  );


  not
  g790
  (
    n1602,
    n306
  );


  not
  g791
  (
    n1503,
    n186
  );


  buf
  g792
  (
    n690,
    n138
  );


  not
  g793
  (
    n905,
    n162
  );


  not
  g794
  (
    n1645,
    n393
  );


  buf
  g795
  (
    n1206,
    n401
  );


  not
  g796
  (
    n737,
    n274
  );


  not
  g797
  (
    n1256,
    n180
  );


  not
  g798
  (
    n446,
    n316
  );


  not
  g799
  (
    n1108,
    n157
  );


  buf
  g800
  (
    n1568,
    n205
  );


  buf
  g801
  (
    n1199,
    n110
  );


  buf
  g802
  (
    n503,
    n296
  );


  not
  g803
  (
    n1227,
    n314
  );


  not
  g804
  (
    n631,
    n344
  );


  not
  g805
  (
    n1070,
    n219
  );


  not
  g806
  (
    n868,
    n147
  );


  not
  g807
  (
    n1622,
    n353
  );


  buf
  g808
  (
    n748,
    n396
  );


  not
  g809
  (
    n510,
    n324
  );


  buf
  g810
  (
    n1412,
    n359
  );


  not
  g811
  (
    n1305,
    n329
  );


  buf
  g812
  (
    n429,
    n266
  );


  buf
  g813
  (
    n887,
    n152
  );


  buf
  g814
  (
    n1389,
    n234
  );


  not
  g815
  (
    n1237,
    n203
  );


  buf
  g816
  (
    n1519,
    n122
  );


  not
  g817
  (
    n628,
    n223
  );


  buf
  g818
  (
    n895,
    n160
  );


  buf
  g819
  (
    n1142,
    n199
  );


  not
  g820
  (
    n1022,
    n364
  );


  not
  g821
  (
    n1145,
    n373
  );


  buf
  g822
  (
    n1410,
    n390
  );


  buf
  g823
  (
    n1260,
    n244
  );


  not
  g824
  (
    n892,
    n418
  );


  buf
  g825
  (
    n878,
    n229
  );


  not
  g826
  (
    n1498,
    n183
  );


  buf
  g827
  (
    n1669,
    n419
  );


  not
  g828
  (
    n616,
    n391
  );


  buf
  g829
  (
    n505,
    n308
  );


  not
  g830
  (
    n1190,
    n313
  );


  not
  g831
  (
    n1269,
    n369
  );


  buf
  g832
  (
    n922,
    n150
  );


  buf
  g833
  (
    n1047,
    n309
  );


  buf
  g834
  (
    n1469,
    n119
  );


  buf
  g835
  (
    n1405,
    n126
  );


  not
  g836
  (
    n436,
    n185
  );


  buf
  g837
  (
    n1524,
    n277
  );


  buf
  g838
  (
    n652,
    n318
  );


  not
  g839
  (
    n1643,
    n334
  );


  not
  g840
  (
    n609,
    n243
  );


  not
  g841
  (
    n1546,
    n188
  );


  not
  g842
  (
    n728,
    n259
  );


  buf
  g843
  (
    n556,
    n216
  );


  not
  g844
  (
    n736,
    n318
  );


  buf
  g845
  (
    n1654,
    n220
  );


  not
  g846
  (
    n1658,
    n412
  );


  not
  g847
  (
    n663,
    n363
  );


  not
  g848
  (
    n1119,
    n188
  );


  buf
  g849
  (
    n1344,
    n398
  );


  buf
  g850
  (
    n717,
    n396
  );


  buf
  g851
  (
    n693,
    n165
  );


  buf
  g852
  (
    n1382,
    n190
  );


  buf
  g853
  (
    n897,
    n339
  );


  buf
  g854
  (
    n466,
    n172
  );


  not
  g855
  (
    n486,
    n257
  );


  not
  g856
  (
    n562,
    n389
  );


  not
  g857
  (
    n945,
    n107
  );


  not
  g858
  (
    n531,
    n135
  );


  buf
  g859
  (
    n1671,
    n372
  );


  buf
  g860
  (
    n937,
    n177
  );


  not
  g861
  (
    n724,
    n329
  );


  not
  g862
  (
    n608,
    n412
  );


  buf
  g863
  (
    n1608,
    n421
  );


  buf
  g864
  (
    KeyWire_0_21,
    n253
  );


  buf
  g865
  (
    n997,
    n238
  );


  not
  g866
  (
    n962,
    n407
  );


  buf
  g867
  (
    n1581,
    n255
  );


  buf
  g868
  (
    n644,
    n139
  );


  buf
  g869
  (
    n790,
    n194
  );


  not
  g870
  (
    n1333,
    n286
  );


  not
  g871
  (
    n1500,
    n147
  );


  buf
  g872
  (
    n1557,
    n180
  );


  buf
  g873
  (
    n1054,
    n291
  );


  not
  g874
  (
    n1378,
    n343
  );


  not
  g875
  (
    n571,
    n168
  );


  not
  g876
  (
    n643,
    n243
  );


  buf
  g877
  (
    n584,
    n345
  );


  not
  g878
  (
    n983,
    n169
  );


  buf
  g879
  (
    n455,
    n319
  );


  not
  g880
  (
    n1587,
    n138
  );


  not
  g881
  (
    n1200,
    n220
  );


  not
  g882
  (
    n704,
    n340
  );


  buf
  g883
  (
    n1248,
    n328
  );


  buf
  g884
  (
    n667,
    n176
  );


  not
  g885
  (
    n1501,
    n211
  );


  not
  g886
  (
    n1173,
    n350
  );


  not
  g887
  (
    n982,
    n151
  );


  not
  g888
  (
    n1046,
    n149
  );


  buf
  g889
  (
    n665,
    n302
  );


  buf
  g890
  (
    n1154,
    n372
  );


  not
  g891
  (
    n1107,
    n175
  );


  not
  g892
  (
    n1452,
    n398
  );


  buf
  g893
  (
    n561,
    n154
  );


  not
  g894
  (
    n1082,
    n210
  );


  not
  g895
  (
    n1506,
    n300
  );


  buf
  g896
  (
    n611,
    n121
  );


  buf
  g897
  (
    n874,
    n333
  );


  buf
  g898
  (
    n1386,
    n315
  );


  buf
  g899
  (
    n474,
    n164
  );


  not
  g900
  (
    n1168,
    n324
  );


  buf
  g901
  (
    n1286,
    n276
  );


  not
  g902
  (
    n1605,
    n323
  );


  buf
  g903
  (
    n735,
    n210
  );


  buf
  g904
  (
    n1444,
    n219
  );


  buf
  g905
  (
    n1084,
    n119
  );


  buf
  g906
  (
    n1507,
    n332
  );


  buf
  g907
  (
    n1069,
    n418
  );


  buf
  g908
  (
    n1617,
    n119
  );


  not
  g909
  (
    n540,
    n303
  );


  not
  g910
  (
    n1613,
    n351
  );


  not
  g911
  (
    n1460,
    n296
  );


  not
  g912
  (
    n1564,
    n306
  );


  not
  g913
  (
    n1267,
    n154
  );


  buf
  g914
  (
    n1028,
    n218
  );


  not
  g915
  (
    n658,
    n144
  );


  not
  g916
  (
    n526,
    n283
  );


  buf
  g917
  (
    n671,
    n260
  );


  buf
  g918
  (
    n1018,
    n265
  );


  buf
  g919
  (
    n1399,
    n346
  );


  not
  g920
  (
    n599,
    n137
  );


  buf
  g921
  (
    n917,
    n143
  );


  buf
  g922
  (
    n1415,
    n337
  );


  not
  g923
  (
    n1158,
    n356
  );


  buf
  g924
  (
    KeyWire_0_17,
    n141
  );


  buf
  g925
  (
    n819,
    n198
  );


  buf
  g926
  (
    n1001,
    n127
  );


  not
  g927
  (
    n1488,
    n144
  );


  not
  g928
  (
    n751,
    n138
  );


  not
  g929
  (
    n1549,
    n248
  );


  not
  g930
  (
    n1160,
    n289
  );


  not
  g931
  (
    n1187,
    n174
  );


  not
  g932
  (
    n1422,
    n354
  );


  not
  g933
  (
    n995,
    n148
  );


  not
  g934
  (
    n933,
    n135
  );


  not
  g935
  (
    n1129,
    n254
  );


  not
  g936
  (
    n1179,
    n183
  );


  not
  g937
  (
    n1426,
    n133
  );


  buf
  g938
  (
    n1105,
    n123
  );


  not
  g939
  (
    n899,
    n332
  );


  buf
  g940
  (
    n1236,
    n270
  );


  not
  g941
  (
    n488,
    n379
  );


  not
  g942
  (
    n793,
    n212
  );


  not
  g943
  (
    n845,
    n375
  );


  buf
  g944
  (
    n876,
    n158
  );


  not
  g945
  (
    n820,
    n264
  );


  not
  g946
  (
    n1420,
    n297
  );


  not
  g947
  (
    n1435,
    n397
  );


  buf
  g948
  (
    n990,
    n294
  );


  not
  g949
  (
    n1577,
    n281
  );


  not
  g950
  (
    n1192,
    n381
  );


  not
  g951
  (
    n843,
    n213
  );


  buf
  g952
  (
    n1651,
    n384
  );


  not
  g953
  (
    n1112,
    n368
  );


  not
  g954
  (
    n430,
    n318
  );


  buf
  g955
  (
    n706,
    n288
  );


  buf
  g956
  (
    n1320,
    n200
  );


  not
  g957
  (
    n1655,
    n239
  );


  buf
  g958
  (
    n1036,
    n360
  );


  not
  g959
  (
    n799,
    n345
  );


  buf
  g960
  (
    n1282,
    n297
  );


  not
  g961
  (
    n858,
    n381
  );


  not
  g962
  (
    n760,
    n208
  );


  not
  g963
  (
    n1570,
    n287
  );


  not
  g964
  (
    n1417,
    n362
  );


  not
  g965
  (
    n763,
    n332
  );


  not
  g966
  (
    n1049,
    n367
  );


  not
  g967
  (
    n1159,
    n120
  );


  buf
  g968
  (
    n437,
    n234
  );


  buf
  g969
  (
    n1311,
    n331
  );


  buf
  g970
  (
    n992,
    n230
  );


  not
  g971
  (
    n925,
    n412
  );


  not
  g972
  (
    n1484,
    n398
  );


  buf
  g973
  (
    n1619,
    n392
  );


  not
  g974
  (
    n1060,
    n310
  );


  not
  g975
  (
    n1352,
    n369
  );


  not
  g976
  (
    n1537,
    n331
  );


  buf
  g977
  (
    n1584,
    n382
  );


  not
  g978
  (
    n1328,
    n342
  );


  buf
  g979
  (
    n1376,
    n388
  );


  not
  g980
  (
    n504,
    n360
  );


  not
  g981
  (
    n1310,
    n271
  );


  buf
  g982
  (
    n1665,
    n408
  );


  not
  g983
  (
    n479,
    n270
  );


  buf
  g984
  (
    n808,
    n152
  );


  buf
  g985
  (
    n750,
    n126
  );


  buf
  g986
  (
    n475,
    n153
  );


  not
  g987
  (
    n1057,
    n279
  );


  buf
  g988
  (
    n1111,
    n137
  );


  not
  g989
  (
    n635,
    n250
  );


  not
  g990
  (
    n1331,
    n386
  );


  buf
  g991
  (
    n1674,
    n170
  );


  buf
  g992
  (
    n835,
    n402
  );


  not
  g993
  (
    n1627,
    n411
  );


  buf
  g994
  (
    n1330,
    n316
  );


  buf
  g995
  (
    n1657,
    n182
  );


  buf
  g996
  (
    n1148,
    n364
  );


  not
  g997
  (
    n1370,
    n333
  );


  buf
  g998
  (
    n1125,
    n294
  );


  buf
  g999
  (
    n955,
    n320
  );


  buf
  g1000
  (
    n1416,
    n342
  );


  not
  g1001
  (
    n1515,
    n289
  );


  not
  g1002
  (
    n1221,
    n260
  );


  not
  g1003
  (
    n1659,
    n189
  );


  not
  g1004
  (
    n1045,
    n201
  );


  buf
  g1005
  (
    n770,
    n317
  );


  not
  g1006
  (
    n492,
    n370
  );


  buf
  g1007
  (
    n782,
    n175
  );


  not
  g1008
  (
    n1670,
    n121
  );


  buf
  g1009
  (
    n521,
    n242
  );


  buf
  g1010
  (
    n931,
    n376
  );


  not
  g1011
  (
    n848,
    n387
  );


  not
  g1012
  (
    n918,
    n153
  );


  not
  g1013
  (
    n773,
    n136
  );


  not
  g1014
  (
    n547,
    n131
  );


  buf
  g1015
  (
    n580,
    n336
  );


  not
  g1016
  (
    n791,
    n336
  );


  not
  g1017
  (
    n424,
    n107
  );


  not
  g1018
  (
    KeyWire_0_6,
    n304
  );


  not
  g1019
  (
    n978,
    n146
  );


  not
  g1020
  (
    n991,
    n379
  );


  not
  g1021
  (
    n685,
    n136
  );


  not
  g1022
  (
    n1122,
    n338
  );


  not
  g1023
  (
    n1458,
    n141
  );


  not
  g1024
  (
    n431,
    n129
  );


  buf
  g1025
  (
    n1242,
    n228
  );


  buf
  g1026
  (
    n1124,
    n281
  );


  not
  g1027
  (
    n1315,
    n272
  );


  buf
  g1028
  (
    n1403,
    n229
  );


  buf
  g1029
  (
    n1401,
    n394
  );


  buf
  g1030
  (
    n1274,
    n320
  );


  not
  g1031
  (
    n1135,
    n400
  );


  buf
  g1032
  (
    n441,
    n422
  );


  buf
  g1033
  (
    n1341,
    n288
  );


  buf
  g1034
  (
    n1323,
    n128
  );


  not
  g1035
  (
    n1629,
    n422
  );


  not
  g1036
  (
    n984,
    n278
  );


  not
  g1037
  (
    n857,
    n289
  );


  not
  g1038
  (
    n1411,
    n122
  );


  buf
  g1039
  (
    n576,
    n285
  );


  not
  g1040
  (
    n564,
    n149
  );


  not
  g1041
  (
    n725,
    n408
  );


  not
  g1042
  (
    n423,
    n359
  );


  not
  g1043
  (
    n877,
    n251
  );


  buf
  g1044
  (
    n537,
    n367
  );


  not
  g1045
  (
    n602,
    n178
  );


  not
  g1046
  (
    n946,
    n358
  );


  buf
  g1047
  (
    n678,
    n420
  );


  buf
  g1048
  (
    n1261,
    n362
  );


  not
  g1049
  (
    n909,
    n196
  );


  buf
  g1050
  (
    n947,
    n118
  );


  not
  g1051
  (
    n478,
    n140
  );


  buf
  g1052
  (
    n731,
    n365
  );


  buf
  g1053
  (
    n1428,
    n235
  );


  buf
  g1054
  (
    n1540,
    n373
  );


  not
  g1055
  (
    n1573,
    n227
  );


  buf
  g1056
  (
    n834,
    n393
  );


  buf
  g1057
  (
    n572,
    n117
  );


  buf
  g1058
  (
    n565,
    n215
  );


  buf
  g1059
  (
    n715,
    n357
  );


  not
  g1060
  (
    n588,
    n178
  );


  buf
  g1061
  (
    n1486,
    n138
  );


  not
  g1062
  (
    n1294,
    n159
  );


  not
  g1063
  (
    n1075,
    n351
  );


  not
  g1064
  (
    n1121,
    n194
  );


  buf
  g1065
  (
    n965,
    n202
  );


  not
  g1066
  (
    n1184,
    n296
  );


  buf
  g1067
  (
    n512,
    n340
  );


  buf
  g1068
  (
    n762,
    n272
  );


  not
  g1069
  (
    n1365,
    n214
  );


  buf
  g1070
  (
    n939,
    n328
  );


  buf
  g1071
  (
    n1120,
    n386
  );


  not
  g1072
  (
    n1118,
    n151
  );


  not
  g1073
  (
    n523,
    n160
  );


  not
  g1074
  (
    n1620,
    n297
  );


  buf
  g1075
  (
    n1576,
    n130
  );


  not
  g1076
  (
    n852,
    n256
  );


  buf
  g1077
  (
    n449,
    n208
  );


  not
  g1078
  (
    n593,
    n403
  );


  not
  g1079
  (
    n502,
    n154
  );


  buf
  g1080
  (
    n489,
    n238
  );


  buf
  g1081
  (
    n575,
    n415
  );


  buf
  g1082
  (
    n1554,
    n295
  );


  not
  g1083
  (
    n653,
    n146
  );


  buf
  g1084
  (
    n944,
    n170
  );


  not
  g1085
  (
    n1361,
    n277
  );


  buf
  g1086
  (
    n769,
    n405
  );


  not
  g1087
  (
    n1116,
    n272
  );


  not
  g1088
  (
    n1117,
    n167
  );


  buf
  g1089
  (
    n1157,
    n249
  );


  buf
  g1090
  (
    n1522,
    n154
  );


  buf
  g1091
  (
    n932,
    n280
  );


  buf
  g1092
  (
    n1137,
    n211
  );


  buf
  g1093
  (
    KeyWire_0_23,
    n349
  );


  buf
  g1094
  (
    n1076,
    n337
  );


  buf
  g1095
  (
    n1343,
    n253
  );


  not
  g1096
  (
    KeyWire_0_5,
    n327
  );


  not
  g1097
  (
    n1141,
    n127
  );


  not
  g1098
  (
    n988,
    n231
  );


  buf
  g1099
  (
    n681,
    n230
  );


  not
  g1100
  (
    n626,
    n305
  );


  buf
  g1101
  (
    n1255,
    n231
  );


  not
  g1102
  (
    n716,
    n191
  );


  buf
  g1103
  (
    n1201,
    n373
  );


  buf
  g1104
  (
    n454,
    n377
  );


  not
  g1105
  (
    n968,
    n330
  );


  not
  g1106
  (
    n1037,
    n123
  );


  buf
  g1107
  (
    n920,
    n143
  );


  buf
  g1108
  (
    n1134,
    n363
  );


  not
  g1109
  (
    n1136,
    n244
  );


  buf
  g1110
  (
    n1388,
    n151
  );


  buf
  g1111
  (
    n660,
    n132
  );


  buf
  g1112
  (
    n1209,
    n218
  );


  buf
  g1113
  (
    n673,
    n262
  );


  buf
  g1114
  (
    n1115,
    n196
  );


  buf
  g1115
  (
    n814,
    n226
  );


  not
  g1116
  (
    n598,
    n296
  );


  buf
  g1117
  (
    n1383,
    n231
  );


  buf
  g1118
  (
    n840,
    n402
  );


  buf
  g1119
  (
    n1326,
    n161
  );


  buf
  g1120
  (
    n587,
    n247
  );


  buf
  g1121
  (
    n1374,
    n406
  );


  not
  g1122
  (
    n1213,
    n394
  );


  not
  g1123
  (
    n1680,
    n260
  );


  buf
  g1124
  (
    n1181,
    n391
  );


  not
  g1125
  (
    n1093,
    n135
  );


  buf
  g1126
  (
    n1099,
    n109
  );


  not
  g1127
  (
    n867,
    n417
  );


  buf
  g1128
  (
    n1650,
    n184
  );


  not
  g1129
  (
    n921,
    n371
  );


  buf
  g1130
  (
    n1625,
    n241
  );


  buf
  g1131
  (
    n1663,
    n245
  );


  buf
  g1132
  (
    KeyWire_0_10,
    n326
  );


  buf
  g1133
  (
    n1423,
    n283
  );


  not
  g1134
  (
    n994,
    n341
  );


  buf
  g1135
  (
    n1565,
    n302
  );


  not
  g1136
  (
    n996,
    n279
  );


  buf
  g1137
  (
    n821,
    n216
  );


  not
  g1138
  (
    n1316,
    n305
  );


  buf
  g1139
  (
    n1147,
    n269
  );


  buf
  g1140
  (
    n710,
    n356
  );


  not
  g1141
  (
    n1170,
    n370
  );


  buf
  g1142
  (
    n1649,
    n380
  );


  not
  g1143
  (
    n1089,
    n202
  );


  buf
  g1144
  (
    n1110,
    n290
  );


  not
  g1145
  (
    n828,
    n148
  );


  not
  g1146
  (
    n794,
    n117
  );


  buf
  g1147
  (
    n815,
    n287
  );


  not
  g1148
  (
    n594,
    n197
  );


  not
  g1149
  (
    n680,
    n383
  );


  not
  g1150
  (
    n755,
    n221
  );


  not
  g1151
  (
    n847,
    n167
  );


  buf
  g1152
  (
    n1586,
    n345
  );


  not
  g1153
  (
    n1155,
    n157
  );


  not
  g1154
  (
    n559,
    n315
  );


  buf
  g1155
  (
    n574,
    n328
  );


  not
  g1156
  (
    n1302,
    n358
  );


  not
  g1157
  (
    n1063,
    n187
  );


  not
  g1158
  (
    n1555,
    n148
  );


  not
  g1159
  (
    n636,
    n116
  );


  not
  g1160
  (
    n1011,
    n193
  );


  buf
  g1161
  (
    n568,
    n181
  );


  buf
  g1162
  (
    n1510,
    n133
  );


  buf
  g1163
  (
    n1594,
    n364
  );


  buf
  g1164
  (
    n1578,
    n292
  );


  not
  g1165
  (
    n558,
    n121
  );


  buf
  g1166
  (
    n1456,
    n261
  );


  not
  g1167
  (
    n1020,
    n255
  );


  not
  g1168
  (
    n456,
    n238
  );


  buf
  g1169
  (
    n875,
    n372
  );


  buf
  g1170
  (
    n830,
    n221
  );


  buf
  g1171
  (
    n1478,
    n187
  );


  buf
  g1172
  (
    n1074,
    n268
  );


  not
  g1173
  (
    n1471,
    n340
  );


  not
  g1174
  (
    n1591,
    n268
  );


  not
  g1175
  (
    n1580,
    n182
  );


  buf
  g1176
  (
    n1349,
    n278
  );


  not
  g1177
  (
    n1485,
    n112
  );


  not
  g1178
  (
    n1667,
    n123
  );


  not
  g1179
  (
    n1676,
    n322
  );


  buf
  g1180
  (
    n637,
    n230
  );


  buf
  g1181
  (
    n1357,
    n118
  );


  not
  g1182
  (
    n1585,
    n386
  );


  not
  g1183
  (
    n902,
    n287
  );


  not
  g1184
  (
    n971,
    n226
  );


  not
  g1185
  (
    n811,
    n267
  );


  not
  g1186
  (
    n1453,
    n169
  );


  not
  g1187
  (
    n1483,
    n210
  );


  buf
  g1188
  (
    n766,
    n285
  );


  buf
  g1189
  (
    n472,
    n136
  );


  buf
  g1190
  (
    n1475,
    n203
  );


  buf
  g1191
  (
    n911,
    n168
  );


  buf
  g1192
  (
    KeyWire_0_0,
    n228
  );


  not
  g1193
  (
    n924,
    n181
  );


  buf
  g1194
  (
    n711,
    n338
  );


  buf
  g1195
  (
    n1166,
    n334
  );


  buf
  g1196
  (
    n1472,
    n356
  );


  buf
  g1197
  (
    n809,
    n182
  );


  not
  g1198
  (
    n707,
    n113
  );


  not
  g1199
  (
    n646,
    n212
  );


  buf
  g1200
  (
    n718,
    n252
  );


  buf
  g1201
  (
    n1424,
    n114
  );


  not
  g1202
  (
    n1288,
    n420
  );


  buf
  g1203
  (
    n500,
    n233
  );


  buf
  g1204
  (
    n1291,
    n262
  );


  buf
  g1205
  (
    n1188,
    n274
  );


  buf
  g1206
  (
    n595,
    n113
  );


  buf
  g1207
  (
    n817,
    n313
  );


  buf
  g1208
  (
    n1290,
    n311
  );


  buf
  g1209
  (
    n1362,
    n382
  );


  buf
  g1210
  (
    n684,
    n341
  );


  buf
  g1211
  (
    n986,
    n299
  );


  not
  g1212
  (
    n1441,
    n298
  );


  buf
  g1213
  (
    n554,
    n118
  );


  buf
  g1214
  (
    n589,
    n388
  );


  buf
  g1215
  (
    n541,
    n312
  );


  buf
  g1216
  (
    n1152,
    n121
  );


  not
  g1217
  (
    n1032,
    n176
  );


  buf
  g1218
  (
    n1238,
    n306
  );


  not
  g1219
  (
    n1220,
    n207
  );


  buf
  g1220
  (
    n1140,
    n127
  );


  not
  g1221
  (
    n535,
    n391
  );


  not
  g1222
  (
    n453,
    n222
  );


  buf
  g1223
  (
    n1132,
    n239
  );


  not
  g1224
  (
    n515,
    n327
  );


  buf
  g1225
  (
    n778,
    n358
  );


  not
  g1226
  (
    n1502,
    n323
  );


  buf
  g1227
  (
    n1520,
    n287
  );


  buf
  g1228
  (
    n703,
    n273
  );


  not
  g1229
  (
    n806,
    n302
  );


  buf
  g1230
  (
    n1660,
    n142
  );


  buf
  g1231
  (
    n846,
    n181
  );


  not
  g1232
  (
    n1631,
    n115
  );


  buf
  g1233
  (
    n686,
    n350
  );


  buf
  g1234
  (
    n539,
    n311
  );


  buf
  g1235
  (
    n607,
    n367
  );


  buf
  g1236
  (
    n1253,
    n127
  );


  buf
  g1237
  (
    n513,
    n321
  );


  buf
  g1238
  (
    KeyWire_0_25,
    n352
  );


  buf
  g1239
  (
    n473,
    n195
  );


  not
  g1240
  (
    n930,
    n376
  );


  buf
  g1241
  (
    n1462,
    n400
  );


  not
  g1242
  (
    n787,
    n284
  );


  buf
  g1243
  (
    n1364,
    n162
  );


  not
  g1244
  (
    n839,
    n266
  );


  not
  g1245
  (
    n1638,
    n217
  );


  not
  g1246
  (
    n816,
    n357
  );


  not
  g1247
  (
    n1257,
    n344
  );


  not
  g1248
  (
    n1308,
    n352
  );


  buf
  g1249
  (
    KeyWire_0_16,
    n223
  );


  buf
  g1250
  (
    n1167,
    n111
  );


  not
  g1251
  (
    n1275,
    n295
  );


  buf
  g1252
  (
    n1262,
    n275
  );


  buf
  g1253
  (
    n1635,
    n187
  );


  not
  g1254
  (
    n481,
    n403
  );


  not
  g1255
  (
    n1218,
    n307
  );


  not
  g1256
  (
    n1247,
    n124
  );


  buf
  g1257
  (
    n563,
    n324
  );


  not
  g1258
  (
    n950,
    n111
  );


  buf
  g1259
  (
    n476,
    n189
  );


  buf
  g1260
  (
    n1525,
    n159
  );


  buf
  g1261
  (
    n1151,
    n149
  );


  not
  g1262
  (
    n527,
    n328
  );


  not
  g1263
  (
    n550,
    n305
  );


  buf
  g1264
  (
    n854,
    n147
  );


  buf
  g1265
  (
    n1492,
    n285
  );


  not
  g1266
  (
    n783,
    n214
  );


  not
  g1267
  (
    n1050,
    n186
  );


  buf
  g1268
  (
    n1626,
    n360
  );


  not
  g1269
  (
    n461,
    n235
  );


  not
  g1270
  (
    n805,
    n155
  );


  not
  g1271
  (
    n1174,
    n342
  );


  buf
  g1272
  (
    n883,
    n414
  );


  not
  g1273
  (
    n1149,
    n267
  );


  not
  g1274
  (
    n777,
    n421
  );


  buf
  g1275
  (
    n493,
    n137
  );


  not
  g1276
  (
    n1055,
    n320
  );


  not
  g1277
  (
    n1487,
    n184
  );


  not
  g1278
  (
    n1392,
    n341
  );


  buf
  g1279
  (
    n1029,
    n249
  );


  buf
  g1280
  (
    n1068,
    n361
  );


  buf
  g1281
  (
    n1385,
    n335
  );


  not
  g1282
  (
    n1180,
    n186
  );


  not
  g1283
  (
    n1544,
    n155
  );


  not
  g1284
  (
    n872,
    n227
  );


  buf
  g1285
  (
    n543,
    n300
  );


  buf
  g1286
  (
    n792,
    n225
  );


  buf
  g1287
  (
    n934,
    n402
  );


  buf
  g1288
  (
    n1015,
    n401
  );


  not
  g1289
  (
    n687,
    n179
  );


  not
  g1290
  (
    n529,
    n172
  );


  not
  g1291
  (
    n1225,
    n190
  );


  buf
  g1292
  (
    n597,
    n153
  );


  not
  g1293
  (
    n634,
    n146
  );


  not
  g1294
  (
    n604,
    n311
  );


  buf
  g1295
  (
    n1301,
    n366
  );


  buf
  g1296
  (
    n1342,
    n390
  );


  not
  g1297
  (
    n1489,
    n318
  );


  not
  g1298
  (
    n1634,
    n322
  );


  not
  g1299
  (
    n566,
    n248
  );


  buf
  g1300
  (
    n941,
    n263
  );


  not
  g1301
  (
    n1346,
    n245
  );


  not
  g1302
  (
    n640,
    n332
  );


  not
  g1303
  (
    n708,
    n398
  );


  buf
  g1304
  (
    n1407,
    n212
  );


  not
  g1305
  (
    n662,
    n412
  );


  not
  g1306
  (
    n689,
    n256
  );


  not
  g1307
  (
    n1406,
    n116
  );


  not
  g1308
  (
    n683,
    n338
  );


  not
  g1309
  (
    n699,
    n411
  );


  not
  g1310
  (
    n1642,
    n302
  );


  not
  g1311
  (
    n1442,
    n387
  );


  not
  g1312
  (
    n1246,
    n411
  );


  buf
  g1313
  (
    n596,
    n301
  );


  buf
  g1314
  (
    n1672,
    n275
  );


  not
  g1315
  (
    n1508,
    n273
  );


  buf
  g1316
  (
    n603,
    n343
  );


  buf
  g1317
  (
    n1516,
    n390
  );


  buf
  g1318
  (
    n862,
    n219
  );


  buf
  g1319
  (
    n1087,
    n173
  );


  not
  g1320
  (
    n1285,
    n246
  );


  not
  g1321
  (
    n914,
    n115
  );


  not
  g1322
  (
    n1434,
    n354
  );


  buf
  g1323
  (
    n818,
    n244
  );


  not
  g1324
  (
    n1596,
    n204
  );


  buf
  g1325
  (
    n1482,
    n267
  );


  not
  g1326
  (
    n1497,
    n368
  );


  buf
  g1327
  (
    n427,
    n301
  );


  not
  g1328
  (
    n825,
    n278
  );


  not
  g1329
  (
    n1012,
    n168
  );


  buf
  g1330
  (
    n1284,
    n132
  );


  buf
  g1331
  (
    n1427,
    n396
  );


  buf
  g1332
  (
    n659,
    n289
  );


  buf
  g1333
  (
    n752,
    n336
  );


  not
  g1334
  (
    n1321,
    n165
  );


  buf
  g1335
  (
    n1224,
    n193
  );


  not
  g1336
  (
    n1080,
    n159
  );


  not
  g1337
  (
    n1447,
    n420
  );


  buf
  g1338
  (
    n448,
    n218
  );


  buf
  g1339
  (
    n928,
    n266
  );


  not
  g1340
  (
    n1526,
    n338
  );


  buf
  g1341
  (
    n509,
    n281
  );


  not
  g1342
  (
    n1465,
    n176
  );


  buf
  g1343
  (
    n583,
    n185
  );


  not
  g1344
  (
    n1567,
    n207
  );


  not
  g1345
  (
    n1641,
    n334
  );


  buf
  g1346
  (
    n1628,
    n190
  );


  buf
  g1347
  (
    n1381,
    n124
  );


  not
  g1348
  (
    n732,
    n254
  );


  buf
  g1349
  (
    n1165,
    n303
  );


  buf
  g1350
  (
    n1681,
    n175
  );


  not
  g1351
  (
    n754,
    n375
  );


  buf
  g1352
  (
    n721,
    n254
  );


  not
  g1353
  (
    n802,
    n361
  );


  buf
  g1354
  (
    n1235,
    n389
  );


  buf
  g1355
  (
    n638,
    n397
  );


  buf
  g1356
  (
    n470,
    n231
  );


  buf
  g1357
  (
    n1325,
    n215
  );


  not
  g1358
  (
    n844,
    n329
  );


  buf
  g1359
  (
    n487,
    n132
  );


  not
  g1360
  (
    n1446,
    n250
  );


  not
  g1361
  (
    n1171,
    n262
  );


  buf
  g1362
  (
    n954,
    n215
  );


  buf
  g1363
  (
    n497,
    n315
  );


  not
  g1364
  (
    n702,
    n208
  );


  not
  g1365
  (
    n1026,
    n330
  );


  buf
  g1366
  (
    n893,
    n221
  );


  buf
  g1367
  (
    n1139,
    n339
  );


  not
  g1368
  (
    n1138,
    n321
  );


  buf
  g1369
  (
    n841,
    n326
  );


  buf
  g1370
  (
    n1336,
    n179
  );


  buf
  g1371
  (
    n1481,
    n293
  );


  not
  g1372
  (
    n629,
    n383
  );


  buf
  g1373
  (
    n891,
    n135
  );


  not
  g1374
  (
    n499,
    n257
  );


  buf
  g1375
  (
    n853,
    n130
  );


  not
  g1376
  (
    n1019,
    n319
  );


  not
  g1377
  (
    n1296,
    n309
  );


  buf
  g1378
  (
    n795,
    n109
  );


  not
  g1379
  (
    n1006,
    n194
  );


  not
  g1380
  (
    n498,
    n420
  );


  buf
  g1381
  (
    n1266,
    n243
  );


  not
  g1382
  (
    n879,
    n249
  );


  not
  g1383
  (
    n1205,
    n130
  );


  buf
  g1384
  (
    n501,
    n155
  );


  buf
  g1385
  (
    n1398,
    n266
  );


  buf
  g1386
  (
    n1010,
    n149
  );


  not
  g1387
  (
    n1400,
    n137
  );


  buf
  g1388
  (
    n1566,
    n355
  );


  not
  g1389
  (
    n1182,
    n246
  );


  not
  g1390
  (
    n1332,
    n330
  );


  not
  g1391
  (
    n1551,
    n258
  );


  buf
  g1392
  (
    n432,
    n173
  );


  buf
  g1393
  (
    n483,
    n383
  );


  not
  g1394
  (
    n980,
    n226
  );


  buf
  g1395
  (
    n1394,
    n271
  );


  not
  g1396
  (
    n1086,
    n240
  );


  buf
  g1397
  (
    n705,
    n352
  );


  buf
  g1398
  (
    n1230,
    n327
  );


  not
  g1399
  (
    n987,
    n199
  );


  buf
  g1400
  (
    n1085,
    n376
  );


  not
  g1401
  (
    n1521,
    n142
  );


  buf
  g1402
  (
    n1590,
    n309
  );


  buf
  g1403
  (
    n1380,
    n369
  );


  buf
  g1404
  (
    n1081,
    n399
  );


  buf
  g1405
  (
    KeyWire_0_2,
    n331
  );


  not
  g1406
  (
    n1340,
    n196
  );


  not
  g1407
  (
    n477,
    n311
  );


  buf
  g1408
  (
    n442,
    n148
  );


  buf
  g1409
  (
    n1161,
    n164
  );


  not
  g1410
  (
    n452,
    n263
  );


  not
  g1411
  (
    n1219,
    n241
  );


  not
  g1412
  (
    n861,
    n213
  );


  not
  g1413
  (
    n800,
    n225
  );


  buf
  g1414
  (
    n460,
    n354
  );


  buf
  g1415
  (
    n959,
    n159
  );


  not
  g1416
  (
    n1530,
    n348
  );


  not
  g1417
  (
    n727,
    n371
  );


  not
  g1418
  (
    n864,
    n325
  );


  buf
  g1419
  (
    n742,
    n278
  );


  not
  g1420
  (
    n1303,
    n286
  );


  buf
  g1421
  (
    n1096,
    n323
  );


  not
  g1422
  (
    n688,
    n242
  );


  buf
  g1423
  (
    n967,
    n171
  );


  not
  g1424
  (
    n426,
    n113
  );


  not
  g1425
  (
    n1588,
    n128
  );


  buf
  g1426
  (
    n1277,
    n280
  );


  buf
  g1427
  (
    n1396,
    n179
  );


  buf
  g1428
  (
    n940,
    n381
  );


  not
  g1429
  (
    n894,
    n156
  );


  not
  g1430
  (
    n1189,
    n339
  );


  not
  g1431
  (
    n1259,
    n375
  );


  not
  g1432
  (
    n1592,
    n224
  );


  buf
  g1433
  (
    n1222,
    n113
  );


  not
  g1434
  (
    n813,
    n409
  );


  buf
  g1435
  (
    n1329,
    n416
  );


  buf
  g1436
  (
    n1644,
    n195
  );


  buf
  g1437
  (
    n963,
    n409
  );


  not
  g1438
  (
    n434,
    n281
  );


  buf
  g1439
  (
    n1556,
    n344
  );


  buf
  g1440
  (
    n679,
    n271
  );


  buf
  g1441
  (
    n1250,
    n122
  );


  not
  g1442
  (
    n838,
    n345
  );


  not
  g1443
  (
    n1327,
    n385
  );


  buf
  g1444
  (
    n1639,
    n399
  );


  not
  g1445
  (
    n1251,
    n273
  );


  buf
  g1446
  (
    n1100,
    n397
  );


  buf
  g1447
  (
    n528,
    n222
  );


  buf
  g1448
  (
    n675,
    n388
  );


  buf
  g1449
  (
    n849,
    n416
  );


  not
  g1450
  (
    n1033,
    n384
  );


  buf
  g1451
  (
    n444,
    n385
  );


  not
  g1452
  (
    n972,
    n355
  );


  buf
  g1453
  (
    n1375,
    n304
  );


  buf
  g1454
  (
    n630,
    n304
  );


  not
  g1455
  (
    n677,
    n392
  );


  not
  g1456
  (
    n1195,
    n402
  );


  not
  g1457
  (
    n606,
    n260
  );


  not
  g1458
  (
    n713,
    n327
  );


  not
  g1459
  (
    n985,
    n223
  );


  not
  g1460
  (
    n1039,
    n115
  );


  buf
  g1461
  (
    n1368,
    n226
  );


  buf
  g1462
  (
    n723,
    n347
  );


  not
  g1463
  (
    n530,
    n117
  );


  buf
  g1464
  (
    n1059,
    n120
  );


  buf
  g1465
  (
    n871,
    n184
  );


  not
  g1466
  (
    n1589,
    n290
  );


  buf
  g1467
  (
    n1348,
    n350
  );


  buf
  g1468
  (
    n1065,
    n298
  );


  not
  g1469
  (
    n534,
    n319
  );


  not
  g1470
  (
    n958,
    n348
  );


  not
  g1471
  (
    n1439,
    n111
  );


  not
  g1472
  (
    n1004,
    n312
  );


  buf
  g1473
  (
    n1527,
    n369
  );


  buf
  g1474
  (
    n1324,
    n214
  );


  buf
  g1475
  (
    n1009,
    n244
  );


  buf
  g1476
  (
    n979,
    n382
  );


  buf
  g1477
  (
    n648,
    n174
  );


  not
  g1478
  (
    n546,
    n220
  );


  buf
  g1479
  (
    n1169,
    n155
  );


  not
  g1480
  (
    n1437,
    n182
  );


  buf
  g1481
  (
    n1464,
    n413
  );


  buf
  g1482
  (
    n1005,
    n163
  );


  buf
  g1483
  (
    n1335,
    n237
  );


  buf
  g1484
  (
    n1661,
    n251
  );


  not
  g1485
  (
    n1528,
    n370
  );


  buf
  g1486
  (
    n1476,
    n271
  );


  not
  g1487
  (
    n1228,
    n264
  );


  not
  g1488
  (
    n860,
    n384
  );


  buf
  g1489
  (
    n1603,
    n139
  );


  buf
  g1490
  (
    n1574,
    n216
  );


  not
  g1491
  (
    n881,
    n141
  );


  buf
  g1492
  (
    n622,
    n192
  );


  not
  g1493
  (
    n1583,
    n191
  );


  buf
  g1494
  (
    n600,
    n150
  );


  not
  g1495
  (
    n1466,
    n306
  );


  not
  g1496
  (
    n906,
    n139
  );


  not
  g1497
  (
    n661,
    n316
  );


  buf
  g1498
  (
    n1146,
    n234
  );


  not
  g1499
  (
    n508,
    n309
  );


  not
  g1500
  (
    n904,
    n144
  );


  buf
  g1501
  (
    n1123,
    n166
  );


  not
  g1502
  (
    n1172,
    n250
  );


  not
  g1503
  (
    n1289,
    n217
  );


  buf
  g1504
  (
    n1393,
    n162
  );


  buf
  g1505
  (
    n964,
    n228
  );


  buf
  g1506
  (
    n1094,
    n204
  );


  not
  g1507
  (
    n786,
    n356
  );


  not
  g1508
  (
    n824,
    n292
  );


  not
  g1509
  (
    n1258,
    n189
  );


  not
  g1510
  (
    n1366,
    n347
  );


  buf
  g1511
  (
    n465,
    n203
  );


  buf
  g1512
  (
    n1071,
    n174
  );


  not
  g1513
  (
    n469,
    n407
  );


  buf
  g1514
  (
    n900,
    n391
  );


  buf
  g1515
  (
    n682,
    n347
  );


  buf
  g1516
  (
    n1106,
    n165
  );


  buf
  g1517
  (
    n837,
    n193
  );


  buf
  g1518
  (
    n1113,
    n126
  );


  buf
  g1519
  (
    n1270,
    n235
  );


  not
  g1520
  (
    n625,
    n129
  );


  not
  g1521
  (
    n552,
    n205
  );


  buf
  g1522
  (
    n577,
    n150
  );


  not
  g1523
  (
    n863,
    n232
  );


  not
  g1524
  (
    n829,
    n349
  );


  buf
  g1525
  (
    n1675,
    n254
  );


  buf
  g1526
  (
    n1552,
    n368
  );


  not
  g1527
  (
    n1101,
    n240
  );


  not
  g1528
  (
    KeyWire_0_22,
    n310
  );


  buf
  g1529
  (
    n804,
    n116
  );


  buf
  g1530
  (
    n1276,
    n343
  );


  buf
  g1531
  (
    n1683,
    n178
  );


  buf
  g1532
  (
    n1384,
    n166
  );


  buf
  g1533
  (
    n1413,
    n233
  );


  buf
  g1534
  (
    n803,
    n178
  );


  buf
  g1535
  (
    n1436,
    n274
  );


  buf
  g1536
  (
    n1632,
    n192
  );


  buf
  g1537
  (
    n519,
    n232
  );


  not
  g1538
  (
    n1061,
    n357
  );


  buf
  g1539
  (
    n696,
    n346
  );


  buf
  g1540
  (
    n1490,
    n404
  );


  not
  g1541
  (
    n612,
    n377
  );


  buf
  g1542
  (
    n645,
    n125
  );


  buf
  g1543
  (
    n1538,
    n225
  );


  not
  g1544
  (
    n1607,
    n399
  );


  not
  g1545
  (
    n1216,
    n334
  );


  not
  g1546
  (
    n1468,
    n381
  );


  buf
  g1547
  (
    n1429,
    n396
  );


  buf
  g1548
  (
    n1679,
    n180
  );


  not
  g1549
  (
    n1599,
    n329
  );


  buf
  g1550
  (
    n451,
    n156
  );


  not
  g1551
  (
    n1212,
    n290
  );


  buf
  g1552
  (
    n506,
    n108
  );


  buf
  g1553
  (
    n1048,
    n112
  );


  buf
  g1554
  (
    n1318,
    n246
  );


  buf
  g1555
  (
    n1505,
    n273
  );


  buf
  g1556
  (
    n974,
    n215
  );


  not
  g1557
  (
    n490,
    n245
  );


  buf
  g1558
  (
    n517,
    n156
  );


  buf
  g1559
  (
    n1395,
    n291
  );


  buf
  g1560
  (
    n697,
    n409
  );


  buf
  g1561
  (
    n961,
    n408
  );


  buf
  g1562
  (
    n1363,
    n312
  );


  buf
  g1563
  (
    n1304,
    n209
  );


  buf
  g1564
  (
    n698,
    n291
  );


  not
  g1565
  (
    n745,
    n276
  );


  not
  g1566
  (
    n765,
    n282
  );


  buf
  g1567
  (
    n1397,
    n199
  );


  not
  g1568
  (
    n1072,
    n417
  );


  buf
  g1569
  (
    n1536,
    n169
  );


  not
  g1570
  (
    n781,
    n251
  );


  buf
  g1571
  (
    n555,
    n349
  );


  not
  g1572
  (
    n1183,
    n419
  );


  buf
  g1573
  (
    n913,
    n291
  );


  buf
  g1574
  (
    n1338,
    n237
  );


  buf
  g1575
  (
    n633,
    n400
  );


  not
  g1576
  (
    n758,
    n141
  );


  not
  g1577
  (
    n969,
    n299
  );


  not
  g1578
  (
    n889,
    n171
  );


  not
  g1579
  (
    n1513,
    n394
  );


  not
  g1580
  (
    n1103,
    n322
  );


  not
  g1581
  (
    n1542,
    n401
  );


  not
  g1582
  (
    n1541,
    n140
  );


  not
  g1583
  (
    n1504,
    n349
  );


  not
  g1584
  (
    n759,
    n354
  );


  buf
  g1585
  (
    n536,
    n134
  );


  buf
  g1586
  (
    n1470,
    n292
  );


  not
  g1587
  (
    n1621,
    n315
  );


  not
  g1588
  (
    n463,
    n219
  );


  not
  g1589
  (
    n1668,
    n410
  );


  buf
  g1590
  (
    n1595,
    n188
  );


  buf
  g1591
  (
    n789,
    n145
  );


  buf
  g1592
  (
    n1319,
    n144
  );


  buf
  g1593
  (
    n927,
    n325
  );


  buf
  g1594
  (
    n740,
    n325
  );


  not
  g1595
  (
    n650,
    n280
  );


  buf
  g1596
  (
    n1090,
    n122
  );


  buf
  g1597
  (
    n774,
    n405
  );


  buf
  g1598
  (
    KeyWire_0_18,
    n147
  );


  buf
  g1599
  (
    n1572,
    n234
  );


  buf
  g1600
  (
    n1127,
    n263
  );


  buf
  g1601
  (
    n1104,
    n172
  );


  not
  g1602
  (
    n1678,
    n191
  );


  buf
  g1603
  (
    n966,
    n393
  );


  not
  g1604
  (
    n1451,
    n124
  );


  buf
  g1605
  (
    n1390,
    n161
  );


  not
  g1606
  (
    n1042,
    n145
  );


  buf
  g1607
  (
    n1459,
    n201
  );


  not
  g1608
  (
    n1322,
    n166
  );


  buf
  g1609
  (
    n1373,
    n129
  );


  buf
  g1610
  (
    n1194,
    n341
  );


  not
  g1611
  (
    n480,
    n177
  );


  not
  g1612
  (
    n1239,
    n200
  );


  buf
  g1613
  (
    n1178,
    n211
  );


  buf
  g1614
  (
    n1007,
    n414
  );


  buf
  g1615
  (
    n1252,
    n374
  );


  buf
  g1616
  (
    n1264,
    n387
  );


  not
  g1617
  (
    n560,
    n257
  );


  not
  g1618
  (
    n613,
    n264
  );


  not
  g1619
  (
    n1043,
    n131
  );


  not
  g1620
  (
    n1509,
    n361
  );


  not
  g1621
  (
    n533,
    n130
  );


  buf
  g1622
  (
    n1495,
    n158
  );


  buf
  g1623
  (
    n1562,
    n418
  );


  buf
  g1624
  (
    n1474,
    n409
  );


  buf
  g1625
  (
    n1611,
    n199
  );


  not
  g1626
  (
    n514,
    n242
  );


  not
  g1627
  (
    n557,
    n197
  );


  not
  g1628
  (
    n1243,
    n263
  );


  buf
  g1629
  (
    n912,
    n404
  );


  not
  g1630
  (
    n468,
    n217
  );


  not
  g1631
  (
    n695,
    n257
  );


  not
  g1632
  (
    n1677,
    n298
  );


  not
  g1633
  (
    n1379,
    n415
  );


  buf
  g1634
  (
    n1499,
    n368
  );


  buf
  g1635
  (
    n1314,
    n275
  );


  buf
  g1636
  (
    n908,
    n282
  );


  not
  g1637
  (
    n507,
    n410
  );


  not
  g1638
  (
    n957,
    n406
  );


  not
  g1639
  (
    n1095,
    n314
  );


  not
  g1640
  (
    n1418,
    n304
  );


  not
  g1641
  (
    n1233,
    n224
  );


  not
  g1642
  (
    n1164,
    n160
  );


  not
  g1643
  (
    n1245,
    n305
  );


  buf
  g1644
  (
    n923,
    n129
  );


  buf
  g1645
  (
    n749,
    n186
  );


  not
  g1646
  (
    n433,
    n206
  );


  buf
  g1647
  (
    n1647,
    n125
  );


  buf
  g1648
  (
    n601,
    n293
  );


  not
  g1649
  (
    n1016,
    n232
  );


  not
  g1650
  (
    n1083,
    n126
  );


  not
  g1651
  (
    n484,
    n343
  );


  buf
  g1652
  (
    n989,
    n188
  );


  buf
  g1653
  (
    n1013,
    n298
  );


  buf
  g1654
  (
    n1317,
    n212
  );


  not
  g1655
  (
    n869,
    n132
  );


  not
  g1656
  (
    n641,
    n283
  );


  not
  g1657
  (
    n1432,
    n230
  );


  buf
  g1658
  (
    n551,
    n403
  );


  nand
  g1659
  (
    n2067,
    n1513,
    n1101,
    n1555,
    n1449
  );


  nor
  g1660
  (
    n1763,
    n1336,
    n1481,
    n1395,
    n465
  );


  or
  g1661
  (
    n1957,
    n1551,
    n1597,
    n1331,
    n1093
  );


  or
  g1662
  (
    n2052,
    n633,
    n1506,
    n1317,
    n1478
  );


  xor
  g1663
  (
    n1887,
    n1167,
    n1548,
    n1504,
    n1480
  );


  and
  g1664
  (
    n1971,
    n1065,
    n1551,
    n1516,
    n651
  );


  and
  g1665
  (
    n1848,
    n1457,
    n1261,
    n1371,
    n1495
  );


  or
  g1666
  (
    n1973,
    n1404,
    n1333,
    n1601,
    n457
  );


  xnor
  g1667
  (
    KeyWire_0_24,
    n935,
    n1554,
    n1530,
    n1348
  );


  xnor
  g1668
  (
    n2054,
    n1016,
    n1351,
    n1339,
    n894
  );


  xnor
  g1669
  (
    n1923,
    n1631,
    n1301,
    n618,
    n479
  );


  nand
  g1670
  (
    n1731,
    n1284,
    n1466,
    n1282,
    n1294
  );


  xor
  g1671
  (
    n1772,
    n1435,
    n1352,
    n1155,
    n1362
  );


  and
  g1672
  (
    n1691,
    n1438,
    n1424,
    n503,
    n1453
  );


  xor
  g1673
  (
    n1719,
    n1073,
    n620,
    n1109,
    n734
  );


  xnor
  g1674
  (
    n1819,
    n1171,
    n1622,
    n1491,
    n1627
  );


  nor
  g1675
  (
    n2198,
    n1268,
    n1546,
    n1088,
    n1349
  );


  nand
  g1676
  (
    n2011,
    n667,
    n548,
    n1587,
    n927
  );


  and
  g1677
  (
    n1916,
    n1531,
    n594,
    n1020,
    n792
  );


  nand
  g1678
  (
    n1889,
    n1486,
    n743,
    n945,
    n1582
  );


  xnor
  g1679
  (
    n1783,
    n552,
    n1454,
    n1527,
    n1453
  );


  nand
  g1680
  (
    n1687,
    n433,
    n1308,
    n1372,
    n1574
  );


  or
  g1681
  (
    n1744,
    n839,
    n900,
    n431,
    n622
  );


  xor
  g1682
  (
    n1801,
    n1503,
    n841,
    n1176,
    n1524
  );


  xor
  g1683
  (
    n2091,
    n1389,
    n1631,
    n933,
    n1406
  );


  or
  g1684
  (
    n1754,
    n1576,
    n1493,
    n753,
    n1314
  );


  and
  g1685
  (
    n2004,
    n1542,
    n1592,
    n1490,
    n1163
  );


  and
  g1686
  (
    n1846,
    n721,
    n1459,
    n1402,
    n1017
  );


  xnor
  g1687
  (
    n2169,
    n492,
    n1427,
    n1080,
    n1495
  );


  nand
  g1688
  (
    n2134,
    n1258,
    n1351,
    n1297,
    n673
  );


  nand
  g1689
  (
    n1758,
    n1518,
    n1461,
    n899,
    n1594
  );


  xnor
  g1690
  (
    n2143,
    n1346,
    n1442,
    n652,
    n1437
  );


  or
  g1691
  (
    n1770,
    n1005,
    n1374,
    n1463,
    n1056
  );


  or
  g1692
  (
    n2020,
    n1226,
    n1476,
    n1002,
    n1429
  );


  nand
  g1693
  (
    n2016,
    n1501,
    n1014,
    n1074,
    n1190
  );


  and
  g1694
  (
    n1990,
    n1561,
    n1558,
    n1424,
    n1347
  );


  xor
  g1695
  (
    n2101,
    n575,
    n1316,
    n807,
    n1436
  );


  nand
  g1696
  (
    n1905,
    n1379,
    n1402,
    n1623,
    n1598
  );


  xor
  g1697
  (
    n1958,
    n1477,
    n504,
    n1616,
    n1330
  );


  xnor
  g1698
  (
    n1824,
    n901,
    n1578,
    n1280,
    n1177
  );


  nand
  g1699
  (
    n1688,
    n1045,
    n1631,
    n1515,
    n885
  );


  nor
  g1700
  (
    n1982,
    n832,
    n1575,
    n1572,
    n1483
  );


  nand
  g1701
  (
    n1978,
    n1090,
    n1390,
    n1417,
    n664
  );


  nor
  g1702
  (
    n2234,
    n775,
    n543,
    n691,
    n1453
  );


  and
  g1703
  (
    n2042,
    n719,
    n1568,
    n876,
    n1299
  );


  nor
  g1704
  (
    n1767,
    n1291,
    n941,
    n1572,
    n1289
  );


  and
  g1705
  (
    n1829,
    n970,
    n1536,
    n1108,
    n973
  );


  or
  g1706
  (
    n2074,
    n1293,
    n1500,
    n1419,
    n1591
  );


  or
  g1707
  (
    n2235,
    n610,
    n1431,
    n1625,
    n1352
  );


  or
  g1708
  (
    n1720,
    n1576,
    n956,
    n1443,
    n1084
  );


  nand
  g1709
  (
    n1791,
    n992,
    n1548,
    n685,
    n1114
  );


  or
  g1710
  (
    n2160,
    n1315,
    n1538,
    n1519,
    n1464
  );


  nand
  g1711
  (
    n1712,
    n1546,
    n1260,
    n924,
    n1218
  );


  nor
  g1712
  (
    n2099,
    n1335,
    n511,
    n451,
    n1486
  );


  or
  g1713
  (
    n2034,
    n1285,
    n1308,
    n704,
    n1530
  );


  nand
  g1714
  (
    n1797,
    n506,
    n1414,
    n1460,
    n1173
  );


  xnor
  g1715
  (
    n2253,
    n1309,
    n650,
    n905,
    n1574
  );


  and
  g1716
  (
    n2210,
    n1158,
    n1488,
    n1192,
    n1474
  );


  nand
  g1717
  (
    n1868,
    n1142,
    n1449,
    n1465,
    n1105
  );


  and
  g1718
  (
    n2216,
    n982,
    n1341,
    n1319,
    n637
  );


  xnor
  g1719
  (
    n2230,
    n1611,
    n1441,
    n442,
    n1492
  );


  or
  g1720
  (
    n1816,
    n1361,
    n1013,
    n1015,
    n1029
  );


  nor
  g1721
  (
    n2113,
    n1363,
    n1254,
    n1450,
    n1301
  );


  and
  g1722
  (
    n1793,
    n1343,
    n1350,
    n1356,
    n874
  );


  or
  g1723
  (
    n2015,
    n1426,
    n1311,
    n484,
    n623
  );


  nand
  g1724
  (
    n2121,
    n1577,
    n1552,
    n1299,
    n1432
  );


  xnor
  g1725
  (
    n2238,
    n564,
    n1011,
    n1312,
    n1574
  );


  or
  g1726
  (
    n2153,
    n1345,
    n1535,
    n1369,
    n1289
  );


  or
  g1727
  (
    n1997,
    n831,
    n1609,
    n1237,
    n801
  );


  nand
  g1728
  (
    n2199,
    n1083,
    n1630,
    n1277,
    n1505
  );


  nand
  g1729
  (
    n1778,
    n1310,
    n436,
    n1387,
    n1570
  );


  nor
  g1730
  (
    n2060,
    n508,
    n1403,
    n1428,
    n1325
  );


  and
  g1731
  (
    n1896,
    n742,
    n953,
    n1514,
    n1304
  );


  or
  g1732
  (
    n1689,
    n425,
    n1554,
    n1532,
    n1327
  );


  nor
  g1733
  (
    n1937,
    n1587,
    n1235,
    n1605,
    n1371
  );


  or
  g1734
  (
    n1922,
    n1308,
    n1354,
    n1434,
    n1496
  );


  or
  g1735
  (
    n2162,
    n1394,
    n1420,
    n1324,
    n1374
  );


  xnor
  g1736
  (
    KeyWire_0_1,
    n1416,
    n556,
    n1531,
    n811
  );


  and
  g1737
  (
    n2028,
    n1502,
    n1041,
    n1606,
    n1497
  );


  xor
  g1738
  (
    n1821,
    n1157,
    n1449,
    n489,
    n1577
  );


  nand
  g1739
  (
    n1912,
    n606,
    n1077,
    n1436,
    n1485
  );


  xnor
  g1740
  (
    n1796,
    n1357,
    n1411,
    n805,
    n1630
  );


  nor
  g1741
  (
    n1962,
    n1225,
    n1297,
    n538,
    n1612
  );


  xnor
  g1742
  (
    n2254,
    n1613,
    n706,
    n1197,
    n1358
  );


  nor
  g1743
  (
    n2148,
    n1599,
    n1344,
    n1170,
    n1443
  );


  nor
  g1744
  (
    n1949,
    n1617,
    n1547,
    n1602,
    n1341
  );


  xor
  g1745
  (
    n2263,
    n1269,
    n1505,
    n454,
    n1509
  );


  nor
  g1746
  (
    n2239,
    n1427,
    n1260,
    n1411,
    n1563
  );


  nor
  g1747
  (
    n1950,
    n1353,
    n1319,
    n1075,
    n946
  );


  nor
  g1748
  (
    n1710,
    n1378,
    n1597,
    n870,
    n1344
  );


  or
  g1749
  (
    n2041,
    n939,
    n1413,
    n1442,
    n1382
  );


  xnor
  g1750
  (
    n2055,
    n1266,
    n1256,
    n452,
    n1447
  );


  xor
  g1751
  (
    n2040,
    n1637,
    n1315,
    n1607,
    n605
  );


  nor
  g1752
  (
    n1959,
    n1407,
    n861,
    n1322,
    n755
  );


  nand
  g1753
  (
    n1968,
    n473,
    n1383,
    n851,
    n1463
  );


  nand
  g1754
  (
    n1795,
    n1595,
    n940,
    n824,
    n1317
  );


  nor
  g1755
  (
    n2140,
    n1524,
    n1184,
    n770,
    n1304
  );


  xor
  g1756
  (
    n2025,
    n1445,
    n1287,
    n1295,
    n1332
  );


  xor
  g1757
  (
    n1882,
    n1541,
    n979,
    n1111,
    n1585
  );


  xnor
  g1758
  (
    n1749,
    n642,
    n972,
    n786,
    n1498
  );


  and
  g1759
  (
    n2069,
    n1568,
    n1362,
    n1551,
    n678
  );


  and
  g1760
  (
    n2137,
    n1421,
    n1470,
    n1624,
    n1346
  );


  xor
  g1761
  (
    n2217,
    n1186,
    n607,
    n1201,
    n1362
  );


  nand
  g1762
  (
    n1727,
    n1276,
    n1286,
    n1498,
    n1486
  );


  nand
  g1763
  (
    n1946,
    n590,
    n1320,
    n1460,
    n1570
  );


  xor
  g1764
  (
    n2264,
    n1459,
    n1321,
    n576,
    n1636
  );


  or
  g1765
  (
    n1713,
    n1472,
    n1396,
    n1366,
    n544
  );


  nand
  g1766
  (
    n1789,
    n1543,
    n1370,
    n1462,
    n1456
  );


  xnor
  g1767
  (
    n1881,
    n1430,
    n1433,
    n1605,
    n891
  );


  and
  g1768
  (
    n2076,
    n539,
    n1343,
    n1553,
    n806
  );


  xnor
  g1769
  (
    n1951,
    n1409,
    n916,
    n1168,
    n1467
  );


  xor
  g1770
  (
    n2065,
    n1281,
    n788,
    n1387,
    n875
  );


  xor
  g1771
  (
    n2211,
    n1004,
    n1602,
    n1421,
    n580
  );


  xor
  g1772
  (
    n2100,
    n1405,
    n1622,
    n1507,
    n1361
  );


  nor
  g1773
  (
    n1876,
    n1489,
    n1347,
    n698,
    n1484
  );


  nand
  g1774
  (
    n2071,
    n493,
    n1390,
    n681,
    n1099
  );


  or
  g1775
  (
    n2173,
    n1538,
    n1307,
    n1613,
    n1559
  );


  nand
  g1776
  (
    n2251,
    n1141,
    n1106,
    n1386,
    n1283
  );


  xnor
  g1777
  (
    n1790,
    n1265,
    n1569,
    n1373,
    n1290
  );


  nor
  g1778
  (
    n2119,
    n553,
    n1546,
    n1418,
    n1007
  );


  nand
  g1779
  (
    n2127,
    n1516,
    n1633,
    n1266,
    n1430
  );


  nand
  g1780
  (
    n1947,
    n1472,
    n1275,
    n991,
    n925
  );


  or
  g1781
  (
    n2064,
    n684,
    n1130,
    n888,
    n1331
  );


  and
  g1782
  (
    n2267,
    n1292,
    n1317,
    n1438,
    n1406
  );


  nor
  g1783
  (
    n2261,
    n1599,
    n1332,
    n1365,
    n817
  );


  and
  g1784
  (
    n2195,
    n1620,
    n1350,
    n877,
    n596
  );


  xnor
  g1785
  (
    n2102,
    n513,
    n1556,
    n1282,
    n1441
  );


  nor
  g1786
  (
    n1836,
    n1326,
    n777,
    n581,
    n579
  );


  xnor
  g1787
  (
    n1804,
    n782,
    n1087,
    n1537,
    n1530
  );


  or
  g1788
  (
    n1705,
    n1471,
    n1224,
    n1351,
    n1464
  );


  nor
  g1789
  (
    n2247,
    n1521,
    n577,
    n1280,
    n993
  );


  xor
  g1790
  (
    n2266,
    n957,
    n1427,
    n774,
    n822
  );


  nor
  g1791
  (
    n2168,
    n1081,
    n1250,
    n1293,
    n922
  );


  nand
  g1792
  (
    n1847,
    n1040,
    n1428,
    n1249,
    n613
  );


  xnor
  g1793
  (
    n2026,
    n522,
    n1439,
    n646,
    n1564
  );


  nand
  g1794
  (
    n2213,
    n920,
    n1274,
    n1466,
    n1603
  );


  xor
  g1795
  (
    n2024,
    n1381,
    n1304,
    n938,
    n1571
  );


  xor
  g1796
  (
    n1835,
    n597,
    n879,
    n441,
    n1323
  );


  nor
  g1797
  (
    n1747,
    n1328,
    n1446,
    n1600,
    n1291
  );


  or
  g1798
  (
    n1808,
    n1259,
    n1589,
    n733,
    n1301
  );


  xor
  g1799
  (
    n2039,
    n1464,
    n1179,
    n1381,
    n591
  );


  and
  g1800
  (
    n1779,
    n1501,
    n668,
    n1631,
    n1588
  );


  and
  g1801
  (
    n1964,
    n1232,
    n448,
    n981,
    n1591
  );


  xnor
  g1802
  (
    n2125,
    n1372,
    n1581,
    n833,
    n1263
  );


  and
  g1803
  (
    n1942,
    n1627,
    n1508,
    n1321,
    n450
  );


  or
  g1804
  (
    n1776,
    n1612,
    n1296,
    n1213,
    n1270
  );


  and
  g1805
  (
    n1817,
    n1510,
    n1431,
    n1586,
    n679
  );


  or
  g1806
  (
    n1883,
    n1009,
    n1583,
    n1104,
    n1220
  );


  nand
  g1807
  (
    n2132,
    n1518,
    n1419,
    n1262,
    n727
  );


  or
  g1808
  (
    n1732,
    n1251,
    n948,
    n1506,
    n1468
  );


  nand
  g1809
  (
    n2077,
    n1455,
    n750,
    n1162,
    n1512
  );


  xor
  g1810
  (
    n1904,
    n1563,
    n1560,
    n752,
    n1608
  );


  or
  g1811
  (
    n1910,
    n1590,
    n793,
    n532,
    n1440
  );


  nor
  g1812
  (
    n2124,
    n1398,
    n1618,
    n796,
    n1502
  );


  or
  g1813
  (
    n2030,
    n1520,
    n1368,
    n1433,
    n1635
  );


  nand
  g1814
  (
    n2059,
    n1128,
    n531,
    n1405,
    n1608
  );


  and
  g1815
  (
    n2237,
    n1469,
    n1615,
    n424,
    n826
  );


  or
  g1816
  (
    n1865,
    n1629,
    n1553,
    n1601,
    n1443
  );


  and
  g1817
  (
    n2104,
    n1551,
    n1324,
    n1449,
    n896
  );


  xnor
  g1818
  (
    n1833,
    n1096,
    n1154,
    n1385,
    n1276
  );


  xor
  g1819
  (
    n1726,
    n558,
    n1578,
    n1288,
    n1301
  );


  nor
  g1820
  (
    n1786,
    n1366,
    n759,
    n1513,
    n440
  );


  xor
  g1821
  (
    n2171,
    n1425,
    n736,
    n1438,
    n1384
  );


  nand
  g1822
  (
    n1806,
    n1542,
    n1422,
    n803,
    n1524
  );


  and
  g1823
  (
    n2110,
    n1493,
    n804,
    n1337,
    n621
  );


  or
  g1824
  (
    n1760,
    n675,
    n1429,
    n1627,
    n1576
  );


  nor
  g1825
  (
    n1730,
    n745,
    n632,
    n760,
    n1606
  );


  xnor
  g1826
  (
    n2009,
    n1501,
    n1438,
    n707,
    n1475
  );


  xor
  g1827
  (
    n1834,
    n1425,
    n789,
    n802,
    n1305
  );


  xor
  g1828
  (
    n1998,
    n1359,
    n855,
    n871,
    n857
  );


  or
  g1829
  (
    n1755,
    n978,
    n820,
    n829,
    n1418
  );


  nor
  g1830
  (
    n2215,
    n1457,
    n1169,
    n1064,
    n1477
  );


  xnor
  g1831
  (
    n1828,
    n1612,
    n819,
    n1461,
    n456
  );


  nand
  g1832
  (
    n1897,
    n1510,
    n1102,
    n1479,
    n1351
  );


  xnor
  g1833
  (
    n1826,
    n971,
    n1352,
    n491,
    n1329
  );


  xnor
  g1834
  (
    n2079,
    n1513,
    n1148,
    n1265,
    n1512
  );


  and
  g1835
  (
    n2192,
    n1478,
    n1472,
    n1454,
    n1327
  );


  nand
  g1836
  (
    n2201,
    n1441,
    n1430,
    n1119,
    n1479
  );


  and
  g1837
  (
    n1850,
    n889,
    n1637,
    n533,
    n1496
  );


  or
  g1838
  (
    n2120,
    n1360,
    n602,
    n914,
    n1620
  );


  and
  g1839
  (
    n1980,
    n1203,
    n1525,
    n1440,
    n986
  );


  xnor
  g1840
  (
    n1707,
    n1318,
    n1429,
    n1393,
    n1604
  );


  nor
  g1841
  (
    n2133,
    n630,
    n604,
    n1537,
    n1223
  );


  xnor
  g1842
  (
    n2174,
    n701,
    n1611,
    n1434,
    n1079
  );


  xor
  g1843
  (
    n1831,
    n917,
    n475,
    n911,
    n969
  );


  or
  g1844
  (
    n2207,
    n1582,
    n1284,
    n1406,
    n497
  );


  or
  g1845
  (
    n1722,
    n1591,
    n1571,
    n1446,
    n1614
  );


  or
  g1846
  (
    n1872,
    n1617,
    n1603,
    n955,
    n1306
  );


  nand
  g1847
  (
    n1827,
    n1393,
    n1413,
    n1404,
    n1422
  );


  xor
  g1848
  (
    n1753,
    n1517,
    n1282,
    n1637,
    n1621
  );


  nand
  g1849
  (
    n1921,
    n1483,
    n868,
    n1069,
    n1497
  );


  or
  g1850
  (
    n1878,
    n1536,
    n1399,
    n1116,
    n1144
  );


  nand
  g1851
  (
    n1953,
    n1423,
    n1019,
    n732,
    n1529
  );


  nor
  g1852
  (
    n1736,
    n674,
    n1435,
    n989,
    n1346
  );


  or
  g1853
  (
    n2172,
    n848,
    n1255,
    n1302,
    n988
  );


  xnor
  g1854
  (
    n2088,
    n1509,
    n1616,
    n1370,
    n1279
  );


  and
  g1855
  (
    n1724,
    n1322,
    n1120,
    n1450,
    n1408
  );


  xnor
  g1856
  (
    n2194,
    n1535,
    n1440,
    n1487,
    n1341
  );


  and
  g1857
  (
    n2033,
    n1473,
    n1389,
    n963,
    n1299
  );


  xor
  g1858
  (
    n2008,
    n740,
    n1420,
    n1295,
    n444
  );


  or
  g1859
  (
    n2051,
    n1630,
    n616,
    n1137,
    n1523
  );


  xnor
  g1860
  (
    n2191,
    n1334,
    n530,
    n514,
    n1611
  );


  nand
  g1861
  (
    n1810,
    n1567,
    n1188,
    n1342,
    n1370
  );


  nand
  g1862
  (
    n1952,
    n731,
    n476,
    n1337,
    n1262
  );


  xor
  g1863
  (
    n1867,
    n747,
    n1284,
    n960,
    n1208
  );


  and
  g1864
  (
    n1870,
    n1609,
    n1624,
    n1596,
    n1474
  );


  xnor
  g1865
  (
    n1812,
    n1364,
    n852,
    n483,
    n1458
  );


  or
  g1866
  (
    n1874,
    n722,
    n542,
    n735,
    n1565
  );


  and
  g1867
  (
    n2188,
    n1348,
    n937,
    n1586,
    n1523
  );


  or
  g1868
  (
    n2094,
    n1594,
    n1476,
    n1550,
    n1303
  );


  or
  g1869
  (
    n1841,
    n561,
    n1433,
    n1451,
    n1487
  );


  nand
  g1870
  (
    n2184,
    n1558,
    n1467,
    n1380,
    n1343
  );


  nand
  g1871
  (
    n2243,
    n1558,
    n1270,
    n1006,
    n611
  );


  nand
  g1872
  (
    n2061,
    n1287,
    n560,
    n994,
    n999
  );


  nand
  g1873
  (
    n2145,
    n1042,
    n1533,
    n1626,
    n429
  );


  nor
  g1874
  (
    n1869,
    n1356,
    n1604,
    n1412
  );


  and
  g1875
  (
    n1879,
    n959,
    n509,
    n1288,
    n1471
  );


  xor
  g1876
  (
    n2129,
    n641,
    n1359,
    n962,
    n1354
  );


  nor
  g1877
  (
    n2111,
    n723,
    n1413,
    n1469,
    n566
  );


  nor
  g1878
  (
    n2106,
    n1561,
    n1423,
    n1509,
    n821
  );


  xnor
  g1879
  (
    n1734,
    n729,
    n1319,
    n1180,
    n1475
  );


  nor
  g1880
  (
    n1764,
    n1396,
    n1480,
    n1085,
    n1635
  );


  nor
  g1881
  (
    n1769,
    n1637,
    n1357,
    n1124,
    n1214
  );


  nor
  g1882
  (
    n1794,
    n1450,
    n1340,
    n884,
    n791
  );


  xor
  g1883
  (
    n2157,
    n1417,
    n1037,
    n694,
    n1428
  );


  and
  g1884
  (
    n2103,
    n1526,
    n485,
    n1602,
    n1187
  );


  nor
  g1885
  (
    n2190,
    n1451,
    n1018,
    n1446,
    n1476
  );


  nor
  g1886
  (
    n2013,
    n1121,
    n463,
    n1579,
    n928
  );


  or
  g1887
  (
    n1774,
    n563,
    n499,
    n1492,
    n699
  );


  and
  g1888
  (
    n1773,
    n1127,
    n1332,
    n1291,
    n1381
  );


  nor
  g1889
  (
    n1860,
    n1543,
    n1508,
    n1557,
    n1525
  );


  nor
  g1890
  (
    n1935,
    n1092,
    n1385,
    n1563,
    n1401
  );


  nor
  g1891
  (
    n1920,
    n1369,
    n1589,
    n1067,
    n1437
  );


  xor
  g1892
  (
    n1977,
    n1425,
    n520,
    n1580,
    n1532
  );


  nor
  g1893
  (
    n2175,
    n682,
    n764,
    n1397,
    n748
  );


  nand
  g1894
  (
    n1924,
    n1262,
    n1526,
    n1385,
    n1593
  );


  xnor
  g1895
  (
    n1994,
    n1397,
    n1269,
    n647,
    n1634
  );


  and
  g1896
  (
    n2115,
    n1624,
    n426,
    n1467,
    n1437
  );


  or
  g1897
  (
    n2268,
    n1598,
    n1529,
    n1383,
    n1518
  );


  nor
  g1898
  (
    n2223,
    n1276,
    n464,
    n1216,
    n1022
  );


  xnor
  g1899
  (
    n1766,
    n1330,
    n1378,
    n1635,
    n1552
  );


  and
  g1900
  (
    n2043,
    n1393,
    n1497,
    n779,
    n1456
  );


  and
  g1901
  (
    n2189,
    n1434,
    n1517,
    n1465,
    n1115
  );


  nand
  g1902
  (
    n1886,
    n1509,
    n1123,
    n1600,
    n1134
  );


  nand
  g1903
  (
    n2149,
    n1375,
    n1089,
    n769,
    n626
  );


  nand
  g1904
  (
    n2056,
    n809,
    n523,
    n1181,
    n1452
  );


  nor
  g1905
  (
    n2108,
    n1524,
    n1363,
    n1447,
    n1361
  );


  nor
  g1906
  (
    n2224,
    n432,
    n1515,
    n1580,
    n625
  );


  and
  g1907
  (
    n1866,
    n1585,
    n1519,
    n893,
    n1200
  );


  and
  g1908
  (
    n1700,
    n1613,
    n1566,
    n1583,
    n818
  );


  and
  g1909
  (
    n1820,
    n1391,
    n460,
    n1481,
    n1444
  );


  xnor
  g1910
  (
    n1785,
    n1588,
    n1610,
    n1194,
    n985
  );


  or
  g1911
  (
    n1792,
    n1335,
    n1071,
    n430,
    n1317
  );


  and
  g1912
  (
    n1961,
    n495,
    n1287,
    n459,
    n1462
  );


  xnor
  g1913
  (
    n1757,
    n980,
    n517,
    n1440,
    n624
  );


  or
  g1914
  (
    n1908,
    n1569,
    n1507,
    n1389,
    n1150
  );


  and
  g1915
  (
    n1803,
    n1139,
    n1554,
    n1532,
    n1283
  );


  xor
  g1916
  (
    n1721,
    n1426,
    n1341,
    n1353,
    n1527
  );


  nand
  g1917
  (
    n2090,
    n741,
    n1270,
    n1451,
    n1054
  );


  xnor
  g1918
  (
    n2236,
    n1277,
    n466,
    n1326,
    n1521
  );


  xnor
  g1919
  (
    n2126,
    n1100,
    n1336,
    n932,
    n1146
  );


  xnor
  g1920
  (
    n2166,
    n1564,
    n669,
    n1183,
    n1435
  );


  and
  g1921
  (
    n1832,
    n1407,
    n1634,
    n1138,
    n1178
  );


  nand
  g1922
  (
    n1902,
    n1366,
    n1136,
    n1307,
    n1582
  );


  and
  g1923
  (
    n1843,
    n1455,
    n800,
    n1242,
    n705
  );


  nand
  g1924
  (
    n1798,
    n1504,
    n1293,
    n1588,
    n1614
  );


  xor
  g1925
  (
    n1740,
    n1319,
    n614,
    n1300,
    n1521
  );


  nand
  g1926
  (
    n1733,
    n1193,
    n1566,
    n1601,
    n1495
  );


  nor
  g1927
  (
    n2142,
    n644,
    n998,
    n1356,
    n1402
  );


  or
  g1928
  (
    n2000,
    n1586,
    n1375,
    n481,
    n1159
  );


  nand
  g1929
  (
    n1884,
    n1633,
    n1373,
    n655,
    n435
  );


  xnor
  g1930
  (
    n1926,
    n1217,
    n1408,
    n1118,
    n1097
  );


  xnor
  g1931
  (
    n1861,
    n968,
    n1313,
    n1472,
    n1269
  );


  xnor
  g1932
  (
    n1984,
    n1394,
    n768,
    n449,
    n1350
  );


  xnor
  g1933
  (
    n2176,
    n648,
    n1161,
    n659,
    n1499
  );


  nand
  g1934
  (
    n1837,
    n1403,
    n1323,
    n907,
    n813
  );


  nand
  g1935
  (
    n1745,
    n665,
    n1247,
    n1326,
    n1629
  );


  nand
  g1936
  (
    n1940,
    n926,
    n850,
    n525,
    n536
  );


  xnor
  g1937
  (
    n1913,
    n1615,
    n1132,
    n825,
    n1542
  );


  nand
  g1938
  (
    n2063,
    n1617,
    n1282,
    n1285,
    n1395
  );


  or
  g1939
  (
    n1989,
    n726,
    n1288,
    n1284,
    n1326
  );


  and
  g1940
  (
    n1856,
    n1596,
    n1231,
    n1129,
    n1547
  );


  or
  g1941
  (
    n2159,
    n1391,
    n1636,
    n1447,
    n662
  );


  or
  g1942
  (
    n1914,
    n1061,
    n562,
    n1415,
    n1576
  );


  nor
  g1943
  (
    n1782,
    n1363,
    n1347,
    n1585,
    n1452
  );


  nand
  g1944
  (
    n1751,
    n1479,
    n1619,
    n1567,
    n1503
  );


  and
  g1945
  (
    n1974,
    n1406,
    n1368,
    n1160,
    n467
  );


  xnor
  g1946
  (
    n2170,
    n1416,
    n930,
    n1327,
    n585
  );


  nor
  g1947
  (
    n1859,
    n814,
    n1377,
    n983,
    n1030
  );


  and
  g1948
  (
    n1943,
    n863,
    n1542,
    n1314,
    n501
  );


  xor
  g1949
  (
    n1741,
    n1210,
    n1052,
    n615,
    n1353
  );


  xnor
  g1950
  (
    n1852,
    n1410,
    n1366,
    n529,
    n1202
  );


  xor
  g1951
  (
    n2087,
    n1523,
    n794,
    n1522,
    n1315
  );


  and
  g1952
  (
    n1871,
    n619,
    n1293,
    n1596,
    n1349
  );


  xnor
  g1953
  (
    n2130,
    n881,
    n1415,
    n1199,
    n943
  );


  or
  g1954
  (
    n2098,
    n1579,
    n1376,
    n695,
    n919
  );


  or
  g1955
  (
    n2155,
    n835,
    n1380,
    n515,
    n510
  );


  nor
  g1956
  (
    n1877,
    n570,
    n1625,
    n1550,
    n1435
  );


  xor
  g1957
  (
    n1988,
    n1055,
    n847,
    n1583,
    n903
  );


  nand
  g1958
  (
    n1919,
    n512,
    n1567,
    n1574,
    n1259
  );


  and
  g1959
  (
    n1761,
    n1318,
    n1309,
    n1489,
    n1605
  );


  xnor
  g1960
  (
    n2123,
    n537,
    n816,
    n1432,
    n1310
  );


  or
  g1961
  (
    n2109,
    n1503,
    n787,
    n1516,
    n1315
  );


  or
  g1962
  (
    n1706,
    n844,
    n1261,
    n1527,
    n1575
  );


  nand
  g1963
  (
    n2032,
    n1414,
    n1590,
    n1264,
    n1484
  );


  xnor
  g1964
  (
    n1701,
    n1593,
    n628,
    n1534,
    n1300
  );


  nand
  g1965
  (
    n1956,
    n1335,
    n798,
    n1174,
    n572
  );


  and
  g1966
  (
    n1742,
    n1555,
    n478,
    n1416,
    n1384
  );


  xor
  g1967
  (
    n1845,
    n573,
    n1444,
    n661,
    n1485
  );


  xor
  g1968
  (
    n2116,
    n1469,
    n1328,
    n1400,
    n1236
  );


  and
  g1969
  (
    n1807,
    n1338,
    n1432,
    n1043,
    n1372
  );


  nor
  g1970
  (
    n2049,
    n1035,
    n1498,
    n1491,
    n1175
  );


  nor
  g1971
  (
    n2227,
    n1329,
    n1454,
    n567,
    n773
  );


  and
  g1972
  (
    n1685,
    n952,
    n1384,
    n1499,
    n587
  );


  and
  g1973
  (
    n1686,
    n589,
    n795,
    n1047,
    n1454
  );


  nor
  g1974
  (
    n2085,
    n1364,
    n490,
    n1404,
    n744
  );


  nor
  g1975
  (
    n1818,
    n1433,
    n1505,
    n1283,
    n1545
  );


  nor
  g1976
  (
    n2163,
    n1484,
    n1588,
    n1482,
    n627
  );


  xnor
  g1977
  (
    n1825,
    n1233,
    n1511,
    n1418,
    n1318
  );


  xor
  g1978
  (
    n2156,
    n1596,
    n1382,
    n540,
    n1526
  );


  and
  g1979
  (
    n1941,
    n810,
    n1613,
    n1620,
    n1303
  );


  nor
  g1980
  (
    n1853,
    n535,
    n1632,
    n1053,
    n672
  );


  nor
  g1981
  (
    n1822,
    n1547,
    n1422,
    n1320,
    n895
  );


  xnor
  g1982
  (
    n2018,
    n1409,
    n737,
    n890,
    n1410
  );


  xor
  g1983
  (
    n1800,
    n1458,
    n1271,
    n1492,
    n1562
  );


  or
  g1984
  (
    n2178,
    n1525,
    n588,
    n1500,
    n471
  );


  and
  g1985
  (
    n1917,
    n645,
    n1280,
    n1488,
    n1389
  );


  nor
  g1986
  (
    n1909,
    n1535,
    n873,
    n1310,
    n1265
  );


  and
  g1987
  (
    n1955,
    n1023,
    n1471,
    n1530,
    n1365
  );


  nand
  g1988
  (
    n2225,
    n1581,
    n1582,
    n1323,
    n1298
  );


  nand
  g1989
  (
    n2057,
    n1367,
    n1275,
    n1632,
    n1415
  );


  xor
  g1990
  (
    n2154,
    n555,
    n1427,
    n1513,
    n1633
  );


  and
  g1991
  (
    n2078,
    n1267,
    n1409,
    n1580,
    n1360
  );


  and
  g1992
  (
    n2053,
    n446,
    n494,
    n853,
    n658
  );


  and
  g1993
  (
    n2081,
    n1522,
    n1514,
    n601,
    n593
  );


  xor
  g1994
  (
    n1934,
    n1473,
    n1541,
    n1448,
    n1535
  );


  nand
  g1995
  (
    n1781,
    n1333,
    n1512,
    n710,
    n987
  );


  xor
  g1996
  (
    n2045,
    n1298,
    n1552,
    n1277,
    n1402
  );


  xor
  g1997
  (
    n2257,
    n686,
    n516,
    n977,
    n996
  );


  nand
  g1998
  (
    n2035,
    n1470,
    n1607,
    n1529,
    n1196
  );


  xor
  g1999
  (
    n1738,
    n1205,
    n1364,
    n1297,
    n1305
  );


  nand
  g2000
  (
    n2062,
    n1559,
    n715,
    n797,
    n683
  );


  nand
  g2001
  (
    n1694,
    n1592,
    n1290,
    n1345,
    n1439
  );


  and
  g2002
  (
    n1892,
    n1424,
    n763,
    n1348,
    n1589
  );


  and
  g2003
  (
    n2246,
    n785,
    n1603,
    n842,
    n1330
  );


  and
  g2004
  (
    n2221,
    n1375,
    n486,
    n1367,
    n1560
  );


  xnor
  g2005
  (
    n2259,
    n1477,
    n912,
    n690,
    n1416
  );


  nor
  g2006
  (
    n1933,
    n1528,
    n1603,
    n638,
    n1278
  );


  xnor
  g2007
  (
    n1901,
    n1539,
    n660,
    n799,
    n1610
  );


  xnor
  g2008
  (
    n1996,
    n1500,
    n1281,
    n1570,
    n1633
  );


  and
  g2009
  (
    n2244,
    n1549,
    n1091,
    n1540,
    n815
  );


  nand
  g2010
  (
    n2075,
    n1520,
    n1384,
    n838,
    n1593
  );


  xor
  g2011
  (
    n2084,
    n966,
    n1621,
    n1325,
    n1622
  );


  or
  g2012
  (
    n2206,
    n428,
    n856,
    n1597,
    n1461
  );


  and
  g2013
  (
    n1750,
    n1595,
    n1273,
    n1514,
    n1333
  );


  nor
  g2014
  (
    n1809,
    n902,
    n1206,
    n670,
    n1300
  );


  or
  g2015
  (
    n2152,
    n906,
    n1605,
    n872,
    n1198
  );


  nand
  g2016
  (
    n2072,
    n1024,
    n1487,
    n830,
    n546
  );


  nor
  g2017
  (
    n1775,
    n1281,
    n964,
    n1609,
    n666
  );


  nand
  g2018
  (
    n2019,
    n1403,
    n1274,
    n1289,
    n689
  );


  nor
  g2019
  (
    n2167,
    n849,
    n1209,
    n1555,
    n1463
  );


  and
  g2020
  (
    n2144,
    n1534,
    n1295,
    n739,
    n559
  );


  nor
  g2021
  (
    n2196,
    n1313,
    n1352,
    n1271,
    n1463
  );


  and
  g2022
  (
    n1802,
    n600,
    n1562,
    n1572,
    n1635
  );


  xnor
  g2023
  (
    n1975,
    n1547,
    n954,
    n1426,
    n1165
  );


  and
  g2024
  (
    n2248,
    n1423,
    n676,
    n1291,
    n1034
  );


  nand
  g2025
  (
    n1788,
    n629,
    n472,
    n1536,
    n1606
  );


  nand
  g2026
  (
    n2023,
    n1117,
    n1240,
    n1344,
    n1541
  );


  or
  g2027
  (
    n1880,
    n1354,
    n639,
    n1339,
    n1468
  );


  nand
  g2028
  (
    n1752,
    n1333,
    n1394,
    n840,
    n1131
  );


  or
  g2029
  (
    n2031,
    n653,
    n1399,
    n1468,
    n761
  );


  or
  g2030
  (
    n1697,
    n1219,
    n1031,
    n1571,
    n1010
  );


  xnor
  g2031
  (
    n2233,
    n1526,
    n934,
    n1307,
    n1257
  );


  and
  g2032
  (
    n1844,
    n1369,
    n1457,
    n1544,
    n1528
  );


  xor
  g2033
  (
    n2105,
    n692,
    n1286,
    n1539,
    n1428
  );


  xor
  g2034
  (
    n1900,
    n1540,
    n1248,
    n1412,
    n1584
  );


  nand
  g2035
  (
    n2262,
    n1149,
    n1488,
    n1336,
    n1044
  );


  and
  g2036
  (
    n2001,
    n843,
    n1628,
    n1338,
    n1365
  );


  xor
  g2037
  (
    n1746,
    n554,
    n1078,
    n1587,
    n1314
  );


  or
  g2038
  (
    n2250,
    n1361,
    n445,
    n1436,
    n1518
  );


  xor
  g2039
  (
    n1711,
    n1556,
    n1057,
    n1381,
    n1355
  );


  or
  g2040
  (
    n1911,
    n1485,
    n1522,
    n1275,
    n1459
  );


  nor
  g2041
  (
    n1890,
    n1368,
    n1398,
    n1618,
    n1479
  );


  xnor
  g2042
  (
    n2029,
    n502,
    n1145,
    n1520,
    n772
  );


  nor
  g2043
  (
    n1979,
    n1182,
    n1422,
    n1172,
    n1424
  );


  and
  g2044
  (
    n1999,
    n557,
    n1471,
    n1358,
    n524
  );


  nor
  g2045
  (
    n2118,
    n1512,
    n1441,
    n974,
    n1459
  );


  nor
  g2046
  (
    n2245,
    n812,
    n1553,
    n1271,
    n1490
  );


  nand
  g2047
  (
    n1759,
    n1221,
    n1540,
    n488,
    n1469
  );


  xnor
  g2048
  (
    n1944,
    n860,
    n915,
    n498,
    n1609
  );


  nor
  g2049
  (
    n1885,
    n1565,
    n1388,
    n1519,
    n1420
  );


  nand
  g2050
  (
    n2017,
    n1355,
    n534,
    n1628,
    n1545
  );


  xor
  g2051
  (
    n2037,
    n865,
    n1417,
    n643,
    n1156
  );


  or
  g2052
  (
    n1851,
    n1545,
    n1355,
    n1374,
    n1133
  );


  xor
  g2053
  (
    n1970,
    n1379,
    n1425,
    n1305,
    n1614
  );


  nor
  g2054
  (
    n1839,
    n671,
    n1296,
    n1230,
    n1227
  );


  nor
  g2055
  (
    n2220,
    n1465,
    n1349,
    n677,
    n1439
  );


  xnor
  g2056
  (
    n2027,
    n1398,
    n1063,
    n738,
    n1443
  );


  and
  g2057
  (
    n2222,
    n714,
    n1458,
    n1126,
    n551
  );


  or
  g2058
  (
    n2046,
    n1046,
    n1277,
    n1272,
    n1460
  );


  nand
  g2059
  (
    n2092,
    n1306,
    n1376,
    n1533,
    n1204
  );


  nand
  g2060
  (
    n2114,
    n1632,
    n862,
    n1616,
    n1280
  );


  nor
  g2061
  (
    n2012,
    n1500,
    n1464,
    n612,
    n1536
  );


  xnor
  g2062
  (
    n2165,
    n1537,
    n1152,
    n474,
    n1539
  );


  nor
  g2063
  (
    n2135,
    n1508,
    n1415,
    n1147,
    n1008
  );


  or
  g2064
  (
    n1893,
    n1303,
    n1570,
    n1094,
    n1332
  );


  xor
  g2065
  (
    KeyWire_0_14,
    n749,
    n1565,
    n1466,
    n1386
  );


  and
  g2066
  (
    n1715,
    n1294,
    n1294,
    n1610,
    n1245
  );


  xnor
  g2067
  (
    n2089,
    n1598,
    n1039,
    n1388,
    n1481
  );


  xnor
  g2068
  (
    n1842,
    n918,
    n1619,
    n1413,
    n1252
  );


  and
  g2069
  (
    n1993,
    n1510,
    n1504,
    n1311,
    n1329
  );


  nand
  g2070
  (
    n1728,
    n1295,
    n1553,
    n711,
    n595
  );


  xor
  g2071
  (
    n1992,
    n1390,
    n1564,
    n1525,
    n1426
  );


  xor
  g2072
  (
    n1954,
    n976,
    n1511,
    n892,
    n1060
  );


  or
  g2073
  (
    n1894,
    n1343,
    n1026,
    n1458,
    n1358
  );


  or
  g2074
  (
    n1976,
    n1281,
    n1334,
    n1001,
    n1408
  );


  or
  g2075
  (
    n1830,
    n1482,
    n586,
    n1501,
    n1452
  );


  xnor
  g2076
  (
    n1864,
    n1495,
    n1586,
    n1571,
    n1215
  );


  nand
  g2077
  (
    n1698,
    n1494,
    n1593,
    n1594,
    n1507
  );


  xor
  g2078
  (
    n2204,
    n1490,
    n1625,
    n921,
    n867
  );


  xor
  g2079
  (
    n2068,
    n1337,
    n1483,
    n1316,
    n1532
  );


  or
  g2080
  (
    n2200,
    n1279,
    n1558,
    n923,
    n469
  );


  nand
  g2081
  (
    n2139,
    n1353,
    n1290,
    n1299,
    n1191
  );


  xor
  g2082
  (
    n1756,
    n1626,
    n1623,
    n1557,
    n584
  );


  or
  g2083
  (
    n2151,
    n1481,
    n1493,
    n582,
    n1380
  );


  and
  g2084
  (
    n1765,
    n931,
    n967,
    n437,
    n1357
  );


  or
  g2085
  (
    n2047,
    n1508,
    n756,
    n1618,
    n780
  );


  xnor
  g2086
  (
    n2208,
    n1400,
    n1385,
    n1401,
    n1334
  );


  or
  g2087
  (
    n1771,
    n1534,
    n521,
    n1275,
    n1268
  );


  and
  g2088
  (
    n1777,
    n1556,
    n1401,
    n1618,
    n720
  );


  xor
  g2089
  (
    n1873,
    n1383,
    n1480,
    n1491,
    n1450
  );


  nand
  g2090
  (
    n1967,
    n913,
    n656,
    n887,
    n1340
  );


  or
  g2091
  (
    n2205,
    n1447,
    n1600,
    n1496,
    n1414
  );


  xor
  g2092
  (
    n1823,
    n1480,
    n1338,
    n1395,
    n1021
  );


  xor
  g2093
  (
    n1704,
    n1316,
    n1595,
    n640,
    n1302
  );


  xor
  g2094
  (
    n2086,
    n1456,
    n1573,
    n1189,
    n1304
  );


  or
  g2095
  (
    n1716,
    n1451,
    n1594,
    n965,
    n990
  );


  or
  g2096
  (
    n2209,
    n1414,
    n878,
    n1461,
    n1246
  );


  and
  g2097
  (
    n1938,
    n1517,
    n1626,
    n1625,
    n1342
  );


  and
  g2098
  (
    n1995,
    n1453,
    n480,
    n1457,
    n1239
  );


  xnor
  g2099
  (
    n1805,
    n1566,
    n1330,
    n598,
    n1604
  );


  nor
  g2100
  (
    n1985,
    n1347,
    n1360,
    n1368,
    n864
  );


  and
  g2101
  (
    n2141,
    n1311,
    n693,
    n1550,
    n725
  );


  nand
  g2102
  (
    n1991,
    n708,
    n1391,
    n1578,
    n1504
  );


  nor
  g2103
  (
    n2229,
    n1392,
    n1411,
    n898,
    n712
  );


  or
  g2104
  (
    n2260,
    n1405,
    n470,
    n1068,
    n1515
  );


  nor
  g2105
  (
    n2038,
    n1541,
    n1544,
    n1511,
    n1288
  );


  xor
  g2106
  (
    n2083,
    n1499,
    n1379,
    n1066,
    n1455
  );


  and
  g2107
  (
    n1936,
    n1322,
    n1485,
    n482,
    n1496
  );


  xor
  g2108
  (
    n2240,
    n1392,
    n1418,
    n1497,
    n1599
  );


  xor
  g2109
  (
    n2212,
    n443,
    n866,
    n1626,
    n1421
  );


  nand
  g2110
  (
    n1799,
    n519,
    n1308,
    n717,
    n599
  );


  and
  g2111
  (
    n1787,
    n1318,
    n950,
    n1430,
    n1483
  );


  and
  g2112
  (
    n1714,
    n578,
    n757,
    n1578,
    n1484
  );


  and
  g2113
  (
    n1702,
    n1569,
    n680,
    n1321,
    n1278
  );


  nor
  g2114
  (
    n2131,
    n1397,
    n1376,
    n1567,
    n1493
  );


  nor
  g2115
  (
    n1849,
    n1475,
    n713,
    n1337,
    n1392
  );


  nand
  g2116
  (
    n1906,
    n1393,
    n949,
    n1573,
    n631
  );


  nor
  g2117
  (
    n1875,
    n1399,
    n434,
    n1462,
    n1456
  );


  xor
  g2118
  (
    n2231,
    n1211,
    n1522,
    n1552,
    n1486
  );


  or
  g2119
  (
    n1903,
    n568,
    n1369,
    n1306,
    n1412
  );


  nor
  g2120
  (
    n1743,
    n1027,
    n1448,
    n1290,
    n500
  );


  xnor
  g2121
  (
    n1895,
    n439,
    n565,
    n1624,
    n702
  );


  nor
  g2122
  (
    n2181,
    n1579,
    n1263,
    n1628,
    n1267
  );


  and
  g2123
  (
    n1929,
    n1587,
    n1620,
    n716,
    n1601
  );


  xor
  g2124
  (
    n2095,
    n1573,
    n1298,
    n1356,
    n1151
  );


  and
  g2125
  (
    n1723,
    n1382,
    n728,
    n1434,
    n1059
  );


  xor
  g2126
  (
    n1925,
    n1533,
    n854,
    n1506,
    n1153
  );


  or
  g2127
  (
    n1855,
    n1348,
    n1357,
    n1610,
    n1494
  );


  nand
  g2128
  (
    n1862,
    n1538,
    n1549,
    n1629,
    n1095
  );


  nor
  g2129
  (
    n2158,
    n1309,
    n1452,
    n1444,
    n1549
  );


  or
  g2130
  (
    n1784,
    n574,
    n1506,
    n1437,
    n1238
  );


  or
  g2131
  (
    n2117,
    n1540,
    n1373,
    n1207,
    n1360
  );


  and
  g2132
  (
    n2249,
    n746,
    n1545,
    n1565,
    n1546
  );


  xor
  g2133
  (
    n2080,
    n1365,
    n1354,
    n1292,
    n1442
  );


  nor
  g2134
  (
    n1703,
    n1329,
    n778,
    n1359,
    n1421
  );


  or
  g2135
  (
    n1972,
    n1488,
    n1498,
    n1607,
    n1564
  );


  nor
  g2136
  (
    n2242,
    n1327,
    n1442,
    n1373,
    n1076
  );


  and
  g2137
  (
    n2180,
    n762,
    n1112,
    n528,
    n1420
  );


  xnor
  g2138
  (
    n2193,
    n1544,
    n1264,
    n1038,
    n1274
  );


  nand
  g2139
  (
    n2138,
    n1579,
    n1260,
    n709,
    n1334
  );


  nor
  g2140
  (
    n1931,
    n751,
    n837,
    n1519,
    n1520
  );


  and
  g2141
  (
    n1768,
    n1561,
    n1432,
    n1185,
    n1627
  );


  xnor
  g2142
  (
    n1930,
    n1289,
    n724,
    n1345,
    n1367
  );


  and
  g2143
  (
    n2147,
    n1589,
    n1279,
    n1473,
    n1229
  );


  and
  g2144
  (
    n2203,
    n462,
    n1363,
    n1272,
    n1263
  );


  nor
  g2145
  (
    n1960,
    n1478,
    n608,
    n1598,
    n781
  );


  or
  g2146
  (
    n2058,
    n1276,
    n1324,
    n1412,
    n1303
  );


  xor
  g2147
  (
    n1854,
    n1487,
    n1387,
    n703,
    n1272
  );


  and
  g2148
  (
    n1735,
    n1516,
    n571,
    n908,
    n1331
  );


  or
  g2149
  (
    n2070,
    n487,
    n1296,
    n1474,
    n1320
  );


  nor
  g2150
  (
    n2128,
    n1342,
    n1062,
    n1244,
    n1409
  );


  nor
  g2151
  (
    n2002,
    n1417,
    n1292,
    n697,
    n1448
  );


  nor
  g2152
  (
    n2093,
    n834,
    n1591,
    n1468,
    n1359
  );


  and
  g2153
  (
    n1928,
    n1377,
    n1378,
    n541,
    n1110
  );


  nand
  g2154
  (
    n1983,
    n808,
    n1241,
    n1419,
    n583
  );


  xor
  g2155
  (
    n2050,
    n1355,
    n758,
    n1475,
    n783
  );


  xor
  g2156
  (
    n1725,
    n1311,
    n1113,
    n995,
    n1367
  );


  nand
  g2157
  (
    n1737,
    n1371,
    n1575,
    n1557,
    n975
  );


  or
  g2158
  (
    n2183,
    n1410,
    n505,
    n1273,
    n1503
  );


  nand
  g2159
  (
    n1981,
    n1375,
    n1572,
    n942,
    n1543
  );


  and
  g2160
  (
    n2010,
    n654,
    n1527,
    n1590,
    n882
  );


  xor
  g2161
  (
    n2177,
    n886,
    n1467,
    n1568,
    n636
  );


  xnor
  g2162
  (
    n1986,
    n1557,
    n1554,
    n1103,
    n1345
  );


  nor
  g2163
  (
    n1780,
    n1510,
    n904,
    n427,
    n823
  );


  nor
  g2164
  (
    n2150,
    n1278,
    n1634,
    n1583,
    n1122
  );


  nand
  g2165
  (
    n2036,
    n827,
    n1405,
    n880,
    n1349
  );


  and
  g2166
  (
    n2003,
    n1548,
    n1445,
    n1028,
    n1600
  );


  xor
  g2167
  (
    n2218,
    n1316,
    n1386,
    n1302,
    n1597
  );


  or
  g2168
  (
    n2082,
    n1344,
    n1636,
    n1592,
    n1608
  );


  or
  g2169
  (
    n2185,
    n1476,
    n569,
    n1602,
    n550
  );


  nand
  g2170
  (
    n1965,
    n1195,
    n1395,
    n1268,
    n1340
  );


  nand
  g2171
  (
    n2097,
    n1297,
    n958,
    n1261,
    n1058
  );


  xnor
  g2172
  (
    n2136,
    n468,
    n1556,
    n1292,
    n1164
  );


  or
  g2173
  (
    n1813,
    n1478,
    n1374,
    n1511,
    n1350
  );


  and
  g2174
  (
    n2066,
    n1364,
    n1531,
    n1577,
    n1489
  );


  or
  g2175
  (
    n1888,
    n910,
    n1302,
    n1372,
    n859
  );


  and
  g2176
  (
    n1898,
    n1234,
    n1377,
    n1439,
    n1555
  );


  xor
  g2177
  (
    n2214,
    n1595,
    n1294,
    n1607,
    n1569
  );


  xor
  g2178
  (
    n1927,
    n730,
    n1323,
    n1462,
    n947
  );


  xor
  g2179
  (
    n2258,
    n518,
    n1346,
    n1537,
    n845
  );


  xnor
  g2180
  (
    n1932,
    n1621,
    n1135,
    n696,
    n1446
  );


  xnor
  g2181
  (
    n1695,
    n1310,
    n461,
    n1531,
    n1383
  );


  and
  g2182
  (
    n2256,
    n1407,
    n1266,
    n1125,
    n1617
  );


  nand
  g2183
  (
    n2241,
    n1392,
    n1328,
    n1621,
    n1382
  );


  and
  g2184
  (
    n2187,
    n1470,
    n1000,
    n1314,
    n1051
  );


  and
  g2185
  (
    n2228,
    n883,
    n1507,
    n1502,
    n1243
  );


  or
  g2186
  (
    n2146,
    n1222,
    n1410,
    n1563,
    n1494
  );


  or
  g2187
  (
    n1815,
    n1036,
    n1575,
    n1505,
    n1490
  );


  nor
  g2188
  (
    n2112,
    n1401,
    n1376,
    n1286,
    n507
  );


  xor
  g2189
  (
    n2096,
    n1253,
    n1499,
    n1400,
    n1273
  );


  and
  g2190
  (
    n2006,
    n1285,
    n1379,
    n1400,
    n1423
  );


  or
  g2191
  (
    n1693,
    n936,
    n657,
    n858,
    n609
  );


  or
  g2192
  (
    n2265,
    n1592,
    n1404,
    n1477,
    n836
  );


  or
  g2193
  (
    n1969,
    n1629,
    n1049,
    n1491,
    n634
  );


  and
  g2194
  (
    n1729,
    n688,
    n1548,
    n1397,
    n1259
  );


  or
  g2195
  (
    n2226,
    n1391,
    n1470,
    n1562,
    n1313
  );


  xor
  g2196
  (
    n1838,
    n1312,
    n1370,
    n1358,
    n1336
  );


  xnor
  g2197
  (
    n2107,
    n1212,
    n1140,
    n1562,
    n951
  );


  nor
  g2198
  (
    n2022,
    n1387,
    n828,
    n1429,
    n1003
  );


  and
  g2199
  (
    n1692,
    n1307,
    n1634,
    n1533,
    n592
  );


  or
  g2200
  (
    KeyWire_0_15,
    n1300,
    n1561,
    n687,
    n1577
  );


  xnor
  g2201
  (
    n1966,
    n1070,
    n1448,
    n766,
    n649
  );


  nor
  g2202
  (
    n2255,
    n1465,
    n547,
    n1632,
    n1581
  );


  nand
  g2203
  (
    n2164,
    n527,
    n1396,
    n1338,
    n1419
  );


  and
  g2204
  (
    n2197,
    n790,
    n1408,
    n869,
    n1528
  );


  and
  g2205
  (
    n2122,
    n1072,
    n718,
    n1538,
    n846
  );


  or
  g2206
  (
    n1696,
    n1298,
    n1584,
    n1616,
    n1544
  );


  xnor
  g2207
  (
    n1899,
    n1573,
    n1313,
    n771,
    n1328
  );


  or
  g2208
  (
    n1708,
    n1466,
    n1445,
    n1528,
    n438
  );


  nor
  g2209
  (
    n1814,
    n1517,
    n1431,
    n477,
    n1407
  );


  nand
  g2210
  (
    n2021,
    n1619,
    n1033,
    n1559,
    n1630
  );


  xor
  g2211
  (
    KeyWire_0_26,
    n663,
    n1390,
    n1585,
    n1568
  );


  or
  g2212
  (
    n2073,
    n1287,
    n1482,
    n1560,
    n1143
  );


  and
  g2213
  (
    n1717,
    n1581,
    n944,
    n1306,
    n1534
  );


  or
  g2214
  (
    n1718,
    n1321,
    n1521,
    n617,
    n1515
  );


  and
  g2215
  (
    n1858,
    n423,
    n1309,
    n767,
    n1482
  );


  xnor
  g2216
  (
    n1840,
    n1331,
    n700,
    n455,
    n1622
  );


  and
  g2217
  (
    n2232,
    n1615,
    n1394,
    n1523,
    n1543
  );


  and
  g2218
  (
    n2179,
    n1098,
    n447,
    n1444,
    n1305
  );


  xnor
  g2219
  (
    n2005,
    n1279,
    n1608,
    n1283,
    n1082
  );


  nor
  g2220
  (
    n1857,
    n1550,
    n784,
    n1339,
    n1050
  );


  xor
  g2221
  (
    n2161,
    n1580,
    n1614,
    n526,
    n1396
  );


  or
  g2222
  (
    n1939,
    n1549,
    n1362,
    n776,
    n1431
  );


  xnor
  g2223
  (
    n1690,
    n1606,
    n1398,
    n1559,
    n1460
  );


  and
  g2224
  (
    n2048,
    n1411,
    n1436,
    n1590,
    n1342
  );


  nand
  g2225
  (
    n1891,
    n1494,
    n1285,
    n1086,
    n1228
  );


  nand
  g2226
  (
    n1987,
    n1399,
    n1584,
    n1386,
    n1012
  );


  nand
  g2227
  (
    n1948,
    n1403,
    n1623,
    n961,
    n1489
  );


  or
  g2228
  (
    n1945,
    n1636,
    n909,
    n1286,
    n1377
  );


  xnor
  g2229
  (
    n2182,
    n1474,
    n458,
    n1048,
    n635
  );


  nand
  g2230
  (
    n2014,
    n603,
    n929,
    n1502,
    n1032
  );


  and
  g2231
  (
    n2219,
    n997,
    n1325,
    n1539,
    n1445
  );


  nand
  g2232
  (
    n1739,
    n1320,
    n1492,
    n1312,
    n453
  );


  nand
  g2233
  (
    n1748,
    n1296,
    n1267,
    n1628,
    n1312
  );


  xnor
  g2234
  (
    n2007,
    n1380,
    n897,
    n1455,
    n1566
  );


  nand
  g2235
  (
    n2252,
    n1612,
    n549,
    n1378,
    n1278
  );


  and
  g2236
  (
    n1811,
    n1584,
    n1340,
    n1325,
    n1514
  );


  xor
  g2237
  (
    n1699,
    n1025,
    n496,
    n754,
    n984
  );


  nand
  g2238
  (
    n1709,
    n1388,
    n1264,
    n1166,
    n545
  );


  or
  g2239
  (
    n2202,
    n1560,
    n1335,
    n1619,
    n1388
  );


  nand
  g2240
  (
    n2044,
    n1324,
    n1599,
    n1623,
    n1529
  );


  and
  g2241
  (
    n1963,
    n1611,
    n1371,
    n1339,
    n1473
  );


  nand
  g2242
  (
    n1918,
    n1107,
    n765,
    n1615,
    n1322
  );


  not
  g2243
  (
    n2275,
    n1736
  );


  not
  g2244
  (
    n2303,
    n1701
  );


  not
  g2245
  (
    n2278,
    n1695
  );


  buf
  g2246
  (
    n2272,
    n1723
  );


  not
  g2247
  (
    n2296,
    n1801
  );


  buf
  g2248
  (
    n2288,
    n1763
  );


  buf
  g2249
  (
    n2313,
    n1714
  );


  buf
  g2250
  (
    n2328,
    n1782
  );


  buf
  g2251
  (
    n2326,
    n1765
  );


  buf
  g2252
  (
    n2289,
    n1848
  );


  buf
  g2253
  (
    n2271,
    n1740
  );


  not
  g2254
  (
    n2323,
    n1775
  );


  buf
  g2255
  (
    n2287,
    n1831
  );


  not
  g2256
  (
    n2314,
    n1692
  );


  buf
  g2257
  (
    n2306,
    n1803
  );


  not
  g2258
  (
    n2305,
    n1724
  );


  not
  g2259
  (
    n2291,
    n1698
  );


  buf
  g2260
  (
    n2317,
    n1757
  );


  buf
  g2261
  (
    n2281,
    n1824
  );


  not
  g2262
  (
    n2297,
    n1716
  );


  not
  g2263
  (
    n2292,
    n1713
  );


  not
  g2264
  (
    n2273,
    n1835
  );


  buf
  g2265
  (
    n2319,
    n1709
  );


  not
  g2266
  (
    n2274,
    n1784
  );


  and
  g2267
  (
    n2283,
    n1794,
    n1762,
    n1727,
    n1797
  );


  xnor
  g2268
  (
    n2312,
    n1753,
    n1838,
    n1821,
    n1845
  );


  nor
  g2269
  (
    n2322,
    n1688,
    n1705,
    n1818,
    n1697
  );


  nand
  g2270
  (
    n2277,
    n1707,
    n1843,
    n1820,
    n1702
  );


  nand
  g2271
  (
    n2325,
    n1844,
    n1770,
    n1777,
    n1706
  );


  xor
  g2272
  (
    n2321,
    n1836,
    n1816,
    n1790,
    n1788
  );


  and
  g2273
  (
    n2316,
    n1834,
    n1850,
    n1754,
    n1822
  );


  xnor
  g2274
  (
    n2285,
    n1833,
    n1800,
    n1729,
    n1718
  );


  xor
  g2275
  (
    n2293,
    n1774,
    n1773,
    n1819,
    n1793
  );


  nand
  g2276
  (
    n2270,
    n1852,
    n1847,
    n1733,
    n1725
  );


  or
  g2277
  (
    n2311,
    n1791,
    n1840,
    n1826,
    n1813
  );


  nand
  g2278
  (
    n2269,
    n1812,
    n1696,
    n1738,
    n1804
  );


  and
  g2279
  (
    n2299,
    n1712,
    n1828,
    n1783,
    n1719
  );


  xnor
  g2280
  (
    n2298,
    n1715,
    n1717,
    n1810,
    n1722
  );


  xnor
  g2281
  (
    n2309,
    n1741,
    n1743,
    n1778,
    n1750
  );


  xnor
  g2282
  (
    n2280,
    n1798,
    n1690,
    n1846,
    n1785
  );


  nor
  g2283
  (
    n2301,
    n1825,
    n1815,
    n1809,
    n1699
  );


  xor
  g2284
  (
    n2294,
    n1689,
    n1787,
    n1829,
    n1772
  );


  and
  g2285
  (
    n2284,
    n1830,
    n1720,
    n1841,
    n1807
  );


  or
  g2286
  (
    n2318,
    n1764,
    n1742,
    n1756,
    n1710
  );


  nand
  g2287
  (
    n2295,
    n1759,
    n1823,
    n1711,
    n1761
  );


  xor
  g2288
  (
    n2324,
    n1817,
    n1795,
    n1769,
    n1731
  );


  nand
  g2289
  (
    n2286,
    n1780,
    n1732,
    n1748,
    n1746
  );


  nor
  g2290
  (
    n2307,
    n1728,
    n1726,
    n1745,
    n1693
  );


  nor
  g2291
  (
    n2282,
    n1708,
    n1694,
    n1839,
    n1849
  );


  or
  g2292
  (
    n2279,
    n1703,
    n1811,
    n1808,
    n1766
  );


  nor
  g2293
  (
    n2320,
    n1751,
    n1827,
    n1771,
    n1832
  );


  or
  g2294
  (
    n2302,
    n1851,
    n1735,
    n1747,
    n1734
  );


  xnor
  g2295
  (
    n2304,
    n1767,
    n1686,
    n1837,
    n1842
  );


  and
  g2296
  (
    n2300,
    n1755,
    n1758,
    n1737,
    n1744
  );


  xnor
  g2297
  (
    n2308,
    n1802,
    n1814,
    n1752,
    n1760
  );


  or
  g2298
  (
    n2276,
    n1749,
    n1691,
    n1776,
    n1768
  );


  nor
  g2299
  (
    n2310,
    n1786,
    n1685,
    n1779,
    n1721
  );


  xnor
  g2300
  (
    n2315,
    n1700,
    n1806,
    n1792,
    n1739
  );


  nor
  g2301
  (
    n2327,
    n1781,
    n1730,
    n1687,
    n1796
  );


  nor
  g2302
  (
    n2290,
    n1805,
    n1704,
    n1789,
    n1799
  );


  not
  g2303
  (
    n2331,
    n2278
  );


  not
  g2304
  (
    KeyWire_0_27,
    n2283
  );


  buf
  g2305
  (
    n2333,
    n2285
  );


  not
  g2306
  (
    n2329,
    n2274
  );


  buf
  g2307
  (
    n2336,
    n2282
  );


  buf
  g2308
  (
    n2334,
    n2275
  );


  and
  g2309
  (
    n2337,
    n2272,
    n2280,
    n2269,
    n2273
  );


  nand
  g2310
  (
    n2332,
    n2276,
    n2271,
    n2279,
    n2270
  );


  or
  g2311
  (
    n2330,
    n2277,
    n2286,
    n2284,
    n2281
  );


  not
  g2312
  (
    n2346,
    n2329
  );


  not
  g2313
  (
    n2347,
    n2332
  );


  not
  g2314
  (
    n2357,
    n2330
  );


  not
  g2315
  (
    n2345,
    n2333
  );


  buf
  g2316
  (
    n2338,
    n2332
  );


  buf
  g2317
  (
    n2355,
    n2329
  );


  buf
  g2318
  (
    n2353,
    n2330
  );


  buf
  g2319
  (
    n2348,
    n2331
  );


  buf
  g2320
  (
    n2352,
    n2331
  );


  buf
  g2321
  (
    n2354,
    n2331
  );


  buf
  g2322
  (
    n2356,
    n2330
  );


  not
  g2323
  (
    n2349,
    n2332
  );


  buf
  g2324
  (
    n2344,
    n2331
  );


  not
  g2325
  (
    n2340,
    n2333
  );


  not
  g2326
  (
    n2341,
    n2329
  );


  not
  g2327
  (
    n2339,
    n2332
  );


  not
  g2328
  (
    n2350,
    n2329
  );


  not
  g2329
  (
    n2351,
    n2330
  );


  not
  g2330
  (
    n2342,
    n2333
  );


  buf
  g2331
  (
    n2343,
    n2333
  );


  buf
  g2332
  (
    n2374,
    n2287
  );


  not
  g2333
  (
    n2359,
    n2356
  );


  buf
  g2334
  (
    n2371,
    n2347
  );


  not
  g2335
  (
    n2372,
    n2350
  );


  xnor
  g2336
  (
    n2375,
    n2336,
    n422
  );


  or
  g2337
  (
    n2363,
    n2345,
    n2348,
    n1638,
    n2336
  );


  and
  g2338
  (
    n2364,
    n2354,
    n21,
    n2335,
    n2334
  );


  nor
  g2339
  (
    n2360,
    n2340,
    n22,
    n2336,
    n2352
  );


  nand
  g2340
  (
    n2365,
    n2355,
    n1853,
    n2342,
    n2341
  );


  xor
  g2341
  (
    n2368,
    n2349,
    n2337,
    n1638,
    n2357
  );


  xnor
  g2342
  (
    n2366,
    n2288,
    n2343,
    n2338,
    n2344
  );


  xnor
  g2343
  (
    n2373,
    n2335,
    n21,
    n2352
  );


  nor
  g2344
  (
    n2361,
    n1639,
    n2335,
    n2339,
    n2351
  );


  nor
  g2345
  (
    n2370,
    n2346,
    n2334,
    n2354,
    n2356
  );


  nand
  g2346
  (
    n2362,
    n2355,
    n1638,
    n2337,
    n22
  );


  xor
  g2347
  (
    n2358,
    n2337,
    n1639,
    n2334
  );


  or
  g2348
  (
    n2367,
    n22,
    n2353,
    n2334
  );


  and
  g2349
  (
    n2369,
    n2357,
    n2335,
    n1638,
    n2336
  );


  buf
  g2350
  (
    n2381,
    n106
  );


  buf
  g2351
  (
    n2384,
    n2373
  );


  buf
  g2352
  (
    n2379,
    n2375
  );


  not
  g2353
  (
    n2383,
    n2368
  );


  buf
  g2354
  (
    n2386,
    n2359
  );


  buf
  g2355
  (
    n2388,
    n2362
  );


  buf
  g2356
  (
    KeyWire_0_12,
    n2372
  );


  buf
  g2357
  (
    n2391,
    n2364
  );


  buf
  g2358
  (
    n2377,
    n2365
  );


  buf
  g2359
  (
    KeyWire_0_3,
    n105
  );


  buf
  g2360
  (
    n2378,
    n2370
  );


  not
  g2361
  (
    n2389,
    n2363
  );


  nand
  g2362
  (
    n2382,
    n2369,
    n2367,
    n106
  );


  and
  g2363
  (
    n2390,
    n2360,
    n2361,
    n105
  );


  xor
  g2364
  (
    n2387,
    n2371,
    n2374,
    n2366
  );


  xnor
  g2365
  (
    n2385,
    n2358,
    n105
  );


  or
  g2366
  (
    n2392,
    n2378,
    n2379,
    n2376,
    n2377
  );


  buf
  g2367
  (
    n2394,
    n2392
  );


  or
  g2368
  (
    n2393,
    n2392,
    n23,
    n22
  );


  not
  g2369
  (
    n2395,
    n2394
  );


  not
  g2370
  (
    n2400,
    n2394
  );


  buf
  g2371
  (
    n2397,
    n2393
  );


  buf
  g2372
  (
    n2398,
    n2394
  );


  not
  g2373
  (
    n2396,
    n2394
  );


  buf
  g2374
  (
    n2399,
    n2393
  );


  not
  g2375
  (
    n2401,
    n2393
  );


  not
  g2376
  (
    n2403,
    n2398
  );


  buf
  g2377
  (
    n2402,
    n2398
  );


  buf
  g2378
  (
    n2407,
    n2396
  );


  not
  g2379
  (
    n2405,
    n2395
  );


  and
  g2380
  (
    n2404,
    n2395,
    n2397,
    n2398
  );


  and
  g2381
  (
    n2406,
    n2397,
    n2396,
    n2395
  );


  not
  g2382
  (
    KeyWire_0_8,
    n1641
  );


  xnor
  g2383
  (
    n2411,
    n2406,
    n1640,
    n2405
  );


  and
  g2384
  (
    n2408,
    n2407,
    n1639,
    n1640,
    n2403
  );


  xnor
  g2385
  (
    n2410,
    n1640,
    n1640,
    n2404,
    n2402
  );


  xor
  g2386
  (
    n2412,
    n1855,
    n1854,
    n1856,
    n2408
  );


  and
  g2387
  (
    n2413,
    n2412,
    n2294,
    n2289,
    n2292
  );


  nor
  g2388
  (
    n2414,
    n2290,
    n2293,
    n2412,
    n2291
  );


  not
  g2389
  (
    n2418,
    n2414
  );


  not
  g2390
  (
    n2415,
    n2413
  );


  not
  g2391
  (
    n2421,
    n2414
  );


  buf
  g2392
  (
    n2422,
    n2414
  );


  buf
  g2393
  (
    n2417,
    n2413
  );


  not
  g2394
  (
    n2416,
    n2413
  );


  not
  g2395
  (
    n2419,
    n2413
  );


  buf
  g2396
  (
    n2420,
    n2414
  );


  nor
  g2397
  (
    n2433,
    n2420,
    n2417
  );


  nor
  g2398
  (
    n2434,
    n1641,
    n25
  );


  xnor
  g2399
  (
    n2435,
    n25,
    n2422
  );


  xnor
  g2400
  (
    n2436,
    n2417,
    n25
  );


  xor
  g2401
  (
    n2439,
    n23,
    n2418
  );


  nand
  g2402
  (
    n2424,
    n2419,
    n2381
  );


  or
  g2403
  (
    n2431,
    n2419,
    n2380
  );


  nor
  g2404
  (
    n2423,
    n2296,
    n2422
  );


  nor
  g2405
  (
    n2425,
    n2295,
    n2415
  );


  xor
  g2406
  (
    n2430,
    n2420,
    n2421
  );


  or
  g2407
  (
    n2428,
    n2297,
    n23
  );


  nand
  g2408
  (
    n2429,
    n24,
    n2422
  );


  xnor
  g2409
  (
    n2437,
    n25,
    n2421
  );


  xnor
  g2410
  (
    n2426,
    n2415,
    n24
  );


  buf
  g2411
  (
    n2440,
    n2416
  );


  nor
  g2412
  (
    n2427,
    n24,
    n1641
  );


  nand
  g2413
  (
    n2438,
    n2418,
    n24
  );


  xnor
  g2414
  (
    n2432,
    n2421,
    n23
  );


  not
  g2415
  (
    n2456,
    n2430
  );


  not
  g2416
  (
    n2449,
    n2434
  );


  buf
  g2417
  (
    n2452,
    n2428
  );


  not
  g2418
  (
    n2446,
    n2431
  );


  not
  g2419
  (
    n2448,
    n2438
  );


  not
  g2420
  (
    n2450,
    n2423
  );


  buf
  g2421
  (
    n2451,
    n2425
  );


  not
  g2422
  (
    n2442,
    n2427
  );


  not
  g2423
  (
    n2455,
    n2437
  );


  not
  g2424
  (
    n2447,
    n2432
  );


  not
  g2425
  (
    n2453,
    n2435
  );


  buf
  g2426
  (
    n2445,
    n2426
  );


  buf
  g2427
  (
    n2441,
    n2433
  );


  not
  g2428
  (
    n2454,
    n2429
  );


  buf
  g2429
  (
    n2443,
    n2436
  );


  buf
  g2430
  (
    n2444,
    n2424
  );


  nor
  g2431
  (
    n2457,
    n2456,
    n2451,
    n2453
  );


  xor
  g2432
  (
    n2465,
    n2451,
    n2456,
    n2454
  );


  xor
  g2433
  (
    n2464,
    n2456,
    n2451,
    n2382,
    n2445
  );


  xor
  g2434
  (
    n2460,
    n2454,
    n2455,
    n2450
  );


  and
  g2435
  (
    n2466,
    n2441,
    n2453,
    n2442,
    n2452
  );


  nor
  g2436
  (
    n2461,
    n2387,
    n2455,
    n2452,
    n2449
  );


  or
  g2437
  (
    n2459,
    n2446,
    n2385,
    n2444,
    n2455
  );


  and
  g2438
  (
    n2458,
    n2454,
    n2383,
    n2386,
    n2453
  );


  or
  g2439
  (
    n2463,
    n2452,
    n2447,
    n2453,
    n2448
  );


  nand
  g2440
  (
    n2462,
    n2454,
    n2384,
    n2452,
    n2443
  );


  buf
  g2441
  (
    n2473,
    n2460
  );


  not
  g2442
  (
    n2474,
    n2463
  );


  buf
  g2443
  (
    n2471,
    n2461
  );


  not
  g2444
  (
    n2468,
    n2398
  );


  buf
  g2445
  (
    n2470,
    n2459
  );


  xor
  g2446
  (
    n2467,
    n2466,
    n1641,
    n1642
  );


  or
  g2447
  (
    n2469,
    n2465,
    n1642,
    n2464
  );


  nand
  g2448
  (
    n2472,
    n2462,
    n2399,
    n1642
  );


  nand
  g2449
  (
    n2483,
    n2472,
    n1870
  );


  xor
  g2450
  (
    n2490,
    n2400,
    n1858
  );


  xor
  g2451
  (
    n2481,
    n2468,
    n2472
  );


  buf
  g2452
  (
    n2486,
    n2469
  );


  xor
  g2453
  (
    n2491,
    n1857,
    n1860
  );


  and
  g2454
  (
    n2494,
    n1866,
    n1859
  );


  or
  g2455
  (
    n2476,
    n1862,
    n1864
  );


  nand
  g2456
  (
    n2493,
    n1868,
    n2401
  );


  nand
  g2457
  (
    n2478,
    n2473,
    n2471
  );


  xnor
  g2458
  (
    n2487,
    n2471,
    n2473
  );


  and
  g2459
  (
    n2480,
    n2474,
    n2468
  );


  buf
  g2460
  (
    n2492,
    n2470
  );


  or
  g2461
  (
    n2489,
    n1865,
    n1863
  );


  nand
  g2462
  (
    n2475,
    n1871,
    n2399
  );


  or
  g2463
  (
    n2479,
    n2470,
    n1867
  );


  nand
  g2464
  (
    n2485,
    n2400,
    n2467
  );


  xor
  g2465
  (
    n2495,
    n2400,
    n2467
  );


  nor
  g2466
  (
    n2482,
    n2399,
    n2472
  );


  xor
  g2467
  (
    n2477,
    n2467,
    n1872
  );


  nand
  g2468
  (
    n2498,
    n2474,
    n2400
  );


  and
  g2469
  (
    n2484,
    n2469,
    n2401
  );


  or
  g2470
  (
    n2488,
    n2473,
    n2471
  );


  nor
  g2471
  (
    n2497,
    n2474,
    n2468
  );


  xnor
  g2472
  (
    n2496,
    n1869,
    n1861
  );


  buf
  g2473
  (
    n2501,
    n2475
  );


  not
  g2474
  (
    n2507,
    n2482
  );


  buf
  g2475
  (
    n2502,
    n2479
  );


  not
  g2476
  (
    n2504,
    n2477
  );


  not
  g2477
  (
    n2500,
    n2481
  );


  not
  g2478
  (
    n2508,
    n2483
  );


  buf
  g2479
  (
    n2499,
    n2480
  );


  not
  g2480
  (
    n2506,
    n2484
  );


  not
  g2481
  (
    n2505,
    n2476
  );


  not
  g2482
  (
    n2503,
    n2478
  );


  xnor
  g2483
  (
    n2521,
    n2504,
    n2500,
    n2501,
    n2320
  );


  nor
  g2484
  (
    n2520,
    n2507,
    n2502,
    n2508,
    n2309
  );


  nor
  g2485
  (
    n2516,
    n2307,
    n2305,
    n2504,
    n2315
  );


  nand
  g2486
  (
    n2525,
    n2501,
    n2501,
    n2505,
    n2324
  );


  xnor
  g2487
  (
    n2524,
    n2507,
    n2500,
    n2298,
    n2505
  );


  xnor
  g2488
  (
    n2515,
    n2303,
    n2505,
    n2302
  );


  xor
  g2489
  (
    n2513,
    n2311,
    n2300,
    n2502,
    n2319
  );


  xnor
  g2490
  (
    n2517,
    n2313,
    n2322,
    n2308,
    n2318
  );


  or
  g2491
  (
    n2522,
    n2299,
    n2503,
    n2506,
    n2314
  );


  and
  g2492
  (
    n2510,
    n2316,
    n2508,
    n2506,
    n2503
  );


  and
  g2493
  (
    KeyWire_0_13,
    n2503,
    n2506,
    n2502,
    n2312
  );


  nand
  g2494
  (
    n2512,
    n2499,
    n2500,
    n2301,
    n2321
  );


  xnor
  g2495
  (
    n2519,
    n2503,
    n2504,
    n2323,
    n2499
  );


  nor
  g2496
  (
    KeyWire_0_20,
    n2500,
    n2325,
    n2317,
    n2502
  );


  xnor
  g2497
  (
    n2511,
    n2507,
    n2506,
    n2310,
    n2499
  );


  xor
  g2498
  (
    n2514,
    n2501,
    n2507,
    n2304,
    n2508
  );


  xnor
  g2499
  (
    n2523,
    n2306,
    n2504,
    n2508,
    n2499
  );


  buf
  g2500
  (
    n2540,
    n1887
  );


  not
  g2501
  (
    n2530,
    n1886
  );


  and
  g2502
  (
    n2532,
    n2328,
    n2408
  );


  nand
  g2503
  (
    n2535,
    n1882,
    n2326,
    n2411,
    n1881
  );


  nand
  g2504
  (
    n2539,
    n2408,
    n2327,
    n2509,
    n2514
  );


  and
  g2505
  (
    n2536,
    n2516,
    n2409,
    n2524,
    n2513
  );


  xor
  g2506
  (
    n2537,
    n1880,
    n2409,
    n2411,
    n2410
  );


  xnor
  g2507
  (
    n2528,
    n1877,
    n2525,
    n2337,
    n1874
  );


  xor
  g2508
  (
    n2529,
    n2410,
    n1879,
    n2515,
    n2522
  );


  nand
  g2509
  (
    n2531,
    n1885,
    n1878,
    n1888,
    n1873
  );


  xnor
  g2510
  (
    n2527,
    n1875,
    n2410,
    n1883,
    n1884
  );


  or
  g2511
  (
    n2534,
    n2411,
    n2510,
    n2521,
    n2511
  );


  nor
  g2512
  (
    n2538,
    n2410,
    n2408,
    n1876,
    n2411
  );


  xnor
  g2513
  (
    n2526,
    n2517,
    n2518,
    n2409
  );


  xnor
  g2514
  (
    n2533,
    n2512,
    n2520,
    n2519,
    n2523
  );


  buf
  g2515
  (
    n2547,
    n1896
  );


  buf
  g2516
  (
    n2543,
    n1901
  );


  buf
  g2517
  (
    n2548,
    n1892
  );


  not
  g2518
  (
    n2542,
    n1890
  );


  buf
  g2519
  (
    n2545,
    n2529
  );


  not
  g2520
  (
    n2556,
    n1893
  );


  not
  g2521
  (
    n2551,
    n2528
  );


  not
  g2522
  (
    n2549,
    n2535
  );


  not
  g2523
  (
    n2555,
    n2536
  );


  nor
  g2524
  (
    n2552,
    n1900,
    n2532,
    n2531,
    n1891
  );


  nand
  g2525
  (
    n2553,
    n1898,
    n2530,
    n2533,
    n1906
  );


  nand
  g2526
  (
    n2554,
    n2537,
    n1902,
    n1905,
    n2540
  );


  and
  g2527
  (
    n2544,
    n1908,
    n1907,
    n1903,
    n2526
  );


  xor
  g2528
  (
    n2546,
    n1895,
    n2527,
    n2538,
    n2539
  );


  xnor
  g2529
  (
    n2541,
    n1904,
    n2534,
    n1894,
    n1889
  );


  nand
  g2530
  (
    n2550,
    n2412,
    n2540,
    n1897,
    n1899
  );


  nor
  g2531
  (
    n2590,
    n2545,
    n1665,
    n1662,
    n1660
  );


  nand
  g2532
  (
    n2587,
    n1672,
    n1659,
    n1683,
    n1649
  );


  xor
  g2533
  (
    n2608,
    n2546,
    n1670,
    n1661
  );


  nor
  g2534
  (
    n2572,
    n1684,
    n1678,
    n1653,
    n1647
  );


  xor
  g2535
  (
    n2581,
    n2547,
    n1651,
    n2552,
    n1678
  );


  xor
  g2536
  (
    n2592,
    n1682,
    n1648,
    n1677,
    n2391
  );


  xnor
  g2537
  (
    n2582,
    n1668,
    n1659,
    n2556,
    n2544
  );


  xor
  g2538
  (
    n2579,
    n1664,
    n1653,
    n2543,
    n1643
  );


  xnor
  g2539
  (
    n2560,
    n1657,
    n1660,
    n1648,
    n1654
  );


  xnor
  g2540
  (
    n2607,
    n1679,
    n1672,
    n1677,
    n1647
  );


  and
  g2541
  (
    n2584,
    n1659,
    n1909,
    n2551,
    n2489
  );


  nor
  g2542
  (
    n2567,
    n1661,
    n2552,
    n1649,
    n1663
  );


  and
  g2543
  (
    n2602,
    n2546,
    n1667,
    n2495,
    n2547
  );


  or
  g2544
  (
    n2586,
    n2550,
    n1680,
    n1651,
    n2556
  );


  xor
  g2545
  (
    n2611,
    n2553,
    n2496,
    n1666,
    n1673
  );


  nor
  g2546
  (
    n2615,
    n1676,
    n2542,
    n1649,
    n1670
  );


  nor
  g2547
  (
    n2594,
    n1684,
    n2553,
    n1666,
    n1650
  );


  xor
  g2548
  (
    n2620,
    n2546,
    n2485,
    n1684,
    n1683
  );


  nand
  g2549
  (
    n2616,
    n2541,
    n1650,
    n2544,
    n2555
  );


  nor
  g2550
  (
    n2565,
    n1680,
    n1674,
    n2545
  );


  nand
  g2551
  (
    n2618,
    n1666,
    n2543,
    n2549,
    n1665
  );


  and
  g2552
  (
    n2617,
    n1681,
    n1653,
    n1676,
    n1663
  );


  xor
  g2553
  (
    n2557,
    n1656,
    n1679,
    n1673,
    n1671
  );


  and
  g2554
  (
    n2561,
    n1643,
    n2494,
    n2556,
    n1652
  );


  or
  g2555
  (
    n2609,
    n2548,
    n1662,
    n1681,
    n2545
  );


  nand
  g2556
  (
    n2596,
    n2551,
    n1652,
    n2553,
    n1653
  );


  or
  g2557
  (
    n2595,
    n1667,
    n1662,
    n1651,
    n1645
  );


  or
  g2558
  (
    n2599,
    n2550,
    n1669,
    n1675,
    n1651
  );


  xor
  g2559
  (
    n2558,
    n1649,
    n1674,
    n2541,
    n1645
  );


  or
  g2560
  (
    n2601,
    n2554,
    n2390,
    n2541,
    n1676
  );


  or
  g2561
  (
    n2604,
    n2555,
    n2548,
    n2486,
    n1660
  );


  xor
  g2562
  (
    n2568,
    n1645,
    n1668,
    n1676,
    n1683
  );


  or
  g2563
  (
    n2570,
    n1658,
    n2550,
    n1657,
    n1674
  );


  nand
  g2564
  (
    n2605,
    n1663,
    n1656,
    n1654,
    n2495
  );


  and
  g2565
  (
    n2563,
    n2547,
    n1667,
    n1657,
    n2552
  );


  xor
  g2566
  (
    n2575,
    n1669,
    n1645,
    n1680,
    n2542
  );


  or
  g2567
  (
    n2610,
    n1654,
    n2544,
    n2554,
    n1660
  );


  nor
  g2568
  (
    n2603,
    n2542,
    n2542,
    n1668,
    n1679
  );


  xnor
  g2569
  (
    n2585,
    n1664,
    n1644,
    n1673,
    n1675
  );


  xnor
  g2570
  (
    n2564,
    n1681,
    n1646,
    n1652,
    n1678
  );


  xor
  g2571
  (
    n2566,
    n1655,
    n2548,
    n1674,
    n2554
  );


  nor
  g2572
  (
    n2574,
    n1671,
    n1654,
    n1661,
    n1683
  );


  xor
  g2573
  (
    n2571,
    n1659,
    n2554,
    n1677,
    n1668
  );


  or
  g2574
  (
    n2562,
    n1666,
    n2552,
    n1664,
    n2496
  );


  nor
  g2575
  (
    n2589,
    n1657,
    n1658,
    n1655,
    n2549
  );


  nor
  g2576
  (
    n2613,
    n1673,
    n2493,
    n1665,
    n1669
  );


  nor
  g2577
  (
    n2600,
    n2495,
    n1647,
    n2488,
    n1682
  );


  or
  g2578
  (
    n2583,
    n1665,
    n2551,
    n1670,
    n1644
  );


  xor
  g2579
  (
    n2614,
    n2492,
    n2548,
    n2551,
    n1643
  );


  or
  g2580
  (
    n2580,
    n1675,
    n1648,
    n1646,
    n1681
  );


  xor
  g2581
  (
    n2606,
    n2543,
    n1663,
    n1643,
    n1650
  );


  xor
  g2582
  (
    n2578,
    n2389,
    n2495,
    n1672
  );


  xnor
  g2583
  (
    n2576,
    n2555,
    n2493,
    n2549,
    n2388
  );


  nand
  g2584
  (
    n2577,
    n2541,
    n1644,
    n1650
  );


  or
  g2585
  (
    n2597,
    n1647,
    n1680,
    n2487,
    n1646
  );


  or
  g2586
  (
    n2588,
    n1682,
    n2549,
    n1655,
    n1678
  );


  xor
  g2587
  (
    n2559,
    n1664,
    n1646,
    n2550,
    n1661
  );


  nand
  g2588
  (
    n2573,
    n2556,
    n1682,
    n1675,
    n2491
  );


  xor
  g2589
  (
    n2591,
    n1671,
    n1655,
    n1656,
    n2555
  );


  xnor
  g2590
  (
    n2612,
    n2543,
    n1671,
    n2544,
    n2490
  );


  nand
  g2591
  (
    n2593,
    n1652,
    n2553,
    n2496,
    n1677
  );


  nor
  g2592
  (
    n2619,
    n1662,
    n1658,
    n1669,
    n2547
  );


  and
  g2593
  (
    n2598,
    n1684,
    n2494,
    n1648,
    n1679
  );


  and
  g2594
  (
    n2569,
    n1656,
    n2546,
    n1667,
    n1658
  );


  or
  g2595
  (
    n2677,
    n2087,
    n2085,
    n1938,
    n2606
  );


  nand
  g2596
  (
    n2622,
    n2594,
    n2044,
    n2221,
    n2176
  );


  xor
  g2597
  (
    n2715,
    n2093,
    n2192,
    n2012,
    n1977
  );


  or
  g2598
  (
    n2638,
    n2143,
    n2051,
    n2108,
    n2572
  );


  nand
  g2599
  (
    n2680,
    n2096,
    n2594,
    n2159,
    n1982
  );


  nand
  g2600
  (
    n2727,
    n2580,
    n2605,
    n2040,
    n2567
  );


  xor
  g2601
  (
    n2707,
    n2614,
    n2147,
    n2042,
    n2039
  );


  and
  g2602
  (
    n2662,
    n2109,
    n2114,
    n2581,
    n2161
  );


  nand
  g2603
  (
    n2722,
    n2239,
    n2223,
    n2617,
    n1966
  );


  or
  g2604
  (
    n2667,
    n2104,
    n2025,
    n2247,
    n2002
  );


  xnor
  g2605
  (
    n2628,
    n2575,
    n2153,
    n2243,
    n1912
  );


  nand
  g2606
  (
    n2669,
    n2217,
    n2257,
    n2615,
    n2244
  );


  xnor
  g2607
  (
    n2639,
    n2105,
    n2057,
    n2584,
    n2035
  );


  nor
  g2608
  (
    n2731,
    n2249,
    n2578,
    n2256,
    n2056
  );


  or
  g2609
  (
    n2718,
    n2082,
    n1994,
    n2194,
    n2053
  );


  nor
  g2610
  (
    n2642,
    n2229,
    n2614,
    n2561,
    n2140
  );


  or
  g2611
  (
    n2655,
    n2066,
    n2148,
    n2033,
    n2260
  );


  or
  g2612
  (
    n2735,
    n2602,
    n2618,
    n2565,
    n2001
  );


  nand
  g2613
  (
    n2635,
    n1942,
    n2185,
    n2052,
    n2571
  );


  nor
  g2614
  (
    n2630,
    n2186,
    n1988,
    n1932,
    n2055
  );


  nor
  g2615
  (
    n2661,
    n2589,
    n1923,
    n2585,
    n2224
  );


  nor
  g2616
  (
    n2656,
    n2162,
    n1975,
    n2157,
    n2058
  );


  xnor
  g2617
  (
    n2621,
    n2102,
    n2582,
    n2592,
    n2599
  );


  or
  g2618
  (
    n2732,
    n2591,
    n2619,
    n1976,
    n2575
  );


  and
  g2619
  (
    n2676,
    n2022,
    n2198,
    n2191,
    n2007
  );


  or
  g2620
  (
    n2721,
    n2015,
    n2258,
    n2596,
    n2567
  );


  xnor
  g2621
  (
    n2706,
    n2240,
    n2227,
    n2248,
    n2602
  );


  or
  g2622
  (
    n2645,
    n2073,
    n2593,
    n2216,
    n2171
  );


  or
  g2623
  (
    n2650,
    n1951,
    n2173,
    n2600,
    n2251
  );


  and
  g2624
  (
    n2685,
    n1998,
    n2078,
    n2094,
    n1979
  );


  xor
  g2625
  (
    n2703,
    n2195,
    n2564,
    n2031,
    n2152
  );


  xor
  g2626
  (
    n2651,
    n2142,
    n2620,
    n2235,
    n2580
  );


  xnor
  g2627
  (
    n2654,
    n2577,
    n2242,
    n2168,
    n2589
  );


  xor
  g2628
  (
    n2710,
    n2010,
    n2156,
    n2180,
    n2061
  );


  and
  g2629
  (
    n2670,
    n2196,
    n2069,
    n2588,
    n1983
  );


  and
  g2630
  (
    n2708,
    n2184,
    n2189,
    n2107,
    n2144
  );


  xnor
  g2631
  (
    n2728,
    n2263,
    n1969,
    n2129,
    n2212
  );


  nor
  g2632
  (
    n2701,
    n1944,
    n2214,
    n2604,
    n2182
  );


  nand
  g2633
  (
    n2647,
    n2219,
    n2027,
    n1913,
    n2136
  );


  or
  g2634
  (
    n2664,
    n2587,
    n2106,
    n1958,
    n2597
  );


  or
  g2635
  (
    n2631,
    n2172,
    n1987,
    n2034,
    n2618
  );


  or
  g2636
  (
    n2657,
    n2588,
    n2097,
    n2111,
    n2193
  );


  nand
  g2637
  (
    n2733,
    n2578,
    n1930,
    n2586,
    n2112
  );


  nor
  g2638
  (
    n2692,
    n2146,
    n2037,
    n2086,
    n2074
  );


  nor
  g2639
  (
    n2713,
    n1949,
    n2201,
    n1963,
    n1939
  );


  or
  g2640
  (
    n2725,
    n2593,
    n2583,
    n2181,
    n2236
  );


  and
  g2641
  (
    n2689,
    n2576,
    n2026,
    n2117,
    n2041
  );


  or
  g2642
  (
    n2720,
    n1972,
    n1943,
    n2200,
    n2590
  );


  xor
  g2643
  (
    n2644,
    n2150,
    n1911,
    n2072,
    n1996
  );


  nand
  g2644
  (
    n2665,
    n2211,
    n2003,
    n2611,
    n2265
  );


  and
  g2645
  (
    n2712,
    n1964,
    n2253,
    n2178,
    n1971
  );


  and
  g2646
  (
    n2729,
    n2579,
    n2127,
    n1992,
    n2563
  );


  xor
  g2647
  (
    n2653,
    n2131,
    n1959,
    n2226,
    n2209
  );


  xnor
  g2648
  (
    n2686,
    n1929,
    n1921,
    n2154,
    n2213
  );


  xor
  g2649
  (
    n2693,
    n2016,
    n2206,
    n2163,
    n1937
  );


  nand
  g2650
  (
    n2632,
    n2067,
    n2014,
    n2017,
    n1981
  );


  or
  g2651
  (
    n2640,
    n2569,
    n1945,
    n2151,
    n2603
  );


  nor
  g2652
  (
    n2698,
    n1985,
    n2177,
    n1956,
    n2116
  );


  and
  g2653
  (
    n2679,
    n2255,
    n2080,
    n2188,
    n2092
  );


  and
  g2654
  (
    n2737,
    n2075,
    n1993,
    n1980,
    n2573
  );


  xor
  g2655
  (
    n2678,
    n2208,
    n2581,
    n2113,
    n1925
  );


  nand
  g2656
  (
    n2682,
    n2230,
    n2081,
    n2128,
    n2098
  );


  nand
  g2657
  (
    n2700,
    n1920,
    n2601,
    n2613,
    n2063
  );


  xor
  g2658
  (
    n2683,
    n1940,
    n1991,
    n2101,
    n2079
  );


  nor
  g2659
  (
    n2624,
    n1933,
    n2124,
    n1955,
    n2577
  );


  and
  g2660
  (
    n2646,
    n2557,
    n2175,
    n2570,
    n2234
  );


  nand
  g2661
  (
    n2658,
    n1990,
    n2076,
    n2570,
    n2254
  );


  nor
  g2662
  (
    n2696,
    n1914,
    n2062,
    n2615,
    n2169
  );


  and
  g2663
  (
    n2716,
    n2077,
    n2245,
    n1968,
    n2585
  );


  xnor
  g2664
  (
    n2740,
    n2220,
    n2103,
    n2586,
    n2558
  );


  and
  g2665
  (
    n2649,
    n2203,
    n2006,
    n2091,
    n1950
  );


  xnor
  g2666
  (
    n2709,
    n2609,
    n2610,
    n2572,
    n2587
  );


  or
  g2667
  (
    n2705,
    n2207,
    n2048,
    n2164,
    n2599
  );


  xor
  g2668
  (
    n2637,
    n2021,
    n2167,
    n2238,
    n2598
  );


  or
  g2669
  (
    n2636,
    n2008,
    n2204,
    n2232,
    n2083
  );


  xor
  g2670
  (
    n2687,
    n2605,
    n2607,
    n2590,
    n2099
  );


  and
  g2671
  (
    n2714,
    n1924,
    n2562,
    n2043,
    n1973
  );


  nor
  g2672
  (
    n2734,
    n2218,
    n2574,
    n1965,
    n2609
  );


  nand
  g2673
  (
    n2626,
    n2011,
    n2046,
    n2582,
    n2250
  );


  xnor
  g2674
  (
    n2668,
    n2134,
    n2612,
    n2210,
    n2559
  );


  xnor
  g2675
  (
    n2726,
    n2122,
    n2174,
    n2613,
    n2120
  );


  nand
  g2676
  (
    n2730,
    n1967,
    n1989,
    n1926,
    n1978
  );


  xor
  g2677
  (
    n2694,
    n2579,
    n2565,
    n2030,
    n1986
  );


  and
  g2678
  (
    n2739,
    n2132,
    n2560,
    n2597,
    n1953
  );


  and
  g2679
  (
    n2697,
    n2619,
    n2133,
    n1960,
    n2566
  );


  xor
  g2680
  (
    n2699,
    n2569,
    n2029,
    n1974,
    n2568
  );


  and
  g2681
  (
    n2695,
    n2205,
    n2050,
    n2600,
    n2024
  );


  and
  g2682
  (
    n2623,
    n2141,
    n2158,
    n1962,
    n2065
  );


  and
  g2683
  (
    n2627,
    n2121,
    n2267,
    n2118,
    n2179
  );


  nor
  g2684
  (
    n2629,
    n2606,
    n2088,
    n2126,
    n2009
  );


  xnor
  g2685
  (
    n2723,
    n1928,
    n2584,
    n1922,
    n1957
  );


  xnor
  g2686
  (
    n2675,
    n2123,
    n1948,
    n2222,
    n2607
  );


  and
  g2687
  (
    KeyWire_0_7,
    n2612,
    n2036,
    n2603,
    n2090
  );


  xor
  g2688
  (
    n2674,
    n2237,
    n2047,
    n2119,
    n2028
  );


  and
  g2689
  (
    n2711,
    n2145,
    n1918,
    n2135,
    n1995
  );


  nand
  g2690
  (
    n2719,
    n2049,
    n2020,
    n2054,
    n2608
  );


  and
  g2691
  (
    n2625,
    n1941,
    n2611,
    n2266,
    n2264
  );


  xor
  g2692
  (
    n2643,
    n2576,
    n2595,
    n2095,
    n2023
  );


  and
  g2693
  (
    n2688,
    n2013,
    n2160,
    n2598,
    n2000
  );


  xnor
  g2694
  (
    KeyWire_0_29,
    n2608,
    n2166,
    n1915,
    n2170
  );


  nor
  g2695
  (
    n2663,
    n2130,
    n2583,
    n1931,
    n2241
  );


  xnor
  g2696
  (
    n2736,
    n2060,
    n2268,
    n1936,
    n2616
  );


  nand
  g2697
  (
    n2724,
    n2591,
    n2610,
    n2592,
    n2125
  );


  xnor
  g2698
  (
    n2704,
    n1916,
    n2138,
    n2573,
    n2620
  );


  xnor
  g2699
  (
    n2648,
    n2604,
    n2089,
    n2616,
    n2262
  );


  nand
  g2700
  (
    n2652,
    n2566,
    n2137,
    n2233,
    n1919
  );


  xor
  g2701
  (
    n2634,
    n1954,
    n2574,
    n1970,
    n2019
  );


  nor
  g2702
  (
    n2672,
    n2190,
    n2202,
    n2068,
    n2004
  );


  xor
  g2703
  (
    n2671,
    n1946,
    n2100,
    n1984,
    n2115
  );


  nor
  g2704
  (
    n2690,
    n2187,
    n2199,
    n2045,
    n2070
  );


  nand
  g2705
  (
    n2684,
    n2231,
    n2246,
    n2571,
    n1934
  );


  xor
  g2706
  (
    n2633,
    n1997,
    n2183,
    n1961,
    n2197
  );


  xnor
  g2707
  (
    n2641,
    n2005,
    n2064,
    n2059,
    n1927
  );


  or
  g2708
  (
    KeyWire_0_11,
    n1999,
    n2568,
    n2071,
    n2617
  );


  nand
  g2709
  (
    n2717,
    n2018,
    n422,
    n2165,
    n2252
  );


  nand
  g2710
  (
    n2681,
    n2596,
    n1952,
    n2215,
    n2155
  );


  nand
  g2711
  (
    n2702,
    n2110,
    n2038,
    n2149,
    n2601
  );


  xor
  g2712
  (
    n2660,
    n2032,
    n2228,
    n1910,
    n2225
  );


  xor
  g2713
  (
    n2666,
    n2139,
    n2259,
    n2084,
    n1917
  );


  nor
  g2714
  (
    n2673,
    n2261,
    n2595,
    n1947,
    n1935
  );


  xnor
  g2715
  (
    n2744,
    n2696,
    n2725,
    n2649,
    n2648
  );


  nor
  g2716
  (
    n2748,
    n2665,
    n2673,
    n2675,
    n2632
  );


  nand
  g2717
  (
    n2742,
    n2656,
    n2726,
    n2623,
    n2722
  );


  or
  g2718
  (
    n2761,
    n2662,
    n2497,
    n2697,
    n2723
  );


  or
  g2719
  (
    n2743,
    n2627,
    n2737,
    n2657,
    n2706
  );


  xor
  g2720
  (
    n2768,
    n2651,
    n2637,
    n2661,
    n2669
  );


  and
  g2721
  (
    n2755,
    n2715,
    n2653,
    n2659,
    n2680
  );


  or
  g2722
  (
    n2766,
    n2672,
    n2695,
    n2644,
    n2497
  );


  xor
  g2723
  (
    n2756,
    n2704,
    n2733,
    n2708,
    n2724
  );


  and
  g2724
  (
    n2759,
    n2686,
    n2688,
    n2711,
    n2727
  );


  nand
  g2725
  (
    n2771,
    n2676,
    n2641,
    n2645,
    n2698
  );


  xor
  g2726
  (
    n2746,
    n2713,
    n2646,
    n2626,
    n2679
  );


  or
  g2727
  (
    n2760,
    n2714,
    n2716,
    n2689,
    n2734
  );


  nand
  g2728
  (
    n2753,
    n2692,
    n2732,
    n2712,
    n2710
  );


  nand
  g2729
  (
    n2770,
    n2701,
    n2498,
    n2643,
    n2684
  );


  xor
  g2730
  (
    n2747,
    n2683,
    n2674,
    n2728,
    n2634
  );


  or
  g2731
  (
    n2752,
    n2658,
    n2631,
    n2736,
    n2666
  );


  xnor
  g2732
  (
    n2763,
    n2670,
    n2630,
    n2622,
    n2735
  );


  xor
  g2733
  (
    n2751,
    n2740,
    n2642,
    n2647,
    n2635
  );


  nor
  g2734
  (
    KeyWire_0_9,
    n2655,
    n2678,
    n2729,
    n2439
  );


  nand
  g2735
  (
    n2741,
    n2738,
    n2731,
    n2694,
    n2633
  );


  and
  g2736
  (
    n2764,
    n2401,
    n2650,
    n2624,
    n2700
  );


  xor
  g2737
  (
    n2774,
    n2730,
    n2639,
    n2690,
    n2628
  );


  nor
  g2738
  (
    n2773,
    n2440,
    n106,
    n2739,
    n2691
  );


  and
  g2739
  (
    n2767,
    n2497,
    n2681,
    n2677,
    n2703
  );


  xor
  g2740
  (
    n2765,
    n2717,
    n2740,
    n2401,
    n2663
  );


  xor
  g2741
  (
    n2754,
    n2496,
    n2707,
    n2654,
    n2660
  );


  xor
  g2742
  (
    n2757,
    n2682,
    n2687,
    n2671,
    n2664
  );


  or
  g2743
  (
    n2745,
    n2497,
    n2699,
    n2702,
    n2640
  );


  or
  g2744
  (
    n2762,
    n2719,
    n2705,
    n2720,
    n2721
  );


  xor
  g2745
  (
    n2758,
    n2440,
    n2668,
    n2638,
    n2625
  );


  xnor
  g2746
  (
    n2769,
    n2709,
    n2685,
    n2636,
    n2629
  );


  and
  g2747
  (
    n2772,
    n2693,
    n2667,
    n2718,
    n2498
  );


  or
  g2748
  (
    KeyWire_0_19,
    n2652,
    n2498,
    n106
  );


  xor
  KeyGate_0_0
  (
    n445,
    keyIn_0_0,
    KeyWire_0_0
  );


  xnor
  KeyGate_0_1
  (
    n2186,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n548,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n2376,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n123,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    n796,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n591,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n2738,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n2409,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n2749,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    n615,
    keyIn_0_10,
    KeyWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    n2659,
    keyIn_0_11,
    KeyWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n2380,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n2518,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1915,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n1863,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1637,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n669,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n1035,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n2750,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n2509,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n647,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n1445,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1203,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n1907,
    keyIn_0_24,
    KeyWire_0_24
  );


  xnor
  KeyGate_0_25
  (
    n1041,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n1762,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n2335,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n729,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    n2691,
    keyIn_0_29,
    KeyWire_0_29
  );


  xor
  KeyGate_0_30
  (
    n393,
    keyIn_0_30,
    KeyWire_0_30
  );


  xnor
  KeyGate_0_31
  (
    n79,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


