// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_1000_104 written by SynthGen on 2021/04/05 11:08:33
module Stat_1000_104( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n731, n623, n637, n649, n677, n718, n675, n616,
 n668, n707, n643, n626, n701, n625, n735, n681,
 n627, n1022, n1020, n1019, n1031, n1026, n1029, n1023,
 n1021, n1024, n1025, n1027, n1030, n1028, n1018, n1032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n731, n623, n637, n649, n677, n718, n675, n616,
 n668, n707, n643, n626, n701, n625, n735, n681,
 n627, n1022, n1020, n1019, n1031, n1026, n1029, n1023,
 n1021, n1024, n1025, n1027, n1030, n1028, n1018, n1032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n442, n443, n444, n445, n446, n447, n448,
 n449, n450, n451, n452, n453, n454, n455, n456,
 n457, n458, n459, n460, n461, n462, n463, n464,
 n465, n466, n467, n468, n469, n470, n471, n472,
 n473, n474, n475, n476, n477, n478, n479, n480,
 n481, n482, n483, n484, n485, n486, n487, n488,
 n489, n490, n491, n492, n493, n494, n495, n496,
 n497, n498, n499, n500, n501, n502, n503, n504,
 n505, n506, n507, n508, n509, n510, n511, n512,
 n513, n514, n515, n516, n517, n518, n519, n520,
 n521, n522, n523, n524, n525, n526, n527, n528,
 n529, n530, n531, n532, n533, n534, n535, n536,
 n537, n538, n539, n540, n541, n542, n543, n544,
 n545, n546, n547, n548, n549, n550, n551, n552,
 n553, n554, n555, n556, n557, n558, n559, n560,
 n561, n562, n563, n564, n565, n566, n567, n568,
 n569, n570, n571, n572, n573, n574, n575, n576,
 n577, n578, n579, n580, n581, n582, n583, n584,
 n585, n586, n587, n588, n589, n590, n591, n592,
 n593, n594, n595, n596, n597, n598, n599, n600,
 n601, n602, n603, n604, n605, n606, n607, n608,
 n609, n610, n611, n612, n613, n614, n615, n617,
 n618, n619, n620, n621, n622, n624, n628, n629,
 n630, n631, n632, n633, n634, n635, n636, n638,
 n639, n640, n641, n642, n644, n645, n646, n647,
 n648, n650, n651, n652, n653, n654, n655, n656,
 n657, n658, n659, n660, n661, n662, n663, n664,
 n665, n666, n667, n669, n670, n671, n672, n673,
 n674, n676, n678, n679, n680, n682, n683, n684,
 n685, n686, n687, n688, n689, n690, n691, n692,
 n693, n694, n695, n696, n697, n698, n699, n700,
 n702, n703, n704, n705, n706, n708, n709, n710,
 n711, n712, n713, n714, n715, n716, n717, n719,
 n720, n721, n722, n723, n724, n725, n726, n727,
 n728, n729, n730, n732, n733, n734, n736, n737,
 n738, n739, n740, n741, n742, n743, n744, n745,
 n746, n747, n748, n749, n750, n751, n752, n753,
 n754, n755, n756, n757, n758, n759, n760, n761,
 n762, n763, n764, n765, n766, n767, n768, n769,
 n770, n771, n772, n773, n774, n775, n776, n777,
 n778, n779, n780, n781, n782, n783, n784, n785,
 n786, n787, n788, n789, n790, n791, n792, n793,
 n794, n795, n796, n797, n798, n799, n800, n801,
 n802, n803, n804, n805, n806, n807, n808, n809,
 n810, n811, n812, n813, n814, n815, n816, n817,
 n818, n819, n820, n821, n822, n823, n824, n825,
 n826, n827, n828, n829, n830, n831, n832, n833,
 n834, n835, n836, n837, n838, n839, n840, n841,
 n842, n843, n844, n845, n846, n847, n848, n849,
 n850, n851, n852, n853, n854, n855, n856, n857,
 n858, n859, n860, n861, n862, n863, n864, n865,
 n866, n867, n868, n869, n870, n871, n872, n873,
 n874, n875, n876, n877, n878, n879, n880, n881,
 n882, n883, n884, n885, n886, n887, n888, n889,
 n890, n891, n892, n893, n894, n895, n896, n897,
 n898, n899, n900, n901, n902, n903, n904, n905,
 n906, n907, n908, n909, n910, n911, n912, n913,
 n914, n915, n916, n917, n918, n919, n920, n921,
 n922, n923, n924, n925, n926, n927, n928, n929,
 n930, n931, n932, n933, n934, n935, n936, n937,
 n938, n939, n940, n941, n942, n943, n944, n945,
 n946, n947, n948, n949, n950, n951, n952, n953,
 n954, n955, n956, n957, n958, n959, n960, n961,
 n962, n963, n964, n965, n966, n967, n968, n969,
 n970, n971, n972, n973, n974, n975, n976, n977,
 n978, n979, n980, n981, n982, n983, n984, n985,
 n986, n987, n988, n989, n990, n991, n992, n993,
 n994, n995, n996, n997, n998, n999, n1000, n1001,
 n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
 n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017;

buf  g0 (n158, n30);
not  g1 (n71, n16);
buf  g2 (n147, n11);
buf  g3 (n101, n22);
not  g4 (n96, n22);
not  g5 (n157, n29);
buf  g6 (n159, n27);
buf  g7 (n37, n10);
buf  g8 (n126, n10);
buf  g9 (n73, n4);
not  g10 (n120, n27);
buf  g11 (n152, n32);
not  g12 (n47, n23);
not  g13 (n41, n8);
buf  g14 (n110, n24);
not  g15 (n90, n13);
buf  g16 (n72, n5);
buf  g17 (n99, n1);
not  g18 (n69, n25);
not  g19 (n145, n26);
buf  g20 (n55, n1);
buf  g21 (n98, n25);
not  g22 (n60, n6);
not  g23 (n116, n3);
buf  g24 (n92, n18);
buf  g25 (n82, n28);
not  g26 (n59, n8);
buf  g27 (n49, n12);
buf  g28 (n61, n15);
buf  g29 (n132, n14);
not  g30 (n58, n16);
buf  g31 (n67, n21);
buf  g32 (n106, n21);
buf  g33 (n144, n6);
not  g34 (n140, n15);
buf  g35 (n93, n19);
not  g36 (n121, n17);
not  g37 (n64, n13);
not  g38 (n115, n18);
not  g39 (n130, n20);
buf  g40 (n112, n5);
buf  g41 (n76, n28);
not  g42 (n156, n7);
buf  g43 (n89, n26);
buf  g44 (n87, n7);
buf  g45 (n46, n26);
buf  g46 (n77, n4);
buf  g47 (n33, n14);
buf  g48 (n80, n18);
not  g49 (n151, n32);
buf  g50 (n108, n31);
buf  g51 (n52, n11);
not  g52 (n48, n17);
not  g53 (n36, n26);
buf  g54 (n128, n12);
not  g55 (n65, n20);
not  g56 (n119, n15);
buf  g57 (n102, n7);
buf  g58 (n153, n12);
buf  g59 (n134, n2);
not  g60 (n114, n7);
buf  g61 (n40, n1);
buf  g62 (n94, n20);
buf  g63 (n74, n19);
buf  g64 (n63, n24);
not  g65 (n154, n31);
buf  g66 (n38, n25);
buf  g67 (n43, n15);
not  g68 (n136, n11);
not  g69 (n113, n22);
not  g70 (n42, n21);
buf  g71 (n44, n10);
not  g72 (n133, n8);
not  g73 (n143, n30);
buf  g74 (n85, n31);
not  g75 (n45, n27);
buf  g76 (n81, n16);
buf  g77 (n57, n3);
not  g78 (n104, n4);
buf  g79 (n111, n24);
not  g80 (n95, n14);
buf  g81 (n68, n19);
buf  g82 (n124, n30);
buf  g83 (n34, n17);
buf  g84 (n100, n9);
not  g85 (n105, n28);
not  g86 (n123, n29);
not  g87 (n53, n29);
buf  g88 (n39, n23);
buf  g89 (n139, n1);
buf  g90 (n125, n13);
buf  g91 (n160, n3);
not  g92 (n131, n21);
buf  g93 (n97, n22);
buf  g94 (n122, n4);
buf  g95 (n138, n32);
not  g96 (n127, n23);
buf  g97 (n84, n14);
buf  g98 (n51, n27);
buf  g99 (n117, n3);
not  g100 (n146, n6);
buf  g101 (n149, n5);
buf  g102 (n141, n2);
buf  g103 (n135, n10);
buf  g104 (n83, n20);
buf  g105 (n142, n9);
buf  g106 (n78, n28);
buf  g107 (n75, n12);
not  g108 (n88, n16);
buf  g109 (n54, n29);
not  g110 (n109, n31);
not  g111 (n155, n2);
buf  g112 (n148, n9);
not  g113 (n86, n8);
buf  g114 (n66, n11);
buf  g115 (n118, n19);
buf  g116 (n137, n18);
not  g117 (n91, n9);
not  g118 (n103, n17);
buf  g119 (n70, n5);
not  g120 (n129, n32);
not  g121 (n56, n23);
buf  g122 (n107, n2);
not  g123 (n62, n13);
buf  g124 (n79, n30);
not  g125 (n35, n24);
buf  g126 (n50, n25);
not  g127 (n150, n6);
xor  g128 (n273, n112, n82);
xor  g129 (n274, n115, n33);
and  g130 (n300, n83, n112);
nor  g131 (n180, n99, n41);
or   g132 (n250, n52, n38);
nand g133 (n181, n80, n77);
nand g134 (n230, n46, n114);
and  g135 (n276, n52, n90);
xnor g136 (n196, n62, n94);
or   g137 (n182, n56, n62);
and  g138 (n167, n84, n91);
and  g139 (n322, n60, n56);
and  g140 (n177, n82, n47);
nand g141 (n261, n122, n98);
xor  g142 (n166, n63, n50);
or   g143 (n169, n124, n115);
xor  g144 (n236, n87, n111);
nand g145 (n282, n100, n77);
nand g146 (n279, n33, n106);
and  g147 (n227, n60, n52);
or   g148 (n268, n44, n106);
and  g149 (n319, n65, n104);
xnor g150 (n259, n126, n46);
nor  g151 (n294, n81, n55);
nor  g152 (n246, n57, n118);
xor  g153 (n321, n86, n65);
and  g154 (n216, n35, n67);
nor  g155 (n314, n43, n58);
nor  g156 (n299, n71, n103);
and  g157 (n239, n70, n117);
or   g158 (n281, n72, n94);
and  g159 (n188, n89, n94);
xnor g160 (n211, n47, n41);
nand g161 (n218, n71, n74);
and  g162 (n286, n87, n69);
xnor g163 (n215, n86, n57);
nand g164 (n290, n104, n46);
or   g165 (n317, n39, n93);
nor  g166 (n307, n108, n81);
nand g167 (n219, n107, n44);
and  g168 (n187, n39, n91);
nand g169 (n285, n61, n92);
or   g170 (n217, n105, n107);
and  g171 (n208, n117, n44);
nand g172 (n309, n86, n97);
or   g173 (n170, n85, n114);
or   g174 (n249, n92, n45);
xor  g175 (n207, n48, n106);
xnor g176 (n256, n73, n60);
nand g177 (n210, n122, n40);
nand g178 (n179, n75, n123);
or   g179 (n238, n68, n85);
xor  g180 (n292, n37, n80);
xor  g181 (n265, n117, n85);
xor  g182 (n229, n73, n113);
nand g183 (n185, n96, n121);
or   g184 (n209, n63, n114);
and  g185 (n260, n45, n102);
xor  g186 (n289, n93, n111);
xnor g187 (n320, n110, n72);
xnor g188 (n164, n72, n71);
xnor g189 (n168, n88, n89);
xnor g190 (n172, n110, n34);
nand g191 (n226, n72, n52);
and  g192 (n306, n78, n67);
nor  g193 (n315, n42, n113);
xnor g194 (n271, n42, n57);
nand g195 (n162, n101, n125);
or   g196 (n241, n119, n122);
or   g197 (n225, n63, n100);
xor  g198 (n310, n83, n89);
xnor g199 (n194, n109, n83);
nand g200 (n221, n62, n86);
xor  g201 (n288, n74, n63);
or   g202 (n308, n88, n110);
xor  g203 (n203, n34, n67);
xnor g204 (n272, n61, n59);
and  g205 (n243, n121, n119);
and  g206 (n312, n36, n74);
and  g207 (n264, n123, n57);
xor  g208 (n206, n68, n116);
or   g209 (n298, n76, n98);
xnor g210 (n220, n101, n118);
and  g211 (n201, n45, n41);
and  g212 (n176, n125, n45);
xor  g213 (n174, n40, n125);
and  g214 (n305, n46, n98);
xor  g215 (n235, n40, n64);
nor  g216 (n200, n53, n66);
xor  g217 (n269, n58, n109);
nand g218 (n171, n38, n74);
or   g219 (n297, n82, n33);
and  g220 (n247, n102, n69);
and  g221 (n237, n107, n34);
xor  g222 (n313, n95, n55);
and  g223 (n301, n61, n38);
nor  g224 (n214, n96, n61);
nand g225 (n280, n59, n44);
and  g226 (n202, n66, n64);
xnor g227 (n253, n114, n65);
nor  g228 (n192, n39, n43);
and  g229 (n223, n37, n64);
and  g230 (n296, n104, n91);
xor  g231 (n233, n49, n108);
xnor g232 (n284, n73, n106);
xnor g233 (n163, n35, n78);
nor  g234 (n267, n59, n81);
xor  g235 (n193, n101, n113);
nand g236 (n303, n121, n105);
xor  g237 (n183, n84, n108);
xnor g238 (n266, n124, n66);
and  g239 (n302, n68, n54);
or   g240 (n191, n89, n95);
nor  g241 (n198, n53, n40);
xnor g242 (n224, n116, n124);
and  g243 (n277, n69, n97);
and  g244 (n287, n48, n92);
nor  g245 (n242, n112, n75);
nand g246 (n189, n85, n33);
nand g247 (n254, n79, n120);
xor  g248 (n234, n87, n35);
and  g249 (n190, n119, n51);
xor  g250 (n318, n94, n104);
nand g251 (n255, n93, n109);
or   g252 (n293, n103, n49);
xor  g253 (n197, n43, n41);
or   g254 (n204, n116, n69);
nand g255 (n252, n111, n48);
or   g256 (n199, n77, n103);
and  g257 (n304, n53, n97);
and  g258 (n262, n36, n120);
nor  g259 (n195, n120, n77);
and  g260 (n175, n98, n67);
nor  g261 (n248, n96, n124);
xor  g262 (n283, n60, n113);
xnor g263 (n173, n62, n50);
and  g264 (n311, n56, n108);
nor  g265 (n228, n64, n51);
xor  g266 (n245, n95, n37);
or   g267 (n258, n120, n88);
nor  g268 (n324, n102, n79);
xor  g269 (n232, n42, n107, n80);
xnor g270 (n275, n58, n122, n79, n84);
nand g271 (n295, n118, n79, n73, n65);
xnor g272 (n244, n84, n78, n93, n54);
nor  g273 (n316, n123, n119, n95, n101);
xnor g274 (n205, n103, n97, n105, n70);
xor  g275 (n186, n111, n88, n109, n55);
nor  g276 (n291, n49, n58, n75, n71);
and  g277 (n257, n48, n91, n110, n121);
and  g278 (n240, n70, n117, n99, n76);
or   g279 (n213, n80, n116, n87, n105);
xor  g280 (n212, n100, n54, n112, n102);
nor  g281 (n278, n56, n82, n38, n118);
xnor g282 (n323, n90, n99, n34, n75);
xnor g283 (n231, n83, n37, n81, n59);
and  g284 (n165, n96, n70, n76, n55);
xnor g285 (n222, n68, n125, n76, n54);
and  g286 (n178, n50, n115, n123, n92);
nand g287 (n270, n47, n42, n39, n90);
nand g288 (n161, n90, n49, n66, n36);
or   g289 (n184, n36, n115, n43, n99);
or   g290 (n251, n47, n78, n51, n100);
and  g291 (n263, n35, n50, n53, n51);
not  g292 (n378, n273);
not  g293 (n463, n191);
buf  g294 (n487, n296);
buf  g295 (n349, n224);
not  g296 (n453, n240);
not  g297 (n383, n201);
buf  g298 (n471, n182);
not  g299 (n454, n209);
not  g300 (n413, n278);
not  g301 (n426, n181);
not  g302 (n470, n288);
not  g303 (n412, n264);
buf  g304 (n386, n258);
buf  g305 (n358, n301);
buf  g306 (n340, n284);
not  g307 (n385, n288);
buf  g308 (n356, n244);
nor  g309 (n394, n255, n251);
nand g310 (n434, n269, n248, n196, n216);
and  g311 (n488, n279, n269, n271, n130);
and  g312 (n457, n280, n210, n282, n135);
or   g313 (n384, n225, n218, n242, n164);
xor  g314 (n351, n260, n278, n205);
nor  g315 (n360, n185, n130, n303, n180);
xor  g316 (n331, n258, n228, n131, n213);
or   g317 (n490, n247, n166, n274, n199);
xnor g318 (n414, n275, n289, n204, n128);
xnor g319 (n461, n255, n166, n215, n201);
xnor g320 (n456, n283, n289, n245, n187);
xor  g321 (n432, n205, n273, n202, n210);
nor  g322 (n447, n287, n236, n127, n231);
xor  g323 (n410, n176, n180, n262, n302);
nor  g324 (n326, n133, n194, n192, n280);
nor  g325 (n425, n169, n236, n244, n276);
nand g326 (n407, n260, n183, n217);
xor  g327 (n485, n229, n199, n261, n162);
nand g328 (n422, n179, n168, n250, n212);
or   g329 (n439, n194, n294, n127, n201);
xnor g330 (n477, n272, n254, n245, n191);
xor  g331 (n372, n163, n251, n190, n184);
or   g332 (n436, n280, n246, n216, n263);
nand g333 (n376, n255, n189, n168, n266);
xnor g334 (n474, n232, n248, n161, n164);
xor  g335 (n341, n135, n185, n178, n212);
nand g336 (n330, n294, n255, n170, n285);
nand g337 (n466, n221, n238, n271, n136);
nor  g338 (n444, n299, n166, n195, n256);
or   g339 (n449, n192, n207, n238, n128);
xor  g340 (n409, n275, n228, n206, n291);
xnor g341 (n482, n173, n130, n259, n186);
nand g342 (n411, n276, n233, n249);
and  g343 (n357, n269, n167, n211, n196);
or   g344 (n421, n239, n232, n198, n191);
nor  g345 (n334, n266, n194, n133, n275);
xor  g346 (n364, n136, n252, n267, n246);
nand g347 (n390, n135, n240, n248, n188);
xor  g348 (n445, n301, n184, n203, n226);
xor  g349 (n489, n177, n247, n281, n165);
or   g350 (n345, n182, n216, n208, n244);
nand g351 (n325, n194, n253, n201, n273);
xnor g352 (n440, n132, n185, n218, n281);
xor  g353 (n458, n263, n298, n294, n174);
xnor g354 (n481, n244, n282, n227, n195);
or   g355 (n479, n293, n189, n130, n268);
xor  g356 (n393, n243, n253, n248, n167);
nand g357 (n327, n284, n241, n256, n212);
xnor g358 (n455, n246, n265, n254, n172);
and  g359 (n374, n173, n241, n131, n285);
and  g360 (n430, n263, n203, n235, n282);
xor  g361 (n438, n219, n290, n198, n170);
and  g362 (n337, n174, n169, n286, n186);
nand g363 (n329, n213, n126, n250, n303);
or   g364 (n348, n209, n275, n261, n163);
nor  g365 (n381, n175, n219, n167, n231);
nor  g366 (n361, n227, n242, n204, n129);
and  g367 (n443, n134, n240, n221, n237);
nand g368 (n366, n258, n279, n226, n289);
nor  g369 (n469, n272, n300, n190, n269);
nor  g370 (n419, n210, n178, n177, n252);
xor  g371 (n408, n220, n268, n128, n242);
xnor g372 (n406, n170, n276, n213, n172);
nor  g373 (n465, n224, n281, n285, n193);
xnor g374 (n459, n227, n170, n206, n203);
nor  g375 (n328, n165, n210, n173, n181);
xnor g376 (n452, n250, n220, n134, n200);
xor  g377 (n427, n291, n270, n245, n274);
or   g378 (n442, n193, n172, n195);
or   g379 (n446, n222, n292, n188, n168);
nor  g380 (n377, n181, n293, n162, n183);
nand g381 (n415, n126, n287, n161, n192);
xor  g382 (n342, n223, n207, n175, n229);
xor  g383 (n335, n225, n249, n287, n265);
or   g384 (n365, n128, n230, n182, n129);
nand g385 (n354, n229, n257, n301, n175);
xnor g386 (n382, n176, n214, n204, n233);
xnor g387 (n373, n277, n230, n208, n184);
or   g388 (n450, n260, n188, n258, n223);
nand g389 (n472, n228, n278, n217, n259);
nand g390 (n387, n203, n234, n214, n131);
xor  g391 (n460, n230, n239, n232, n133);
nand g392 (n424, n192, n266, n298, n129);
nand g393 (n401, n302, n250, n221, n256);
nand g394 (n433, n205, n190, n171, n289);
nor  g395 (n346, n178, n207, n165, n209);
xnor g396 (n375, n300, n221, n284, n297);
nor  g397 (n431, n131, n199, n240, n161);
or   g398 (n350, n232, n126, n268, n237);
or   g399 (n429, n259, n164, n222, n162);
or   g400 (n362, n223, n202, n283, n264);
and  g401 (n396, n288, n163, n286, n291);
and  g402 (n451, n197, n296, n283, n247);
and  g403 (n403, n127, n174, n290, n206);
nand g404 (n391, n241, n134, n185, n299);
or   g405 (n435, n177, n271, n163);
or   g406 (n473, n292, n231, n219, n272);
or   g407 (n347, n169, n245, n277, n179);
xor  g408 (n476, n287, n279, n295, n189);
nand g409 (n344, n263, n206, n300, n261);
nor  g410 (n417, n262, n186, n236, n195);
nand g411 (n416, n251, n173, n270, n252);
nor  g412 (n448, n297, n183, n268, n257);
nor  g413 (n486, n270, n225, n175, n299);
nand g414 (n395, n267, n292, n181, n246);
xor  g415 (n338, n187, n234, n238, n243);
nand g416 (n462, n298, n276, n217, n171);
and  g417 (n389, n134, n262, n197, n238);
nor  g418 (n353, n215, n296, n171, n252);
or   g419 (n336, n233, n296, n298, n236);
nand g420 (n428, n212, n198, n174, n264);
or   g421 (n437, n167, n234, n282, n227);
nand g422 (n355, n189, n202, n237, n253);
nor  g423 (n467, n253, n229, n198, n215);
xor  g424 (n370, n135, n292, n274, n171);
and  g425 (n369, n211, n211, n224, n294);
xnor g426 (n398, n290, n265, n165, n247);
and  g427 (n468, n168, n286, n205, n235);
or   g428 (n483, n211, n200, n295, n272);
and  g429 (n359, n230, n196, n200);
xor  g430 (n363, n132, n226, n166, n207);
xnor g431 (n402, n164, n184, n214, n179);
nor  g432 (n423, n277, n213, n267, n182);
xnor g433 (n388, n243, n169, n235, n237);
and  g434 (n405, n228, n266, n187, n265);
and  g435 (n480, n133, n239, n204, n127);
nand g436 (n464, n302, n286, n279, n193);
nand g437 (n399, n257, n262, n270, n225);
and  g438 (n484, n176, n220, n178, n186);
xnor g439 (n397, n299, n235, n233, n188);
and  g440 (n339, n297, n197, n301, n293);
xnor g441 (n392, n177, n241, n231, n216);
xor  g442 (n333, n256, n254, n234, n214);
nor  g443 (n332, n226, n187, n239, n222);
and  g444 (n441, n223, n191, n220, n260);
nand g445 (n379, n215, n293, n300, n190);
nor  g446 (n371, n297, n281, n285, n257);
xor  g447 (n420, n302, n199, n242, n295);
xnor g448 (n475, n129, n288, n208, n274);
xnor g449 (n367, n180, n180, n273, n219);
nand g450 (n400, n291, n222, n161, n218);
and  g451 (n343, n283, n259, n208, n249);
xor  g452 (n352, n218, n209, n132, n295);
nand g453 (n368, n290, n267, n132, n196);
xor  g454 (n478, n197, n280, n251, n254);
nor  g455 (n418, n179, n277, n261, n162);
nand g456 (n380, n264, n176, n284, n224);
nor  g457 (n404, n243, n193, n202, n217);
xnor g458 (n491, n330, n339, n336, n326);
and  g459 (n504, n331, n339, n334, n328);
xor  g460 (n501, n326, n327, n330, n332);
xor  g461 (n493, n338, n331, n341, n333);
and  g462 (n499, n332, n334, n331, n338);
or   g463 (n505, n340, n329, n339);
xor  g464 (n497, n336, n332, n333);
or   g465 (n495, n333, n335, n340);
xnor g466 (n502, n327, n341);
or   g467 (n498, n329, n326, n328, n337);
nand g468 (n500, n330, n334, n335, n331);
nand g469 (n492, n327, n340, n330, n337);
and  g470 (n506, n337, n326, n338);
xnor g471 (n496, n329, n341, n339, n335);
nor  g472 (n494, n334, n328, n337);
nand g473 (n503, n340, n336, n332);
buf  g474 (n509, n496);
buf  g475 (n511, n501);
buf  g476 (n515, n504);
buf  g477 (n512, n497);
buf  g478 (n528, n501);
buf  g479 (n508, n506);
buf  g480 (n524, n493);
buf  g481 (n510, n503);
not  g482 (n514, n502);
buf  g483 (n526, n506);
not  g484 (n518, n505);
not  g485 (n519, n504);
not  g486 (n523, n500);
not  g487 (n507, n491);
buf  g488 (n527, n492);
not  g489 (n522, n495);
buf  g490 (n521, n499);
buf  g491 (n516, n503);
buf  g492 (n513, n502);
buf  g493 (n517, n505);
not  g494 (n525, n494);
not  g495 (n520, n498);
nand g496 (n539, n359, n384, n361, n377);
xnor g497 (n541, n366, n525, n516, n141);
xnor g498 (n578, n352, n364, n513, n142);
nor  g499 (n604, n520, n350, n515, n347);
or   g500 (n582, n523, n521, n364, n385);
xor  g501 (n542, n382, n523, n365, n142);
xnor g502 (n581, n512, n140, n357, n511);
or   g503 (n580, n143, n352, n521, n353);
xor  g504 (n546, n356, n362, n345, n368);
xnor g505 (n571, n374, n381, n369, n520);
or   g506 (n559, n368, n151, n376, n511);
xnor g507 (n577, n526, n362, n146, n350);
xor  g508 (n595, n377, n507, n140, n347);
xor  g509 (n574, n344, n524, n148, n510);
nor  g510 (n566, n375, n508, n140, n520);
xor  g511 (n588, n522, n383, n517, n142);
or   g512 (n589, n136, n150, n382, n377);
or   g513 (n548, n138, n146, n344, n515);
xnor g514 (n600, n375, n371, n342, n142);
xnor g515 (n573, n345, n374, n382, n358);
nor  g516 (n596, n378, n373, n342, n374);
or   g517 (n602, n525, n373, n511, n517);
xor  g518 (n547, n516, n346, n378, n141);
xor  g519 (n556, n518, n526, n350, n381);
xor  g520 (n562, n372, n523, n347, n371);
nor  g521 (n530, n360, n521, n371, n348);
xor  g522 (n572, n507, n150, n526, n370);
and  g523 (n545, n527, n138, n139, n363);
nand g524 (n532, n349, n373, n375, n147);
xor  g525 (n607, n383, n342, n139, n145);
and  g526 (n586, n517, n510, n144, n379);
nor  g527 (n585, n357, n379, n514, n360);
xnor g528 (n557, n149, n152, n145, n513);
or   g529 (n553, n147, n362, n366, n376);
xor  g530 (n584, n151, n380, n385, n508);
nand g531 (n533, n345, n357, n141, n368);
xnor g532 (n540, n513, n152, n144, n524);
and  g533 (n558, n522, n522, n361, n360);
nand g534 (n565, n149, n514, n355, n508);
and  g535 (n603, n380, n348, n346, n507);
and  g536 (n590, n521, n152, n355, n377);
or   g537 (n583, n352, n526, n149, n358);
xnor g538 (n576, n520, n375, n356, n516);
xnor g539 (n606, n145, n363, n376, n349);
nand g540 (n592, n378, n510, n148, n508);
or   g541 (n608, n347, n381, n518, n354);
nor  g542 (n555, n380, n352, n145, n140);
and  g543 (n579, n514, n137, n365, n362);
or   g544 (n598, n354, n371, n382, n343);
xnor g545 (n552, n370, n150, n512, n137);
or   g546 (n550, n146, n374, n345, n381);
xor  g547 (n609, n523, n512, n364, n148);
and  g548 (n531, n525, n144, n346, n343);
nor  g549 (n551, n141, n517, n363, n139);
nor  g550 (n605, n385, n376, n379, n518);
nor  g551 (n594, n510, n366, n351);
nor  g552 (n599, n509, n369, n357, n519);
and  g553 (n568, n370, n151, n384, n380);
and  g554 (n601, n372, n370, n348, n358);
nand g555 (n554, n355, n136, n515, n361);
xor  g556 (n543, n509, n348, n369, n356);
and  g557 (n567, n353, n151, n378, n139);
or   g558 (n538, n153, n137, n372, n356);
or   g559 (n569, n519, n149, n351, n150);
xnor g560 (n570, n519, n346, n518, n359);
or   g561 (n561, n509, n358, n351, n350);
xor  g562 (n537, n367, n524, n355);
or   g563 (n535, n379, n383, n367);
xor  g564 (n597, n148, n384, n138, n519);
xnor g565 (n564, n147, n143, n361, n369);
xor  g566 (n560, n513, n515, n509, n344);
xor  g567 (n544, n516, n144, n368, n143);
nor  g568 (n549, n365, n360, n364, n343);
xor  g569 (n529, n365, n359, n349, n512);
xor  g570 (n587, n511, n351, n514, n138);
or   g571 (n593, n147, n143, n525, n367);
and  g572 (n563, n146, n137, n363, n385);
and  g573 (n591, n367, n522, n353, n384);
xor  g574 (n536, n353, n372, n354, n507);
nor  g575 (n575, n152, n342, n359, n349);
nand g576 (n534, n343, n344, n373, n354);
not  g577 (n624, n574);
buf  g578 (n636, n552);
not  g579 (n685, n570);
buf  g580 (n639, n533);
buf  g581 (n680, n553);
not  g582 (n659, n528);
buf  g583 (n627, n311);
not  g584 (n629, n420);
or   g585 (n679, n403, n562, n429, n425);
xnor g586 (n737, n576, n399, n557, n542);
nand g587 (n697, n571, n405, n569, n418);
xor  g588 (n653, n423, n538, n561, n319);
and  g589 (n692, n542, n319, n404, n153);
and  g590 (n654, n541, n569, n316, n320);
xor  g591 (n700, n530, n427, n155, n408);
or   g592 (n615, n406, n571, n155, n555);
and  g593 (n704, n573, n157, n564, n558);
xnor g594 (n670, n430, n321, n407);
xnor g595 (n610, n321, n533, n547, n426);
xnor g596 (n727, n578, n323, n572, n389);
nand g597 (n613, n569, n413, n540, n318);
and  g598 (n709, n424, n552, n309, n417);
or   g599 (n681, n154, n323, n420, n401);
nand g600 (n663, n318, n321, n315, n409);
and  g601 (n725, n565, n417, n309, n429);
xor  g602 (n626, n156, n414, n399, n548);
and  g603 (n675, n540, n576, n553, n570);
xnor g604 (n733, n552, n393, n426, n391);
and  g605 (n688, n567, n559, n532, n527);
and  g606 (n694, n530, n427, n551, n418);
xnor g607 (n631, n546, n548, n306, n391);
and  g608 (n635, n534, n306, n533, n550);
and  g609 (n650, n547, n566, n306, n549);
xnor g610 (n705, n397, n566, n396, n569);
xnor g611 (n662, n316, n428, n580, n390);
or   g612 (n655, n411, n532, n393, n539);
nand g613 (n721, n431, n529, n560, n538);
and  g614 (n652, n397, n420, n419, n579);
nor  g615 (n728, n554, n546, n529, n310);
nor  g616 (n684, n578, n560, n535, n318);
nand g617 (n634, n578, n406, n537, n309);
and  g618 (n637, n547, n571, n398, n317);
nor  g619 (n646, n568, n531, n416, n408);
and  g620 (n690, n403, n531, n555, n395);
nand g621 (n644, n323, n415, n389, n423);
xnor g622 (n642, n410, n577, n430, n386);
or   g623 (n656, n554, n403, n536, n424);
nand g624 (n730, n154, n407, n320, n315);
nand g625 (n630, n535, n426, n549, n539);
nand g626 (n643, n401, n541, n554, n422);
or   g627 (n726, n574, n303, n539, n552);
nor  g628 (n710, n556, n561, n306, n425);
xnor g629 (n625, n404, n565, n413, n392);
or   g630 (n689, n422, n153, n429, n304);
nor  g631 (n638, n545, n559, n412, n536);
or   g632 (n683, n431, n407, n528, n413);
or   g633 (n723, n315, n551, n402, n400);
xnor g634 (n648, n316, n540, n421, n533);
and  g635 (n686, n402, n393, n430, n406);
and  g636 (n735, n568, n421, n551, n317);
and  g637 (n671, n410, n308, n419, n563);
xnor g638 (n701, n314, n576, n418, n313);
and  g639 (n677, n544, n425, n570, n314);
nand g640 (n687, n546, n317, n388, n556);
nand g641 (n696, n537, n313, n156, n558);
nand g642 (n695, n398, n312, n402, n553);
nand g643 (n693, n153, n155, n577, n311);
nand g644 (n645, n547, n415, n538, n412);
or   g645 (n706, n565, n568, n391, n555);
nor  g646 (n738, n527, n409, n579, n570);
xnor g647 (n658, n428, n558, n539, n531);
nor  g648 (n729, n541, n572, n558, n307);
nor  g649 (n665, n549, n529, n577, n550);
nand g650 (n707, n392, n412, n553, n556);
nor  g651 (n703, n398, n554, n312, n424);
xnor g652 (n673, n394, n304, n534, n423);
xnor g653 (n647, n575, n408, n560, n534);
nand g654 (n660, n154, n308, n557, n420);
and  g655 (n736, n305, n308, n312, n572);
xnor g656 (n708, n395, n317, n387, n562);
or   g657 (n672, n398, n312, n561, n154);
nor  g658 (n611, n536, n397, n405, n411);
nor  g659 (n714, n563, n322, n562, n542);
xnor g660 (n612, n564, n572, n422, n313);
xnor g661 (n712, n396, n386, n417, n401);
or   g662 (n640, n545, n548, n405, n426);
nor  g663 (n702, n557, n573, n571, n544);
or   g664 (n716, n409, n425, n390, n305);
and  g665 (n732, n549, n575, n528, n431);
xnor g666 (n682, n532, n156, n559, n556);
xor  g667 (n657, n419, n565, n395, n403);
nand g668 (n678, n555, n411, n563, n416);
and  g669 (n616, n307, n396, n427, n527);
nor  g670 (n623, n545, n394, n577, n406);
nand g671 (n632, n396, n307, n575, n546);
xor  g672 (n641, n416, n537, n566, n389);
xor  g673 (n731, n395, n404, n580, n305);
xnor g674 (n699, n324, n568, n315, n532);
or   g675 (n619, n562, n404, n388, n544);
nor  g676 (n628, n400, n540, n544, n430);
xor  g677 (n667, n543, n431, n576, n399);
or   g678 (n633, n566, n538, n316, n402);
or   g679 (n691, n543, n387, n559, n310);
nand g680 (n676, n414, n543, n567, n400);
and  g681 (n666, n543, n407, n394, n542);
xor  g682 (n649, n550, n564, n392, n531);
xor  g683 (n614, n310, n319, n416, n389);
xnor g684 (n722, n567, n388, n390, n320);
and  g685 (n720, n415, n412, n541, n319);
and  g686 (n621, n573, n564, n417, n308);
xor  g687 (n661, n535, n423, n529, n307);
nor  g688 (n734, n418, n422, n397, n563);
nand g689 (n664, n427, n311, n415, n303);
xor  g690 (n668, n537, n155, n387, n424);
nor  g691 (n711, n392, n414, n567);
or   g692 (n715, n322, n386, n318, n388);
nor  g693 (n724, n387, n400, n310, n530);
and  g694 (n698, n530, n573, n386, n419);
xor  g695 (n674, n534, n313, n579, n575);
and  g696 (n620, n428, n560, n323, n535);
nand g697 (n713, n391, n401, n428, n390);
xnor g698 (n617, n304, n561, n410, n421);
and  g699 (n618, n393, n574, n309, n408);
xnor g700 (n718, n304, n409, n413, n394);
nand g701 (n651, n156, n320, n574, n548);
xor  g702 (n622, n314, n551, n536, n399);
xor  g703 (n719, n305, n528, n579, n557);
and  g704 (n739, n311, n322, n410, n578);
xor  g705 (n669, n550, n421, n545, n411);
xor  g706 (n717, n314, n405, n429, n322);
nand g707 (n784, n476, n717, n471, n599);
and  g708 (n813, n658, n462, n736, n437);
and  g709 (n824, n619, n478, n615, n584);
nand g710 (n956, n669, n604, n725, n629);
xor  g711 (n918, n679, n159, n718, n651);
nand g712 (n752, n717, n693, n683, n684);
and  g713 (n929, n586, n460, n665, n733);
and  g714 (n838, n682, n646, n457, n664);
and  g715 (n923, n600, n461, n724, n693);
xnor g716 (n879, n665, n444, n659, n607);
and  g717 (n859, n650, n704, n456, n652);
or   g718 (n753, n601, n675, n720, n725);
and  g719 (n863, n721, n478, n581, n714);
xor  g720 (n846, n620, n448, n724, n726);
nand g721 (n827, n450, n725, n625, n443);
or   g722 (n869, n680, n477, n604, n489);
and  g723 (n819, n721, n483, n607, n713);
xnor g724 (n772, n696, n667, n457, n676);
or   g725 (n804, n728, n594, n709, n676);
xnor g726 (n886, n617, n702, n605, n634);
or   g727 (n945, n655, n463, n476, n643);
nor  g728 (n925, n617, n667, n588, n683);
nor  g729 (n820, n485, n721, n690, n583);
nand g730 (n759, n695, n641, n642, n451);
xor  g731 (n877, n606, n682, n635, n704);
and  g732 (n816, n587, n592, n705, n619);
xnor g733 (n791, n593, n616, n454, n601);
nor  g734 (n950, n435, n701, n641, n636);
nand g735 (n740, n597, n632, n662, n681);
xor  g736 (n851, n727, n608, n638, n702);
and  g737 (n912, n657, n633, n732, n157);
xnor g738 (n774, n719, n447, n437, n470);
and  g739 (n832, n722, n688, n643, n697);
and  g740 (n953, n588, n697, n466, n660);
or   g741 (n903, n631, n454, n666, n738);
or   g742 (n823, n622, n720, n624, n672);
or   g743 (n775, n475, n694, n686, n636);
nand g744 (n814, n690, n490, n446, n689);
nand g745 (n907, n451, n590, n719, n685);
xnor g746 (n882, n635, n432, n644, n734);
xnor g747 (n921, n677, n626, n600, n478);
nor  g748 (n788, n471, n598, n490, n673);
nor  g749 (n857, n604, n475, n631, n589);
xor  g750 (n761, n588, n732, n451, n484);
xor  g751 (n856, n645, n484, n728, n480);
xnor g752 (n942, n590, n620, n488, n443);
xor  g753 (n811, n611, n623, n657, n690);
or   g754 (n762, n653, n442, n463, n458);
xor  g755 (n828, n692, n664, n643, n609);
and  g756 (n826, n580, n662, n658, n617);
nor  g757 (n890, n472, n731, n640, n614);
xor  g758 (n944, n613, n433, n472, n597);
or   g759 (n906, n699, n686, n587, n729);
xor  g760 (n871, n598, n730, n639, n695);
nor  g761 (n795, n649, n665, n630, n706);
and  g762 (n936, n463, n607, n731, n643);
nor  g763 (n798, n618, n656, n446, n603);
xnor g764 (n924, n436, n735, n733, n585);
or   g765 (n755, n699, n652, n472, n677);
nand g766 (n872, n698, n159, n662, n605);
nor  g767 (n742, n631, n680, n661, n648);
xnor g768 (n931, n658, n622, n713, n451);
nor  g769 (n844, n585, n669, n735, n639);
xor  g770 (n778, n458, n440, n645, n456);
and  g771 (n951, n481, n690, n487, n594);
nor  g772 (n747, n649, n630, n593, n638);
nand g773 (n852, n652, n473, n470, n589);
xor  g774 (n881, n473, n723, n625, n734);
nand g775 (n917, n675, n660, n640, n635);
xor  g776 (n947, n687, n739, n447, n621);
xor  g777 (n938, n478, n629, n476, n461);
nor  g778 (n803, n472, n648, n602);
nand g779 (n941, n482, n632, n437, n646);
or   g780 (n901, n461, n465, n582, n659);
xor  g781 (n770, n632, n455, n474, n623);
xnor g782 (n905, n461, n488, n730, n669);
nor  g783 (n751, n474, n726, n711, n668);
or   g784 (n922, n708, n710, n722, n467);
xor  g785 (n842, n682, n468, n584, n712);
nand g786 (n861, n608, n678, n696, n433);
and  g787 (n833, n701, n609, n466, n624);
and  g788 (n900, n666, n444, n489, n160);
nand g789 (n948, n675, n606, n637, n670);
nor  g790 (n930, n678, n160, n674, n599);
and  g791 (n949, n434, n696, n453, n645);
xnor g792 (n836, n732, n704, n734, n606);
nand g793 (n760, n716, n698, n679, n673);
xor  g794 (n766, n452, n600, n691, n708);
xnor g795 (n800, n598, n700, n449, n738);
nand g796 (n779, n710, n586, n441, n696);
and  g797 (n777, n455, n441, n629, n703);
nand g798 (n909, n585, n674, n490, n626);
nand g799 (n837, n160, n625, n483);
nor  g800 (n904, n444, n439, n459, n638);
nand g801 (n867, n464, n691, n723, n581);
nand g802 (n815, n469, n605, n738, n636);
xnor g803 (n865, n477, n597, n709, n716);
nor  g804 (n939, n708, n644, n669, n589);
nor  g805 (n932, n718, n440, n714, n583);
xnor g806 (n785, n651, n449, n655, n694);
nand g807 (n749, n606, n432, n730, n677);
and  g808 (n802, n710, n468, n707, n477);
and  g809 (n822, n468, n456, n440, n641);
and  g810 (n748, n703, n453, n434, n432);
xnor g811 (n843, n436, n450, n595, n712);
or   g812 (n792, n627, n485, n452, n474);
and  g813 (n817, n628, n726, n596, n729);
nor  g814 (n758, n700, n158, n716, n602);
nand g815 (n873, n705, n434, n462, n654);
or   g816 (n896, n444, n435, n436, n642);
nor  g817 (n794, n637, n620, n724, n583);
or   g818 (n887, n706, n589, n692, n694);
and  g819 (n864, n657, n682, n640, n590);
nor  g820 (n831, n474, n439, n660, n647);
and  g821 (n916, n450, n596, n672, n693);
or   g822 (n850, n486, n720, n630, n469);
xor  g823 (n952, n157, n728, n717, n442);
and  g824 (n888, n442, n157, n699, n443);
xnor g825 (n889, n653, n678, n679, n623);
xnor g826 (n883, n477, n595, n715, n707);
and  g827 (n809, n628, n702, n686, n637);
xnor g828 (n913, n603, n487, n612, n645);
nand g829 (n899, n698, n715, n473, n686);
or   g830 (n845, n667, n455, n650, n711);
nand g831 (n744, n731, n612, n688, n448);
and  g832 (n866, n593, n703, n483, n449);
or   g833 (n765, n714, n619, n691, n471);
xnor g834 (n825, n588, n615, n159, n694);
xnor g835 (n767, n432, n666, n622, n445);
nor  g836 (n935, n711, n621, n618, n446);
xor  g837 (n875, n734, n460, n674, n727);
nor  g838 (n781, n433, n722, n582, n616);
xor  g839 (n847, n663, n739, n633, n490);
nor  g840 (n898, n608, n688, n698, n596);
xnor g841 (n928, n158, n159, n678, n695);
xor  g842 (n943, n603, n671, n475, n470);
and  g843 (n926, n482, n624, n460, n715);
nor  g844 (n764, n700, n464, n626, n673);
and  g845 (n839, n658, n685, n707, n729);
and  g846 (n745, n654, n158, n597, n467);
nor  g847 (n884, n668, n656, n701, n726);
and  g848 (n915, n458, n663, n709, n731);
and  g849 (n750, n459, n466, n446, n644);
nor  g850 (n920, n656, n609, n708, n685);
xnor g851 (n829, n445, n438, n621, n634);
nand g852 (n893, n651, n719, n725, n652);
or   g853 (n927, n480, n691, n634, n668);
xor  g854 (n911, n622, n706, n650, n671);
or   g855 (n880, n604, n627, n633, n479);
xnor g856 (n937, n650, n685, n480, n590);
and  g857 (n955, n466, n661, n687, n448);
nand g858 (n853, n485, n671, n445, n627);
xor  g859 (n854, n659, n733, n719, n594);
xnor g860 (n754, n489, n467, n628, n692);
nand g861 (n855, n602, n443, n692, n670);
xor  g862 (n946, n587, n663, n601, n651);
or   g863 (n768, n720, n448, n716, n687);
xnor g864 (n796, n469, n591, n624, n482);
xor  g865 (n862, n664, n617, n614, n482);
xnor g866 (n786, n677, n647, n437, n735);
nand g867 (n806, n450, n459, n739, n586);
or   g868 (n858, n592, n605, n632, n736);
xnor g869 (n835, n438, n736, n584, n681);
xor  g870 (n940, n457, n465, n456, n712);
nand g871 (n776, n641, n637, n689, n681);
xnor g872 (n780, n683, n705, n663, n638);
nor  g873 (n849, n462, n598, n656, n438);
xnor g874 (n756, n486, n675, n697, n458);
nand g875 (n810, n667, n724, n647, n661);
nand g876 (n910, n654, n676, n439, n592);
and  g877 (n801, n618, n581, n706, n653);
xor  g878 (n746, n462, n486, n728, n680);
xnor g879 (n790, n619, n487, n479, n488);
nand g880 (n895, n730, n608, n160, n649);
xnor g881 (n773, n704, n665, n584, n657);
xnor g882 (n821, n441, n631, n599, n435);
nand g883 (n805, n666, n591, n627, n435);
nor  g884 (n902, n648, n596, n447, n683);
xnor g885 (n763, n487, n693, n737, n646);
and  g886 (n954, n712, n459, n463, n460);
xnor g887 (n757, n595, n684, n445, n473);
or   g888 (n892, n626, n697, n469, n452);
xnor g889 (n818, n713, n736, n722, n738);
xor  g890 (n897, n727, n486, n737, n464);
nor  g891 (n885, n707, n436, n639, n479);
and  g892 (n782, n587, n453, n684, n702);
and  g893 (n769, n705, n684, n471, n653);
and  g894 (n840, n628, n672, n709, n465);
or   g895 (n812, n648, n636, n618, n735);
and  g896 (n808, n452, n673, n635, n455);
nand g897 (n874, n732, n672, n642, n733);
xnor g898 (n807, n674, n454, n467, n687);
and  g899 (n894, n639, n670, n601, n158);
nor  g900 (n848, n689, n642, n620, n703);
xor  g901 (n876, n649, n655, n454, n464);
nand g902 (n891, n668, n438, n442, n433);
and  g903 (n741, n723, n583, n727, n591);
nor  g904 (n834, n644, n646, n447, n481);
xor  g905 (n934, n721, n713, n470, n623);
and  g906 (n793, n457, n679, n489, n655);
or   g907 (n860, n586, n465, n485, n661);
and  g908 (n919, n441, n449, n599, n592);
or   g909 (n783, n634, n481, n591, n711);
or   g910 (n933, n585, n613, n654, n609);
xnor g911 (n830, n593, n700, n737, n600);
xor  g912 (n957, n681, n710, n715, n714);
xnor g913 (n799, n660, n488, n671, n676);
nor  g914 (n878, n737, n603, n607, n475);
and  g915 (n771, n453, n699, n439, n484);
nand g916 (n797, n594, n580, n595, n582);
and  g917 (n908, n689, n662, n659, n479);
or   g918 (n789, n476, n633, n664, n581);
xor  g919 (n870, n630, n480, n647, n688);
xnor g920 (n868, n670, n625, n629, n484);
nand g921 (n787, n640, n718, n717, n729);
or   g922 (n841, n440, n701, n723, n621);
and  g923 (n743, n468, n434, n718, n582);
and  g924 (n914, n680, n739, n695, n481);
and  g925 (n983, n824, n767, n928, n868);
and  g926 (n979, n799, n895, n893, n952);
xor  g927 (n973, n810, n942, n936, n919);
or   g928 (n960, n842, n807, n778, n918);
nor  g929 (n1013, n814, n782, n945, n948);
nor  g930 (n964, n761, n836, n950, n941);
or   g931 (n971, n780, n932, n917, n774);
nor  g932 (n965, n783, n884, n921, n853);
xor  g933 (n997, n852, n813, n869, n896);
xor  g934 (n989, n792, n885, n907, n944);
nor  g935 (n966, n832, n851, n950, n938);
and  g936 (n975, n882, n881, n771, n891);
nor  g937 (n990, n957, n759, n887, n827);
nor  g938 (n995, n945, n826, n935, n812);
xnor g939 (n976, n776, n809, n946, n784);
or   g940 (n1011, n841, n937, n769, n837);
xor  g941 (n982, n954, n899, n839, n931);
xnor g942 (n1004, n788, n828, n930, n938);
nand g943 (n968, n875, n324, n956, n903);
nor  g944 (n998, n858, n889, n805, n900);
or   g945 (n980, n855, n872, n854, n905);
xnor g946 (n963, n946, n864, n949, n951);
xor  g947 (n999, n927, n867, n877, n796);
or   g948 (n1000, n838, n890, n932, n870);
nor  g949 (n1010, n781, n791, n760, n808);
or   g950 (n981, n862, n848, n786, n873);
xnor g951 (n967, n821, n910, n806, n940);
nand g952 (n986, n772, n789, n757, n324);
nor  g953 (n970, n888, n770, n795, n787);
xor  g954 (n1002, n755, n897, n941, n947);
nor  g955 (n969, n880, n871, n861, n804);
xor  g956 (n988, n816, n773, n825, n785);
xnor g957 (n984, n798, n777, n878, n811);
or   g958 (n978, n925, n765, n764, n833);
and  g959 (n1015, n859, n819, n883, n803);
xnor g960 (n1008, n955, n956, n797, n834);
nor  g961 (n961, n860, n914, n754, n953);
xnor g962 (n991, n840, n763, n911, n944);
or   g963 (n972, n955, n902, n845, n324);
or   g964 (n977, n779, n915, n904, n879);
or   g965 (n996, n857, n892, n898, n913);
or   g966 (n1003, n933, n766, n849, n912);
or   g967 (n974, n934, n802, n758, n943);
nor  g968 (n1007, n909, n957, n906, n937);
nand g969 (n962, n936, n790, n843, n948);
and  g970 (n993, n929, n924, n822, n947);
xor  g971 (n959, n863, n876, n856, n866);
nand g972 (n958, n931, n927, n952, n916);
nor  g973 (n1001, n957, n901, n933, n942);
or   g974 (n985, n847, n823, n835, n886);
xnor g975 (n1017, n926, n844, n831, n928);
nor  g976 (n1009, n939, n954, n850, n957);
nand g977 (n987, n930, n756, n951, n815);
or   g978 (n1006, n768, n920, n940, n846);
and  g979 (n992, n801, n953, n817, n820);
nor  g980 (n1005, n934, n894, n818, n935);
xor  g981 (n1016, n908, n794, n923, n874);
nor  g982 (n1012, n929, n829, n800, n775);
xor  g983 (n1014, n949, n830, n793, n922);
and  g984 (n994, n865, n939, n943, n762);
or   g985 (n1025, n1007, n1003, n981, n982);
nand g986 (n1028, n972, n1002, n975, n971);
and  g987 (n1019, n979, n1006, n994, n985);
nor  g988 (n1030, n1001, n1015, n1010, n966);
xor  g989 (n1032, n973, n987, n1017, n1012);
or   g990 (n1027, n963, n977, n1014, n978);
xnor g991 (n1023, n980, n1008, n961, n988);
and  g992 (n1020, n960, n1004, n1005, n990);
nand g993 (n1024, n1016, n969, n995, n970);
xnor g994 (n1018, n1000, n984, n958, n967);
nor  g995 (n1031, n1009, n976, n991, n999);
nand g996 (n1029, n992, n989, n983, n959);
or   g997 (n1021, n965, n968, n996, n962);
or   g998 (n1026, n986, n1013, n974, n997);
xor  g999 (n1022, n964, n1011, n998, n993);
endmodule
