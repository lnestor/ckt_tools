

module Stat_1000_108
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n983,
  n995,
  n984,
  n974,
  n967,
  n1008,
  n962,
  n965,
  n1015,
  n993,
  n988,
  n981,
  n1003,
  n973,
  n989,
  n970,
  n1021,
  n1029,
  n1025,
  n1023,
  n1026,
  n1032,
  n1022,
  n1020,
  n1027,
  n1017,
  n1024,
  n1030,
  n1019,
  n1018,
  n1028,
  n1031,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  output n983;
  output n995;
  output n984;
  output n974;
  output n967;
  output n1008;
  output n962;
  output n965;
  output n1015;
  output n993;
  output n988;
  output n981;
  output n1003;
  output n973;
  output n989;
  output n970;
  output n1021;
  output n1029;
  output n1025;
  output n1023;
  output n1026;
  output n1032;
  output n1022;
  output n1020;
  output n1027;
  output n1017;
  output n1024;
  output n1030;
  output n1019;
  output n1018;
  output n1028;
  output n1031;
  wire n33;
  wire n34;
  wire n35;
  wire n36;
  wire n37;
  wire n38;
  wire n39;
  wire n40;
  wire n41;
  wire n42;
  wire n43;
  wire n44;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n925;
  wire n926;
  wire n927;
  wire n928;
  wire n929;
  wire n930;
  wire n931;
  wire n932;
  wire n933;
  wire n934;
  wire n935;
  wire n936;
  wire n937;
  wire n938;
  wire n939;
  wire n940;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n963;
  wire n964;
  wire n966;
  wire n968;
  wire n969;
  wire n971;
  wire n972;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n982;
  wire n985;
  wire n986;
  wire n987;
  wire n990;
  wire n991;
  wire n992;
  wire n994;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1016;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyNOTWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyNOTWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyNOTWire_0_15;

  not
  g0
  (
    n138,
    n7
  );


  not
  g1
  (
    n109,
    n13
  );


  buf
  g2
  (
    n79,
    n2
  );


  buf
  g3
  (
    n64,
    n25
  );


  buf
  g4
  (
    n99,
    n25
  );


  not
  g5
  (
    n56,
    n4
  );


  not
  g6
  (
    n67,
    n17
  );


  buf
  g7
  (
    n40,
    n12
  );


  buf
  g8
  (
    n103,
    n2
  );


  buf
  g9
  (
    n121,
    n3
  );


  buf
  g10
  (
    n115,
    n16
  );


  buf
  g11
  (
    n135,
    n11
  );


  not
  g12
  (
    n89,
    n27
  );


  not
  g13
  (
    n52,
    n21
  );


  not
  g14
  (
    n33,
    n17
  );


  not
  g15
  (
    n133,
    n13
  );


  buf
  g16
  (
    KeyWire_0_0,
    n11
  );


  not
  g17
  (
    n119,
    n5
  );


  buf
  g18
  (
    n141,
    n9
  );


  buf
  g19
  (
    n134,
    n20
  );


  not
  g20
  (
    n118,
    n18
  );


  buf
  g21
  (
    n108,
    n15
  );


  not
  g22
  (
    n49,
    n19
  );


  not
  g23
  (
    n57,
    n8
  );


  not
  g24
  (
    n102,
    n7
  );


  not
  g25
  (
    n116,
    n24
  );


  buf
  g26
  (
    n75,
    n10
  );


  buf
  g27
  (
    n36,
    n14
  );


  not
  g28
  (
    n53,
    n1
  );


  buf
  g29
  (
    n94,
    n6
  );


  not
  g30
  (
    n85,
    n22
  );


  buf
  g31
  (
    n107,
    n24
  );


  not
  g32
  (
    n101,
    n15
  );


  buf
  g33
  (
    n58,
    n10
  );


  buf
  g34
  (
    n87,
    n15
  );


  not
  g35
  (
    n143,
    n21
  );


  not
  g36
  (
    n106,
    n14
  );


  not
  g37
  (
    n100,
    n27
  );


  buf
  g38
  (
    n93,
    n26
  );


  not
  g39
  (
    n44,
    n6
  );


  buf
  g40
  (
    n105,
    n18
  );


  not
  g41
  (
    n110,
    n8
  );


  buf
  g42
  (
    n111,
    n22
  );


  buf
  g43
  (
    n77,
    n13
  );


  buf
  g44
  (
    KeyWire_0_12,
    n5
  );


  not
  g45
  (
    n66,
    n2
  );


  buf
  g46
  (
    n139,
    n28
  );


  not
  g47
  (
    n114,
    n17
  );


  not
  g48
  (
    n80,
    n1
  );


  buf
  g49
  (
    n144,
    n25
  );


  not
  g50
  (
    n126,
    n1
  );


  buf
  g51
  (
    n54,
    n16
  );


  buf
  g52
  (
    n86,
    n22
  );


  not
  g53
  (
    n129,
    n23
  );


  not
  g54
  (
    n39,
    n5
  );


  buf
  g55
  (
    n62,
    n10
  );


  not
  g56
  (
    n45,
    n15
  );


  buf
  g57
  (
    n117,
    n24
  );


  not
  g58
  (
    n69,
    n25
  );


  not
  g59
  (
    n124,
    n21
  );


  buf
  g60
  (
    n51,
    n2
  );


  buf
  g61
  (
    n78,
    n26
  );


  not
  g62
  (
    n43,
    n6
  );


  not
  g63
  (
    n55,
    n8
  );


  buf
  g64
  (
    n84,
    n6
  );


  buf
  g65
  (
    n35,
    n18
  );


  buf
  g66
  (
    n73,
    n27
  );


  buf
  g67
  (
    n96,
    n16
  );


  not
  g68
  (
    n104,
    n24
  );


  buf
  g69
  (
    n70,
    n28
  );


  not
  g70
  (
    n81,
    n10
  );


  buf
  g71
  (
    n98,
    n14
  );


  buf
  g72
  (
    n130,
    n22
  );


  buf
  g73
  (
    n38,
    n26
  );


  not
  g74
  (
    n48,
    n3
  );


  not
  g75
  (
    n74,
    n9
  );


  buf
  g76
  (
    n59,
    n3
  );


  buf
  g77
  (
    n92,
    n8
  );


  buf
  g78
  (
    n131,
    n4
  );


  buf
  g79
  (
    n97,
    n17
  );


  not
  g80
  (
    n60,
    n28
  );


  not
  g81
  (
    n65,
    n12
  );


  buf
  g82
  (
    n136,
    n12
  );


  not
  g83
  (
    n132,
    n4
  );


  not
  g84
  (
    n112,
    n12
  );


  not
  g85
  (
    n137,
    n20
  );


  not
  g86
  (
    n91,
    n11
  );


  buf
  g87
  (
    n122,
    n4
  );


  not
  g88
  (
    n127,
    n18
  );


  not
  g89
  (
    n71,
    n13
  );


  buf
  g90
  (
    n95,
    n20
  );


  not
  g91
  (
    n123,
    n19
  );


  not
  g92
  (
    n113,
    n9
  );


  not
  g93
  (
    n42,
    n5
  );


  not
  g94
  (
    n125,
    n14
  );


  not
  g95
  (
    n47,
    n19
  );


  buf
  g96
  (
    n140,
    n21
  );


  not
  g97
  (
    n76,
    n1
  );


  buf
  g98
  (
    KeyWire_0_8,
    n23
  );


  buf
  g99
  (
    n128,
    n11
  );


  not
  g100
  (
    n41,
    n23
  );


  buf
  g101
  (
    n142,
    n9
  );


  buf
  g102
  (
    n72,
    n19
  );


  buf
  g103
  (
    n61,
    n23
  );


  not
  g104
  (
    n63,
    n26
  );


  not
  g105
  (
    n46,
    n20
  );


  buf
  g106
  (
    n120,
    n28
  );


  buf
  g107
  (
    n88,
    n7
  );


  buf
  g108
  (
    n90,
    n16
  );


  not
  g109
  (
    n83,
    n7
  );


  buf
  g110
  (
    n82,
    n27
  );


  not
  g111
  (
    n50,
    n3
  );


  buf
  g112
  (
    n236,
    n56
  );


  buf
  g113
  (
    n201,
    n74
  );


  not
  g114
  (
    n248,
    n58
  );


  not
  g115
  (
    n149,
    n70
  );


  not
  g116
  (
    n309,
    n75
  );


  not
  g117
  (
    n184,
    n36
  );


  buf
  g118
  (
    n209,
    n57
  );


  buf
  g119
  (
    n171,
    n31
  );


  buf
  g120
  (
    n163,
    n71
  );


  buf
  g121
  (
    n237,
    n50
  );


  buf
  g122
  (
    n241,
    n34
  );


  not
  g123
  (
    n294,
    n52
  );


  buf
  g124
  (
    n207,
    n64
  );


  not
  g125
  (
    n316,
    n42
  );


  buf
  g126
  (
    n159,
    n70
  );


  not
  g127
  (
    n203,
    n45
  );


  buf
  g128
  (
    n175,
    n49
  );


  buf
  g129
  (
    n273,
    n39
  );


  not
  g130
  (
    n205,
    n65
  );


  buf
  g131
  (
    n307,
    n60
  );


  not
  g132
  (
    n177,
    n29
  );


  buf
  g133
  (
    n188,
    n66
  );


  not
  g134
  (
    n311,
    n45
  );


  not
  g135
  (
    n225,
    n41
  );


  buf
  g136
  (
    n257,
    n60
  );


  buf
  g137
  (
    n280,
    n62
  );


  not
  g138
  (
    n252,
    n73
  );


  buf
  g139
  (
    n187,
    n56
  );


  buf
  g140
  (
    n238,
    n46
  );


  not
  g141
  (
    n293,
    n61
  );


  not
  g142
  (
    n224,
    n57
  );


  buf
  g143
  (
    n227,
    n37
  );


  not
  g144
  (
    n310,
    n44
  );


  not
  g145
  (
    n290,
    n67
  );


  buf
  g146
  (
    n214,
    n44
  );


  not
  g147
  (
    n189,
    n34
  );


  not
  g148
  (
    n244,
    n51
  );


  not
  g149
  (
    n253,
    n65
  );


  not
  g150
  (
    n314,
    n59
  );


  not
  g151
  (
    n308,
    n50
  );


  buf
  g152
  (
    n176,
    n76
  );


  buf
  g153
  (
    n160,
    n36
  );


  buf
  g154
  (
    n234,
    n44
  );


  buf
  g155
  (
    n165,
    n72
  );


  not
  g156
  (
    n230,
    n33
  );


  not
  g157
  (
    n301,
    n35
  );


  not
  g158
  (
    n212,
    n47
  );


  buf
  g159
  (
    n157,
    n52
  );


  buf
  g160
  (
    n202,
    n30
  );


  buf
  g161
  (
    n170,
    n72
  );


  not
  g162
  (
    n256,
    n59
  );


  not
  g163
  (
    n263,
    n39
  );


  not
  g164
  (
    n276,
    n48
  );


  not
  g165
  (
    n279,
    n61
  );


  not
  g166
  (
    n194,
    n69
  );


  not
  g167
  (
    n216,
    n67
  );


  buf
  g168
  (
    n195,
    n47
  );


  not
  g169
  (
    n180,
    n70
  );


  not
  g170
  (
    n231,
    n53
  );


  not
  g171
  (
    n318,
    n66
  );


  not
  g172
  (
    n199,
    n49
  );


  buf
  g173
  (
    n173,
    n66
  );


  not
  g174
  (
    n261,
    n40
  );


  buf
  g175
  (
    n191,
    n69
  );


  buf
  g176
  (
    n283,
    n68
  );


  buf
  g177
  (
    n197,
    n68
  );


  not
  g178
  (
    n255,
    n38
  );


  not
  g179
  (
    n267,
    n49
  );


  buf
  g180
  (
    n303,
    n37
  );


  not
  g181
  (
    n297,
    n67
  );


  not
  g182
  (
    n218,
    n31
  );


  buf
  g183
  (
    n233,
    n55
  );


  not
  g184
  (
    n295,
    n49
  );


  not
  g185
  (
    n221,
    n30
  );


  not
  g186
  (
    n240,
    n75
  );


  not
  g187
  (
    n287,
    n68
  );


  buf
  g188
  (
    n245,
    n43
  );


  buf
  g189
  (
    n161,
    n34
  );


  not
  g190
  (
    n289,
    n44
  );


  not
  g191
  (
    n152,
    n37
  );


  not
  g192
  (
    n148,
    n63
  );


  buf
  g193
  (
    n223,
    n43
  );


  buf
  g194
  (
    n264,
    n29
  );


  not
  g195
  (
    n243,
    n33
  );


  not
  g196
  (
    n168,
    n55
  );


  buf
  g197
  (
    n247,
    n40
  );


  not
  g198
  (
    n217,
    n74
  );


  buf
  g199
  (
    n196,
    n46
  );


  not
  g200
  (
    n183,
    n39
  );


  buf
  g201
  (
    n271,
    n63
  );


  not
  g202
  (
    n312,
    n47
  );


  not
  g203
  (
    n299,
    n29
  );


  not
  g204
  (
    n185,
    n41
  );


  not
  g205
  (
    n158,
    n42
  );


  not
  g206
  (
    n246,
    n62
  );


  buf
  g207
  (
    n210,
    n62
  );


  buf
  g208
  (
    n304,
    n73
  );


  not
  g209
  (
    n296,
    n40
  );


  not
  g210
  (
    n153,
    n38
  );


  not
  g211
  (
    n292,
    n41
  );


  not
  g212
  (
    n319,
    n60
  );


  not
  g213
  (
    n146,
    n56
  );


  buf
  g214
  (
    n232,
    n33
  );


  not
  g215
  (
    n239,
    n69
  );


  buf
  g216
  (
    n288,
    n64
  );


  not
  g217
  (
    n269,
    n48
  );


  not
  g218
  (
    n154,
    n38
  );


  buf
  g219
  (
    n174,
    n41
  );


  buf
  g220
  (
    n222,
    n71
  );


  not
  g221
  (
    n182,
    n57
  );


  buf
  g222
  (
    n250,
    n35
  );


  buf
  g223
  (
    n274,
    n63
  );


  not
  g224
  (
    KeyWire_0_7,
    n51
  );


  buf
  g225
  (
    n155,
    n58
  );


  not
  g226
  (
    n179,
    n64
  );


  not
  g227
  (
    n249,
    n74
  );


  not
  g228
  (
    n313,
    n58
  );


  not
  g229
  (
    n198,
    n34
  );


  not
  g230
  (
    n254,
    n75
  );


  not
  g231
  (
    n164,
    n76
  );


  not
  g232
  (
    n204,
    n60
  );


  buf
  g233
  (
    n228,
    n52
  );


  not
  g234
  (
    n172,
    n58
  );


  buf
  g235
  (
    n260,
    n55
  );


  not
  g236
  (
    n282,
    n71
  );


  not
  g237
  (
    n285,
    n54
  );


  not
  g238
  (
    n259,
    n33
  );


  not
  g239
  (
    n192,
    n55
  );


  buf
  g240
  (
    n162,
    n59
  );


  not
  g241
  (
    n178,
    n36
  );


  buf
  g242
  (
    n278,
    n69
  );


  buf
  g243
  (
    n169,
    n56
  );


  buf
  g244
  (
    n281,
    n63
  );


  buf
  g245
  (
    n229,
    n54
  );


  not
  g246
  (
    n242,
    n45
  );


  buf
  g247
  (
    n147,
    n50
  );


  not
  g248
  (
    n150,
    n57
  );


  buf
  g249
  (
    n206,
    n66
  );


  not
  g250
  (
    n181,
    n75
  );


  not
  g251
  (
    n235,
    n72
  );


  not
  g252
  (
    n300,
    n48
  );


  not
  g253
  (
    n302,
    n30
  );


  not
  g254
  (
    n272,
    n53
  );


  not
  g255
  (
    n305,
    n73
  );


  buf
  g256
  (
    n298,
    n42
  );


  not
  g257
  (
    n213,
    n53
  );


  buf
  g258
  (
    KeyWire_0_11,
    n61
  );


  buf
  g259
  (
    n275,
    n71
  );


  buf
  g260
  (
    n190,
    n76
  );


  buf
  g261
  (
    n211,
    n48
  );


  buf
  g262
  (
    n186,
    n46
  );


  buf
  g263
  (
    n317,
    n61
  );


  buf
  g264
  (
    n219,
    n35
  );


  not
  g265
  (
    n167,
    n54
  );


  buf
  g266
  (
    n268,
    n51
  );


  not
  g267
  (
    n265,
    n67
  );


  buf
  g268
  (
    n262,
    n62
  );


  not
  g269
  (
    n277,
    n68
  );


  not
  g270
  (
    n215,
    n35
  );


  not
  g271
  (
    n270,
    n29
  );


  not
  g272
  (
    n156,
    n70
  );


  not
  g273
  (
    n258,
    n51
  );


  buf
  g274
  (
    n145,
    n54
  );


  buf
  g275
  (
    n284,
    n46
  );


  buf
  g276
  (
    n266,
    n30
  );


  not
  g277
  (
    n200,
    n53
  );


  not
  g278
  (
    n291,
    n37
  );


  not
  g279
  (
    n226,
    n74
  );


  buf
  g280
  (
    n208,
    n39
  );


  not
  g281
  (
    n251,
    n65
  );


  not
  g282
  (
    n286,
    n31
  );


  xor
  g283
  (
    n306,
    n65,
    n50,
    n47,
    n43
  );


  or
  g284
  (
    n220,
    n38,
    n40,
    n45,
    n64
  );


  and
  g285
  (
    n193,
    n52,
    n42,
    n31,
    n36
  );


  and
  g286
  (
    n315,
    n73,
    n72,
    n43,
    n59
  );


  buf
  g287
  (
    n326,
    n76
  );


  not
  g288
  (
    n340,
    n89
  );


  buf
  g289
  (
    n341,
    n32
  );


  buf
  g290
  (
    n372,
    n82
  );


  buf
  g291
  (
    n373,
    n153
  );


  not
  g292
  (
    n338,
    n79
  );


  not
  g293
  (
    n351,
    n83
  );


  not
  g294
  (
    n357,
    n147
  );


  not
  g295
  (
    n347,
    n148
  );


  buf
  g296
  (
    n324,
    n85
  );


  buf
  g297
  (
    n344,
    n80
  );


  buf
  g298
  (
    n364,
    n147
  );


  buf
  g299
  (
    n366,
    n150
  );


  buf
  g300
  (
    n361,
    n146
  );


  buf
  g301
  (
    n321,
    n80
  );


  buf
  g302
  (
    n348,
    n90
  );


  buf
  g303
  (
    n331,
    n152
  );


  buf
  g304
  (
    n355,
    n148
  );


  not
  g305
  (
    n346,
    n157
  );


  not
  g306
  (
    n328,
    n150
  );


  buf
  g307
  (
    n354,
    n158
  );


  not
  g308
  (
    n369,
    n155
  );


  buf
  g309
  (
    n362,
    n90
  );


  not
  g310
  (
    n332,
    n84
  );


  not
  g311
  (
    n322,
    n87
  );


  not
  g312
  (
    n345,
    n149
  );


  not
  g313
  (
    n367,
    n145
  );


  not
  g314
  (
    n336,
    n152
  );


  not
  g315
  (
    n333,
    n147
  );


  buf
  g316
  (
    n356,
    n87
  );


  buf
  g317
  (
    n334,
    n84
  );


  not
  g318
  (
    n323,
    n88
  );


  not
  g319
  (
    n327,
    n77
  );


  buf
  g320
  (
    n353,
    n83
  );


  xor
  g321
  (
    n339,
    n78,
    n85,
    n157,
    n82
  );


  xor
  g322
  (
    n350,
    n86,
    n85,
    n90,
    n78
  );


  or
  g323
  (
    n370,
    n153,
    n78,
    n149,
    n151
  );


  or
  g324
  (
    n360,
    n152,
    n86,
    n158,
    n154
  );


  nor
  g325
  (
    n337,
    n88,
    n79,
    n146,
    n150
  );


  nor
  g326
  (
    n330,
    n77,
    n79,
    n89,
    n146
  );


  and
  g327
  (
    n329,
    n150,
    n86,
    n148,
    n82
  );


  nand
  g328
  (
    n363,
    n149,
    n156,
    n32,
    n80
  );


  xor
  g329
  (
    n371,
    n85,
    n87,
    n155,
    n156
  );


  xnor
  g330
  (
    n365,
    n151,
    n153,
    n82,
    n32
  );


  xor
  g331
  (
    n352,
    n157,
    n87,
    n84,
    n86
  );


  or
  g332
  (
    n359,
    n156,
    n80,
    n81,
    n153
  );


  nor
  g333
  (
    n342,
    n83,
    n155,
    n88,
    n157
  );


  xnor
  g334
  (
    n358,
    n145,
    n151,
    n79,
    n89
  );


  nand
  g335
  (
    n349,
    n155,
    n146,
    n84,
    n154
  );


  xnor
  g336
  (
    n368,
    n77,
    n32,
    n152,
    n83
  );


  and
  g337
  (
    n320,
    n154,
    n145
  );


  and
  g338
  (
    n343,
    n149,
    n147,
    n81,
    n89
  );


  nand
  g339
  (
    n325,
    n148,
    n77,
    n88,
    n78
  );


  or
  g340
  (
    n335,
    n151,
    n156,
    n81
  );


  nor
  g341
  (
    n392,
    n231,
    n98,
    n286,
    n287
  );


  nor
  g342
  (
    n466,
    n163,
    n367,
    n162,
    n263
  );


  nor
  g343
  (
    n563,
    n252,
    n105,
    n279,
    n221
  );


  xor
  g344
  (
    n494,
    n344,
    n320,
    n208,
    n197
  );


  and
  g345
  (
    n385,
    n187,
    n301,
    n221,
    n322
  );


  nand
  g346
  (
    n401,
    n235,
    n160,
    n90,
    n335
  );


  nor
  g347
  (
    n537,
    n214,
    n338,
    n168,
    n202
  );


  and
  g348
  (
    n398,
    n356,
    n342,
    n159,
    n222
  );


  and
  g349
  (
    KeyWire_0_3,
    n188,
    n363,
    n258,
    n230
  );


  xor
  g350
  (
    n473,
    n242,
    n300,
    n262,
    n299
  );


  nand
  g351
  (
    n582,
    n266,
    n284,
    n228,
    n257
  );


  xnor
  g352
  (
    n439,
    n359,
    n271,
    n246,
    n362
  );


  xor
  g353
  (
    n569,
    n297,
    n358,
    n189,
    n343
  );


  xor
  g354
  (
    n574,
    n256,
    n371,
    n205,
    n234
  );


  nor
  g355
  (
    n374,
    n161,
    n244,
    n238,
    n357
  );


  xor
  g356
  (
    n476,
    n225,
    n221,
    n170,
    n208
  );


  xnor
  g357
  (
    n549,
    n101,
    n333,
    n327,
    n366
  );


  and
  g358
  (
    n532,
    n335,
    n345,
    n185
  );


  xnor
  g359
  (
    n454,
    n293,
    n211,
    n162,
    n183
  );


  or
  g360
  (
    n554,
    n339,
    n234,
    n175,
    n344
  );


  xnor
  g361
  (
    n397,
    n220,
    n341,
    n257,
    n95
  );


  xnor
  g362
  (
    n464,
    n260,
    n293,
    n165,
    n249
  );


  and
  g363
  (
    n526,
    n254,
    n282,
    n189,
    n372
  );


  and
  g364
  (
    n493,
    n92,
    n104,
    n172,
    n325
  );


  xnor
  g365
  (
    n424,
    n265,
    n279,
    n270,
    n367
  );


  or
  g366
  (
    n479,
    n283,
    n216,
    n351,
    n366
  );


  nor
  g367
  (
    n525,
    n273,
    n203,
    n268,
    n289
  );


  xor
  g368
  (
    n390,
    n263,
    n250,
    n99,
    n321
  );


  and
  g369
  (
    n492,
    n286,
    n104,
    n255,
    n222
  );


  nand
  g370
  (
    n465,
    n295,
    n227,
    n324,
    n235
  );


  nor
  g371
  (
    n380,
    n249,
    n373,
    n360,
    n351
  );


  xor
  g372
  (
    n410,
    n277,
    n354,
    n326
  );


  nor
  g373
  (
    n429,
    n176,
    n103,
    n178,
    n274
  );


  nor
  g374
  (
    n388,
    n256,
    n217,
    n227,
    n94
  );


  or
  g375
  (
    n575,
    n240,
    n286,
    n201,
    n190
  );


  nor
  g376
  (
    n520,
    n252,
    n184,
    n201,
    n244
  );


  nand
  g377
  (
    n470,
    n249,
    n176,
    n167,
    n334
  );


  xor
  g378
  (
    n430,
    n344,
    n92,
    n327,
    n196
  );


  xnor
  g379
  (
    KeyWire_0_10,
    n187,
    n204,
    n279,
    n224
  );


  nor
  g380
  (
    n522,
    n206,
    n241,
    n220,
    n356
  );


  xnor
  g381
  (
    n431,
    n358,
    n196,
    n233,
    n212
  );


  xor
  g382
  (
    n440,
    n263,
    n264,
    n239,
    n329
  );


  xnor
  g383
  (
    n584,
    n260,
    n336,
    n178,
    n331
  );


  nor
  g384
  (
    n434,
    n237,
    n202,
    n222,
    n219
  );


  nor
  g385
  (
    KeyWire_0_1,
    n238,
    n96,
    n171,
    n170
  );


  and
  g386
  (
    n571,
    n100,
    n191,
    n371,
    n203
  );


  nor
  g387
  (
    n472,
    n351,
    n192,
    n173,
    n199
  );


  xnor
  g388
  (
    n428,
    n105,
    n247,
    n365,
    n91
  );


  and
  g389
  (
    n435,
    n371,
    n161,
    n207,
    n367
  );


  or
  g390
  (
    KeyWire_0_4,
    n162,
    n170,
    n248,
    n195
  );


  xnor
  g391
  (
    n417,
    n171,
    n355,
    n220,
    n227
  );


  or
  g392
  (
    n394,
    n203,
    n100,
    n209,
    n350
  );


  nor
  g393
  (
    n450,
    n96,
    n237,
    n101,
    n182
  );


  xor
  g394
  (
    n572,
    n172,
    n360,
    n253,
    n273
  );


  xnor
  g395
  (
    n409,
    n186,
    n196,
    n370,
    n177
  );


  xnor
  g396
  (
    n570,
    n176,
    n210,
    n357,
    n213
  );


  nand
  g397
  (
    n540,
    n229,
    n93,
    n365,
    n176
  );


  and
  g398
  (
    n497,
    n165,
    n99,
    n197,
    n181
  );


  xnor
  g399
  (
    n521,
    n188,
    n369,
    n248,
    n95
  );


  xor
  g400
  (
    n421,
    n186,
    n321,
    n161,
    n267
  );


  or
  g401
  (
    n527,
    n352,
    n253,
    n267,
    n167
  );


  nor
  g402
  (
    n416,
    n288,
    n369,
    n229,
    n234
  );


  or
  g403
  (
    n517,
    n270,
    n186,
    n329,
    n350
  );


  nand
  g404
  (
    n391,
    n213,
    n326,
    n246,
    n245
  );


  nand
  g405
  (
    n542,
    n241,
    n104,
    n197,
    n274
  );


  and
  g406
  (
    n523,
    n357,
    n215,
    n206,
    n180
  );


  xor
  g407
  (
    n568,
    n194,
    n179,
    n183,
    n331
  );


  and
  g408
  (
    n487,
    n218,
    n284,
    n246,
    n223
  );


  xor
  g409
  (
    n550,
    n216,
    n234,
    n262,
    n291
  );


  nor
  g410
  (
    n387,
    n362,
    n361,
    n285,
    n298
  );


  or
  g411
  (
    n507,
    n293,
    n346,
    n279,
    n189
  );


  xnor
  g412
  (
    n448,
    n183,
    n260,
    n103,
    n254
  );


  nand
  g413
  (
    n469,
    n338,
    n160,
    n295,
    n353
  );


  nor
  g414
  (
    KeyWire_0_5,
    n373,
    n275,
    n244,
    n247
  );


  or
  g415
  (
    n412,
    n102,
    n102,
    n290,
    n297
  );


  xnor
  g416
  (
    n580,
    n226,
    n328,
    n200,
    n294
  );


  nand
  g417
  (
    n406,
    n106,
    n214,
    n293,
    n345
  );


  or
  g418
  (
    n559,
    n240,
    n205,
    n213,
    n360
  );


  nand
  g419
  (
    n471,
    n182,
    n272,
    n276,
    n246
  );


  xor
  g420
  (
    n558,
    n94,
    n327,
    n188,
    n259
  );


  nor
  g421
  (
    n567,
    n186,
    n211,
    n350,
    n212
  );


  nor
  g422
  (
    n411,
    n359,
    n265,
    n347,
    n276
  );


  and
  g423
  (
    n415,
    n97,
    n353,
    n323
  );


  nor
  g424
  (
    n543,
    n93,
    n320,
    n366,
    n262
  );


  xnor
  g425
  (
    n403,
    n332,
    n348,
    n273,
    n191
  );


  or
  g426
  (
    n395,
    n346,
    n94,
    n248,
    n187
  );


  xor
  g427
  (
    n578,
    n105,
    n261,
    n300
  );


  xnor
  g428
  (
    n566,
    n332,
    n237,
    n290,
    n236
  );


  or
  g429
  (
    n586,
    n301,
    n224,
    n280,
    n294
  );


  xor
  g430
  (
    n452,
    n93,
    n251,
    n165,
    n265
  );


  or
  g431
  (
    n505,
    n269,
    n214,
    n288,
    n171
  );


  nand
  g432
  (
    n478,
    n177,
    n212,
    n240,
    n289
  );


  xnor
  g433
  (
    n519,
    n292,
    n256,
    n96,
    n209
  );


  and
  g434
  (
    n539,
    n201,
    n251,
    n250,
    n180
  );


  xnor
  g435
  (
    n536,
    n289,
    n290,
    n258,
    n340
  );


  xnor
  g436
  (
    n457,
    n193,
    n181,
    n199,
    n368
  );


  nor
  g437
  (
    n474,
    n239,
    n298,
    n178,
    n275
  );


  and
  g438
  (
    n534,
    n346,
    n339,
    n277,
    n329
  );


  nand
  g439
  (
    n538,
    n292,
    n181,
    n320,
    n198
  );


  xnor
  g440
  (
    n496,
    n339,
    n103,
    n98,
    n324
  );


  xnor
  g441
  (
    KeyWire_0_13,
    n224,
    n294,
    n288,
    n166
  );


  xor
  g442
  (
    n477,
    n224,
    n231,
    n256,
    n207
  );


  and
  g443
  (
    n407,
    n183,
    n171,
    n349,
    n282
  );


  xor
  g444
  (
    n425,
    n272,
    n92,
    n239,
    n228
  );


  xnor
  g445
  (
    n515,
    n369,
    n164,
    n322,
    n163
  );


  and
  g446
  (
    n581,
    n349,
    n335,
    n255,
    n269
  );


  xnor
  g447
  (
    n544,
    n91,
    n258,
    n361,
    n286
  );


  and
  g448
  (
    n462,
    n221,
    n210,
    n295,
    n329
  );


  nand
  g449
  (
    n418,
    n179,
    n362,
    n225,
    n175
  );


  nand
  g450
  (
    n502,
    n218,
    n217,
    n258,
    n347
  );


  xor
  g451
  (
    n548,
    n287,
    n164,
    n185,
    n91
  );


  or
  g452
  (
    n447,
    n164,
    n352,
    n185,
    n95
  );


  xnor
  g453
  (
    n486,
    n346,
    n337,
    n267,
    n349
  );


  or
  g454
  (
    n458,
    n344,
    n355,
    n188,
    n321
  );


  or
  g455
  (
    n404,
    n297,
    n247,
    n202,
    n322
  );


  nand
  g456
  (
    n500,
    n252,
    n231,
    n208,
    n326
  );


  xnor
  g457
  (
    n400,
    n219,
    n98,
    n291,
    n184
  );


  nand
  g458
  (
    n378,
    n276,
    n97,
    n334,
    n338
  );


  xnor
  g459
  (
    n432,
    n101,
    n285,
    n358,
    n158
  );


  or
  g460
  (
    n463,
    n217,
    n247,
    n180,
    n271
  );


  nor
  g461
  (
    n459,
    n238,
    n206,
    n174,
    n324
  );


  xnor
  g462
  (
    n451,
    n349,
    n348,
    n193
  );


  and
  g463
  (
    n414,
    n193,
    n323,
    n233,
    n200
  );


  and
  g464
  (
    n511,
    n292,
    n264,
    n174,
    n260
  );


  and
  g465
  (
    n506,
    n205,
    n225,
    n235,
    n105
  );


  or
  g466
  (
    n490,
    n190,
    n272,
    n360,
    n270
  );


  nand
  g467
  (
    n579,
    n162,
    n160,
    n253,
    n191
  );


  xnor
  g468
  (
    n530,
    n177,
    n181,
    n274
  );


  xor
  g469
  (
    n446,
    n192,
    n211,
    n275,
    n330
  );


  and
  g470
  (
    n510,
    n368,
    n354,
    n259,
    n170
  );


  nand
  g471
  (
    n484,
    n180,
    n194,
    n354,
    n284
  );


  nor
  g472
  (
    n485,
    n160,
    n270,
    n198,
    n169
  );


  xor
  g473
  (
    n438,
    n241,
    n333,
    n331,
    n97
  );


  xnor
  g474
  (
    n442,
    n323,
    n253,
    n262,
    n372
  );


  xnor
  g475
  (
    n443,
    n348,
    n242,
    n281,
    n163
  );


  or
  g476
  (
    n528,
    n192,
    n175,
    n216,
    n248
  );


  and
  g477
  (
    n565,
    n207,
    n328,
    n332,
    n354
  );


  xnor
  g478
  (
    n386,
    n223,
    n353,
    n236,
    n102
  );


  or
  g479
  (
    n557,
    n91,
    n226,
    n290,
    n163
  );


  nand
  g480
  (
    n503,
    n268,
    n272,
    n266,
    n365
  );


  or
  g481
  (
    n427,
    n347,
    n284,
    n172,
    n254
  );


  nand
  g482
  (
    n408,
    n300,
    n194,
    n363,
    n100
  );


  xor
  g483
  (
    n545,
    n366,
    n257,
    n294,
    n351
  );


  or
  g484
  (
    n489,
    n343,
    n327,
    n371,
    n97
  );


  nor
  g485
  (
    n501,
    n227,
    n191,
    n352,
    n177
  );


  nor
  g486
  (
    n468,
    n232,
    n341,
    n277,
    n335
  );


  xnor
  g487
  (
    n504,
    n238,
    n173,
    n207,
    n276
  );


  xnor
  g488
  (
    n551,
    n337,
    n261,
    n356,
    n243
  );


  nand
  g489
  (
    n541,
    n363,
    n336,
    n198,
    n261
  );


  xor
  g490
  (
    n512,
    n330,
    n340,
    n215,
    n295
  );


  xnor
  g491
  (
    n455,
    n242,
    n169,
    n283,
    n243
  );


  or
  g492
  (
    n513,
    n209,
    n340,
    n266,
    n252
  );


  and
  g493
  (
    n547,
    n325,
    n250,
    n179,
    n282
  );


  xnor
  g494
  (
    n377,
    n178,
    n300,
    n196,
    n245
  );


  or
  g495
  (
    n482,
    n370,
    n368,
    n166,
    n299
  );


  and
  g496
  (
    n382,
    n218,
    n232,
    n159,
    n211
  );


  nand
  g497
  (
    n585,
    n333,
    n231,
    n165,
    n195
  );


  nor
  g498
  (
    n402,
    n357,
    n277,
    n330
  );


  xnor
  g499
  (
    n381,
    n283,
    n291,
    n200,
    n219
  );


  nor
  g500
  (
    n546,
    n369,
    n159,
    n158,
    n278
  );


  xor
  g501
  (
    n560,
    n265,
    n239,
    n102,
    n220
  );


  nor
  g502
  (
    n552,
    n334,
    n200,
    n251,
    n223
  );


  xnor
  g503
  (
    n467,
    n281,
    n184,
    n208,
    n273
  );


  xnor
  g504
  (
    n524,
    n190,
    n296,
    n269,
    n99
  );


  nor
  g505
  (
    n422,
    n280,
    n103,
    n267,
    n361
  );


  xnor
  g506
  (
    n498,
    n166,
    n331,
    n362,
    n278
  );


  nor
  g507
  (
    n426,
    n226,
    n98,
    n337,
    n336
  );


  or
  g508
  (
    n475,
    n218,
    n259,
    n281,
    n167
  );


  nor
  g509
  (
    n413,
    n356,
    n347,
    n214,
    n199
  );


  or
  g510
  (
    n583,
    n100,
    n343,
    n268,
    n249
  );


  and
  g511
  (
    n531,
    n325,
    n182,
    n280,
    n301
  );


  xor
  g512
  (
    n445,
    n173,
    n264,
    n228,
    n199
  );


  and
  g513
  (
    n576,
    n106,
    n297,
    n202,
    n169
  );


  and
  g514
  (
    n437,
    n350,
    n161,
    n174,
    n324
  );


  nor
  g515
  (
    n379,
    n92,
    n187,
    n245,
    n296
  );


  and
  g516
  (
    n556,
    n189,
    n298,
    n195,
    n179
  );


  xor
  g517
  (
    n514,
    n332,
    n325,
    n172,
    n285
  );


  xor
  g518
  (
    n553,
    n255,
    n225,
    n233,
    n264
  );


  nor
  g519
  (
    n375,
    n278,
    n368,
    n203,
    n230
  );


  nand
  g520
  (
    n499,
    n341,
    n195,
    n372,
    n339
  );


  nor
  g521
  (
    KeyWire_0_9,
    n204,
    n345,
    n283,
    n173
  );


  and
  g522
  (
    n577,
    n287,
    n242,
    n244,
    n229
  );


  nor
  g523
  (
    n495,
    n93,
    n358,
    n359,
    n230
  );


  and
  g524
  (
    n561,
    n323,
    n222,
    n226,
    n223
  );


  xnor
  g525
  (
    n433,
    n237,
    n299,
    n168
  );


  nor
  g526
  (
    n420,
    n219,
    n321,
    n359,
    n236
  );


  or
  g527
  (
    n516,
    n174,
    n182,
    n204,
    n250
  );


  or
  g528
  (
    n376,
    n210,
    n287,
    n340,
    n99
  );


  nand
  g529
  (
    n396,
    n257,
    n328,
    n296,
    n301
  );


  or
  g530
  (
    n384,
    n278,
    n236,
    n167,
    n291
  );


  xnor
  g531
  (
    n488,
    n364,
    n370,
    n210,
    n212
  );


  and
  g532
  (
    n555,
    n364,
    n254,
    n104,
    n245
  );


  and
  g533
  (
    n436,
    n363,
    n296,
    n343,
    n367
  );


  and
  g534
  (
    n562,
    n280,
    n215,
    n201,
    n289
  );


  or
  g535
  (
    n449,
    n364,
    n336,
    n164,
    n361
  );


  and
  g536
  (
    n481,
    n342,
    n240,
    n185,
    n285
  );


  xnor
  g537
  (
    n441,
    n228,
    n204,
    n275,
    n190
  );


  nor
  g538
  (
    n419,
    n230,
    n229,
    n106,
    n266
  );


  xor
  g539
  (
    n405,
    n166,
    n251,
    n193,
    n235
  );


  or
  g540
  (
    n480,
    n355,
    n334,
    n282,
    n106
  );


  nand
  g541
  (
    n508,
    n365,
    n168,
    n328,
    n213
  );


  xnor
  g542
  (
    n453,
    n184,
    n341,
    n271,
    n255
  );


  or
  g543
  (
    n483,
    n232,
    n95,
    n281,
    n259
  );


  nand
  g544
  (
    n535,
    n370,
    n205,
    n337,
    n352
  );


  xor
  g545
  (
    n564,
    n243,
    n192,
    n342,
    n241
  );


  and
  g546
  (
    n389,
    n209,
    n197,
    n96,
    n269
  );


  xor
  g547
  (
    n399,
    n159,
    n263,
    n292,
    n215
  );


  and
  g548
  (
    n393,
    n271,
    n342,
    n338,
    n355
  );


  xor
  g549
  (
    n444,
    n288,
    n243,
    n364,
    n168
  );


  xnor
  g550
  (
    n423,
    n217,
    n268,
    n94,
    n194
  );


  nand
  g551
  (
    n383,
    n175,
    n333,
    n322,
    n233
  );


  and
  g552
  (
    n529,
    n169,
    n232,
    n216,
    n206
  );


  xor
  g553
  (
    n491,
    n198,
    n298,
    n372,
    n101
  );


  and
  g554
  (
    n588,
    n137,
    n123,
    n117,
    n107
  );


  xnor
  g555
  (
    n601,
    n140,
    n303,
    n138,
    n111
  );


  xor
  g556
  (
    n634,
    n141,
    n142,
    n389,
    n388
  );


  nor
  g557
  (
    n626,
    n118,
    n107,
    n378
  );


  nor
  g558
  (
    n631,
    n374,
    n108,
    n139,
    n124
  );


  nand
  g559
  (
    n627,
    n308,
    n379,
    n113,
    n133
  );


  xnor
  g560
  (
    n608,
    n123,
    n136,
    n384
  );


  xor
  g561
  (
    n617,
    n118,
    n130,
    n121,
    n132
  );


  nand
  g562
  (
    n600,
    n109,
    n117,
    n114,
    n144
  );


  xor
  g563
  (
    n611,
    n119,
    n114,
    n115,
    n377
  );


  and
  g564
  (
    n612,
    n383,
    n381,
    n129,
    n387
  );


  xor
  g565
  (
    n591,
    n387,
    n389,
    n132,
    n382
  );


  or
  g566
  (
    n622,
    n141,
    n122,
    n143,
    n134
  );


  or
  g567
  (
    n638,
    n120,
    n113,
    n116
  );


  or
  g568
  (
    n610,
    n373,
    n121,
    n141,
    n143
  );


  xnor
  g569
  (
    n596,
    n117,
    n381,
    n127,
    n302
  );


  and
  g570
  (
    n616,
    n124,
    n390,
    n119,
    n111
  );


  or
  g571
  (
    n615,
    n142,
    n378,
    n130,
    n144
  );


  and
  g572
  (
    n613,
    n142,
    n120,
    n121,
    n375
  );


  xnor
  g573
  (
    n633,
    n380,
    n131,
    n109,
    n140
  );


  nor
  g574
  (
    n614,
    n122,
    n127,
    n125,
    n120
  );


  or
  g575
  (
    n603,
    n139,
    n382,
    n140,
    n129
  );


  and
  g576
  (
    n624,
    n135,
    n304,
    n134
  );


  xnor
  g577
  (
    n595,
    n388,
    n305,
    n375,
    n306
  );


  nor
  g578
  (
    n589,
    n379,
    n125,
    n138,
    n112
  );


  xor
  g579
  (
    n618,
    n111,
    n376,
    n385,
    n108
  );


  nor
  g580
  (
    n597,
    n140,
    n133,
    n387,
    n380
  );


  nor
  g581
  (
    n598,
    n377,
    n116,
    n386,
    n118
  );


  or
  g582
  (
    n635,
    n109,
    n304,
    n137,
    n302
  );


  nor
  g583
  (
    n630,
    n131,
    n112,
    n136,
    n144
  );


  and
  g584
  (
    n628,
    n128,
    n391,
    n118,
    n133
  );


  xor
  g585
  (
    n606,
    n123,
    n133,
    n125,
    n115
  );


  or
  g586
  (
    n623,
    n385,
    n114,
    n374,
    n143
  );


  xor
  g587
  (
    n594,
    n392,
    n393,
    n109,
    n381
  );


  or
  g588
  (
    n599,
    n135,
    n379,
    n386,
    n107
  );


  or
  g589
  (
    n639,
    n302,
    n136,
    n305,
    n385
  );


  nand
  g590
  (
    n625,
    n113,
    n303,
    n115,
    n139
  );


  nor
  g591
  (
    n643,
    n306,
    n134,
    n131,
    n121
  );


  and
  g592
  (
    n632,
    n306,
    n127,
    n108,
    n117
  );


  or
  g593
  (
    n605,
    n122,
    n384,
    n138,
    n391
  );


  nor
  g594
  (
    n641,
    n393,
    n129,
    n144,
    n120
  );


  nand
  g595
  (
    n646,
    n123,
    n134,
    n124,
    n125
  );


  and
  g596
  (
    n590,
    n374,
    n391,
    n305,
    n110
  );


  nand
  g597
  (
    n619,
    n132,
    n128,
    n384,
    n122
  );


  or
  g598
  (
    n609,
    n138,
    n110
  );


  xor
  g599
  (
    n587,
    n137,
    n130,
    n143,
    n111
  );


  and
  g600
  (
    n604,
    n129,
    n141,
    n135,
    n132
  );


  xnor
  g601
  (
    n593,
    n377,
    n130,
    n142,
    n376
  );


  nor
  g602
  (
    n620,
    n373,
    n128,
    n126,
    n107
  );


  nor
  g603
  (
    n621,
    n112,
    n302,
    n392,
    n393
  );


  and
  g604
  (
    n640,
    n306,
    n308,
    n376,
    n139
  );


  nor
  g605
  (
    n602,
    n303,
    n116,
    n392
  );


  and
  g606
  (
    n636,
    n307,
    n390,
    n112,
    n388
  );


  nor
  g607
  (
    n637,
    n137,
    n108,
    n307,
    n126
  );


  or
  g608
  (
    n642,
    n386,
    n380,
    n375,
    n115
  );


  xor
  g609
  (
    n645,
    n127,
    n126,
    n128,
    n114
  );


  xor
  g610
  (
    n607,
    n119,
    n307,
    n124
  );


  or
  g611
  (
    n629,
    n304,
    n383,
    n135,
    n126
  );


  xnor
  g612
  (
    n644,
    n131,
    n119,
    n383,
    n303
  );


  nand
  g613
  (
    n592,
    n389,
    n305,
    n382,
    n390
  );


  nor
  g614
  (
    n689,
    n506,
    n514,
    n641,
    n423
  );


  and
  g615
  (
    n647,
    n471,
    n637,
    n483,
    n486
  );


  and
  g616
  (
    n685,
    n414,
    n513,
    n638,
    n642
  );


  nand
  g617
  (
    n738,
    n473,
    n636,
    n618,
    n489
  );


  and
  g618
  (
    n713,
    n631,
    n474,
    n587,
    n427
  );


  nor
  g619
  (
    n711,
    n515,
    n415,
    n465,
    n495
  );


  xnor
  g620
  (
    n660,
    n466,
    n618,
    n460,
    n424
  );


  and
  g621
  (
    n722,
    n615,
    n458,
    n400,
    n473
  );


  nor
  g622
  (
    n726,
    n403,
    n441,
    n635,
    n447
  );


  xnor
  g623
  (
    n690,
    n628,
    n477,
    n482,
    n509
  );


  nand
  g624
  (
    n661,
    n512,
    n439,
    n508,
    n499
  );


  xnor
  g625
  (
    n762,
    n462,
    n402,
    n638,
    n454
  );


  nand
  g626
  (
    n686,
    n419,
    n504,
    n453,
    n628
  );


  nor
  g627
  (
    n761,
    n644,
    n625,
    n433,
    n426
  );


  or
  g628
  (
    n696,
    n401,
    n453,
    n633,
    n498
  );


  and
  g629
  (
    n694,
    n626,
    n500,
    n408,
    n627
  );


  nor
  g630
  (
    n702,
    n469,
    n631,
    n430,
    n496
  );


  and
  g631
  (
    n718,
    n400,
    n398,
    n639,
    n600
  );


  nand
  g632
  (
    n715,
    n413,
    n616,
    n442,
    n395
  );


  nor
  g633
  (
    n723,
    n466,
    n399,
    n487,
    n451
  );


  xor
  g634
  (
    n719,
    n407,
    n437,
    n462,
    n409
  );


  xor
  g635
  (
    n740,
    n633,
    n436,
    n416,
    n445
  );


  and
  g636
  (
    n763,
    n414,
    n426,
    n646,
    n644
  );


  or
  g637
  (
    n697,
    n464,
    n624,
    n427,
    n404
  );


  or
  g638
  (
    n766,
    n462,
    n641,
    n629,
    n609
  );


  xnor
  g639
  (
    n760,
    n481,
    n464,
    n453,
    n411
  );


  nand
  g640
  (
    n683,
    n632,
    n514,
    n415,
    n399
  );


  xor
  g641
  (
    n649,
    n505,
    n616,
    n633,
    n620
  );


  nor
  g642
  (
    n650,
    n396,
    n405,
    n459,
    n408
  );


  and
  g643
  (
    n730,
    n447,
    n505,
    n469,
    n606
  );


  and
  g644
  (
    n734,
    n607,
    n611,
    n623,
    n429
  );


  xnor
  g645
  (
    n751,
    n412,
    n403,
    n442,
    n404
  );


  nor
  g646
  (
    n669,
    n512,
    n394,
    n631,
    n448
  );


  nor
  g647
  (
    n755,
    n455,
    n634,
    n470,
    n485
  );


  xnor
  g648
  (
    n680,
    n438,
    n417,
    n479,
    n461
  );


  xnor
  g649
  (
    n752,
    n646,
    n625,
    n424,
    n457
  );


  nand
  g650
  (
    n674,
    n490,
    n397,
    n604,
    n488
  );


  or
  g651
  (
    n666,
    n446,
    n591,
    n449,
    n396
  );


  xor
  g652
  (
    n733,
    n481,
    n640,
    n617,
    n509
  );


  and
  g653
  (
    n692,
    n413,
    n494,
    n460,
    n467
  );


  xor
  g654
  (
    n677,
    n418,
    n636,
    n610,
    n406
  );


  or
  g655
  (
    n678,
    n439,
    n623,
    n498,
    n450
  );


  nor
  g656
  (
    n721,
    n416,
    n460,
    n424,
    n643
  );


  or
  g657
  (
    n758,
    n602,
    n507,
    n425,
    n464
  );


  nand
  g658
  (
    n743,
    n494,
    n411,
    n500,
    n432
  );


  and
  g659
  (
    KeyWire_0_14,
    n401,
    n456,
    n511,
    n399
  );


  xor
  g660
  (
    n746,
    n434,
    n645,
    n478,
    n632
  );


  nand
  g661
  (
    n662,
    n430,
    n494,
    n440,
    n638
  );


  xnor
  g662
  (
    n684,
    n501,
    n483,
    n410,
    n403
  );


  and
  g663
  (
    n695,
    n485,
    n476,
    n468,
    n472
  );


  and
  g664
  (
    n732,
    n496,
    n489,
    n446,
    n415
  );


  xnor
  g665
  (
    n672,
    n433,
    n433,
    n506,
    n612
  );


  nand
  g666
  (
    n745,
    n432,
    n476,
    n640,
    n405
  );


  or
  g667
  (
    n741,
    n617,
    n510,
    n469,
    n468
  );


  or
  g668
  (
    n720,
    n482,
    n411,
    n475,
    n445
  );


  nor
  g669
  (
    n705,
    n628,
    n637,
    n435,
    n630
  );


  or
  g670
  (
    n747,
    n465,
    n436,
    n484,
    n430
  );


  nand
  g671
  (
    KeyWire_0_15,
    n452,
    n402,
    n467,
    n438
  );


  xor
  g672
  (
    n664,
    n620,
    n400,
    n452,
    n503
  );


  and
  g673
  (
    n652,
    n497,
    n501,
    n639,
    n398
  );


  xnor
  g674
  (
    n671,
    n511,
    n467,
    n488,
    n624
  );


  and
  g675
  (
    n725,
    n479,
    n444,
    n629,
    n515
  );


  xnor
  g676
  (
    n691,
    n429,
    n420,
    n491,
    n488
  );


  or
  g677
  (
    n765,
    n414,
    n509,
    n504,
    n608
  );


  or
  g678
  (
    n693,
    n613,
    n445,
    n443,
    n601
  );


  and
  g679
  (
    n744,
    n419,
    n479,
    n629,
    n448
  );


  and
  g680
  (
    n703,
    n404,
    n468,
    n642,
    n426
  );


  nand
  g681
  (
    n710,
    n487,
    n486,
    n471,
    n437
  );


  nand
  g682
  (
    n748,
    n508,
    n492,
    n420,
    n619
  );


  nor
  g683
  (
    n735,
    n431,
    n417,
    n461,
    n475
  );


  and
  g684
  (
    n653,
    n407,
    n487,
    n621,
    n425
  );


  or
  g685
  (
    n727,
    n422,
    n516,
    n459,
    n496
  );


  nand
  g686
  (
    n739,
    n605,
    n478,
    n434,
    n410
  );


  and
  g687
  (
    n708,
    n428,
    n484,
    n427,
    n497
  );


  nand
  g688
  (
    n731,
    n594,
    n474,
    n639,
    n499
  );


  xnor
  g689
  (
    n750,
    n516,
    n418,
    n480,
    n417
  );


  nand
  g690
  (
    n756,
    n626,
    n437,
    n413,
    n444
  );


  xnor
  g691
  (
    n757,
    n513,
    n431,
    n593,
    n483
  );


  nor
  g692
  (
    n709,
    n428,
    n412,
    n635,
    n456
  );


  and
  g693
  (
    n728,
    n492,
    n634,
    n420,
    n477
  );


  xor
  g694
  (
    n753,
    n457,
    n472,
    n423,
    n493
  );


  nor
  g695
  (
    n724,
    n441,
    n616,
    n619,
    n463
  );


  xor
  g696
  (
    n673,
    n621,
    n595,
    n603,
    n480
  );


  xor
  g697
  (
    n742,
    n407,
    n406,
    n397
  );


  and
  g698
  (
    KeyWire_0_2,
    n588,
    n421,
    n481,
    n627
  );


  or
  g699
  (
    n670,
    n421,
    n449,
    n644,
    n475
  );


  xnor
  g700
  (
    n736,
    n642,
    n457,
    n500,
    n592
  );


  and
  g701
  (
    n657,
    n508,
    n408,
    n435,
    n422
  );


  xnor
  g702
  (
    n767,
    n416,
    n598,
    n451,
    n432
  );


  or
  g703
  (
    n679,
    n458,
    n491,
    n516,
    n625
  );


  xor
  g704
  (
    n699,
    n503,
    n590,
    n472,
    n597
  );


  xnor
  g705
  (
    n648,
    n514,
    n515,
    n482,
    n440
  );


  xnor
  g706
  (
    n754,
    n495,
    n409,
    n618,
    n643
  );


  and
  g707
  (
    n700,
    n505,
    n476,
    n627,
    n645
  );


  xnor
  g708
  (
    n704,
    n434,
    n645,
    n634,
    n635
  );


  nand
  g709
  (
    n769,
    n495,
    n619,
    n513,
    n493
  );


  nand
  g710
  (
    n681,
    n507,
    n589,
    n614,
    n395
  );


  xor
  g711
  (
    n768,
    n470,
    n492,
    n622,
    n412
  );


  and
  g712
  (
    n682,
    n405,
    n471,
    n502,
    n474
  );


  nor
  g713
  (
    n701,
    n478,
    n466,
    n623,
    n396
  );


  and
  g714
  (
    n712,
    n438,
    n461,
    n501,
    n439
  );


  xor
  g715
  (
    n729,
    n443,
    n410,
    n621,
    n498
  );


  and
  g716
  (
    n749,
    n441,
    n418,
    n463,
    n422
  );


  nand
  g717
  (
    n656,
    n506,
    n452,
    n394,
    n443
  );


  xor
  g718
  (
    n698,
    n401,
    n473,
    n486,
    n429
  );


  xor
  g719
  (
    n716,
    n599,
    n448,
    n491,
    n502
  );


  xnor
  g720
  (
    n668,
    n455,
    n409,
    n450,
    n398
  );


  xnor
  g721
  (
    n759,
    n512,
    n397,
    n626,
    n636
  );


  xor
  g722
  (
    n737,
    n447,
    n622,
    n630
  );


  or
  g723
  (
    n706,
    n449,
    n436,
    n395,
    n402
  );


  or
  g724
  (
    n717,
    n641,
    n503,
    n423,
    n480
  );


  nor
  g725
  (
    n651,
    n394,
    n510,
    n477,
    n490
  );


  nor
  g726
  (
    n658,
    n643,
    n620,
    n617,
    n428
  );


  xor
  g727
  (
    n675,
    n640,
    n507,
    n596,
    n450
  );


  nor
  g728
  (
    n676,
    n630,
    n425,
    n490,
    n470
  );


  nor
  g729
  (
    n655,
    n624,
    n419,
    n463,
    n431
  );


  or
  g730
  (
    n667,
    n510,
    n502,
    n646,
    n485
  );


  and
  g731
  (
    n665,
    n454,
    n465,
    n444,
    n440
  );


  and
  g732
  (
    n714,
    n459,
    n435,
    n504,
    n637
  );


  or
  g733
  (
    n663,
    n455,
    n451,
    n456,
    n632
  );


  or
  g734
  (
    n707,
    n493,
    n489,
    n454,
    n446
  );


  nand
  g735
  (
    n659,
    n458,
    n497,
    n499,
    n646
  );


  and
  g736
  (
    n687,
    n484,
    n442,
    n511,
    n421
  );


  xnor
  g737
  (
    n803,
    n662,
    n652,
    n550,
    n539
  );


  and
  g738
  (
    n786,
    n656,
    n530,
    n544,
    n312
  );


  xnor
  g739
  (
    n770,
    n550,
    n525,
    n542,
    n310
  );


  nand
  g740
  (
    n814,
    n659,
    n309,
    n523,
    n539
  );


  and
  g741
  (
    n798,
    n546,
    n657,
    n522,
    n553
  );


  xor
  g742
  (
    n808,
    n532,
    n531,
    n310,
    n309
  );


  xnor
  g743
  (
    n774,
    n315,
    n546,
    n658,
    n653
  );


  and
  g744
  (
    n818,
    n649,
    n311,
    n543,
    n538
  );


  xnor
  g745
  (
    n797,
    n318,
    n313,
    n517,
    n663
  );


  nor
  g746
  (
    n791,
    n527,
    n656,
    n650,
    n318
  );


  nand
  g747
  (
    n776,
    n314,
    n521,
    n548,
    n522
  );


  nor
  g748
  (
    n813,
    n548,
    n533,
    n524,
    n654
  );


  or
  g749
  (
    n822,
    n551,
    n312,
    n533,
    n660
  );


  xor
  g750
  (
    n821,
    n656,
    n520,
    n527,
    n537
  );


  nand
  g751
  (
    n800,
    n655,
    n316,
    n313,
    n518
  );


  nand
  g752
  (
    n819,
    n317,
    n316,
    n524,
    n526
  );


  xnor
  g753
  (
    n804,
    n552,
    n526,
    n535,
    n524
  );


  xnor
  g754
  (
    n795,
    n534,
    n521,
    n319,
    n529
  );


  xnor
  g755
  (
    n805,
    n540,
    n317,
    n517,
    n664
  );


  nor
  g756
  (
    n809,
    n536,
    n310,
    n552,
    n663
  );


  nor
  g757
  (
    n778,
    n309,
    n553,
    n542,
    n319
  );


  nor
  g758
  (
    n772,
    n554,
    n552,
    n529,
    n541
  );


  nand
  g759
  (
    n801,
    n531,
    n523,
    n537,
    n659
  );


  nand
  g760
  (
    n812,
    n521,
    n314,
    n313,
    n317
  );


  and
  g761
  (
    n815,
    n652,
    n527,
    n651,
    n543
  );


  xor
  g762
  (
    n784,
    n538,
    n530,
    n650,
    n534
  );


  nor
  g763
  (
    n782,
    n311,
    n551,
    n519,
    n663
  );


  xor
  g764
  (
    n806,
    n548,
    n649,
    n523,
    n525
  );


  xnor
  g765
  (
    n777,
    n648,
    n313,
    n658,
    n517
  );


  xor
  g766
  (
    n771,
    n520,
    n549,
    n661,
    n651
  );


  xor
  g767
  (
    n810,
    n315,
    n551,
    n518,
    n664
  );


  xnor
  g768
  (
    n794,
    n547,
    n653,
    n309,
    n540
  );


  or
  g769
  (
    n773,
    n647,
    n545,
    n314,
    n652
  );


  or
  g770
  (
    n817,
    n531,
    n544,
    n519,
    n532
  );


  or
  g771
  (
    n781,
    n650,
    n314,
    n648,
    n536
  );


  nor
  g772
  (
    n799,
    n554,
    n311,
    n661,
    n310
  );


  xor
  g773
  (
    n788,
    n541,
    n537,
    n520,
    n315
  );


  nand
  g774
  (
    n780,
    n528,
    n660,
    n544,
    n522
  );


  xor
  g775
  (
    n787,
    n549,
    n662,
    n539,
    n533
  );


  nand
  g776
  (
    n796,
    n319,
    n316,
    n662,
    n317
  );


  or
  g777
  (
    n775,
    n648,
    n664,
    n532,
    n545
  );


  nand
  g778
  (
    n807,
    n538,
    n655,
    n553,
    n312
  );


  nor
  g779
  (
    n820,
    n655,
    n653,
    n316,
    n312
  );


  xnor
  g780
  (
    n802,
    n651,
    n542,
    n658,
    n545
  );


  xor
  g781
  (
    n792,
    n308,
    n543,
    n525,
    n535
  );


  or
  g782
  (
    n789,
    n536,
    n529,
    n318,
    n550
  );


  xnor
  g783
  (
    n793,
    n649,
    n540,
    n319,
    n530
  );


  and
  g784
  (
    n816,
    n528,
    n547,
    n654,
    n519
  );


  xnor
  g785
  (
    n779,
    n534,
    n654,
    n549,
    n660
  );


  xor
  g786
  (
    n785,
    n535,
    n308,
    n518,
    n657
  );


  xnor
  g787
  (
    n811,
    n659,
    n661,
    n318,
    n528
  );


  xnor
  g788
  (
    n783,
    n657,
    n547,
    n663,
    n541
  );


  xor
  g789
  (
    n790,
    n546,
    n526,
    n315,
    n311
  );


  or
  g790
  (
    n879,
    n756,
    n722,
    n686,
    n735
  );


  or
  g791
  (
    n922,
    n666,
    n667,
    n745,
    n754
  );


  or
  g792
  (
    n849,
    n708,
    n675,
    n792,
    n724
  );


  and
  g793
  (
    n915,
    n787,
    n735,
    n786,
    n716
  );


  nor
  g794
  (
    n888,
    n703,
    n708,
    n810,
    n681
  );


  nand
  g795
  (
    n917,
    n811,
    n687,
    n802,
    n715
  );


  nor
  g796
  (
    n826,
    n698,
    n712,
    n711,
    n741
  );


  xnor
  g797
  (
    n855,
    n700,
    n698,
    n744,
    n799
  );


  xnor
  g798
  (
    n844,
    n797,
    n712,
    n739,
    n702
  );


  xor
  g799
  (
    n851,
    n717,
    n733,
    n689,
    n696
  );


  xor
  g800
  (
    n884,
    n741,
    n694,
    n690,
    n743
  );


  and
  g801
  (
    n839,
    n780,
    n742,
    n665,
    n788
  );


  nand
  g802
  (
    n918,
    n674,
    n797,
    n677,
    n748
  );


  xor
  g803
  (
    n951,
    n731,
    n822,
    n718,
    n805
  );


  xnor
  g804
  (
    n927,
    n796,
    n696,
    n693,
    n677
  );


  or
  g805
  (
    n906,
    n821,
    n682,
    n758,
    n805
  );


  xor
  g806
  (
    n866,
    n781,
    n756,
    n777,
    n740
  );


  nand
  g807
  (
    n882,
    n692,
    n794,
    n755,
    n723
  );


  xnor
  g808
  (
    n897,
    n697,
    n690,
    n692,
    n706
  );


  xnor
  g809
  (
    n824,
    n785,
    n750,
    n682,
    n678
  );


  nor
  g810
  (
    n827,
    n750,
    n739,
    n734,
    n670
  );


  nand
  g811
  (
    n860,
    n707,
    n694,
    n708,
    n716
  );


  xnor
  g812
  (
    n935,
    n807,
    n797,
    n688,
    n668
  );


  and
  g813
  (
    n941,
    n707,
    n729,
    n746,
    n820
  );


  nand
  g814
  (
    n905,
    n778,
    n816,
    n757,
    n722
  );


  or
  g815
  (
    n853,
    n686,
    n758,
    n677,
    n554
  );


  xnor
  g816
  (
    n904,
    n808,
    n685,
    n720,
    n669
  );


  xnor
  g817
  (
    n894,
    n694,
    n714,
    n812,
    n735
  );


  xor
  g818
  (
    n942,
    n725,
    n740,
    n822,
    n732
  );


  nand
  g819
  (
    n889,
    n686,
    n728,
    n802,
    n714
  );


  xor
  g820
  (
    n933,
    n809,
    n679,
    n742
  );


  nor
  g821
  (
    n911,
    n817,
    n807,
    n757,
    n753
  );


  nor
  g822
  (
    n890,
    n748,
    n711,
    n710,
    n707
  );


  xor
  g823
  (
    n937,
    n691,
    n677,
    n741,
    n814
  );


  xnor
  g824
  (
    n925,
    n761,
    n685,
    n759,
    n813
  );


  xor
  g825
  (
    n896,
    n740,
    n770,
    n702,
    n795
  );


  nand
  g826
  (
    n945,
    n692,
    n819,
    n690,
    n801
  );


  nor
  g827
  (
    n847,
    n743,
    n685,
    n681,
    n729
  );


  xnor
  g828
  (
    KeyWire_0_6,
    n800,
    n712,
    n678
  );


  xnor
  g829
  (
    n932,
    n665,
    n753,
    n791,
    n754
  );


  and
  g830
  (
    n944,
    n747,
    n700,
    n816,
    n775
  );


  nor
  g831
  (
    n862,
    n808,
    n667,
    n799,
    n692
  );


  xor
  g832
  (
    n828,
    n806,
    n708,
    n744,
    n805
  );


  nor
  g833
  (
    n833,
    n798,
    n705,
    n714,
    n737
  );


  and
  g834
  (
    n863,
    n752,
    n784,
    n710,
    n727
  );


  or
  g835
  (
    n861,
    n671,
    n743,
    n820,
    n693
  );


  or
  g836
  (
    n881,
    n815,
    n793,
    n666,
    n691
  );


  nand
  g837
  (
    n841,
    n796,
    n683,
    n666,
    n681
  );


  nand
  g838
  (
    n946,
    n738,
    n703,
    n801,
    n748
  );


  nor
  g839
  (
    n876,
    n757,
    n710,
    n693,
    n745
  );


  and
  g840
  (
    n920,
    n786,
    n670,
    n815,
    n725
  );


  nand
  g841
  (
    n830,
    n701,
    n746,
    n814,
    n713
  );


  or
  g842
  (
    n891,
    n711,
    n789,
    n684,
    n822
  );


  nor
  g843
  (
    n899,
    n814,
    n739,
    n785,
    n751
  );


  and
  g844
  (
    n923,
    n734,
    n746,
    n803,
    n679
  );


  xor
  g845
  (
    n865,
    n745,
    n779,
    n737,
    n756
  );


  and
  g846
  (
    n854,
    n705,
    n720,
    n809,
    n678
  );


  nor
  g847
  (
    n910,
    n718,
    n732,
    n706,
    n680
  );


  xnor
  g848
  (
    n936,
    n749,
    n690,
    n724,
    n803
  );


  and
  g849
  (
    n838,
    n671,
    n761,
    n676,
    n701
  );


  xor
  g850
  (
    n872,
    n669,
    n711,
    n792,
    n732
  );


  or
  g851
  (
    n869,
    n821,
    n790,
    n689,
    n753
  );


  and
  g852
  (
    n950,
    n800,
    n730,
    n746,
    n736
  );


  xor
  g853
  (
    n870,
    n700,
    n725,
    n758,
    n670
  );


  nand
  g854
  (
    n850,
    n717,
    n669,
    n674,
    n703
  );


  xor
  g855
  (
    n939,
    n697,
    n817,
    n705,
    n715
  );


  nand
  g856
  (
    n878,
    n666,
    n680,
    n817,
    n750
  );


  or
  g857
  (
    n908,
    n713,
    n749,
    n790,
    n729
  );


  xor
  g858
  (
    n912,
    n721,
    n723,
    n806,
    n755
  );


  and
  g859
  (
    n947,
    n706,
    n678,
    n693,
    n731
  );


  nor
  g860
  (
    n931,
    n796,
    n675,
    n757,
    n722
  );


  nand
  g861
  (
    n914,
    n755,
    n754,
    n813,
    n738
  );


  xor
  g862
  (
    n929,
    n747,
    n799,
    n721,
    n774
  );


  xor
  g863
  (
    n840,
    n679,
    n720,
    n758,
    n773
  );


  xor
  g864
  (
    n864,
    n667,
    n696,
    n689,
    n819
  );


  nand
  g865
  (
    n856,
    n731,
    n810,
    n804,
    n709
  );


  nand
  g866
  (
    n832,
    n725,
    n728,
    n804,
    n760
  );


  nand
  g867
  (
    n877,
    n742,
    n710,
    n782,
    n680
  );


  and
  g868
  (
    n919,
    n760,
    n787,
    n812,
    n815
  );


  xor
  g869
  (
    n940,
    n555,
    n731,
    n719,
    n822
  );


  nor
  g870
  (
    n857,
    n809,
    n751,
    n674,
    n795
  );


  xor
  g871
  (
    n835,
    n668,
    n673,
    n709,
    n719
  );


  and
  g872
  (
    n867,
    n801,
    n695,
    n776,
    n738
  );


  xnor
  g873
  (
    n949,
    n737,
    n730,
    n689,
    n771
  );


  or
  g874
  (
    n837,
    n681,
    n787,
    n798,
    n716
  );


  xor
  g875
  (
    n952,
    n740,
    n687,
    n807,
    n818
  );


  nor
  g876
  (
    n842,
    n783,
    n688,
    n751,
    n744
  );


  nand
  g877
  (
    n825,
    n811,
    n716,
    n726,
    n680
  );


  and
  g878
  (
    n934,
    n697,
    n672,
    n732,
    n727
  );


  nand
  g879
  (
    n913,
    n736,
    n700,
    n750,
    n794
  );


  nand
  g880
  (
    n858,
    n722,
    n713,
    n759,
    n715
  );


  xnor
  g881
  (
    n938,
    n811,
    n709,
    n726,
    n734
  );


  nand
  g882
  (
    n868,
    n791,
    n818,
    n738,
    n671
  );


  xor
  g883
  (
    n901,
    n724,
    n672,
    n703,
    n682
  );


  xnor
  g884
  (
    n880,
    n793,
    n726,
    n665,
    n743
  );


  xnor
  g885
  (
    n895,
    n699,
    n694,
    n715,
    n792
  );


  xnor
  g886
  (
    n916,
    n676,
    n759,
    n679,
    n705
  );


  nand
  g887
  (
    n875,
    n665,
    n749,
    n686,
    n685
  );


  and
  g888
  (
    n898,
    n744,
    n752,
    n719,
    n747
  );


  nor
  g889
  (
    n836,
    n667,
    n727,
    n741,
    n795
  );


  nor
  g890
  (
    n909,
    n816,
    n676,
    n752,
    n727
  );


  or
  g891
  (
    n921,
    n687,
    n721,
    n723,
    n719
  );


  xnor
  g892
  (
    n883,
    n669,
    n818,
    n699,
    n674
  );


  xnor
  g893
  (
    n831,
    n704,
    n760,
    n672,
    n737
  );


  xor
  g894
  (
    n924,
    n745,
    n684,
    n804,
    n736
  );


  and
  g895
  (
    n885,
    n684,
    n717,
    n751,
    n696
  );


  xor
  g896
  (
    n903,
    n709,
    n683,
    n707,
    n736
  );


  xor
  g897
  (
    n874,
    n810,
    n726,
    n683,
    n701
  );


  or
  g898
  (
    n902,
    n675,
    n733,
    n670,
    n739
  );


  and
  g899
  (
    n859,
    n788,
    n793,
    n806,
    n704
  );


  xor
  g900
  (
    n893,
    n794,
    n668,
    n821,
    n747
  );


  or
  g901
  (
    n892,
    n702,
    n812,
    n756,
    n691
  );


  xor
  g902
  (
    n846,
    n717,
    n672,
    n730,
    n706
  );


  xor
  g903
  (
    n900,
    n668,
    n673,
    n555,
    n788
  );


  xor
  g904
  (
    n907,
    n683,
    n753,
    n728,
    n760
  );


  or
  g905
  (
    n871,
    n704,
    n755,
    n688,
    n759
  );


  xor
  g906
  (
    n926,
    n664,
    n728,
    n704,
    n673
  );


  xnor
  g907
  (
    n948,
    n798,
    n718,
    n695,
    n721
  );


  and
  g908
  (
    n829,
    n673,
    n702,
    n688,
    n808
  );


  or
  g909
  (
    n823,
    n682,
    n733,
    n698,
    n752
  );


  and
  g910
  (
    n873,
    n733,
    n803,
    n791,
    n800
  );


  and
  g911
  (
    n928,
    n687,
    n713,
    n730,
    n749
  );


  xor
  g912
  (
    n843,
    n684,
    n734,
    n714,
    n813
  );


  xor
  g913
  (
    n930,
    n675,
    n695,
    n785,
    n697
  );


  nand
  g914
  (
    n943,
    n701,
    n790,
    n720,
    n786
  );


  nor
  g915
  (
    n852,
    n729,
    n698,
    n699,
    n754
  );


  or
  g916
  (
    n845,
    n789,
    n735,
    n819,
    n802
  );


  xor
  g917
  (
    n848,
    n718,
    n691,
    n772,
    n724
  );


  nand
  g918
  (
    n887,
    n820,
    n723,
    n676,
    n695
  );


  and
  g919
  (
    n834,
    n699,
    n789,
    n671,
    n748
  );


  or
  g920
  (
    n986,
    n884,
    n846,
    n575,
    n870
  );


  xnor
  g921
  (
    n981,
    n570,
    n873,
    n574,
    n921
  );


  nand
  g922
  (
    n953,
    n557,
    n876,
    n887,
    n575
  );


  and
  g923
  (
    n977,
    n583,
    n563,
    n561,
    n558
  );


  or
  g924
  (
    n985,
    n569,
    n564,
    n582,
    n907
  );


  and
  g925
  (
    n1016,
    n826,
    n577,
    n845,
    n561
  );


  nor
  g926
  (
    n956,
    n575,
    n581,
    n933,
    n926
  );


  or
  g927
  (
    n976,
    n763,
    n573,
    n909,
    n766
  );


  and
  g928
  (
    n961,
    n901,
    n761,
    n769,
    n763
  );


  and
  g929
  (
    n1015,
    n567,
    n580,
    n857,
    n934
  );


  or
  g930
  (
    n975,
    n881,
    n922,
    n848,
    n912
  );


  xnor
  g931
  (
    n994,
    n880,
    n915,
    n584,
    n823
  );


  xor
  g932
  (
    n968,
    n571,
    n866,
    n556,
    n768
  );


  and
  g933
  (
    n1009,
    n847,
    n856,
    n767,
    n898
  );


  nand
  g934
  (
    n960,
    n904,
    n763,
    n581,
    n906
  );


  xor
  g935
  (
    n969,
    n919,
    n852,
    n854,
    n829
  );


  xor
  g936
  (
    n989,
    n916,
    n562,
    n878,
    n563
  );


  nor
  g937
  (
    n963,
    n570,
    n578,
    n566,
    n894
  );


  xnor
  g938
  (
    n1012,
    n576,
    n902,
    n570,
    n765
  );


  nand
  g939
  (
    n980,
    n929,
    n564,
    n580,
    n882
  );


  xor
  g940
  (
    n990,
    n763,
    n872,
    n889,
    n582
  );


  nand
  g941
  (
    n979,
    n581,
    n762,
    n936,
    n557
  );


  or
  g942
  (
    n1003,
    n890,
    n908,
    n555,
    n586
  );


  xor
  g943
  (
    n971,
    n913,
    n858,
    n865,
    n877
  );


  and
  g944
  (
    n959,
    n874,
    n580,
    n843,
    n892
  );


  and
  g945
  (
    n999,
    n766,
    n838,
    n582,
    n769
  );


  xor
  g946
  (
    n972,
    n769,
    n886,
    n585,
    n861
  );


  or
  g947
  (
    n974,
    n832,
    n840,
    n584,
    n879
  );


  nand
  g948
  (
    n1001,
    n565,
    n580,
    n576,
    n572
  );


  or
  g949
  (
    n962,
    n769,
    n569,
    n911,
    n577
  );


  nand
  g950
  (
    n987,
    n577,
    n825,
    n574,
    n568
  );


  nor
  g951
  (
    n992,
    n585,
    n875,
    n851,
    n841
  );


  xnor
  g952
  (
    n998,
    n586,
    n565,
    n867,
    n561
  );


  nand
  g953
  (
    n1014,
    n566,
    n583,
    n584,
    n850
  );


  or
  g954
  (
    n1010,
    n920,
    n828,
    n765,
    n925
  );


  xor
  g955
  (
    n983,
    n918,
    n842,
    n930,
    n579
  );


  xor
  g956
  (
    n1000,
    n837,
    n849,
    n571,
    n556
  );


  nand
  g957
  (
    n993,
    n768,
    n905,
    n836,
    n834
  );


  and
  g958
  (
    n973,
    n559,
    n869,
    n899,
    n768
  );


  or
  g959
  (
    n1007,
    n917,
    n910,
    n578,
    n927
  );


  or
  g960
  (
    n978,
    n827,
    n833,
    n764,
    n563
  );


  xor
  g961
  (
    n958,
    n575,
    n767,
    n895,
    n853
  );


  or
  g962
  (
    n982,
    n572,
    n762,
    n574,
    n585
  );


  xnor
  g963
  (
    n954,
    n583,
    n900,
    n767,
    n577
  );


  or
  g964
  (
    n1008,
    n839,
    n871,
    n766,
    n562
  );


  and
  g965
  (
    n964,
    n573,
    n558,
    n574,
    n893
  );


  xor
  g966
  (
    n1013,
    n935,
    n585,
    n579,
    n573
  );


  or
  g967
  (
    n1006,
    n560,
    n914,
    n924,
    n764
  );


  xor
  g968
  (
    n984,
    n579,
    n586,
    n565,
    n923
  );


  or
  g969
  (
    n996,
    n557,
    n768,
    n564,
    n576
  );


  xor
  g970
  (
    n995,
    n888,
    n883,
    n859,
    n568
  );


  nand
  g971
  (
    n966,
    n566,
    n568,
    n558,
    n855
  );


  nand
  g972
  (
    n988,
    n560,
    n560,
    n762,
    n582
  );


  and
  g973
  (
    n955,
    n586,
    n862,
    n864,
    n567
  );


  xor
  g974
  (
    n1011,
    n824,
    n559,
    n860,
    n569
  );


  and
  g975
  (
    n1005,
    n830,
    n584,
    n761,
    n767
  );


  and
  g976
  (
    n1002,
    n764,
    n765,
    n932,
    n559
  );


  and
  g977
  (
    n957,
    n903,
    n578,
    n572,
    n579
  );


  or
  g978
  (
    n965,
    n571,
    n891,
    n765,
    n576
  );


  xor
  g979
  (
    n1004,
    n844,
    n931,
    n764,
    n578
  );


  and
  g980
  (
    n991,
    n567,
    n766,
    n573,
    n863
  );


  nor
  g981
  (
    n997,
    n885,
    n581,
    n556,
    n868
  );


  and
  g982
  (
    n970,
    n762,
    n928,
    n562,
    n896
  );


  xor
  g983
  (
    n967,
    n897,
    n835,
    n831,
    n583
  );


  xnor
  g984
  (
    n1029,
    n1009,
    n943,
    n997,
    n972
  );


  xnor
  g985
  (
    n1028,
    n1005,
    n948,
    n940,
    n983
  );


  nand
  g986
  (
    n1021,
    n949,
    n992,
    n985,
    n971
  );


  and
  g987
  (
    n1017,
    n952,
    n1002,
    n1012,
    n1010
  );


  xor
  g988
  (
    n1022,
    n1000,
    n1013,
    n991,
    n1003
  );


  and
  g989
  (
    n1025,
    n947,
    n976,
    n1016,
    n939
  );


  xnor
  g990
  (
    n1024,
    n979,
    n974,
    n1008,
    n998
  );


  xnor
  g991
  (
    n1020,
    n993,
    n975,
    n945,
    n987
  );


  nor
  g992
  (
    n1027,
    n981,
    n951,
    n1015,
    n990
  );


  xor
  g993
  (
    n1023,
    n1001,
    n946,
    n950,
    n984
  );


  xor
  g994
  (
    n1018,
    n977,
    n1004,
    n986,
    n978
  );


  or
  g995
  (
    n1032,
    n1014,
    n982,
    n995,
    n969
  );


  or
  g996
  (
    n1031,
    n996,
    n989,
    n944,
    n988
  );


  and
  g997
  (
    n1019,
    n999,
    n938,
    n942,
    n941
  );


  and
  g998
  (
    n1026,
    n973,
    n994,
    n980,
    n1006
  );


  nor
  g999
  (
    n1030,
    n1011,
    n937,
    n1007,
    n970
  );


  xnor
  KeyGate_0_0
  (
    n34,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n509,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n654,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n460,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n518,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n573,
    KeyNOTWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n886,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n151,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n37,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n533,
    KeyNOTWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n461,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n166,
    KeyNOTWire_0_11
  );


  xor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n68,
    KeyNOTWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    n456,
    keyIn_0_13,
    KeyWire_0_13
  );


  xor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n688,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n764,
    KeyNOTWire_0_15
  );


endmodule

