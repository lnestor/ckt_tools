

module Stat_2540_401
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n33,
  n34,
  n35,
  n36,
  n37,
  n38,
  n39,
  n40,
  n41,
  n42,
  n43,
  n44,
  n940,
  n933,
  n939,
  n937,
  n926,
  n932,
  n938,
  n925,
  n935,
  n936,
  n931,
  n930,
  n929,
  n934,
  n2453,
  n2482,
  n2525,
  n2526,
  n2523,
  n2524,
  n2521,
  n2557,
  n2581,
  n2580,
  n2570,
  n2579,
  n2553,
  n2559,
  n2584,
  n2573,
  n2571,
  n2558,
  n2577,
  n2562,
  n2572,
  n2560,
  n2569,
  n2576,
  n2568,
  n2567,
  n2564,
  n2574,
  n2583,
  n2561,
  n2554,
  n2563,
  n2582,
  n2555,
  n2575,
  n2566,
  n2578,
  n2556,
  n2565,
  keyIn_0_0,
  keyIn_0_1,
  keyIn_0_2,
  keyIn_0_3,
  keyIn_0_4,
  keyIn_0_5,
  keyIn_0_6,
  keyIn_0_7,
  keyIn_0_8,
  keyIn_0_9,
  keyIn_0_10,
  keyIn_0_11,
  keyIn_0_12,
  keyIn_0_13,
  keyIn_0_14,
  keyIn_0_15,
  keyIn_0_16,
  keyIn_0_17,
  keyIn_0_18,
  keyIn_0_19,
  keyIn_0_20,
  keyIn_0_21,
  keyIn_0_22,
  keyIn_0_23,
  keyIn_0_24,
  keyIn_0_25,
  keyIn_0_26,
  keyIn_0_27,
  keyIn_0_28,
  keyIn_0_29,
  keyIn_0_30,
  keyIn_0_31,
  keyIn_0_32,
  keyIn_0_33,
  keyIn_0_34,
  keyIn_0_35,
  keyIn_0_36,
  keyIn_0_37,
  keyIn_0_38,
  keyIn_0_39,
  keyIn_0_40,
  keyIn_0_41,
  keyIn_0_42,
  keyIn_0_43,
  keyIn_0_44,
  keyIn_0_45,
  keyIn_0_46,
  keyIn_0_47,
  keyIn_0_48,
  keyIn_0_49,
  keyIn_0_50,
  keyIn_0_51,
  keyIn_0_52,
  keyIn_0_53,
  keyIn_0_54,
  keyIn_0_55,
  keyIn_0_56,
  keyIn_0_57,
  keyIn_0_58,
  keyIn_0_59,
  keyIn_0_60,
  keyIn_0_61,
  keyIn_0_62,
  keyIn_0_63
);

  input n1;
  input n2;
  input n3;
  input n4;
  input n5;
  input n6;
  input n7;
  input n8;
  input n9;
  input n10;
  input n11;
  input n12;
  input n13;
  input n14;
  input n15;
  input n16;
  input n17;
  input n18;
  input n19;
  input n20;
  input n21;
  input n22;
  input n23;
  input n24;
  input n25;
  input n26;
  input n27;
  input n28;
  input n29;
  input n30;
  input n31;
  input n32;
  input n33;
  input n34;
  input n35;
  input n36;
  input n37;
  input n38;
  input n39;
  input n40;
  input n41;
  input n42;
  input n43;
  input n44;
  input keyIn_0_0;
  input keyIn_0_1;
  input keyIn_0_2;
  input keyIn_0_3;
  input keyIn_0_4;
  input keyIn_0_5;
  input keyIn_0_6;
  input keyIn_0_7;
  input keyIn_0_8;
  input keyIn_0_9;
  input keyIn_0_10;
  input keyIn_0_11;
  input keyIn_0_12;
  input keyIn_0_13;
  input keyIn_0_14;
  input keyIn_0_15;
  input keyIn_0_16;
  input keyIn_0_17;
  input keyIn_0_18;
  input keyIn_0_19;
  input keyIn_0_20;
  input keyIn_0_21;
  input keyIn_0_22;
  input keyIn_0_23;
  input keyIn_0_24;
  input keyIn_0_25;
  input keyIn_0_26;
  input keyIn_0_27;
  input keyIn_0_28;
  input keyIn_0_29;
  input keyIn_0_30;
  input keyIn_0_31;
  input keyIn_0_32;
  input keyIn_0_33;
  input keyIn_0_34;
  input keyIn_0_35;
  input keyIn_0_36;
  input keyIn_0_37;
  input keyIn_0_38;
  input keyIn_0_39;
  input keyIn_0_40;
  input keyIn_0_41;
  input keyIn_0_42;
  input keyIn_0_43;
  input keyIn_0_44;
  input keyIn_0_45;
  input keyIn_0_46;
  input keyIn_0_47;
  input keyIn_0_48;
  input keyIn_0_49;
  input keyIn_0_50;
  input keyIn_0_51;
  input keyIn_0_52;
  input keyIn_0_53;
  input keyIn_0_54;
  input keyIn_0_55;
  input keyIn_0_56;
  input keyIn_0_57;
  input keyIn_0_58;
  input keyIn_0_59;
  input keyIn_0_60;
  input keyIn_0_61;
  input keyIn_0_62;
  input keyIn_0_63;
  output n940;
  output n933;
  output n939;
  output n937;
  output n926;
  output n932;
  output n938;
  output n925;
  output n935;
  output n936;
  output n931;
  output n930;
  output n929;
  output n934;
  output n2453;
  output n2482;
  output n2525;
  output n2526;
  output n2523;
  output n2524;
  output n2521;
  output n2557;
  output n2581;
  output n2580;
  output n2570;
  output n2579;
  output n2553;
  output n2559;
  output n2584;
  output n2573;
  output n2571;
  output n2558;
  output n2577;
  output n2562;
  output n2572;
  output n2560;
  output n2569;
  output n2576;
  output n2568;
  output n2567;
  output n2564;
  output n2574;
  output n2583;
  output n2561;
  output n2554;
  output n2563;
  output n2582;
  output n2555;
  output n2575;
  output n2566;
  output n2578;
  output n2556;
  output n2565;
  wire n45;
  wire n46;
  wire n47;
  wire n48;
  wire n49;
  wire n50;
  wire n51;
  wire n52;
  wire n53;
  wire n54;
  wire n55;
  wire n56;
  wire n57;
  wire n58;
  wire n59;
  wire n60;
  wire n61;
  wire n62;
  wire n63;
  wire n64;
  wire n65;
  wire n66;
  wire n67;
  wire n68;
  wire n69;
  wire n70;
  wire n71;
  wire n72;
  wire n73;
  wire n74;
  wire n75;
  wire n76;
  wire n77;
  wire n78;
  wire n79;
  wire n80;
  wire n81;
  wire n82;
  wire n83;
  wire n84;
  wire n85;
  wire n86;
  wire n87;
  wire n88;
  wire n89;
  wire n90;
  wire n91;
  wire n92;
  wire n93;
  wire n94;
  wire n95;
  wire n96;
  wire n97;
  wire n98;
  wire n99;
  wire n100;
  wire n101;
  wire n102;
  wire n103;
  wire n104;
  wire n105;
  wire n106;
  wire n107;
  wire n108;
  wire n109;
  wire n110;
  wire n111;
  wire n112;
  wire n113;
  wire n114;
  wire n115;
  wire n116;
  wire n117;
  wire n118;
  wire n119;
  wire n120;
  wire n121;
  wire n122;
  wire n123;
  wire n124;
  wire n125;
  wire n126;
  wire n127;
  wire n128;
  wire n129;
  wire n130;
  wire n131;
  wire n132;
  wire n133;
  wire n134;
  wire n135;
  wire n136;
  wire n137;
  wire n138;
  wire n139;
  wire n140;
  wire n141;
  wire n142;
  wire n143;
  wire n144;
  wire n145;
  wire n146;
  wire n147;
  wire n148;
  wire n149;
  wire n150;
  wire n151;
  wire n152;
  wire n153;
  wire n154;
  wire n155;
  wire n156;
  wire n157;
  wire n158;
  wire n159;
  wire n160;
  wire n161;
  wire n162;
  wire n163;
  wire n164;
  wire n165;
  wire n166;
  wire n167;
  wire n168;
  wire n169;
  wire n170;
  wire n171;
  wire n172;
  wire n173;
  wire n174;
  wire n175;
  wire n176;
  wire n177;
  wire n178;
  wire n179;
  wire n180;
  wire n181;
  wire n182;
  wire n183;
  wire n184;
  wire n185;
  wire n186;
  wire n187;
  wire n188;
  wire n189;
  wire n190;
  wire n191;
  wire n192;
  wire n193;
  wire n194;
  wire n195;
  wire n196;
  wire n197;
  wire n198;
  wire n199;
  wire n200;
  wire n201;
  wire n202;
  wire n203;
  wire n204;
  wire n205;
  wire n206;
  wire n207;
  wire n208;
  wire n209;
  wire n210;
  wire n211;
  wire n212;
  wire n213;
  wire n214;
  wire n215;
  wire n216;
  wire n217;
  wire n218;
  wire n219;
  wire n220;
  wire n221;
  wire n222;
  wire n223;
  wire n224;
  wire n225;
  wire n226;
  wire n227;
  wire n228;
  wire n229;
  wire n230;
  wire n231;
  wire n232;
  wire n233;
  wire n234;
  wire n235;
  wire n236;
  wire n237;
  wire n238;
  wire n239;
  wire n240;
  wire n241;
  wire n242;
  wire n243;
  wire n244;
  wire n245;
  wire n246;
  wire n247;
  wire n248;
  wire n249;
  wire n250;
  wire n251;
  wire n252;
  wire n253;
  wire n254;
  wire n255;
  wire n256;
  wire n257;
  wire n258;
  wire n259;
  wire n260;
  wire n261;
  wire n262;
  wire n263;
  wire n264;
  wire n265;
  wire n266;
  wire n267;
  wire n268;
  wire n269;
  wire n270;
  wire n271;
  wire n272;
  wire n273;
  wire n274;
  wire n275;
  wire n276;
  wire n277;
  wire n278;
  wire n279;
  wire n280;
  wire n281;
  wire n282;
  wire n283;
  wire n284;
  wire n285;
  wire n286;
  wire n287;
  wire n288;
  wire n289;
  wire n290;
  wire n291;
  wire n292;
  wire n293;
  wire n294;
  wire n295;
  wire n296;
  wire n297;
  wire n298;
  wire n299;
  wire n300;
  wire n301;
  wire n302;
  wire n303;
  wire n304;
  wire n305;
  wire n306;
  wire n307;
  wire n308;
  wire n309;
  wire n310;
  wire n311;
  wire n312;
  wire n313;
  wire n314;
  wire n315;
  wire n316;
  wire n317;
  wire n318;
  wire n319;
  wire n320;
  wire n321;
  wire n322;
  wire n323;
  wire n324;
  wire n325;
  wire n326;
  wire n327;
  wire n328;
  wire n329;
  wire n330;
  wire n331;
  wire n332;
  wire n333;
  wire n334;
  wire n335;
  wire n336;
  wire n337;
  wire n338;
  wire n339;
  wire n340;
  wire n341;
  wire n342;
  wire n343;
  wire n344;
  wire n345;
  wire n346;
  wire n347;
  wire n348;
  wire n349;
  wire n350;
  wire n351;
  wire n352;
  wire n353;
  wire n354;
  wire n355;
  wire n356;
  wire n357;
  wire n358;
  wire n359;
  wire n360;
  wire n361;
  wire n362;
  wire n363;
  wire n364;
  wire n365;
  wire n366;
  wire n367;
  wire n368;
  wire n369;
  wire n370;
  wire n371;
  wire n372;
  wire n373;
  wire n374;
  wire n375;
  wire n376;
  wire n377;
  wire n378;
  wire n379;
  wire n380;
  wire n381;
  wire n382;
  wire n383;
  wire n384;
  wire n385;
  wire n386;
  wire n387;
  wire n388;
  wire n389;
  wire n390;
  wire n391;
  wire n392;
  wire n393;
  wire n394;
  wire n395;
  wire n396;
  wire n397;
  wire n398;
  wire n399;
  wire n400;
  wire n401;
  wire n402;
  wire n403;
  wire n404;
  wire n405;
  wire n406;
  wire n407;
  wire n408;
  wire n409;
  wire n410;
  wire n411;
  wire n412;
  wire n413;
  wire n414;
  wire n415;
  wire n416;
  wire n417;
  wire n418;
  wire n419;
  wire n420;
  wire n421;
  wire n422;
  wire n423;
  wire n424;
  wire n425;
  wire n426;
  wire n427;
  wire n428;
  wire n429;
  wire n430;
  wire n431;
  wire n432;
  wire n433;
  wire n434;
  wire n435;
  wire n436;
  wire n437;
  wire n438;
  wire n439;
  wire n440;
  wire n441;
  wire n442;
  wire n443;
  wire n444;
  wire n445;
  wire n446;
  wire n447;
  wire n448;
  wire n449;
  wire n450;
  wire n451;
  wire n452;
  wire n453;
  wire n454;
  wire n455;
  wire n456;
  wire n457;
  wire n458;
  wire n459;
  wire n460;
  wire n461;
  wire n462;
  wire n463;
  wire n464;
  wire n465;
  wire n466;
  wire n467;
  wire n468;
  wire n469;
  wire n470;
  wire n471;
  wire n472;
  wire n473;
  wire n474;
  wire n475;
  wire n476;
  wire n477;
  wire n478;
  wire n479;
  wire n480;
  wire n481;
  wire n482;
  wire n483;
  wire n484;
  wire n485;
  wire n486;
  wire n487;
  wire n488;
  wire n489;
  wire n490;
  wire n491;
  wire n492;
  wire n493;
  wire n494;
  wire n495;
  wire n496;
  wire n497;
  wire n498;
  wire n499;
  wire n500;
  wire n501;
  wire n502;
  wire n503;
  wire n504;
  wire n505;
  wire n506;
  wire n507;
  wire n508;
  wire n509;
  wire n510;
  wire n511;
  wire n512;
  wire n513;
  wire n514;
  wire n515;
  wire n516;
  wire n517;
  wire n518;
  wire n519;
  wire n520;
  wire n521;
  wire n522;
  wire n523;
  wire n524;
  wire n525;
  wire n526;
  wire n527;
  wire n528;
  wire n529;
  wire n530;
  wire n531;
  wire n532;
  wire n533;
  wire n534;
  wire n535;
  wire n536;
  wire n537;
  wire n538;
  wire n539;
  wire n540;
  wire n541;
  wire n542;
  wire n543;
  wire n544;
  wire n545;
  wire n546;
  wire n547;
  wire n548;
  wire n549;
  wire n550;
  wire n551;
  wire n552;
  wire n553;
  wire n554;
  wire n555;
  wire n556;
  wire n557;
  wire n558;
  wire n559;
  wire n560;
  wire n561;
  wire n562;
  wire n563;
  wire n564;
  wire n565;
  wire n566;
  wire n567;
  wire n568;
  wire n569;
  wire n570;
  wire n571;
  wire n572;
  wire n573;
  wire n574;
  wire n575;
  wire n576;
  wire n577;
  wire n578;
  wire n579;
  wire n580;
  wire n581;
  wire n582;
  wire n583;
  wire n584;
  wire n585;
  wire n586;
  wire n587;
  wire n588;
  wire n589;
  wire n590;
  wire n591;
  wire n592;
  wire n593;
  wire n594;
  wire n595;
  wire n596;
  wire n597;
  wire n598;
  wire n599;
  wire n600;
  wire n601;
  wire n602;
  wire n603;
  wire n604;
  wire n605;
  wire n606;
  wire n607;
  wire n608;
  wire n609;
  wire n610;
  wire n611;
  wire n612;
  wire n613;
  wire n614;
  wire n615;
  wire n616;
  wire n617;
  wire n618;
  wire n619;
  wire n620;
  wire n621;
  wire n622;
  wire n623;
  wire n624;
  wire n625;
  wire n626;
  wire n627;
  wire n628;
  wire n629;
  wire n630;
  wire n631;
  wire n632;
  wire n633;
  wire n634;
  wire n635;
  wire n636;
  wire n637;
  wire n638;
  wire n639;
  wire n640;
  wire n641;
  wire n642;
  wire n643;
  wire n644;
  wire n645;
  wire n646;
  wire n647;
  wire n648;
  wire n649;
  wire n650;
  wire n651;
  wire n652;
  wire n653;
  wire n654;
  wire n655;
  wire n656;
  wire n657;
  wire n658;
  wire n659;
  wire n660;
  wire n661;
  wire n662;
  wire n663;
  wire n664;
  wire n665;
  wire n666;
  wire n667;
  wire n668;
  wire n669;
  wire n670;
  wire n671;
  wire n672;
  wire n673;
  wire n674;
  wire n675;
  wire n676;
  wire n677;
  wire n678;
  wire n679;
  wire n680;
  wire n681;
  wire n682;
  wire n683;
  wire n684;
  wire n685;
  wire n686;
  wire n687;
  wire n688;
  wire n689;
  wire n690;
  wire n691;
  wire n692;
  wire n693;
  wire n694;
  wire n695;
  wire n696;
  wire n697;
  wire n698;
  wire n699;
  wire n700;
  wire n701;
  wire n702;
  wire n703;
  wire n704;
  wire n705;
  wire n706;
  wire n707;
  wire n708;
  wire n709;
  wire n710;
  wire n711;
  wire n712;
  wire n713;
  wire n714;
  wire n715;
  wire n716;
  wire n717;
  wire n718;
  wire n719;
  wire n720;
  wire n721;
  wire n722;
  wire n723;
  wire n724;
  wire n725;
  wire n726;
  wire n727;
  wire n728;
  wire n729;
  wire n730;
  wire n731;
  wire n732;
  wire n733;
  wire n734;
  wire n735;
  wire n736;
  wire n737;
  wire n738;
  wire n739;
  wire n740;
  wire n741;
  wire n742;
  wire n743;
  wire n744;
  wire n745;
  wire n746;
  wire n747;
  wire n748;
  wire n749;
  wire n750;
  wire n751;
  wire n752;
  wire n753;
  wire n754;
  wire n755;
  wire n756;
  wire n757;
  wire n758;
  wire n759;
  wire n760;
  wire n761;
  wire n762;
  wire n763;
  wire n764;
  wire n765;
  wire n766;
  wire n767;
  wire n768;
  wire n769;
  wire n770;
  wire n771;
  wire n772;
  wire n773;
  wire n774;
  wire n775;
  wire n776;
  wire n777;
  wire n778;
  wire n779;
  wire n780;
  wire n781;
  wire n782;
  wire n783;
  wire n784;
  wire n785;
  wire n786;
  wire n787;
  wire n788;
  wire n789;
  wire n790;
  wire n791;
  wire n792;
  wire n793;
  wire n794;
  wire n795;
  wire n796;
  wire n797;
  wire n798;
  wire n799;
  wire n800;
  wire n801;
  wire n802;
  wire n803;
  wire n804;
  wire n805;
  wire n806;
  wire n807;
  wire n808;
  wire n809;
  wire n810;
  wire n811;
  wire n812;
  wire n813;
  wire n814;
  wire n815;
  wire n816;
  wire n817;
  wire n818;
  wire n819;
  wire n820;
  wire n821;
  wire n822;
  wire n823;
  wire n824;
  wire n825;
  wire n826;
  wire n827;
  wire n828;
  wire n829;
  wire n830;
  wire n831;
  wire n832;
  wire n833;
  wire n834;
  wire n835;
  wire n836;
  wire n837;
  wire n838;
  wire n839;
  wire n840;
  wire n841;
  wire n842;
  wire n843;
  wire n844;
  wire n845;
  wire n846;
  wire n847;
  wire n848;
  wire n849;
  wire n850;
  wire n851;
  wire n852;
  wire n853;
  wire n854;
  wire n855;
  wire n856;
  wire n857;
  wire n858;
  wire n859;
  wire n860;
  wire n861;
  wire n862;
  wire n863;
  wire n864;
  wire n865;
  wire n866;
  wire n867;
  wire n868;
  wire n869;
  wire n870;
  wire n871;
  wire n872;
  wire n873;
  wire n874;
  wire n875;
  wire n876;
  wire n877;
  wire n878;
  wire n879;
  wire n880;
  wire n881;
  wire n882;
  wire n883;
  wire n884;
  wire n885;
  wire n886;
  wire n887;
  wire n888;
  wire n889;
  wire n890;
  wire n891;
  wire n892;
  wire n893;
  wire n894;
  wire n895;
  wire n896;
  wire n897;
  wire n898;
  wire n899;
  wire n900;
  wire n901;
  wire n902;
  wire n903;
  wire n904;
  wire n905;
  wire n906;
  wire n907;
  wire n908;
  wire n909;
  wire n910;
  wire n911;
  wire n912;
  wire n913;
  wire n914;
  wire n915;
  wire n916;
  wire n917;
  wire n918;
  wire n919;
  wire n920;
  wire n921;
  wire n922;
  wire n923;
  wire n924;
  wire n927;
  wire n928;
  wire n941;
  wire n942;
  wire n943;
  wire n944;
  wire n945;
  wire n946;
  wire n947;
  wire n948;
  wire n949;
  wire n950;
  wire n951;
  wire n952;
  wire n953;
  wire n954;
  wire n955;
  wire n956;
  wire n957;
  wire n958;
  wire n959;
  wire n960;
  wire n961;
  wire n962;
  wire n963;
  wire n964;
  wire n965;
  wire n966;
  wire n967;
  wire n968;
  wire n969;
  wire n970;
  wire n971;
  wire n972;
  wire n973;
  wire n974;
  wire n975;
  wire n976;
  wire n977;
  wire n978;
  wire n979;
  wire n980;
  wire n981;
  wire n982;
  wire n983;
  wire n984;
  wire n985;
  wire n986;
  wire n987;
  wire n988;
  wire n989;
  wire n990;
  wire n991;
  wire n992;
  wire n993;
  wire n994;
  wire n995;
  wire n996;
  wire n997;
  wire n998;
  wire n999;
  wire n1000;
  wire n1001;
  wire n1002;
  wire n1003;
  wire n1004;
  wire n1005;
  wire n1006;
  wire n1007;
  wire n1008;
  wire n1009;
  wire n1010;
  wire n1011;
  wire n1012;
  wire n1013;
  wire n1014;
  wire n1015;
  wire n1016;
  wire n1017;
  wire n1018;
  wire n1019;
  wire n1020;
  wire n1021;
  wire n1022;
  wire n1023;
  wire n1024;
  wire n1025;
  wire n1026;
  wire n1027;
  wire n1028;
  wire n1029;
  wire n1030;
  wire n1031;
  wire n1032;
  wire n1033;
  wire n1034;
  wire n1035;
  wire n1036;
  wire n1037;
  wire n1038;
  wire n1039;
  wire n1040;
  wire n1041;
  wire n1042;
  wire n1043;
  wire n1044;
  wire n1045;
  wire n1046;
  wire n1047;
  wire n1048;
  wire n1049;
  wire n1050;
  wire n1051;
  wire n1052;
  wire n1053;
  wire n1054;
  wire n1055;
  wire n1056;
  wire n1057;
  wire n1058;
  wire n1059;
  wire n1060;
  wire n1061;
  wire n1062;
  wire n1063;
  wire n1064;
  wire n1065;
  wire n1066;
  wire n1067;
  wire n1068;
  wire n1069;
  wire n1070;
  wire n1071;
  wire n1072;
  wire n1073;
  wire n1074;
  wire n1075;
  wire n1076;
  wire n1077;
  wire n1078;
  wire n1079;
  wire n1080;
  wire n1081;
  wire n1082;
  wire n1083;
  wire n1084;
  wire n1085;
  wire n1086;
  wire n1087;
  wire n1088;
  wire n1089;
  wire n1090;
  wire n1091;
  wire n1092;
  wire n1093;
  wire n1094;
  wire n1095;
  wire n1096;
  wire n1097;
  wire n1098;
  wire n1099;
  wire n1100;
  wire n1101;
  wire n1102;
  wire n1103;
  wire n1104;
  wire n1105;
  wire n1106;
  wire n1107;
  wire n1108;
  wire n1109;
  wire n1110;
  wire n1111;
  wire n1112;
  wire n1113;
  wire n1114;
  wire n1115;
  wire n1116;
  wire n1117;
  wire n1118;
  wire n1119;
  wire n1120;
  wire n1121;
  wire n1122;
  wire n1123;
  wire n1124;
  wire n1125;
  wire n1126;
  wire n1127;
  wire n1128;
  wire n1129;
  wire n1130;
  wire n1131;
  wire n1132;
  wire n1133;
  wire n1134;
  wire n1135;
  wire n1136;
  wire n1137;
  wire n1138;
  wire n1139;
  wire n1140;
  wire n1141;
  wire n1142;
  wire n1143;
  wire n1144;
  wire n1145;
  wire n1146;
  wire n1147;
  wire n1148;
  wire n1149;
  wire n1150;
  wire n1151;
  wire n1152;
  wire n1153;
  wire n1154;
  wire n1155;
  wire n1156;
  wire n1157;
  wire n1158;
  wire n1159;
  wire n1160;
  wire n1161;
  wire n1162;
  wire n1163;
  wire n1164;
  wire n1165;
  wire n1166;
  wire n1167;
  wire n1168;
  wire n1169;
  wire n1170;
  wire n1171;
  wire n1172;
  wire n1173;
  wire n1174;
  wire n1175;
  wire n1176;
  wire n1177;
  wire n1178;
  wire n1179;
  wire n1180;
  wire n1181;
  wire n1182;
  wire n1183;
  wire n1184;
  wire n1185;
  wire n1186;
  wire n1187;
  wire n1188;
  wire n1189;
  wire n1190;
  wire n1191;
  wire n1192;
  wire n1193;
  wire n1194;
  wire n1195;
  wire n1196;
  wire n1197;
  wire n1198;
  wire n1199;
  wire n1200;
  wire n1201;
  wire n1202;
  wire n1203;
  wire n1204;
  wire n1205;
  wire n1206;
  wire n1207;
  wire n1208;
  wire n1209;
  wire n1210;
  wire n1211;
  wire n1212;
  wire n1213;
  wire n1214;
  wire n1215;
  wire n1216;
  wire n1217;
  wire n1218;
  wire n1219;
  wire n1220;
  wire n1221;
  wire n1222;
  wire n1223;
  wire n1224;
  wire n1225;
  wire n1226;
  wire n1227;
  wire n1228;
  wire n1229;
  wire n1230;
  wire n1231;
  wire n1232;
  wire n1233;
  wire n1234;
  wire n1235;
  wire n1236;
  wire n1237;
  wire n1238;
  wire n1239;
  wire n1240;
  wire n1241;
  wire n1242;
  wire n1243;
  wire n1244;
  wire n1245;
  wire n1246;
  wire n1247;
  wire n1248;
  wire n1249;
  wire n1250;
  wire n1251;
  wire n1252;
  wire n1253;
  wire n1254;
  wire n1255;
  wire n1256;
  wire n1257;
  wire n1258;
  wire n1259;
  wire n1260;
  wire n1261;
  wire n1262;
  wire n1263;
  wire n1264;
  wire n1265;
  wire n1266;
  wire n1267;
  wire n1268;
  wire n1269;
  wire n1270;
  wire n1271;
  wire n1272;
  wire n1273;
  wire n1274;
  wire n1275;
  wire n1276;
  wire n1277;
  wire n1278;
  wire n1279;
  wire n1280;
  wire n1281;
  wire n1282;
  wire n1283;
  wire n1284;
  wire n1285;
  wire n1286;
  wire n1287;
  wire n1288;
  wire n1289;
  wire n1290;
  wire n1291;
  wire n1292;
  wire n1293;
  wire n1294;
  wire n1295;
  wire n1296;
  wire n1297;
  wire n1298;
  wire n1299;
  wire n1300;
  wire n1301;
  wire n1302;
  wire n1303;
  wire n1304;
  wire n1305;
  wire n1306;
  wire n1307;
  wire n1308;
  wire n1309;
  wire n1310;
  wire n1311;
  wire n1312;
  wire n1313;
  wire n1314;
  wire n1315;
  wire n1316;
  wire n1317;
  wire n1318;
  wire n1319;
  wire n1320;
  wire n1321;
  wire n1322;
  wire n1323;
  wire n1324;
  wire n1325;
  wire n1326;
  wire n1327;
  wire n1328;
  wire n1329;
  wire n1330;
  wire n1331;
  wire n1332;
  wire n1333;
  wire n1334;
  wire n1335;
  wire n1336;
  wire n1337;
  wire n1338;
  wire n1339;
  wire n1340;
  wire n1341;
  wire n1342;
  wire n1343;
  wire n1344;
  wire n1345;
  wire n1346;
  wire n1347;
  wire n1348;
  wire n1349;
  wire n1350;
  wire n1351;
  wire n1352;
  wire n1353;
  wire n1354;
  wire n1355;
  wire n1356;
  wire n1357;
  wire n1358;
  wire n1359;
  wire n1360;
  wire n1361;
  wire n1362;
  wire n1363;
  wire n1364;
  wire n1365;
  wire n1366;
  wire n1367;
  wire n1368;
  wire n1369;
  wire n1370;
  wire n1371;
  wire n1372;
  wire n1373;
  wire n1374;
  wire n1375;
  wire n1376;
  wire n1377;
  wire n1378;
  wire n1379;
  wire n1380;
  wire n1381;
  wire n1382;
  wire n1383;
  wire n1384;
  wire n1385;
  wire n1386;
  wire n1387;
  wire n1388;
  wire n1389;
  wire n1390;
  wire n1391;
  wire n1392;
  wire n1393;
  wire n1394;
  wire n1395;
  wire n1396;
  wire n1397;
  wire n1398;
  wire n1399;
  wire n1400;
  wire n1401;
  wire n1402;
  wire n1403;
  wire n1404;
  wire n1405;
  wire n1406;
  wire n1407;
  wire n1408;
  wire n1409;
  wire n1410;
  wire n1411;
  wire n1412;
  wire n1413;
  wire n1414;
  wire n1415;
  wire n1416;
  wire n1417;
  wire n1418;
  wire n1419;
  wire n1420;
  wire n1421;
  wire n1422;
  wire n1423;
  wire n1424;
  wire n1425;
  wire n1426;
  wire n1427;
  wire n1428;
  wire n1429;
  wire n1430;
  wire n1431;
  wire n1432;
  wire n1433;
  wire n1434;
  wire n1435;
  wire n1436;
  wire n1437;
  wire n1438;
  wire n1439;
  wire n1440;
  wire n1441;
  wire n1442;
  wire n1443;
  wire n1444;
  wire n1445;
  wire n1446;
  wire n1447;
  wire n1448;
  wire n1449;
  wire n1450;
  wire n1451;
  wire n1452;
  wire n1453;
  wire n1454;
  wire n1455;
  wire n1456;
  wire n1457;
  wire n1458;
  wire n1459;
  wire n1460;
  wire n1461;
  wire n1462;
  wire n1463;
  wire n1464;
  wire n1465;
  wire n1466;
  wire n1467;
  wire n1468;
  wire n1469;
  wire n1470;
  wire n1471;
  wire n1472;
  wire n1473;
  wire n1474;
  wire n1475;
  wire n1476;
  wire n1477;
  wire n1478;
  wire n1479;
  wire n1480;
  wire n1481;
  wire n1482;
  wire n1483;
  wire n1484;
  wire n1485;
  wire n1486;
  wire n1487;
  wire n1488;
  wire n1489;
  wire n1490;
  wire n1491;
  wire n1492;
  wire n1493;
  wire n1494;
  wire n1495;
  wire n1496;
  wire n1497;
  wire n1498;
  wire n1499;
  wire n1500;
  wire n1501;
  wire n1502;
  wire n1503;
  wire n1504;
  wire n1505;
  wire n1506;
  wire n1507;
  wire n1508;
  wire n1509;
  wire n1510;
  wire n1511;
  wire n1512;
  wire n1513;
  wire n1514;
  wire n1515;
  wire n1516;
  wire n1517;
  wire n1518;
  wire n1519;
  wire n1520;
  wire n1521;
  wire n1522;
  wire n1523;
  wire n1524;
  wire n1525;
  wire n1526;
  wire n1527;
  wire n1528;
  wire n1529;
  wire n1530;
  wire n1531;
  wire n1532;
  wire n1533;
  wire n1534;
  wire n1535;
  wire n1536;
  wire n1537;
  wire n1538;
  wire n1539;
  wire n1540;
  wire n1541;
  wire n1542;
  wire n1543;
  wire n1544;
  wire n1545;
  wire n1546;
  wire n1547;
  wire n1548;
  wire n1549;
  wire n1550;
  wire n1551;
  wire n1552;
  wire n1553;
  wire n1554;
  wire n1555;
  wire n1556;
  wire n1557;
  wire n1558;
  wire n1559;
  wire n1560;
  wire n1561;
  wire n1562;
  wire n1563;
  wire n1564;
  wire n1565;
  wire n1566;
  wire n1567;
  wire n1568;
  wire n1569;
  wire n1570;
  wire n1571;
  wire n1572;
  wire n1573;
  wire n1574;
  wire n1575;
  wire n1576;
  wire n1577;
  wire n1578;
  wire n1579;
  wire n1580;
  wire n1581;
  wire n1582;
  wire n1583;
  wire n1584;
  wire n1585;
  wire n1586;
  wire n1587;
  wire n1588;
  wire n1589;
  wire n1590;
  wire n1591;
  wire n1592;
  wire n1593;
  wire n1594;
  wire n1595;
  wire n1596;
  wire n1597;
  wire n1598;
  wire n1599;
  wire n1600;
  wire n1601;
  wire n1602;
  wire n1603;
  wire n1604;
  wire n1605;
  wire n1606;
  wire n1607;
  wire n1608;
  wire n1609;
  wire n1610;
  wire n1611;
  wire n1612;
  wire n1613;
  wire n1614;
  wire n1615;
  wire n1616;
  wire n1617;
  wire n1618;
  wire n1619;
  wire n1620;
  wire n1621;
  wire n1622;
  wire n1623;
  wire n1624;
  wire n1625;
  wire n1626;
  wire n1627;
  wire n1628;
  wire n1629;
  wire n1630;
  wire n1631;
  wire n1632;
  wire n1633;
  wire n1634;
  wire n1635;
  wire n1636;
  wire n1637;
  wire n1638;
  wire n1639;
  wire n1640;
  wire n1641;
  wire n1642;
  wire n1643;
  wire n1644;
  wire n1645;
  wire n1646;
  wire n1647;
  wire n1648;
  wire n1649;
  wire n1650;
  wire n1651;
  wire n1652;
  wire n1653;
  wire n1654;
  wire n1655;
  wire n1656;
  wire n1657;
  wire n1658;
  wire n1659;
  wire n1660;
  wire n1661;
  wire n1662;
  wire n1663;
  wire n1664;
  wire n1665;
  wire n1666;
  wire n1667;
  wire n1668;
  wire n1669;
  wire n1670;
  wire n1671;
  wire n1672;
  wire n1673;
  wire n1674;
  wire n1675;
  wire n1676;
  wire n1677;
  wire n1678;
  wire n1679;
  wire n1680;
  wire n1681;
  wire n1682;
  wire n1683;
  wire n1684;
  wire n1685;
  wire n1686;
  wire n1687;
  wire n1688;
  wire n1689;
  wire n1690;
  wire n1691;
  wire n1692;
  wire n1693;
  wire n1694;
  wire n1695;
  wire n1696;
  wire n1697;
  wire n1698;
  wire n1699;
  wire n1700;
  wire n1701;
  wire n1702;
  wire n1703;
  wire n1704;
  wire n1705;
  wire n1706;
  wire n1707;
  wire n1708;
  wire n1709;
  wire n1710;
  wire n1711;
  wire n1712;
  wire n1713;
  wire n1714;
  wire n1715;
  wire n1716;
  wire n1717;
  wire n1718;
  wire n1719;
  wire n1720;
  wire n1721;
  wire n1722;
  wire n1723;
  wire n1724;
  wire n1725;
  wire n1726;
  wire n1727;
  wire n1728;
  wire n1729;
  wire n1730;
  wire n1731;
  wire n1732;
  wire n1733;
  wire n1734;
  wire n1735;
  wire n1736;
  wire n1737;
  wire n1738;
  wire n1739;
  wire n1740;
  wire n1741;
  wire n1742;
  wire n1743;
  wire n1744;
  wire n1745;
  wire n1746;
  wire n1747;
  wire n1748;
  wire n1749;
  wire n1750;
  wire n1751;
  wire n1752;
  wire n1753;
  wire n1754;
  wire n1755;
  wire n1756;
  wire n1757;
  wire n1758;
  wire n1759;
  wire n1760;
  wire n1761;
  wire n1762;
  wire n1763;
  wire n1764;
  wire n1765;
  wire n1766;
  wire n1767;
  wire n1768;
  wire n1769;
  wire n1770;
  wire n1771;
  wire n1772;
  wire n1773;
  wire n1774;
  wire n1775;
  wire n1776;
  wire n1777;
  wire n1778;
  wire n1779;
  wire n1780;
  wire n1781;
  wire n1782;
  wire n1783;
  wire n1784;
  wire n1785;
  wire n1786;
  wire n1787;
  wire n1788;
  wire n1789;
  wire n1790;
  wire n1791;
  wire n1792;
  wire n1793;
  wire n1794;
  wire n1795;
  wire n1796;
  wire n1797;
  wire n1798;
  wire n1799;
  wire n1800;
  wire n1801;
  wire n1802;
  wire n1803;
  wire n1804;
  wire n1805;
  wire n1806;
  wire n1807;
  wire n1808;
  wire n1809;
  wire n1810;
  wire n1811;
  wire n1812;
  wire n1813;
  wire n1814;
  wire n1815;
  wire n1816;
  wire n1817;
  wire n1818;
  wire n1819;
  wire n1820;
  wire n1821;
  wire n1822;
  wire n1823;
  wire n1824;
  wire n1825;
  wire n1826;
  wire n1827;
  wire n1828;
  wire n1829;
  wire n1830;
  wire n1831;
  wire n1832;
  wire n1833;
  wire n1834;
  wire n1835;
  wire n1836;
  wire n1837;
  wire n1838;
  wire n1839;
  wire n1840;
  wire n1841;
  wire n1842;
  wire n1843;
  wire n1844;
  wire n1845;
  wire n1846;
  wire n1847;
  wire n1848;
  wire n1849;
  wire n1850;
  wire n1851;
  wire n1852;
  wire n1853;
  wire n1854;
  wire n1855;
  wire n1856;
  wire n1857;
  wire n1858;
  wire n1859;
  wire n1860;
  wire n1861;
  wire n1862;
  wire n1863;
  wire n1864;
  wire n1865;
  wire n1866;
  wire n1867;
  wire n1868;
  wire n1869;
  wire n1870;
  wire n1871;
  wire n1872;
  wire n1873;
  wire n1874;
  wire n1875;
  wire n1876;
  wire n1877;
  wire n1878;
  wire n1879;
  wire n1880;
  wire n1881;
  wire n1882;
  wire n1883;
  wire n1884;
  wire n1885;
  wire n1886;
  wire n1887;
  wire n1888;
  wire n1889;
  wire n1890;
  wire n1891;
  wire n1892;
  wire n1893;
  wire n1894;
  wire n1895;
  wire n1896;
  wire n1897;
  wire n1898;
  wire n1899;
  wire n1900;
  wire n1901;
  wire n1902;
  wire n1903;
  wire n1904;
  wire n1905;
  wire n1906;
  wire n1907;
  wire n1908;
  wire n1909;
  wire n1910;
  wire n1911;
  wire n1912;
  wire n1913;
  wire n1914;
  wire n1915;
  wire n1916;
  wire n1917;
  wire n1918;
  wire n1919;
  wire n1920;
  wire n1921;
  wire n1922;
  wire n1923;
  wire n1924;
  wire n1925;
  wire n1926;
  wire n1927;
  wire n1928;
  wire n1929;
  wire n1930;
  wire n1931;
  wire n1932;
  wire n1933;
  wire n1934;
  wire n1935;
  wire n1936;
  wire n1937;
  wire n1938;
  wire n1939;
  wire n1940;
  wire n1941;
  wire n1942;
  wire n1943;
  wire n1944;
  wire n1945;
  wire n1946;
  wire n1947;
  wire n1948;
  wire n1949;
  wire n1950;
  wire n1951;
  wire n1952;
  wire n1953;
  wire n1954;
  wire n1955;
  wire n1956;
  wire n1957;
  wire n1958;
  wire n1959;
  wire n1960;
  wire n1961;
  wire n1962;
  wire n1963;
  wire n1964;
  wire n1965;
  wire n1966;
  wire n1967;
  wire n1968;
  wire n1969;
  wire n1970;
  wire n1971;
  wire n1972;
  wire n1973;
  wire n1974;
  wire n1975;
  wire n1976;
  wire n1977;
  wire n1978;
  wire n1979;
  wire n1980;
  wire n1981;
  wire n1982;
  wire n1983;
  wire n1984;
  wire n1985;
  wire n1986;
  wire n1987;
  wire n1988;
  wire n1989;
  wire n1990;
  wire n1991;
  wire n1992;
  wire n1993;
  wire n1994;
  wire n1995;
  wire n1996;
  wire n1997;
  wire n1998;
  wire n1999;
  wire n2000;
  wire n2001;
  wire n2002;
  wire n2003;
  wire n2004;
  wire n2005;
  wire n2006;
  wire n2007;
  wire n2008;
  wire n2009;
  wire n2010;
  wire n2011;
  wire n2012;
  wire n2013;
  wire n2014;
  wire n2015;
  wire n2016;
  wire n2017;
  wire n2018;
  wire n2019;
  wire n2020;
  wire n2021;
  wire n2022;
  wire n2023;
  wire n2024;
  wire n2025;
  wire n2026;
  wire n2027;
  wire n2028;
  wire n2029;
  wire n2030;
  wire n2031;
  wire n2032;
  wire n2033;
  wire n2034;
  wire n2035;
  wire n2036;
  wire n2037;
  wire n2038;
  wire n2039;
  wire n2040;
  wire n2041;
  wire n2042;
  wire n2043;
  wire n2044;
  wire n2045;
  wire n2046;
  wire n2047;
  wire n2048;
  wire n2049;
  wire n2050;
  wire n2051;
  wire n2052;
  wire n2053;
  wire n2054;
  wire n2055;
  wire n2056;
  wire n2057;
  wire n2058;
  wire n2059;
  wire n2060;
  wire n2061;
  wire n2062;
  wire n2063;
  wire n2064;
  wire n2065;
  wire n2066;
  wire n2067;
  wire n2068;
  wire n2069;
  wire n2070;
  wire n2071;
  wire n2072;
  wire n2073;
  wire n2074;
  wire n2075;
  wire n2076;
  wire n2077;
  wire n2078;
  wire n2079;
  wire n2080;
  wire n2081;
  wire n2082;
  wire n2083;
  wire n2084;
  wire n2085;
  wire n2086;
  wire n2087;
  wire n2088;
  wire n2089;
  wire n2090;
  wire n2091;
  wire n2092;
  wire n2093;
  wire n2094;
  wire n2095;
  wire n2096;
  wire n2097;
  wire n2098;
  wire n2099;
  wire n2100;
  wire n2101;
  wire n2102;
  wire n2103;
  wire n2104;
  wire n2105;
  wire n2106;
  wire n2107;
  wire n2108;
  wire n2109;
  wire n2110;
  wire n2111;
  wire n2112;
  wire n2113;
  wire n2114;
  wire n2115;
  wire n2116;
  wire n2117;
  wire n2118;
  wire n2119;
  wire n2120;
  wire n2121;
  wire n2122;
  wire n2123;
  wire n2124;
  wire n2125;
  wire n2126;
  wire n2127;
  wire n2128;
  wire n2129;
  wire n2130;
  wire n2131;
  wire n2132;
  wire n2133;
  wire n2134;
  wire n2135;
  wire n2136;
  wire n2137;
  wire n2138;
  wire n2139;
  wire n2140;
  wire n2141;
  wire n2142;
  wire n2143;
  wire n2144;
  wire n2145;
  wire n2146;
  wire n2147;
  wire n2148;
  wire n2149;
  wire n2150;
  wire n2151;
  wire n2152;
  wire n2153;
  wire n2154;
  wire n2155;
  wire n2156;
  wire n2157;
  wire n2158;
  wire n2159;
  wire n2160;
  wire n2161;
  wire n2162;
  wire n2163;
  wire n2164;
  wire n2165;
  wire n2166;
  wire n2167;
  wire n2168;
  wire n2169;
  wire n2170;
  wire n2171;
  wire n2172;
  wire n2173;
  wire n2174;
  wire n2175;
  wire n2176;
  wire n2177;
  wire n2178;
  wire n2179;
  wire n2180;
  wire n2181;
  wire n2182;
  wire n2183;
  wire n2184;
  wire n2185;
  wire n2186;
  wire n2187;
  wire n2188;
  wire n2189;
  wire n2190;
  wire n2191;
  wire n2192;
  wire n2193;
  wire n2194;
  wire n2195;
  wire n2196;
  wire n2197;
  wire n2198;
  wire n2199;
  wire n2200;
  wire n2201;
  wire n2202;
  wire n2203;
  wire n2204;
  wire n2205;
  wire n2206;
  wire n2207;
  wire n2208;
  wire n2209;
  wire n2210;
  wire n2211;
  wire n2212;
  wire n2213;
  wire n2214;
  wire n2215;
  wire n2216;
  wire n2217;
  wire n2218;
  wire n2219;
  wire n2220;
  wire n2221;
  wire n2222;
  wire n2223;
  wire n2224;
  wire n2225;
  wire n2226;
  wire n2227;
  wire n2228;
  wire n2229;
  wire n2230;
  wire n2231;
  wire n2232;
  wire n2233;
  wire n2234;
  wire n2235;
  wire n2236;
  wire n2237;
  wire n2238;
  wire n2239;
  wire n2240;
  wire n2241;
  wire n2242;
  wire n2243;
  wire n2244;
  wire n2245;
  wire n2246;
  wire n2247;
  wire n2248;
  wire n2249;
  wire n2250;
  wire n2251;
  wire n2252;
  wire n2253;
  wire n2254;
  wire n2255;
  wire n2256;
  wire n2257;
  wire n2258;
  wire n2259;
  wire n2260;
  wire n2261;
  wire n2262;
  wire n2263;
  wire n2264;
  wire n2265;
  wire n2266;
  wire n2267;
  wire n2268;
  wire n2269;
  wire n2270;
  wire n2271;
  wire n2272;
  wire n2273;
  wire n2274;
  wire n2275;
  wire n2276;
  wire n2277;
  wire n2278;
  wire n2279;
  wire n2280;
  wire n2281;
  wire n2282;
  wire n2283;
  wire n2284;
  wire n2285;
  wire n2286;
  wire n2287;
  wire n2288;
  wire n2289;
  wire n2290;
  wire n2291;
  wire n2292;
  wire n2293;
  wire n2294;
  wire n2295;
  wire n2296;
  wire n2297;
  wire n2298;
  wire n2299;
  wire n2300;
  wire n2301;
  wire n2302;
  wire n2303;
  wire n2304;
  wire n2305;
  wire n2306;
  wire n2307;
  wire n2308;
  wire n2309;
  wire n2310;
  wire n2311;
  wire n2312;
  wire n2313;
  wire n2314;
  wire n2315;
  wire n2316;
  wire n2317;
  wire n2318;
  wire n2319;
  wire n2320;
  wire n2321;
  wire n2322;
  wire n2323;
  wire n2324;
  wire n2325;
  wire n2326;
  wire n2327;
  wire n2328;
  wire n2329;
  wire n2330;
  wire n2331;
  wire n2332;
  wire n2333;
  wire n2334;
  wire n2335;
  wire n2336;
  wire n2337;
  wire n2338;
  wire n2339;
  wire n2340;
  wire n2341;
  wire n2342;
  wire n2343;
  wire n2344;
  wire n2345;
  wire n2346;
  wire n2347;
  wire n2348;
  wire n2349;
  wire n2350;
  wire n2351;
  wire n2352;
  wire n2353;
  wire n2354;
  wire n2355;
  wire n2356;
  wire n2357;
  wire n2358;
  wire n2359;
  wire n2360;
  wire n2361;
  wire n2362;
  wire n2363;
  wire n2364;
  wire n2365;
  wire n2366;
  wire n2367;
  wire n2368;
  wire n2369;
  wire n2370;
  wire n2371;
  wire n2372;
  wire n2373;
  wire n2374;
  wire n2375;
  wire n2376;
  wire n2377;
  wire n2378;
  wire n2379;
  wire n2380;
  wire n2381;
  wire n2382;
  wire n2383;
  wire n2384;
  wire n2385;
  wire n2386;
  wire n2387;
  wire n2388;
  wire n2389;
  wire n2390;
  wire n2391;
  wire n2392;
  wire n2393;
  wire n2394;
  wire n2395;
  wire n2396;
  wire n2397;
  wire n2398;
  wire n2399;
  wire n2400;
  wire n2401;
  wire n2402;
  wire n2403;
  wire n2404;
  wire n2405;
  wire n2406;
  wire n2407;
  wire n2408;
  wire n2409;
  wire n2410;
  wire n2411;
  wire n2412;
  wire n2413;
  wire n2414;
  wire n2415;
  wire n2416;
  wire n2417;
  wire n2418;
  wire n2419;
  wire n2420;
  wire n2421;
  wire n2422;
  wire n2423;
  wire n2424;
  wire n2425;
  wire n2426;
  wire n2427;
  wire n2428;
  wire n2429;
  wire n2430;
  wire n2431;
  wire n2432;
  wire n2433;
  wire n2434;
  wire n2435;
  wire n2436;
  wire n2437;
  wire n2438;
  wire n2439;
  wire n2440;
  wire n2441;
  wire n2442;
  wire n2443;
  wire n2444;
  wire n2445;
  wire n2446;
  wire n2447;
  wire n2448;
  wire n2449;
  wire n2450;
  wire n2451;
  wire n2452;
  wire n2454;
  wire n2455;
  wire n2456;
  wire n2457;
  wire n2458;
  wire n2459;
  wire n2460;
  wire n2461;
  wire n2462;
  wire n2463;
  wire n2464;
  wire n2465;
  wire n2466;
  wire n2467;
  wire n2468;
  wire n2469;
  wire n2470;
  wire n2471;
  wire n2472;
  wire n2473;
  wire n2474;
  wire n2475;
  wire n2476;
  wire n2477;
  wire n2478;
  wire n2479;
  wire n2480;
  wire n2481;
  wire n2483;
  wire n2484;
  wire n2485;
  wire n2486;
  wire n2487;
  wire n2488;
  wire n2489;
  wire n2490;
  wire n2491;
  wire n2492;
  wire n2493;
  wire n2494;
  wire n2495;
  wire n2496;
  wire n2497;
  wire n2498;
  wire n2499;
  wire n2500;
  wire n2501;
  wire n2502;
  wire n2503;
  wire n2504;
  wire n2505;
  wire n2506;
  wire n2507;
  wire n2508;
  wire n2509;
  wire n2510;
  wire n2511;
  wire n2512;
  wire n2513;
  wire n2514;
  wire n2515;
  wire n2516;
  wire n2517;
  wire n2518;
  wire n2519;
  wire n2520;
  wire n2522;
  wire n2527;
  wire n2528;
  wire n2529;
  wire n2530;
  wire n2531;
  wire n2532;
  wire n2533;
  wire n2534;
  wire n2535;
  wire n2536;
  wire n2537;
  wire n2538;
  wire n2539;
  wire n2540;
  wire n2541;
  wire n2542;
  wire n2543;
  wire n2544;
  wire n2545;
  wire n2546;
  wire n2547;
  wire n2548;
  wire n2549;
  wire n2550;
  wire n2551;
  wire n2552;
  wire KeyWire_0_0;
  wire KeyWire_0_1;
  wire KeyWire_0_2;
  wire KeyNOTWire_0_2;
  wire KeyWire_0_3;
  wire KeyNOTWire_0_3;
  wire KeyWire_0_4;
  wire KeyWire_0_5;
  wire KeyNOTWire_0_5;
  wire KeyWire_0_6;
  wire KeyWire_0_7;
  wire KeyWire_0_8;
  wire KeyNOTWire_0_8;
  wire KeyWire_0_9;
  wire KeyWire_0_10;
  wire KeyNOTWire_0_10;
  wire KeyWire_0_11;
  wire KeyNOTWire_0_11;
  wire KeyWire_0_12;
  wire KeyNOTWire_0_12;
  wire KeyWire_0_13;
  wire KeyWire_0_14;
  wire KeyNOTWire_0_14;
  wire KeyWire_0_15;
  wire KeyWire_0_16;
  wire KeyWire_0_17;
  wire KeyWire_0_18;
  wire KeyNOTWire_0_18;
  wire KeyWire_0_19;
  wire KeyWire_0_20;
  wire KeyWire_0_21;
  wire KeyNOTWire_0_21;
  wire KeyWire_0_22;
  wire KeyWire_0_23;
  wire KeyNOTWire_0_23;
  wire KeyWire_0_24;
  wire KeyWire_0_25;
  wire KeyNOTWire_0_25;
  wire KeyWire_0_26;
  wire KeyNOTWire_0_26;
  wire KeyWire_0_27;
  wire KeyNOTWire_0_27;
  wire KeyWire_0_28;
  wire KeyWire_0_29;
  wire KeyNOTWire_0_29;
  wire KeyWire_0_30;
  wire KeyNOTWire_0_30;
  wire KeyWire_0_31;
  wire KeyNOTWire_0_31;
  wire KeyWire_0_32;
  wire KeyWire_0_33;
  wire KeyNOTWire_0_33;
  wire KeyWire_0_34;
  wire KeyWire_0_35;
  wire KeyWire_0_36;
  wire KeyWire_0_37;
  wire KeyWire_0_38;
  wire KeyNOTWire_0_38;
  wire KeyWire_0_39;
  wire KeyWire_0_40;
  wire KeyWire_0_41;
  wire KeyWire_0_42;
  wire KeyNOTWire_0_42;
  wire KeyWire_0_43;
  wire KeyWire_0_44;
  wire KeyNOTWire_0_44;
  wire KeyWire_0_45;
  wire KeyWire_0_46;
  wire KeyNOTWire_0_46;
  wire KeyWire_0_47;
  wire KeyNOTWire_0_47;
  wire KeyWire_0_48;
  wire KeyNOTWire_0_48;
  wire KeyWire_0_49;
  wire KeyWire_0_50;
  wire KeyNOTWire_0_50;
  wire KeyWire_0_51;
  wire KeyWire_0_52;
  wire KeyNOTWire_0_52;
  wire KeyWire_0_53;
  wire KeyNOTWire_0_53;
  wire KeyWire_0_54;
  wire KeyWire_0_55;
  wire KeyWire_0_56;
  wire KeyNOTWire_0_56;
  wire KeyWire_0_57;
  wire KeyWire_0_58;
  wire KeyNOTWire_0_58;
  wire KeyWire_0_59;
  wire KeyNOTWire_0_59;
  wire KeyWire_0_60;
  wire KeyNOTWire_0_60;
  wire KeyWire_0_61;
  wire KeyNOTWire_0_61;
  wire KeyWire_0_62;
  wire KeyWire_0_63;

  buf
  g0
  (
    n206,
    n33
  );


  not
  g1
  (
    n174,
    n33
  );


  buf
  g2
  (
    n53,
    n4
  );


  not
  g3
  (
    n186,
    n24
  );


  not
  g4
  (
    n175,
    n19
  );


  not
  g5
  (
    n69,
    n39
  );


  not
  g6
  (
    n161,
    n15
  );


  buf
  g7
  (
    n201,
    n39
  );


  buf
  g8
  (
    n97,
    n15
  );


  not
  g9
  (
    n103,
    n23
  );


  buf
  g10
  (
    n105,
    n35
  );


  not
  g11
  (
    n200,
    n26
  );


  not
  g12
  (
    n57,
    n29
  );


  buf
  g13
  (
    n124,
    n3
  );


  buf
  g14
  (
    n156,
    n34
  );


  not
  g15
  (
    n169,
    n6
  );


  not
  g16
  (
    n157,
    n4
  );


  buf
  g17
  (
    n94,
    n35
  );


  not
  g18
  (
    n195,
    n42
  );


  not
  g19
  (
    n77,
    n12
  );


  not
  g20
  (
    n134,
    n36
  );


  buf
  g21
  (
    n179,
    n12
  );


  not
  g22
  (
    n80,
    n22
  );


  buf
  g23
  (
    n145,
    n7
  );


  not
  g24
  (
    n135,
    n44
  );


  not
  g25
  (
    n99,
    n23
  );


  buf
  g26
  (
    n146,
    n31
  );


  not
  g27
  (
    n55,
    n8
  );


  not
  g28
  (
    n81,
    n14
  );


  not
  g29
  (
    KeyWire_0_37,
    n10
  );


  buf
  g30
  (
    n108,
    n23
  );


  buf
  g31
  (
    n216,
    n5
  );


  not
  g32
  (
    n117,
    n35
  );


  buf
  g33
  (
    n164,
    n18
  );


  buf
  g34
  (
    n180,
    n19
  );


  not
  g35
  (
    n190,
    n11
  );


  not
  g36
  (
    n49,
    n41
  );


  not
  g37
  (
    KeyWire_0_34,
    n20
  );


  not
  g38
  (
    n155,
    n25
  );


  buf
  g39
  (
    n126,
    n11
  );


  buf
  g40
  (
    n88,
    n39
  );


  buf
  g41
  (
    n170,
    n27
  );


  buf
  g42
  (
    n107,
    n14
  );


  buf
  g43
  (
    n65,
    n2
  );


  buf
  g44
  (
    n106,
    n10
  );


  not
  g45
  (
    n158,
    n17
  );


  not
  g46
  (
    n139,
    n43
  );


  not
  g47
  (
    n220,
    n8
  );


  buf
  g48
  (
    n79,
    n9
  );


  buf
  g49
  (
    n178,
    n36
  );


  not
  g50
  (
    n185,
    n38
  );


  buf
  g51
  (
    n149,
    n38
  );


  not
  g52
  (
    n148,
    n8
  );


  not
  g53
  (
    n151,
    n20
  );


  not
  g54
  (
    n188,
    n31
  );


  buf
  g55
  (
    n165,
    n17
  );


  buf
  g56
  (
    n93,
    n41
  );


  not
  g57
  (
    n120,
    n40
  );


  buf
  g58
  (
    n127,
    n22
  );


  buf
  g59
  (
    n109,
    n10
  );


  not
  g60
  (
    n172,
    n33
  );


  buf
  g61
  (
    n160,
    n26
  );


  buf
  g62
  (
    n152,
    n40
  );


  not
  g63
  (
    n154,
    n13
  );


  not
  g64
  (
    n136,
    n6
  );


  buf
  g65
  (
    n193,
    n19
  );


  buf
  g66
  (
    n219,
    n17
  );


  buf
  g67
  (
    n52,
    n11
  );


  buf
  g68
  (
    n202,
    n9
  );


  buf
  g69
  (
    n75,
    n16
  );


  not
  g70
  (
    n101,
    n21
  );


  not
  g71
  (
    n47,
    n34
  );


  buf
  g72
  (
    n64,
    n8
  );


  buf
  g73
  (
    n67,
    n14
  );


  buf
  g74
  (
    n138,
    n43
  );


  buf
  g75
  (
    n153,
    n25
  );


  not
  g76
  (
    n45,
    n10
  );


  not
  g77
  (
    n144,
    n44
  );


  buf
  g78
  (
    n111,
    n19
  );


  buf
  g79
  (
    n210,
    n18
  );


  buf
  g80
  (
    n192,
    n15
  );


  buf
  g81
  (
    n209,
    n7
  );


  buf
  g82
  (
    n159,
    n32
  );


  buf
  g83
  (
    n184,
    n38
  );


  buf
  g84
  (
    n114,
    n6
  );


  not
  g85
  (
    n133,
    n24
  );


  not
  g86
  (
    n68,
    n21
  );


  buf
  g87
  (
    n205,
    n25
  );


  not
  g88
  (
    n62,
    n13
  );


  buf
  g89
  (
    n95,
    n44
  );


  buf
  g90
  (
    n168,
    n24
  );


  not
  g91
  (
    n96,
    n35
  );


  buf
  g92
  (
    n87,
    n1
  );


  buf
  g93
  (
    n183,
    n18
  );


  buf
  g94
  (
    n167,
    n29
  );


  buf
  g95
  (
    n121,
    n41
  );


  buf
  g96
  (
    n171,
    n4
  );


  buf
  g97
  (
    n91,
    n5
  );


  not
  g98
  (
    n177,
    n16
  );


  not
  g99
  (
    n66,
    n44
  );


  buf
  g100
  (
    n83,
    n21
  );


  buf
  g101
  (
    KeyWire_0_39,
    n2
  );


  not
  g102
  (
    n60,
    n28
  );


  buf
  g103
  (
    n58,
    n41
  );


  buf
  g104
  (
    n74,
    n30
  );


  buf
  g105
  (
    n50,
    n37
  );


  buf
  g106
  (
    n173,
    n26
  );


  not
  g107
  (
    n214,
    n39
  );


  buf
  g108
  (
    n213,
    n40
  );


  buf
  g109
  (
    n181,
    n42
  );


  not
  g110
  (
    n56,
    n36
  );


  not
  g111
  (
    n76,
    n11
  );


  buf
  g112
  (
    n182,
    n13
  );


  not
  g113
  (
    n116,
    n22
  );


  buf
  g114
  (
    n54,
    n9
  );


  buf
  g115
  (
    n208,
    n1
  );


  not
  g116
  (
    n51,
    n23
  );


  not
  g117
  (
    n166,
    n3
  );


  buf
  g118
  (
    n85,
    n42
  );


  buf
  g119
  (
    n217,
    n40
  );


  buf
  g120
  (
    n199,
    n43
  );


  not
  g121
  (
    n46,
    n15
  );


  not
  g122
  (
    n113,
    n20
  );


  buf
  g123
  (
    n78,
    n43
  );


  not
  g124
  (
    n176,
    n1
  );


  buf
  g125
  (
    n131,
    n2
  );


  not
  g126
  (
    n84,
    n3
  );


  not
  g127
  (
    n82,
    n30
  );


  buf
  g128
  (
    n72,
    n27
  );


  not
  g129
  (
    n204,
    n34
  );


  buf
  g130
  (
    n104,
    n37
  );


  not
  g131
  (
    KeyWire_0_8,
    n7
  );


  buf
  g132
  (
    n129,
    n32
  );


  not
  g133
  (
    n141,
    n4
  );


  not
  g134
  (
    n102,
    n29
  );


  not
  g135
  (
    n147,
    n12
  );


  buf
  g136
  (
    n163,
    n30
  );


  buf
  g137
  (
    n196,
    n36
  );


  not
  g138
  (
    n90,
    n38
  );


  not
  g139
  (
    n197,
    n21
  );


  not
  g140
  (
    n137,
    n20
  );


  not
  g141
  (
    n118,
    n16
  );


  buf
  g142
  (
    n140,
    n28
  );


  buf
  g143
  (
    n86,
    n18
  );


  not
  g144
  (
    n73,
    n9
  );


  buf
  g145
  (
    n189,
    n7
  );


  buf
  g146
  (
    n122,
    n26
  );


  not
  g147
  (
    n119,
    n3
  );


  buf
  g148
  (
    n130,
    n28
  );


  buf
  g149
  (
    n71,
    n16
  );


  buf
  g150
  (
    n194,
    n17
  );


  buf
  g151
  (
    n100,
    n32
  );


  not
  g152
  (
    n48,
    n27
  );


  buf
  g153
  (
    n92,
    n24
  );


  not
  g154
  (
    n211,
    n33
  );


  not
  g155
  (
    n150,
    n34
  );


  buf
  g156
  (
    n198,
    n14
  );


  not
  g157
  (
    KeyWire_0_26,
    n37
  );


  buf
  g158
  (
    n212,
    n31
  );


  not
  g159
  (
    n203,
    n32
  );


  buf
  g160
  (
    n162,
    n37
  );


  buf
  g161
  (
    n89,
    n27
  );


  not
  g162
  (
    n123,
    n6
  );


  buf
  g163
  (
    n215,
    n25
  );


  not
  g164
  (
    n218,
    n13
  );


  buf
  g165
  (
    n112,
    n12
  );


  not
  g166
  (
    n132,
    n5
  );


  buf
  g167
  (
    n125,
    n28
  );


  not
  g168
  (
    n98,
    n2
  );


  not
  g169
  (
    n115,
    n42
  );


  buf
  g170
  (
    n110,
    n31
  );


  not
  g171
  (
    n142,
    n29
  );


  not
  g172
  (
    n191,
    n30
  );


  buf
  g173
  (
    n187,
    n5
  );


  not
  g174
  (
    n61,
    n22
  );


  not
  g175
  (
    n143,
    n1
  );


  not
  g176
  (
    n779,
    n125
  );


  not
  g177
  (
    n431,
    n102
  );


  buf
  g178
  (
    n577,
    n133
  );


  buf
  g179
  (
    n556,
    n194
  );


  not
  g180
  (
    n870,
    n101
  );


  not
  g181
  (
    n254,
    n59
  );


  not
  g182
  (
    n402,
    n176
  );


  buf
  g183
  (
    n253,
    n178
  );


  not
  g184
  (
    n524,
    n157
  );


  buf
  g185
  (
    n643,
    n70
  );


  buf
  g186
  (
    n889,
    n209
  );


  not
  g187
  (
    n351,
    n86
  );


  not
  g188
  (
    KeyWire_0_10,
    n179
  );


  not
  g189
  (
    n442,
    n158
  );


  not
  g190
  (
    n589,
    n48
  );


  not
  g191
  (
    n644,
    n152
  );


  buf
  g192
  (
    n356,
    n170
  );


  not
  g193
  (
    n774,
    n171
  );


  buf
  g194
  (
    n624,
    n71
  );


  buf
  g195
  (
    n848,
    n54
  );


  not
  g196
  (
    n382,
    n182
  );


  buf
  g197
  (
    n464,
    n100
  );


  not
  g198
  (
    n626,
    n56
  );


  buf
  g199
  (
    n830,
    n126
  );


  buf
  g200
  (
    n560,
    n140
  );


  not
  g201
  (
    n623,
    n167
  );


  buf
  g202
  (
    n318,
    n200
  );


  buf
  g203
  (
    n581,
    n76
  );


  not
  g204
  (
    n437,
    n60
  );


  not
  g205
  (
    n653,
    n98
  );


  buf
  g206
  (
    n518,
    n77
  );


  buf
  g207
  (
    n855,
    n86
  );


  not
  g208
  (
    n270,
    n146
  );


  not
  g209
  (
    n882,
    n52
  );


  not
  g210
  (
    n311,
    n81
  );


  buf
  g211
  (
    n479,
    n220
  );


  buf
  g212
  (
    n233,
    n53
  );


  buf
  g213
  (
    n664,
    n89
  );


  buf
  g214
  (
    n591,
    n143
  );


  not
  g215
  (
    n923,
    n85
  );


  buf
  g216
  (
    n618,
    n170
  );


  buf
  g217
  (
    n521,
    n197
  );


  buf
  g218
  (
    n338,
    n70
  );


  buf
  g219
  (
    n661,
    n101
  );


  not
  g220
  (
    n527,
    n205
  );


  not
  g221
  (
    n459,
    n168
  );


  buf
  g222
  (
    n497,
    n99
  );


  buf
  g223
  (
    n597,
    n94
  );


  not
  g224
  (
    n908,
    n85
  );


  not
  g225
  (
    n328,
    n73
  );


  not
  g226
  (
    n612,
    n63
  );


  buf
  g227
  (
    n826,
    n161
  );


  not
  g228
  (
    n852,
    n218
  );


  buf
  g229
  (
    n388,
    n164
  );


  buf
  g230
  (
    n666,
    n45
  );


  buf
  g231
  (
    n236,
    n219
  );


  not
  g232
  (
    n372,
    n183
  );


  buf
  g233
  (
    n821,
    n104
  );


  not
  g234
  (
    n566,
    n214
  );


  not
  g235
  (
    n361,
    n198
  );


  not
  g236
  (
    n456,
    n83
  );


  not
  g237
  (
    n244,
    n83
  );


  not
  g238
  (
    n801,
    n140
  );


  not
  g239
  (
    n829,
    n174
  );


  not
  g240
  (
    n895,
    n47
  );


  not
  g241
  (
    n691,
    n46
  );


  buf
  g242
  (
    n627,
    n51
  );


  buf
  g243
  (
    n711,
    n88
  );


  buf
  g244
  (
    n505,
    n158
  );


  not
  g245
  (
    n540,
    n96
  );


  buf
  g246
  (
    n645,
    n175
  );


  buf
  g247
  (
    n400,
    n79
  );


  buf
  g248
  (
    n884,
    n104
  );


  buf
  g249
  (
    n632,
    n53
  );


  buf
  g250
  (
    n559,
    n169
  );


  not
  g251
  (
    n552,
    n194
  );


  buf
  g252
  (
    n547,
    n81
  );


  buf
  g253
  (
    n381,
    n86
  );


  not
  g254
  (
    n704,
    n217
  );


  buf
  g255
  (
    n648,
    n57
  );


  not
  g256
  (
    n256,
    n204
  );


  buf
  g257
  (
    KeyWire_0_2,
    n219
  );


  buf
  g258
  (
    n385,
    n60
  );


  not
  g259
  (
    n708,
    n193
  );


  buf
  g260
  (
    n777,
    n197
  );


  buf
  g261
  (
    n323,
    n72
  );


  not
  g262
  (
    n823,
    n164
  );


  not
  g263
  (
    n384,
    n191
  );


  buf
  g264
  (
    n430,
    n82
  );


  buf
  g265
  (
    n657,
    n67
  );


  buf
  g266
  (
    n476,
    n142
  );


  buf
  g267
  (
    n449,
    n106
  );


  buf
  g268
  (
    n322,
    n93
  );


  buf
  g269
  (
    n425,
    n50
  );


  buf
  g270
  (
    n592,
    n184
  );


  buf
  g271
  (
    n865,
    n177
  );


  not
  g272
  (
    n825,
    n182
  );


  not
  g273
  (
    n668,
    n71
  );


  buf
  g274
  (
    n802,
    n210
  );


  not
  g275
  (
    n791,
    n216
  );


  buf
  g276
  (
    n881,
    n80
  );


  not
  g277
  (
    n788,
    n132
  );


  not
  g278
  (
    n488,
    n118
  );


  buf
  g279
  (
    n490,
    n127
  );


  not
  g280
  (
    n421,
    n84
  );


  not
  g281
  (
    n371,
    n161
  );


  not
  g282
  (
    n506,
    n103
  );


  not
  g283
  (
    n586,
    n220
  );


  buf
  g284
  (
    n780,
    n187
  );


  not
  g285
  (
    n611,
    n81
  );


  buf
  g286
  (
    n641,
    n149
  );


  buf
  g287
  (
    n733,
    n92
  );


  buf
  g288
  (
    n416,
    n94
  );


  buf
  g289
  (
    n266,
    n207
  );


  not
  g290
  (
    n501,
    n84
  );


  not
  g291
  (
    n575,
    n48
  );


  buf
  g292
  (
    n580,
    n186
  );


  not
  g293
  (
    n241,
    n55
  );


  buf
  g294
  (
    n740,
    n73
  );


  not
  g295
  (
    n271,
    n163
  );


  buf
  g296
  (
    n637,
    n123
  );


  buf
  g297
  (
    n665,
    n155
  );


  buf
  g298
  (
    n463,
    n216
  );


  not
  g299
  (
    n550,
    n149
  );


  not
  g300
  (
    n346,
    n55
  );


  not
  g301
  (
    n427,
    n201
  );


  not
  g302
  (
    n681,
    n106
  );


  buf
  g303
  (
    n498,
    n85
  );


  not
  g304
  (
    n485,
    n109
  );


  buf
  g305
  (
    n594,
    n180
  );


  buf
  g306
  (
    n838,
    n133
  );


  buf
  g307
  (
    n538,
    n200
  );


  buf
  g308
  (
    n806,
    n63
  );


  buf
  g309
  (
    n844,
    n187
  );


  buf
  g310
  (
    n869,
    n165
  );


  not
  g311
  (
    n370,
    n66
  );


  not
  g312
  (
    n342,
    n103
  );


  buf
  g313
  (
    n707,
    n47
  );


  not
  g314
  (
    n755,
    n87
  );


  not
  g315
  (
    n878,
    n63
  );


  buf
  g316
  (
    n794,
    n151
  );


  not
  g317
  (
    n900,
    n185
  );


  buf
  g318
  (
    n348,
    n54
  );


  buf
  g319
  (
    n268,
    n167
  );


  buf
  g320
  (
    n763,
    n208
  );


  buf
  g321
  (
    n819,
    n200
  );


  buf
  g322
  (
    n365,
    n108
  );


  not
  g323
  (
    n354,
    n195
  );


  not
  g324
  (
    n562,
    n100
  );


  buf
  g325
  (
    n746,
    n99
  );


  not
  g326
  (
    n689,
    n145
  );


  not
  g327
  (
    n719,
    n196
  );


  buf
  g328
  (
    n533,
    n52
  );


  not
  g329
  (
    n724,
    n213
  );


  not
  g330
  (
    n451,
    n53
  );


  not
  g331
  (
    n263,
    n153
  );


  buf
  g332
  (
    n678,
    n189
  );


  not
  g333
  (
    n636,
    n56
  );


  not
  g334
  (
    n658,
    n209
  );


  not
  g335
  (
    n810,
    n115
  );


  buf
  g336
  (
    n532,
    n214
  );


  buf
  g337
  (
    n894,
    n49
  );


  buf
  g338
  (
    n410,
    n117
  );


  buf
  g339
  (
    n396,
    n188
  );


  buf
  g340
  (
    n906,
    n58
  );


  not
  g341
  (
    n325,
    n134
  );


  not
  g342
  (
    n745,
    n140
  );


  not
  g343
  (
    n567,
    n99
  );


  not
  g344
  (
    n776,
    n82
  );


  not
  g345
  (
    n863,
    n67
  );


  not
  g346
  (
    n907,
    n116
  );


  buf
  g347
  (
    n287,
    n212
  );


  buf
  g348
  (
    n602,
    n168
  );


  buf
  g349
  (
    n883,
    n71
  );


  not
  g350
  (
    n734,
    n152
  );


  not
  g351
  (
    n903,
    n195
  );


  buf
  g352
  (
    n548,
    n138
  );


  not
  g353
  (
    n500,
    n189
  );


  not
  g354
  (
    n234,
    n71
  );


  buf
  g355
  (
    n748,
    n171
  );


  not
  g356
  (
    n596,
    n87
  );


  buf
  g357
  (
    n905,
    n105
  );


  not
  g358
  (
    n625,
    n121
  );


  not
  g359
  (
    n327,
    n164
  );


  buf
  g360
  (
    n433,
    n208
  );


  not
  g361
  (
    n712,
    n115
  );


  not
  g362
  (
    n670,
    n88
  );


  not
  g363
  (
    n753,
    n55
  );


  not
  g364
  (
    n549,
    n215
  );


  not
  g365
  (
    n605,
    n80
  );


  not
  g366
  (
    n687,
    n75
  );


  buf
  g367
  (
    n909,
    n175
  );


  buf
  g368
  (
    n457,
    n59
  );


  buf
  g369
  (
    n230,
    n72
  );


  buf
  g370
  (
    n887,
    n60
  );


  not
  g371
  (
    n781,
    n176
  );


  buf
  g372
  (
    n474,
    n141
  );


  not
  g373
  (
    n531,
    n145
  );


  buf
  g374
  (
    n555,
    n145
  );


  buf
  g375
  (
    n293,
    n215
  );


  not
  g376
  (
    n279,
    n188
  );


  not
  g377
  (
    n335,
    n50
  );


  not
  g378
  (
    n713,
    n183
  );


  buf
  g379
  (
    n699,
    n139
  );


  buf
  g380
  (
    n743,
    n215
  );


  buf
  g381
  (
    n758,
    n141
  );


  buf
  g382
  (
    n303,
    n211
  );


  buf
  g383
  (
    n697,
    n203
  );


  not
  g384
  (
    n873,
    n159
  );


  not
  g385
  (
    n890,
    n179
  );


  buf
  g386
  (
    n285,
    n165
  );


  buf
  g387
  (
    n647,
    n191
  );


  buf
  g388
  (
    n579,
    n129
  );


  not
  g389
  (
    n493,
    n201
  );


  not
  g390
  (
    n248,
    n96
  );


  buf
  g391
  (
    n675,
    n75
  );


  buf
  g392
  (
    n616,
    n148
  );


  not
  g393
  (
    n920,
    n138
  );


  not
  g394
  (
    n496,
    n127
  );


  buf
  g395
  (
    n423,
    n64
  );


  not
  g396
  (
    n811,
    n82
  );


  buf
  g397
  (
    n332,
    n165
  );


  buf
  g398
  (
    n409,
    n82
  );


  buf
  g399
  (
    n642,
    n181
  );


  buf
  g400
  (
    n470,
    n186
  );


  not
  g401
  (
    n720,
    n192
  );


  buf
  g402
  (
    n911,
    n109
  );


  not
  g403
  (
    n314,
    n68
  );


  not
  g404
  (
    n320,
    n113
  );


  buf
  g405
  (
    n854,
    n157
  );


  not
  g406
  (
    n761,
    n174
  );


  not
  g407
  (
    KeyWire_0_63,
    n168
  );


  not
  g408
  (
    n765,
    n120
  );


  buf
  g409
  (
    n558,
    n62
  );


  not
  g410
  (
    n366,
    n48
  );


  buf
  g411
  (
    n390,
    n182
  );


  buf
  g412
  (
    n565,
    n144
  );


  buf
  g413
  (
    n759,
    n113
  );


  buf
  g414
  (
    n630,
    n114
  );


  not
  g415
  (
    n570,
    n52
  );


  buf
  g416
  (
    n918,
    n151
  );


  not
  g417
  (
    n585,
    n159
  );


  not
  g418
  (
    n462,
    n147
  );


  not
  g419
  (
    n897,
    n217
  );


  not
  g420
  (
    n526,
    n93
  );


  buf
  g421
  (
    n688,
    n132
  );


  buf
  g422
  (
    n291,
    n148
  );


  not
  g423
  (
    n917,
    n129
  );


  not
  g424
  (
    n726,
    n183
  );


  not
  g425
  (
    n814,
    n122
  );


  not
  g426
  (
    n730,
    n79
  );


  not
  g427
  (
    n676,
    n108
  );


  buf
  g428
  (
    n795,
    n106
  );


  not
  g429
  (
    n617,
    n163
  );


  buf
  g430
  (
    n387,
    n206
  );


  buf
  g431
  (
    n503,
    n182
  );


  buf
  g432
  (
    n242,
    n198
  );


  buf
  g433
  (
    n283,
    n119
  );


  buf
  g434
  (
    n329,
    n208
  );


  buf
  g435
  (
    n317,
    n199
  );


  not
  g436
  (
    n252,
    n130
  );


  not
  g437
  (
    n334,
    n65
  );


  buf
  g438
  (
    n709,
    n197
  );


  buf
  g439
  (
    n672,
    n47
  );


  not
  g440
  (
    n715,
    n136
  );


  buf
  g441
  (
    n249,
    n126
  );


  not
  g442
  (
    n614,
    n55
  );


  not
  g443
  (
    n340,
    n59
  );


  not
  g444
  (
    n921,
    n50
  );


  buf
  g445
  (
    n621,
    n147
  );


  not
  g446
  (
    n478,
    n62
  );


  buf
  g447
  (
    n404,
    n169
  );


  not
  g448
  (
    n519,
    n74
  );


  not
  g449
  (
    n834,
    n73
  );


  not
  g450
  (
    n510,
    n61
  );


  not
  g451
  (
    n640,
    n138
  );


  buf
  g452
  (
    n770,
    n154
  );


  not
  g453
  (
    n523,
    n137
  );


  not
  g454
  (
    n288,
    n104
  );


  not
  g455
  (
    n495,
    n207
  );


  buf
  g456
  (
    n662,
    n70
  );


  not
  g457
  (
    n359,
    n49
  );


  not
  g458
  (
    n835,
    n213
  );


  not
  g459
  (
    n245,
    n216
  );


  buf
  g460
  (
    n888,
    n131
  );


  not
  g461
  (
    n786,
    n173
  );


  not
  g462
  (
    n696,
    n210
  );


  buf
  g463
  (
    n654,
    n95
  );


  not
  g464
  (
    n871,
    n75
  );


  buf
  g465
  (
    n259,
    n168
  );


  not
  g466
  (
    n362,
    n172
  );


  buf
  g467
  (
    n557,
    n131
  );


  buf
  g468
  (
    n480,
    n48
  );


  buf
  g469
  (
    n729,
    n87
  );


  not
  g470
  (
    n435,
    n73
  );


  buf
  g471
  (
    n635,
    n180
  );


  buf
  g472
  (
    n899,
    n101
  );


  not
  g473
  (
    n751,
    n123
  );


  buf
  g474
  (
    n756,
    n119
  );


  buf
  g475
  (
    n564,
    n205
  );


  not
  g476
  (
    n659,
    n104
  );


  buf
  g477
  (
    n492,
    n187
  );


  buf
  g478
  (
    n828,
    n136
  );


  buf
  g479
  (
    n554,
    n170
  );


  buf
  g480
  (
    n536,
    n61
  );


  buf
  g481
  (
    n639,
    n109
  );


  buf
  g482
  (
    n469,
    n97
  );


  not
  g483
  (
    n284,
    n167
  );


  buf
  g484
  (
    n764,
    n112
  );


  buf
  g485
  (
    n273,
    n214
  );


  not
  g486
  (
    n376,
    n200
  );


  buf
  g487
  (
    n880,
    n181
  );


  not
  g488
  (
    n842,
    n75
  );


  buf
  g489
  (
    n484,
    n204
  );


  buf
  g490
  (
    n534,
    n126
  );


  not
  g491
  (
    n750,
    n157
  );


  buf
  g492
  (
    n595,
    n91
  );


  buf
  g493
  (
    n299,
    n151
  );


  buf
  g494
  (
    n649,
    n164
  );


  not
  g495
  (
    n762,
    n173
  );


  not
  g496
  (
    n238,
    n141
  );


  not
  g497
  (
    n336,
    n202
  );


  not
  g498
  (
    KeyWire_0_61,
    n115
  );


  not
  g499
  (
    n778,
    n118
  );


  buf
  g500
  (
    n491,
    n143
  );


  not
  g501
  (
    n306,
    n83
  );


  buf
  g502
  (
    n913,
    n155
  );


  buf
  g503
  (
    n584,
    n120
  );


  not
  g504
  (
    n267,
    n45
  );


  not
  g505
  (
    n784,
    n72
  );


  buf
  g506
  (
    n783,
    n57
  );


  not
  g507
  (
    n403,
    n85
  );


  buf
  g508
  (
    n282,
    n74
  );


  buf
  g509
  (
    n298,
    n163
  );


  not
  g510
  (
    n374,
    n215
  );


  not
  g511
  (
    n415,
    n100
  );


  buf
  g512
  (
    n448,
    n64
  );


  buf
  g513
  (
    n467,
    n203
  );


  buf
  g514
  (
    n544,
    n68
  );


  buf
  g515
  (
    n603,
    n185
  );


  buf
  g516
  (
    n789,
    n155
  );


  not
  g517
  (
    KeyWire_0_20,
    n177
  );


  not
  g518
  (
    n693,
    n197
  );


  not
  g519
  (
    n465,
    n63
  );


  buf
  g520
  (
    n773,
    n188
  );


  buf
  g521
  (
    n702,
    n172
  );


  not
  g522
  (
    n680,
    n51
  );


  not
  g523
  (
    n551,
    n84
  );


  not
  g524
  (
    n700,
    n149
  );


  buf
  g525
  (
    n766,
    n179
  );


  not
  g526
  (
    n772,
    n190
  );


  not
  g527
  (
    n226,
    n84
  );


  not
  g528
  (
    n522,
    n95
  );


  not
  g529
  (
    n604,
    n91
  );


  buf
  g530
  (
    n578,
    n146
  );


  not
  g531
  (
    n669,
    n125
  );


  not
  g532
  (
    n486,
    n190
  );


  not
  g533
  (
    n331,
    n207
  );


  buf
  g534
  (
    n915,
    n112
  );


  buf
  g535
  (
    n429,
    n144
  );


  buf
  g536
  (
    n414,
    n134
  );


  not
  g537
  (
    n378,
    n133
  );


  buf
  g538
  (
    n235,
    n122
  );


  buf
  g539
  (
    n258,
    n132
  );


  not
  g540
  (
    n877,
    n111
  );


  buf
  g541
  (
    n228,
    n122
  );


  not
  g542
  (
    n754,
    n94
  );


  buf
  g543
  (
    n651,
    n132
  );


  not
  g544
  (
    n695,
    n46
  );


  not
  g545
  (
    n481,
    n142
  );


  buf
  g546
  (
    n296,
    n125
  );


  buf
  g547
  (
    n598,
    n201
  );


  not
  g548
  (
    n512,
    n169
  );


  not
  g549
  (
    n701,
    n66
  );


  not
  g550
  (
    n265,
    n119
  );


  not
  g551
  (
    n922,
    n120
  );


  buf
  g552
  (
    n817,
    n177
  );


  not
  g553
  (
    n418,
    n78
  );


  buf
  g554
  (
    n309,
    n80
  );


  buf
  g555
  (
    n790,
    n51
  );


  not
  g556
  (
    n482,
    n66
  );


  buf
  g557
  (
    n793,
    n89
  );


  buf
  g558
  (
    n326,
    n96
  );


  not
  g559
  (
    KeyWire_0_3,
    n181
  );


  buf
  g560
  (
    n816,
    n128
  );


  buf
  g561
  (
    n694,
    n118
  );


  not
  g562
  (
    n760,
    n174
  );


  not
  g563
  (
    n721,
    n97
  );


  not
  g564
  (
    n441,
    n195
  );


  buf
  g565
  (
    n440,
    n136
  );


  buf
  g566
  (
    n407,
    n86
  );


  not
  g567
  (
    n477,
    n188
  );


  not
  g568
  (
    n568,
    n191
  );


  buf
  g569
  (
    n910,
    n61
  );


  not
  g570
  (
    n690,
    n176
  );


  not
  g571
  (
    n445,
    n165
  );


  not
  g572
  (
    n472,
    n134
  );


  buf
  g573
  (
    n247,
    n95
  );


  buf
  g574
  (
    n833,
    n100
  );


  not
  g575
  (
    n898,
    n193
  );


  buf
  g576
  (
    n847,
    n206
  );


  buf
  g577
  (
    n798,
    n156
  );


  not
  g578
  (
    n892,
    n107
  );


  buf
  g579
  (
    n367,
    n64
  );


  buf
  g580
  (
    n237,
    n76
  );


  buf
  g581
  (
    n741,
    n114
  );


  buf
  g582
  (
    n785,
    n184
  );


  buf
  g583
  (
    n227,
    n147
  );


  not
  g584
  (
    n674,
    n169
  );


  not
  g585
  (
    n804,
    n159
  );


  not
  g586
  (
    n861,
    n64
  );


  not
  g587
  (
    n858,
    n139
  );


  not
  g588
  (
    n539,
    n166
  );


  not
  g589
  (
    n722,
    n98
  );


  not
  g590
  (
    n446,
    n107
  );


  buf
  g591
  (
    n357,
    n160
  );


  not
  g592
  (
    n737,
    n78
  );


  not
  g593
  (
    n671,
    n123
  );


  not
  g594
  (
    n269,
    n68
  );


  buf
  g595
  (
    n358,
    n199
  );


  not
  g596
  (
    n677,
    n56
  );


  not
  g597
  (
    n364,
    n202
  );


  not
  g598
  (
    n633,
    n49
  );


  buf
  g599
  (
    n638,
    n162
  );


  buf
  g600
  (
    n800,
    n192
  );


  not
  g601
  (
    n412,
    n90
  );


  buf
  g602
  (
    n663,
    n152
  );


  buf
  g603
  (
    n321,
    n116
  );


  not
  g604
  (
    n885,
    n126
  );


  not
  g605
  (
    n489,
    n208
  );


  not
  g606
  (
    n525,
    n51
  );


  buf
  g607
  (
    n386,
    n119
  );


  not
  g608
  (
    n432,
    n108
  );


  not
  g609
  (
    n276,
    n212
  );


  not
  g610
  (
    n593,
    n91
  );


  buf
  g611
  (
    n839,
    n202
  );


  not
  g612
  (
    n347,
    n191
  );


  not
  g613
  (
    n901,
    n130
  );


  buf
  g614
  (
    n406,
    n151
  );


  buf
  g615
  (
    n319,
    n128
  );


  buf
  g616
  (
    n822,
    n130
  );


  not
  g617
  (
    n391,
    n149
  );


  not
  g618
  (
    n727,
    n220
  );


  buf
  g619
  (
    n808,
    n76
  );


  not
  g620
  (
    n454,
    n74
  );


  buf
  g621
  (
    n243,
    n66
  );


  buf
  g622
  (
    n812,
    n184
  );


  not
  g623
  (
    n514,
    n158
  );


  buf
  g624
  (
    n373,
    n88
  );


  not
  g625
  (
    n608,
    n62
  );


  buf
  g626
  (
    n845,
    n120
  );


  not
  g627
  (
    KeyWire_0_25,
    n83
  );


  buf
  g628
  (
    n535,
    n199
  );


  buf
  g629
  (
    n606,
    n56
  );


  buf
  g630
  (
    n316,
    n178
  );


  not
  g631
  (
    n718,
    n203
  );


  buf
  g632
  (
    n458,
    n190
  );


  not
  g633
  (
    n893,
    n156
  );


  buf
  g634
  (
    n511,
    n45
  );


  not
  g635
  (
    n389,
    n105
  );


  not
  g636
  (
    n420,
    n58
  );


  not
  g637
  (
    n260,
    n217
  );


  buf
  g638
  (
    n221,
    n72
  );


  not
  g639
  (
    n424,
    n102
  );


  not
  g640
  (
    n301,
    n87
  );


  buf
  g641
  (
    n286,
    n212
  );


  buf
  g642
  (
    n582,
    n113
  );


  buf
  g643
  (
    n857,
    n98
  );


  buf
  g644
  (
    n747,
    n144
  );


  buf
  g645
  (
    n428,
    n118
  );


  not
  g646
  (
    n815,
    n47
  );


  not
  g647
  (
    n600,
    n160
  );


  not
  g648
  (
    n613,
    n65
  );


  buf
  g649
  (
    n652,
    n65
  );


  buf
  g650
  (
    n588,
    n111
  );


  not
  g651
  (
    n343,
    n124
  );


  not
  g652
  (
    n629,
    n127
  );


  buf
  g653
  (
    n239,
    n124
  );


  not
  g654
  (
    n601,
    n213
  );


  not
  g655
  (
    n487,
    n115
  );


  not
  g656
  (
    n300,
    n57
  );


  not
  g657
  (
    n703,
    n74
  );


  not
  g658
  (
    n546,
    n198
  );


  buf
  g659
  (
    n914,
    n198
  );


  buf
  g660
  (
    n438,
    n194
  );


  buf
  g661
  (
    n820,
    n181
  );


  buf
  g662
  (
    n450,
    n144
  );


  not
  g663
  (
    n257,
    n163
  );


  buf
  g664
  (
    n561,
    n99
  );


  buf
  g665
  (
    n516,
    n219
  );


  not
  g666
  (
    n660,
    n136
  );


  not
  g667
  (
    n609,
    n205
  );


  buf
  g668
  (
    n867,
    n187
  );


  buf
  g669
  (
    n509,
    n117
  );


  not
  g670
  (
    n728,
    n97
  );


  not
  g671
  (
    KeyWire_0_50,
    n219
  );


  buf
  g672
  (
    n836,
    n220
  );


  not
  g673
  (
    n411,
    n199
  );


  not
  g674
  (
    n813,
    n186
  );


  buf
  g675
  (
    n231,
    n79
  );


  buf
  g676
  (
    n818,
    n107
  );


  not
  g677
  (
    n380,
    n121
  );


  not
  g678
  (
    n471,
    n159
  );


  buf
  g679
  (
    KeyWire_0_22,
    n138
  );


  not
  g680
  (
    n856,
    n111
  );


  buf
  g681
  (
    n650,
    n210
  );


  buf
  g682
  (
    n307,
    n141
  );


  buf
  g683
  (
    n573,
    n192
  );


  not
  g684
  (
    n732,
    n69
  );


  not
  g685
  (
    n655,
    n173
  );


  buf
  g686
  (
    n851,
    n171
  );


  buf
  g687
  (
    n792,
    n171
  );


  buf
  g688
  (
    n731,
    n79
  );


  buf
  g689
  (
    n530,
    n93
  );


  not
  g690
  (
    n912,
    n117
  );


  buf
  g691
  (
    n305,
    n58
  );


  buf
  g692
  (
    n902,
    n112
  );


  buf
  g693
  (
    n853,
    n150
  );


  buf
  g694
  (
    n809,
    n94
  );


  not
  g695
  (
    n513,
    n54
  );


  buf
  g696
  (
    n543,
    n90
  );


  not
  g697
  (
    n735,
    n150
  );


  buf
  g698
  (
    n916,
    n93
  );


  buf
  g699
  (
    n872,
    n78
  );


  buf
  g700
  (
    n736,
    n209
  );


  not
  g701
  (
    n308,
    n175
  );


  not
  g702
  (
    n686,
    n196
  );


  buf
  g703
  (
    n345,
    n114
  );


  buf
  g704
  (
    n904,
    n175
  );


  not
  g705
  (
    n274,
    n123
  );


  not
  g706
  (
    n831,
    n192
  );


  buf
  g707
  (
    n222,
    n77
  );


  not
  g708
  (
    n744,
    n166
  );


  buf
  g709
  (
    n864,
    n189
  );


  buf
  g710
  (
    n483,
    n92
  );


  not
  g711
  (
    n698,
    n140
  );


  buf
  g712
  (
    n607,
    n69
  );


  not
  g713
  (
    KeyWire_0_1,
    n97
  );


  not
  g714
  (
    n837,
    n166
  );


  buf
  g715
  (
    n827,
    n46
  );


  buf
  g716
  (
    n310,
    n76
  );


  buf
  g717
  (
    n769,
    n217
  );


  not
  g718
  (
    n599,
    n162
  );


  buf
  g719
  (
    n896,
    n112
  );


  buf
  g720
  (
    n290,
    n194
  );


  not
  g721
  (
    n859,
    n189
  );


  not
  g722
  (
    n355,
    n213
  );


  buf
  g723
  (
    n504,
    n113
  );


  buf
  g724
  (
    n466,
    n210
  );


  buf
  g725
  (
    n280,
    n203
  );


  not
  g726
  (
    n710,
    n67
  );


  not
  g727
  (
    n443,
    n90
  );


  not
  g728
  (
    n537,
    n161
  );


  not
  g729
  (
    n297,
    n110
  );


  buf
  g730
  (
    n807,
    n124
  );


  not
  g731
  (
    n225,
    n129
  );


  not
  g732
  (
    n337,
    n162
  );


  not
  g733
  (
    KeyWire_0_41,
    n135
  );


  buf
  g734
  (
    n520,
    n176
  );


  not
  g735
  (
    n344,
    n135
  );


  not
  g736
  (
    n460,
    n205
  );


  buf
  g737
  (
    n315,
    n206
  );


  buf
  g738
  (
    n405,
    n185
  );


  not
  g739
  (
    n545,
    n160
  );


  buf
  g740
  (
    n368,
    n178
  );


  buf
  g741
  (
    n393,
    n135
  );


  not
  g742
  (
    n352,
    n110
  );


  buf
  g743
  (
    n379,
    n90
  );


  not
  g744
  (
    n333,
    n161
  );


  not
  g745
  (
    n574,
    n125
  );


  not
  g746
  (
    n294,
    n172
  );


  not
  g747
  (
    n563,
    n172
  );


  not
  g748
  (
    n330,
    n214
  );


  not
  g749
  (
    n875,
    n167
  );


  not
  g750
  (
    n289,
    n59
  );


  buf
  g751
  (
    n886,
    n105
  );


  not
  g752
  (
    n716,
    n142
  );


  not
  g753
  (
    n706,
    n178
  );


  not
  g754
  (
    n313,
    n180
  );


  buf
  g755
  (
    n725,
    n158
  );


  buf
  g756
  (
    n656,
    n102
  );


  not
  g757
  (
    n796,
    n49
  );


  not
  g758
  (
    n787,
    n154
  );


  not
  g759
  (
    n646,
    n177
  );


  buf
  g760
  (
    n277,
    n154
  );


  not
  g761
  (
    n508,
    n131
  );


  not
  g762
  (
    n246,
    n143
  );


  not
  g763
  (
    n705,
    n146
  );


  not
  g764
  (
    KeyWire_0_9,
    n150
  );


  buf
  g765
  (
    n395,
    n130
  );


  buf
  g766
  (
    n860,
    n128
  );


  buf
  g767
  (
    n583,
    n69
  );


  buf
  g768
  (
    n324,
    n134
  );


  not
  g769
  (
    n667,
    n218
  );


  buf
  g770
  (
    n302,
    n62
  );


  not
  g771
  (
    n576,
    n70
  );


  buf
  g772
  (
    n717,
    n101
  );


  not
  g773
  (
    n541,
    n68
  );


  buf
  g774
  (
    n281,
    n77
  );


  not
  g775
  (
    n223,
    n81
  );


  not
  g776
  (
    n620,
    n139
  );


  not
  g777
  (
    n874,
    n170
  );


  not
  g778
  (
    n507,
    n186
  );


  not
  g779
  (
    n419,
    n216
  );


  buf
  g780
  (
    n742,
    n179
  );


  not
  g781
  (
    n862,
    n92
  );


  buf
  g782
  (
    n797,
    n122
  );


  not
  g783
  (
    n590,
    n92
  );


  not
  g784
  (
    n615,
    n160
  );


  not
  g785
  (
    n517,
    n153
  );


  not
  g786
  (
    n803,
    n103
  );


  buf
  g787
  (
    n846,
    n148
  );


  buf
  g788
  (
    n240,
    n80
  );


  not
  g789
  (
    n292,
    n61
  );


  not
  g790
  (
    n312,
    n109
  );


  buf
  g791
  (
    n455,
    n204
  );


  buf
  g792
  (
    n866,
    n65
  );


  buf
  g793
  (
    n229,
    n190
  );


  not
  g794
  (
    n569,
    n206
  );


  buf
  g795
  (
    n383,
    n193
  );


  not
  g796
  (
    n444,
    n155
  );


  buf
  g797
  (
    n679,
    n209
  );


  buf
  g798
  (
    n377,
    n98
  );


  buf
  g799
  (
    n752,
    n116
  );


  not
  g800
  (
    n473,
    n121
  );


  not
  g801
  (
    n439,
    n212
  );


  buf
  g802
  (
    n587,
    n147
  );


  buf
  g803
  (
    n397,
    n148
  );


  not
  g804
  (
    n502,
    n89
  );


  not
  g805
  (
    n394,
    n143
  );


  not
  g806
  (
    n261,
    n67
  );


  buf
  g807
  (
    KeyWire_0_30,
    n46
  );


  buf
  g808
  (
    n684,
    n78
  );


  not
  g809
  (
    n553,
    n105
  );


  buf
  g810
  (
    n571,
    n180
  );


  buf
  g811
  (
    n275,
    n89
  );


  buf
  g812
  (
    n255,
    n121
  );


  not
  g813
  (
    n891,
    n91
  );


  buf
  g814
  (
    n749,
    n201
  );


  buf
  g815
  (
    n232,
    n102
  );


  buf
  g816
  (
    n841,
    n207
  );


  not
  g817
  (
    n628,
    n145
  );


  not
  g818
  (
    KeyWire_0_18,
    n139
  );


  buf
  g819
  (
    n622,
    n137
  );


  buf
  g820
  (
    n879,
    n106
  );


  not
  g821
  (
    n634,
    n166
  );


  buf
  g822
  (
    n673,
    n173
  );


  buf
  g823
  (
    n775,
    n60
  );


  not
  g824
  (
    n434,
    n117
  );


  not
  g825
  (
    n876,
    n114
  );


  not
  g826
  (
    n919,
    n108
  );


  buf
  g827
  (
    n461,
    n50
  );


  not
  g828
  (
    n529,
    n116
  );


  not
  g829
  (
    n264,
    n195
  );


  buf
  g830
  (
    n251,
    n57
  );


  not
  g831
  (
    n843,
    n153
  );


  not
  g832
  (
    n417,
    n135
  );


  not
  g833
  (
    n452,
    n193
  );


  buf
  g834
  (
    n542,
    n77
  );


  buf
  g835
  (
    n447,
    n146
  );


  buf
  g836
  (
    n369,
    n103
  );


  not
  g837
  (
    n341,
    n204
  );


  buf
  g838
  (
    n224,
    n54
  );


  buf
  g839
  (
    n360,
    n183
  );


  buf
  g840
  (
    n692,
    n45
  );


  buf
  g841
  (
    n849,
    n196
  );


  not
  g842
  (
    n924,
    n128
  );


  not
  g843
  (
    n631,
    n52
  );


  not
  g844
  (
    n350,
    n129
  );


  not
  g845
  (
    n832,
    n142
  );


  buf
  g846
  (
    n757,
    n150
  );


  buf
  g847
  (
    n295,
    n218
  );


  not
  g848
  (
    n250,
    n162
  );


  not
  g849
  (
    n426,
    n107
  );


  buf
  g850
  (
    n685,
    n184
  );


  buf
  g851
  (
    n408,
    n202
  );


  buf
  g852
  (
    n353,
    n110
  );


  buf
  g853
  (
    n475,
    n69
  );


  buf
  g854
  (
    n398,
    n111
  );


  not
  g855
  (
    n401,
    n174
  );


  buf
  g856
  (
    n868,
    n154
  );


  buf
  g857
  (
    n619,
    n127
  );


  buf
  g858
  (
    n682,
    n156
  );


  not
  g859
  (
    n739,
    n137
  );


  not
  g860
  (
    n453,
    n131
  );


  buf
  g861
  (
    KeyWire_0_17,
    n152
  );


  not
  g862
  (
    n349,
    n88
  );


  not
  g863
  (
    n468,
    n137
  );


  buf
  g864
  (
    n436,
    n110
  );


  not
  g865
  (
    n714,
    n211
  );


  buf
  g866
  (
    n363,
    n58
  );


  not
  g867
  (
    n272,
    n53
  );


  buf
  g868
  (
    n683,
    n185
  );


  buf
  g869
  (
    n767,
    n157
  );


  not
  g870
  (
    n413,
    n124
  );


  not
  g871
  (
    n850,
    n153
  );


  not
  g872
  (
    n771,
    n133
  );


  buf
  g873
  (
    n494,
    n211
  );


  not
  g874
  (
    n515,
    n96
  );


  not
  g875
  (
    n262,
    n196
  );


  buf
  g876
  (
    n304,
    n218
  );


  buf
  g877
  (
    n528,
    n211
  );


  not
  g878
  (
    n339,
    n95
  );


  buf
  g879
  (
    n278,
    n156
  );


  xor
  g880
  (
    n931,
    n234,
    n238,
    n242,
    n221
  );


  xnor
  g881
  (
    n930,
    n252,
    n248,
    n249,
    n233
  );


  xnor
  g882
  (
    n936,
    n245,
    n234,
    n240,
    n228
  );


  xnor
  g883
  (
    n929,
    n227,
    n230,
    n241,
    n248
  );


  nor
  g884
  (
    n938,
    n246,
    n251,
    n229,
    n244
  );


  xor
  g885
  (
    n935,
    n246,
    n229,
    n231,
    n240
  );


  nand
  g886
  (
    n933,
    n232,
    n237,
    n247,
    n223
  );


  and
  g887
  (
    n937,
    n236,
    n250,
    n252
  );


  xnor
  g888
  (
    n934,
    n239,
    n241,
    n245,
    n224
  );


  nor
  g889
  (
    n939,
    n228,
    n236,
    n226,
    n235
  );


  and
  g890
  (
    n940,
    n242,
    n233,
    n226,
    n247
  );


  and
  g891
  (
    n932,
    n249,
    n243,
    n224,
    n238
  );


  xnor
  g892
  (
    n928,
    n243,
    n223,
    n221,
    n231
  );


  and
  g893
  (
    n925,
    n230,
    n244,
    n222
  );


  and
  g894
  (
    n926,
    n237,
    n225,
    n232,
    n227
  );


  nor
  g895
  (
    n927,
    n235,
    n239,
    n251,
    n225
  );


  not
  g896
  (
    n941,
    n939
  );


  buf
  g897
  (
    n942,
    n940
  );


  buf
  g898
  (
    n943,
    n942
  );


  buf
  g899
  (
    n944,
    n942
  );


  not
  g900
  (
    n945,
    n942
  );


  not
  g901
  (
    n947,
    n942
  );


  not
  g902
  (
    n950,
    n941
  );


  not
  g903
  (
    n948,
    n941
  );


  buf
  g904
  (
    n946,
    n941
  );


  not
  g905
  (
    n949,
    n941
  );


  not
  g906
  (
    n954,
    n944
  );


  not
  g907
  (
    n953,
    n943
  );


  buf
  g908
  (
    n955,
    n943
  );


  buf
  g909
  (
    n951,
    n943
  );


  not
  g910
  (
    n952,
    n943
  );


  nor
  g911
  (
    n957,
    n944,
    n955,
    n945,
    n954
  );


  nor
  g912
  (
    n956,
    n256,
    n256,
    n955,
    n255
  );


  xnor
  g913
  (
    n963,
    n947,
    n945,
    n953
  );


  or
  g914
  (
    n958,
    n257,
    n945,
    n954,
    n952
  );


  and
  g915
  (
    n959,
    n254,
    n254,
    n944,
    n952
  );


  nor
  g916
  (
    n960,
    n253,
    n255,
    n944,
    n946
  );


  or
  g917
  (
    n961,
    n953,
    n951,
    n946,
    n253
  );


  nor
  g918
  (
    n962,
    n257,
    n946,
    n951
  );


  not
  g919
  (
    n968,
    n961
  );


  buf
  g920
  (
    n973,
    n963
  );


  buf
  g921
  (
    n971,
    n959
  );


  buf
  g922
  (
    n967,
    n956
  );


  not
  g923
  (
    n965,
    n958
  );


  not
  g924
  (
    n970,
    n960
  );


  buf
  g925
  (
    n966,
    n962
  );


  buf
  g926
  (
    n969,
    n957
  );


  not
  g927
  (
    KeyWire_0_62,
    n962
  );


  not
  g928
  (
    n972,
    n963
  );


  xnor
  g929
  (
    n979,
    n969,
    n264,
    n276,
    n291
  );


  or
  g930
  (
    n977,
    n296,
    n273,
    n259,
    n279
  );


  nand
  g931
  (
    n982,
    n281,
    n293,
    n270,
    n966
  );


  and
  g932
  (
    n989,
    n971,
    n288,
    n966,
    n264
  );


  nand
  g933
  (
    n978,
    n278,
    n296,
    n275,
    n277
  );


  or
  g934
  (
    n994,
    n290,
    n276,
    n294,
    n277
  );


  xor
  g935
  (
    n976,
    n267,
    n971,
    n283,
    n299
  );


  and
  g936
  (
    n992,
    n287,
    n269,
    n289,
    n279
  );


  nor
  g937
  (
    n983,
    n295,
    n268,
    n272,
    n266
  );


  and
  g938
  (
    n988,
    n263,
    n964,
    n274,
    n265
  );


  xnor
  g939
  (
    n999,
    n299,
    n967,
    n965
  );


  xor
  g940
  (
    n991,
    n968,
    n259,
    n290,
    n289
  );


  nand
  g941
  (
    KeyWire_0_60,
    n292,
    n970,
    n273,
    n964
  );


  or
  g942
  (
    n1003,
    n260,
    n285,
    n965,
    n291
  );


  xor
  g943
  (
    n985,
    n293,
    n292,
    n297,
    n301
  );


  or
  g944
  (
    n1000,
    n262,
    n258,
    n969,
    n298
  );


  xnor
  g945
  (
    n998,
    n280,
    n300,
    n287,
    n970
  );


  xor
  g946
  (
    n1002,
    n261,
    n969,
    n284,
    n274
  );


  xnor
  g947
  (
    n984,
    n272,
    n280,
    n966,
    n269
  );


  and
  g948
  (
    n990,
    n278,
    n268,
    n286,
    n263
  );


  or
  g949
  (
    n980,
    n275,
    n266,
    n260,
    n285
  );


  nor
  g950
  (
    n1001,
    n286,
    n282,
    n967
  );


  xnor
  g951
  (
    n986,
    n968,
    n294,
    n964,
    n261
  );


  or
  g952
  (
    n974,
    n265,
    n965,
    n281,
    n283
  );


  xor
  g953
  (
    n997,
    n302,
    n295,
    n301,
    n297
  );


  nor
  g954
  (
    n987,
    n271,
    n298,
    n968,
    n288
  );


  nand
  g955
  (
    n995,
    n965,
    n300,
    n271,
    n969
  );


  nor
  g956
  (
    n996,
    n282,
    n270,
    n970,
    n966
  );


  or
  g957
  (
    n993,
    n284,
    n258,
    n262,
    n968
  );


  or
  g958
  (
    n981,
    n302,
    n964,
    n267,
    n970
  );


  not
  g959
  (
    n1014,
    n977
  );


  buf
  g960
  (
    n1005,
    n975
  );


  not
  g961
  (
    n1012,
    n974
  );


  buf
  g962
  (
    n1007,
    n979
  );


  not
  g963
  (
    n1013,
    n981
  );


  not
  g964
  (
    KeyWire_0_11,
    n981
  );


  buf
  g965
  (
    n1006,
    n978
  );


  not
  g966
  (
    n1015,
    n976
  );


  not
  g967
  (
    KeyWire_0_27,
    n976
  );


  not
  g968
  (
    KeyWire_0_15,
    n978
  );


  nand
  g969
  (
    n1011,
    n974,
    n979
  );


  and
  g970
  (
    n1009,
    n975,
    n980,
    n977
  );


  not
  g971
  (
    n1024,
    n1004
  );


  buf
  g972
  (
    n1021,
    n1005
  );


  not
  g973
  (
    n1031,
    n1005
  );


  buf
  g974
  (
    n1017,
    n1004
  );


  not
  g975
  (
    n1030,
    n1007
  );


  buf
  g976
  (
    n1023,
    n1005
  );


  buf
  g977
  (
    n1019,
    n1007
  );


  buf
  g978
  (
    n1022,
    n1006
  );


  buf
  g979
  (
    n1016,
    n1006
  );


  not
  g980
  (
    n1028,
    n1004
  );


  buf
  g981
  (
    n1025,
    n1004
  );


  buf
  g982
  (
    n1029,
    n1007
  );


  not
  g983
  (
    n1020,
    n1005
  );


  not
  g984
  (
    n1027,
    n1007
  );


  not
  g985
  (
    n1026,
    n1006
  );


  not
  g986
  (
    n1018,
    n1006
  );


  buf
  g987
  (
    n1033,
    n1016
  );


  not
  g988
  (
    n1032,
    n1016
  );


  xnor
  g989
  (
    n1040,
    n1032,
    n1017,
    n1033
  );


  or
  g990
  (
    n1034,
    n1025,
    n1021,
    n304,
    n1020
  );


  xnor
  g991
  (
    n1035,
    n1022,
    n1017,
    n1024
  );


  or
  g992
  (
    n1039,
    n1019,
    n303,
    n1018,
    n1023
  );


  nor
  g993
  (
    n1036,
    n1026,
    n1032,
    n1033,
    n1023
  );


  and
  g994
  (
    n1038,
    n1032,
    n1019,
    n1033,
    n947
  );


  xnor
  g995
  (
    n1041,
    n303,
    n1032,
    n1021,
    n1025
  );


  and
  g996
  (
    n1037,
    n304,
    n1020,
    n1022,
    n1018
  );


  not
  g997
  (
    n1050,
    n982
  );


  not
  g998
  (
    n1043,
    n1040
  );


  not
  g999
  (
    n1053,
    n305
  );


  not
  g1000
  (
    n1047,
    n973
  );


  not
  g1001
  (
    n1049,
    n1034
  );


  not
  g1002
  (
    n1045,
    n1041
  );


  not
  g1003
  (
    n1044,
    n972
  );


  or
  g1004
  (
    n1042,
    n1037,
    n1040,
    n972
  );


  and
  g1005
  (
    n1048,
    n1036,
    n1039,
    n971,
    n1038
  );


  xnor
  g1006
  (
    n1051,
    n982,
    n972,
    n983,
    n306
  );


  nor
  g1007
  (
    n1052,
    n1038,
    n1041,
    n971,
    n305
  );


  nor
  g1008
  (
    n1046,
    n973,
    n1039,
    n1035,
    n972
  );


  not
  g1009
  (
    n1066,
    n1048
  );


  buf
  g1010
  (
    n1074,
    n1051
  );


  buf
  g1011
  (
    n1069,
    n1049
  );


  buf
  g1012
  (
    n1060,
    n1047
  );


  buf
  g1013
  (
    n1063,
    n1049
  );


  not
  g1014
  (
    n1081,
    n1047
  );


  buf
  g1015
  (
    n1070,
    n1050
  );


  not
  g1016
  (
    n1078,
    n1045
  );


  not
  g1017
  (
    n1073,
    n1044
  );


  not
  g1018
  (
    n1064,
    n1043
  );


  not
  g1019
  (
    n1079,
    n1044
  );


  buf
  g1020
  (
    n1075,
    n1048
  );


  not
  g1021
  (
    n1080,
    n1045
  );


  not
  g1022
  (
    n1077,
    n1042
  );


  not
  g1023
  (
    n1059,
    n1043
  );


  buf
  g1024
  (
    n1067,
    n1044
  );


  not
  g1025
  (
    n1056,
    n1046
  );


  buf
  g1026
  (
    n1072,
    n1050
  );


  not
  g1027
  (
    n1054,
    n1046
  );


  not
  g1028
  (
    n1062,
    n1051
  );


  buf
  g1029
  (
    n1068,
    n1042
  );


  buf
  g1030
  (
    n1061,
    n1048
  );


  not
  g1031
  (
    n1055,
    n1049
  );


  buf
  g1032
  (
    n1065,
    n1045
  );


  buf
  g1033
  (
    n1057,
    n1046
  );


  buf
  g1034
  (
    n1071,
    n1047
  );


  buf
  g1035
  (
    n1076,
    n1050
  );


  buf
  g1036
  (
    n1058,
    n1043
  );


  not
  g1037
  (
    n1137,
    n1057
  );


  not
  g1038
  (
    n1149,
    n1064
  );


  buf
  g1039
  (
    n1127,
    n1074
  );


  buf
  g1040
  (
    n1131,
    n1075
  );


  not
  g1041
  (
    n1155,
    n1009
  );


  not
  g1042
  (
    n1083,
    n1014
  );


  not
  g1043
  (
    KeyWire_0_43,
    n1013
  );


  not
  g1044
  (
    n1090,
    n1000
  );


  buf
  g1045
  (
    n1092,
    n1057
  );


  not
  g1046
  (
    n1128,
    n1071
  );


  not
  g1047
  (
    n1104,
    n1067
  );


  not
  g1048
  (
    n1160,
    n1065
  );


  not
  g1049
  (
    n1101,
    n987
  );


  buf
  g1050
  (
    n1157,
    n1080
  );


  not
  g1051
  (
    n1165,
    n1012
  );


  buf
  g1052
  (
    n1088,
    n1064
  );


  buf
  g1053
  (
    n1141,
    n1075
  );


  buf
  g1054
  (
    n1097,
    n1013
  );


  buf
  g1055
  (
    n1122,
    n1055
  );


  buf
  g1056
  (
    n1188,
    n1009
  );


  buf
  g1057
  (
    n1171,
    n1079
  );


  buf
  g1058
  (
    n1173,
    n1071
  );


  not
  g1059
  (
    n1093,
    n1061
  );


  not
  g1060
  (
    KeyWire_0_35,
    n1081
  );


  buf
  g1061
  (
    n1106,
    n990
  );


  not
  g1062
  (
    n1145,
    n1012
  );


  not
  g1063
  (
    n1151,
    n1063
  );


  buf
  g1064
  (
    n1189,
    n1011
  );


  not
  g1065
  (
    n1094,
    n1070
  );


  buf
  g1066
  (
    n1182,
    n1014
  );


  buf
  g1067
  (
    n1191,
    n985
  );


  not
  g1068
  (
    n1169,
    n1077
  );


  not
  g1069
  (
    KeyWire_0_38,
    n994
  );


  buf
  g1070
  (
    n1193,
    n1069
  );


  buf
  g1071
  (
    n1132,
    n1080
  );


  not
  g1072
  (
    n1111,
    n1054
  );


  buf
  g1073
  (
    n1146,
    n991
  );


  buf
  g1074
  (
    n1087,
    n1008
  );


  not
  g1075
  (
    n1129,
    n1072
  );


  not
  g1076
  (
    n1139,
    n1002
  );


  not
  g1077
  (
    n1161,
    n1060
  );


  not
  g1078
  (
    n1109,
    n1081
  );


  buf
  g1079
  (
    n1159,
    n1063
  );


  not
  g1080
  (
    n1192,
    n1062
  );


  not
  g1081
  (
    n1110,
    n1059
  );


  not
  g1082
  (
    n1130,
    n1061
  );


  buf
  g1083
  (
    n1095,
    n1081
  );


  not
  g1084
  (
    n1086,
    n991
  );


  not
  g1085
  (
    n1153,
    n1078
  );


  buf
  g1086
  (
    n1140,
    n1070
  );


  buf
  g1087
  (
    n1150,
    n1062
  );


  not
  g1088
  (
    n1098,
    n1055
  );


  buf
  g1089
  (
    n1120,
    n1002
  );


  not
  g1090
  (
    n1183,
    n1073
  );


  buf
  g1091
  (
    n1180,
    n1071
  );


  not
  g1092
  (
    n1099,
    n1015
  );


  buf
  g1093
  (
    n1158,
    n1070
  );


  buf
  g1094
  (
    n1112,
    n1057
  );


  not
  g1095
  (
    n1166,
    n1067
  );


  buf
  g1096
  (
    n1142,
    n1080
  );


  buf
  g1097
  (
    n1163,
    n1073
  );


  not
  g1098
  (
    n1176,
    n1059
  );


  not
  g1099
  (
    n1103,
    n992
  );


  buf
  g1100
  (
    n1156,
    n1062
  );


  not
  g1101
  (
    n1118,
    n1059
  );


  buf
  g1102
  (
    n1134,
    n1068
  );


  not
  g1103
  (
    n1108,
    n1076
  );


  buf
  g1104
  (
    n1154,
    n1008
  );


  buf
  g1105
  (
    n1167,
    n1011
  );


  buf
  g1106
  (
    n1121,
    n997
  );


  not
  g1107
  (
    n1187,
    n1011
  );


  buf
  g1108
  (
    n1172,
    n1073
  );


  buf
  g1109
  (
    n1102,
    n989
  );


  buf
  g1110
  (
    n1190,
    n1054
  );


  not
  g1111
  (
    n1175,
    n990
  );


  buf
  g1112
  (
    n1136,
    n1079
  );


  buf
  g1113
  (
    n1089,
    n987
  );


  not
  g1114
  (
    n1105,
    n988
  );


  not
  g1115
  (
    n1174,
    n996
  );


  buf
  g1116
  (
    n1082,
    n985
  );


  not
  g1117
  (
    n1135,
    n1061
  );


  buf
  g1118
  (
    KeyWire_0_0,
    n1067
  );


  buf
  g1119
  (
    n1152,
    n993
  );


  buf
  g1120
  (
    n1186,
    n1081
  );


  buf
  g1121
  (
    KeyWire_0_28,
    n1078
  );


  not
  g1122
  (
    n1144,
    n1056
  );


  buf
  g1123
  (
    n1107,
    n1068
  );


  not
  g1124
  (
    n1117,
    n1058
  );


  not
  g1125
  (
    n1133,
    n988
  );


  or
  g1126
  (
    n1177,
    n1064,
    n1066,
    n1001,
    n1071
  );


  nand
  g1127
  (
    n1168,
    n1065,
    n995,
    n1010,
    n1068
  );


  or
  g1128
  (
    n1162,
    n983,
    n1056,
    n1078
  );


  xor
  g1129
  (
    n1126,
    n1054,
    n1069,
    n1070,
    n1075
  );


  xor
  g1130
  (
    n1164,
    n1013,
    n1079,
    n1010,
    n1000
  );


  nor
  g1131
  (
    n1185,
    n1079,
    n1060,
    n1015,
    n1058
  );


  and
  g1132
  (
    n1123,
    n1066,
    n1074,
    n1065,
    n1063
  );


  or
  g1133
  (
    n1124,
    n1008,
    n989,
    n992,
    n1056
  );


  xnor
  g1134
  (
    n1116,
    n1014,
    n995,
    n1009,
    n1069
  );


  xnor
  g1135
  (
    n1170,
    n1077,
    n1060,
    n1054,
    n1008
  );


  nor
  g1136
  (
    n1096,
    n1072,
    n1065,
    n1080,
    n1009
  );


  xor
  g1137
  (
    n1113,
    n1055,
    n1058
  );


  nor
  g1138
  (
    n1138,
    n1061,
    n1010,
    n1059,
    n1011
  );


  xor
  g1139
  (
    n1178,
    n1062,
    n984,
    n1063
  );


  nand
  g1140
  (
    n1148,
    n1074,
    n994,
    n1001,
    n1067
  );


  xor
  g1141
  (
    n1114,
    n999,
    n1077,
    n1076,
    n998
  );


  xnor
  g1142
  (
    n1119,
    n999,
    n996,
    n1060,
    n1077
  );


  xor
  g1143
  (
    n1084,
    n1074,
    n998,
    n1073,
    n986
  );


  and
  g1144
  (
    n1125,
    n1076,
    n1075,
    n993,
    n1069
  );


  xnor
  g1145
  (
    n1179,
    n997,
    n1076,
    n1066,
    n1068
  );


  xnor
  g1146
  (
    n1184,
    n1072,
    n986,
    n1010,
    n1066
  );


  xor
  g1147
  (
    n1085,
    n1012,
    n1014,
    n1056,
    n1064
  );


  xor
  g1148
  (
    n1181,
    n1072,
    n1012,
    n1057,
    n1013
  );


  xor
  g1149
  (
    n1208,
    n623,
    n559,
    n562,
    n658
  );


  nor
  g1150
  (
    n1332,
    n1144,
    n351,
    n695,
    n347
  );


  and
  g1151
  (
    n1444,
    n599,
    n650,
    n1098,
    n364
  );


  xnor
  g1152
  (
    n1634,
    n1088,
    n556,
    n377,
    n561
  );


  and
  g1153
  (
    n1238,
    n535,
    n625,
    n611,
    n643
  );


  xor
  g1154
  (
    n1350,
    n666,
    n1127,
    n1137,
    n550
  );


  nor
  g1155
  (
    n1380,
    n440,
    n568,
    n550,
    n655
  );


  nand
  g1156
  (
    n1612,
    n527,
    n630,
    n1146,
    n679
  );


  and
  g1157
  (
    n1475,
    n654,
    n680,
    n1103,
    n595
  );


  nor
  g1158
  (
    n1225,
    n431,
    n1165,
    n691,
    n1126
  );


  nand
  g1159
  (
    n1462,
    n395,
    n649,
    n583,
    n481
  );


  and
  g1160
  (
    n1284,
    n340,
    n564,
    n523,
    n463
  );


  xor
  g1161
  (
    n1546,
    n713,
    n500,
    n346,
    n1145
  );


  nor
  g1162
  (
    n1430,
    n1131,
    n501,
    n651,
    n641
  );


  nand
  g1163
  (
    n1469,
    n1170,
    n499,
    n629,
    n1147
  );


  and
  g1164
  (
    n1236,
    n306,
    n509,
    n712,
    n611
  );


  xnor
  g1165
  (
    n1479,
    n360,
    n644,
    n598,
    n630
  );


  nor
  g1166
  (
    n1484,
    n526,
    n1148,
    n380,
    n1121
  );


  and
  g1167
  (
    n1261,
    n609,
    n666,
    n569,
    n659
  );


  xor
  g1168
  (
    n1221,
    n1084,
    n651,
    n459,
    n566
  );


  nor
  g1169
  (
    n1386,
    n1175,
    n486,
    n1120,
    n553
  );


  and
  g1170
  (
    n1521,
    n522,
    n397,
    n578,
    n390
  );


  xor
  g1171
  (
    n1579,
    n644,
    n724,
    n693,
    n530
  );


  xnor
  g1172
  (
    n1533,
    n361,
    n1126,
    n1125,
    n1110
  );


  nor
  g1173
  (
    n1200,
    n430,
    n632,
    n667,
    n564
  );


  nor
  g1174
  (
    n1424,
    n607,
    n425,
    n522,
    n400
  );


  xor
  g1175
  (
    n1381,
    n369,
    n680,
    n665,
    n1107
  );


  or
  g1176
  (
    KeyWire_0_36,
    n617,
    n1090,
    n623,
    n535
  );


  xnor
  g1177
  (
    n1576,
    n528,
    n545,
    n506,
    n422
  );


  xnor
  g1178
  (
    n1405,
    n578,
    n683,
    n625,
    n433
  );


  nand
  g1179
  (
    n1325,
    n525,
    n515,
    n617,
    n701
  );


  xor
  g1180
  (
    KeyWire_0_6,
    n602,
    n649,
    n1111,
    n546
  );


  nor
  g1181
  (
    n1594,
    n396,
    n1186,
    n1161,
    n1136
  );


  xnor
  g1182
  (
    n1529,
    n578,
    n718,
    n653,
    n668
  );


  xnor
  g1183
  (
    n1624,
    n1029,
    n693,
    n457,
    n1171
  );


  and
  g1184
  (
    n1467,
    n1137,
    n728,
    n637,
    n594
  );


  xor
  g1185
  (
    n1361,
    n684,
    n570,
    n1158,
    n647
  );


  xor
  g1186
  (
    n1440,
    n498,
    n1105,
    n460,
    n1136
  );


  xor
  g1187
  (
    n1548,
    n1102,
    n363,
    n461,
    n343
  );


  and
  g1188
  (
    n1447,
    n373,
    n541,
    n1193,
    n596
  );


  xor
  g1189
  (
    n1500,
    n514,
    n538,
    n1112,
    n661
  );


  nand
  g1190
  (
    KeyWire_0_33,
    n626,
    n1113,
    n1156,
    n609
  );


  and
  g1191
  (
    n1297,
    n540,
    n540,
    n1094,
    n491
  );


  or
  g1192
  (
    n1404,
    n669,
    n585,
    n561,
    n640
  );


  xor
  g1193
  (
    n1436,
    n551,
    n1138,
    n335,
    n1127
  );


  and
  g1194
  (
    n1491,
    n485,
    n326,
    n566,
    n1127
  );


  and
  g1195
  (
    n1626,
    n647,
    n1127,
    n648,
    n589
  );


  nor
  g1196
  (
    n1274,
    n579,
    n533,
    n430,
    n322
  );


  nand
  g1197
  (
    n1555,
    n1145,
    n308,
    n419,
    n646
  );


  nand
  g1198
  (
    n1618,
    n603,
    n344,
    n539,
    n1160
  );


  xor
  g1199
  (
    n1566,
    n358,
    n362,
    n502,
    n313
  );


  nor
  g1200
  (
    n1291,
    n451,
    n1192,
    n1181,
    n472
  );


  and
  g1201
  (
    KeyWire_0_5,
    n530,
    n644,
    n513,
    n1093
  );


  and
  g1202
  (
    n1453,
    n622,
    n705,
    n670,
    n460
  );


  xor
  g1203
  (
    KeyWire_0_56,
    n723,
    n1161,
    n578,
    n1092
  );


  nand
  g1204
  (
    n1636,
    n1164,
    n434,
    n1097,
    n1136
  );


  nand
  g1205
  (
    KeyWire_0_49,
    n481,
    n1188,
    n478,
    n495
  );


  nand
  g1206
  (
    n1222,
    n1107,
    n1130,
    n449,
    n532
  );


  xor
  g1207
  (
    n1329,
    n1135,
    n649,
    n714,
    n1097
  );


  nand
  g1208
  (
    n1226,
    n1128,
    n456,
    n703,
    n608
  );


  and
  g1209
  (
    n1206,
    n1189,
    n610,
    n433,
    n728
  );


  nor
  g1210
  (
    n1232,
    n615,
    n630,
    n649,
    n565
  );


  nor
  g1211
  (
    n1316,
    n553,
    n499,
    n331,
    n597
  );


  or
  g1212
  (
    n1330,
    n428,
    n720,
    n1139,
    n608
  );


  nand
  g1213
  (
    n1421,
    n711,
    n548,
    n1189,
    n628
  );


  or
  g1214
  (
    n1408,
    n1028,
    n720,
    n678,
    n725
  );


  xor
  g1215
  (
    n1627,
    n632,
    n379,
    n375,
    n691
  );


  xnor
  g1216
  (
    n1456,
    n1123,
    n432,
    n549,
    n658
  );


  xnor
  g1217
  (
    n1582,
    n531,
    n1135,
    n501,
    n539
  );


  xnor
  g1218
  (
    n1287,
    n626,
    n1086,
    n583,
    n554
  );


  nand
  g1219
  (
    n1270,
    n528,
    n1157,
    n557,
    n478
  );


  nor
  g1220
  (
    n1610,
    n516,
    n1146,
    n595,
    n669
  );


  xnor
  g1221
  (
    n1459,
    n1135,
    n1119,
    n1124,
    n1095
  );


  or
  g1222
  (
    n1292,
    n614,
    n662,
    n414,
    n1154
  );


  or
  g1223
  (
    n1517,
    n1170,
    n650,
    n681,
    n359
  );


  xor
  g1224
  (
    n1464,
    n314,
    n708,
    n704,
    n657
  );


  xnor
  g1225
  (
    n1488,
    n1087,
    n319,
    n489,
    n628
  );


  xnor
  g1226
  (
    n1277,
    n1104,
    n1028,
    n1107,
    n508
  );


  xnor
  g1227
  (
    n1558,
    n418,
    n1156,
    n387,
    n495
  );


  nor
  g1228
  (
    n1543,
    n1083,
    n556,
    n409,
    n507
  );


  xor
  g1229
  (
    n1617,
    n549,
    n612,
    n1144,
    n575
  );


  nand
  g1230
  (
    n1468,
    n431,
    n1184,
    n654,
    n546
  );


  nor
  g1231
  (
    n1472,
    n463,
    n661,
    n682,
    n459
  );


  nand
  g1232
  (
    n1333,
    n1185,
    n576,
    n1118,
    n1188
  );


  or
  g1233
  (
    n1429,
    n332,
    n593,
    n1096,
    n629
  );


  or
  g1234
  (
    n1389,
    n311,
    n675,
    n1156,
    n1153
  );


  and
  g1235
  (
    n1514,
    n524,
    n612,
    n688,
    n510
  );


  xor
  g1236
  (
    n1253,
    n568,
    n707,
    n685,
    n598
  );


  or
  g1237
  (
    n1375,
    n718,
    n601,
    n1093,
    n1182
  );


  nand
  g1238
  (
    n1229,
    n648,
    n542,
    n646,
    n602
  );


  xnor
  g1239
  (
    n1283,
    n613,
    n450,
    n1187,
    n597
  );


  or
  g1240
  (
    n1512,
    n1093,
    n468,
    n504,
    n469
  );


  and
  g1241
  (
    n1476,
    n446,
    n385,
    n389,
    n1097
  );


  nor
  g1242
  (
    n1262,
    n355,
    n636,
    n639,
    n562
  );


  xor
  g1243
  (
    n1390,
    n1122,
    n692,
    n404,
    n1094
  );


  xnor
  g1244
  (
    n1377,
    n422,
    n452,
    n516,
    n1193
  );


  nor
  g1245
  (
    n1527,
    n582,
    n333,
    n585,
    n711
  );


  or
  g1246
  (
    n1557,
    n1120,
    n717,
    n328,
    n329
  );


  xnor
  g1247
  (
    n1489,
    n1145,
    n1144,
    n1142,
    n693
  );


  xor
  g1248
  (
    n1511,
    n650,
    n1177,
    n654,
    n560
  );


  or
  g1249
  (
    n1591,
    n1182,
    n310,
    n1151,
    n706
  );


  nor
  g1250
  (
    n1535,
    n594,
    n1114,
    n1176,
    n715
  );


  xnor
  g1251
  (
    n1526,
    n1154,
    n523,
    n1166,
    n1191
  );


  or
  g1252
  (
    n1347,
    n697,
    n712,
    n620,
    n595
  );


  nor
  g1253
  (
    n1311,
    n547,
    n572,
    n670,
    n592
  );


  nor
  g1254
  (
    n1205,
    n1176,
    n331,
    n574,
    n666
  );


  xnor
  g1255
  (
    n1321,
    n1118,
    n494,
    n624,
    n1115
  );


  nand
  g1256
  (
    n1379,
    n642,
    n502,
    n584,
    n456
  );


  or
  g1257
  (
    n1231,
    n577,
    n1193,
    n621,
    n309
  );


  nand
  g1258
  (
    n1368,
    n1129,
    n585,
    n1112,
    n634
  );


  and
  g1259
  (
    n1528,
    n1150,
    n1087,
    n637,
    n669
  );


  xor
  g1260
  (
    n1412,
    n542,
    n546,
    n462,
    n379
  );


  nor
  g1261
  (
    n1267,
    n671,
    n337,
    n548,
    n1162
  );


  nor
  g1262
  (
    n1493,
    n443,
    n634,
    n1099,
    n703
  );


  or
  g1263
  (
    n1196,
    n349,
    n448,
    n635,
    n442
  );


  xnor
  g1264
  (
    n1595,
    n1158,
    n487,
    n634,
    n382
  );


  nand
  g1265
  (
    n1217,
    n687,
    n1152,
    n371,
    n537
  );


  and
  g1266
  (
    n1400,
    n558,
    n1110,
    n607,
    n727
  );


  xor
  g1267
  (
    n1230,
    n412,
    n1125,
    n1112,
    n686
  );


  nor
  g1268
  (
    n1631,
    n370,
    n678,
    n416,
    n708
  );


  or
  g1269
  (
    n1531,
    n1083,
    n535,
    n582,
    n673
  );


  nand
  g1270
  (
    n1248,
    n1083,
    n333,
    n678,
    n1161
  );


  xor
  g1271
  (
    n1490,
    n381,
    n1169,
    n643,
    n633
  );


  or
  g1272
  (
    n1289,
    n397,
    n643,
    n616,
    n324
  );


  and
  g1273
  (
    n1417,
    n1166,
    n694,
    n708,
    n1147
  );


  or
  g1274
  (
    n1411,
    n590,
    n481,
    n683,
    n1102
  );


  xnor
  g1275
  (
    n1515,
    n615,
    n374,
    n707,
    n599
  );


  nand
  g1276
  (
    n1346,
    n548,
    n700,
    n668,
    n437
  );


  xor
  g1277
  (
    n1265,
    n627,
    n493,
    n581,
    n694
  );


  xor
  g1278
  (
    n1483,
    n536,
    n670,
    n659,
    n671
  );


  nand
  g1279
  (
    n1194,
    n525,
    n698,
    n590,
    n699
  );


  nand
  g1280
  (
    n1499,
    n1193,
    n678,
    n606,
    n629
  );


  nand
  g1281
  (
    n1420,
    n512,
    n601,
    n500,
    n544
  );


  or
  g1282
  (
    n1240,
    n658,
    n1139,
    n1118,
    n312
  );


  nor
  g1283
  (
    n1498,
    n365,
    n1108,
    n1164,
    n372
  );


  nand
  g1284
  (
    n1207,
    n497,
    n621,
    n1088,
    n567
  );


  xnor
  g1285
  (
    n1621,
    n538,
    n1168,
    n1092,
    n1091
  );


  nand
  g1286
  (
    n1245,
    n698,
    n1099,
    n639,
    n577
  );


  and
  g1287
  (
    n1536,
    n502,
    n1103,
    n1152,
    n482
  );


  xnor
  g1288
  (
    n1427,
    n420,
    n1148,
    n606,
    n1104
  );


  xor
  g1289
  (
    n1562,
    n1138,
    n472,
    n684,
    n378
  );


  nor
  g1290
  (
    n1314,
    n672,
    n386,
    n700,
    n532
  );


  xnor
  g1291
  (
    n1278,
    n512,
    n1116,
    n718,
    n1155
  );


  nand
  g1292
  (
    n1598,
    n539,
    n1106,
    n339,
    n1087
  );


  or
  g1293
  (
    n1426,
    n1188,
    n1185,
    n517,
    n1174
  );


  nand
  g1294
  (
    n1423,
    n1166,
    n1181,
    n1105,
    n690
  );


  xnor
  g1295
  (
    n1622,
    n487,
    n522,
    n620,
    n605
  );


  xnor
  g1296
  (
    n1435,
    n1121,
    n468,
    n1140,
    n656
  );


  nor
  g1297
  (
    n1252,
    n537,
    n450,
    n497,
    n611
  );


  and
  g1298
  (
    n1446,
    n1095,
    n528,
    n447,
    n497
  );


  or
  g1299
  (
    n1606,
    n376,
    n435,
    n617,
    n458
  );


  or
  g1300
  (
    n1506,
    n519,
    n645,
    n565,
    n1149
  );


  and
  g1301
  (
    n1603,
    n587,
    n675,
    n464,
    n677
  );


  xor
  g1302
  (
    n1549,
    n520,
    n417,
    n601,
    n663
  );


  nor
  g1303
  (
    n1522,
    n567,
    n471,
    n661,
    n625
  );


  nand
  g1304
  (
    n1286,
    n361,
    n514,
    n1176,
    n348
  );


  or
  g1305
  (
    n1471,
    n496,
    n1156,
    n582,
    n1119
  );


  nand
  g1306
  (
    n1224,
    n554,
    n1134,
    n367,
    n513
  );


  nor
  g1307
  (
    n1353,
    n723,
    n413,
    n475,
    n653
  );


  or
  g1308
  (
    n1369,
    n525,
    n1147,
    n715,
    n543
  );


  nand
  g1309
  (
    n1215,
    n662,
    n320,
    n574,
    n1175
  );


  xor
  g1310
  (
    n1586,
    n1117,
    n543,
    n527,
    n493
  );


  and
  g1311
  (
    n1313,
    n664,
    n338,
    n1139,
    n618
  );


  nor
  g1312
  (
    n1349,
    n1092,
    n624,
    n708,
    n628
  );


  or
  g1313
  (
    n1384,
    n480,
    n571,
    n636,
    n517
  );


  or
  g1314
  (
    n1524,
    n1133,
    n489,
    n408,
    n351
  );


  and
  g1315
  (
    n1233,
    n470,
    n695,
    n551,
    n1176
  );


  xor
  g1316
  (
    n1373,
    n455,
    n321,
    n439,
    n383
  );


  or
  g1317
  (
    n1338,
    n1189,
    n1110,
    n660,
    n694
  );


  or
  g1318
  (
    n1520,
    n659,
    n727,
    n1126,
    n512
  );


  xor
  g1319
  (
    n1320,
    n1094,
    n545,
    n1027,
    n642
  );


  xnor
  g1320
  (
    n1538,
    n1171,
    n686,
    n1147,
    n634
  );


  xor
  g1321
  (
    n1395,
    n381,
    n660,
    n631,
    n715
  );


  xnor
  g1322
  (
    n1388,
    n488,
    n1115,
    n1146,
    n591
  );


  and
  g1323
  (
    n1319,
    n663,
    n562,
    n537,
    n608
  );


  nor
  g1324
  (
    n1448,
    n490,
    n707,
    n1167,
    n545
  );


  and
  g1325
  (
    n1441,
    n321,
    n524,
    n562,
    n1186
  );


  and
  g1326
  (
    n1590,
    n716,
    n676,
    n1160,
    n508
  );


  or
  g1327
  (
    n1281,
    n596,
    n668,
    n1151,
    n676
  );


  nand
  g1328
  (
    n1303,
    n590,
    n1101,
    n1186,
    n551
  );


  or
  g1329
  (
    n1326,
    n1086,
    n511,
    n1164,
    n690
  );


  and
  g1330
  (
    n1492,
    n656,
    n587,
    n689,
    n444
  );


  nor
  g1331
  (
    n1523,
    n552,
    n507,
    n633,
    n581
  );


  or
  g1332
  (
    n1630,
    n688,
    n507,
    n445,
    n665
  );


  and
  g1333
  (
    n1615,
    n584,
    n490,
    n696,
    n511
  );


  and
  g1334
  (
    n1415,
    n549,
    n580,
    n1150,
    n457
  );


  and
  g1335
  (
    n1561,
    n1129,
    n710,
    n1132
  );


  and
  g1336
  (
    n1628,
    n1152,
    n1181,
    n438,
    n1099
  );


  nand
  g1337
  (
    n1596,
    n705,
    n336,
    n672,
    n491
  );


  and
  g1338
  (
    n1366,
    n664,
    n543,
    n636,
    n363
  );


  and
  g1339
  (
    n1431,
    n489,
    n684,
    n488,
    n1188
  );


  nand
  g1340
  (
    n1308,
    n559,
    n1151,
    n538,
    n467
  );


  or
  g1341
  (
    n1547,
    n610,
    n1155,
    n1111,
    n1150
  );


  nor
  g1342
  (
    n1530,
    n346,
    n1085,
    n546,
    n652
  );


  or
  g1343
  (
    n1478,
    n645,
    n327,
    n657,
    n650
  );


  or
  g1344
  (
    n1604,
    n1148,
    n670,
    n622,
    n602
  );


  xor
  g1345
  (
    n1541,
    n721,
    n311,
    n685,
    n336
  );


  nor
  g1346
  (
    n1195,
    n1029,
    n620,
    n492,
    n721
  );


  nor
  g1347
  (
    n1363,
    n335,
    n1168,
    n576,
    n721
  );


  nand
  g1348
  (
    n1495,
    n687,
    n635,
    n591,
    n555
  );


  xnor
  g1349
  (
    n1199,
    n709,
    n1166,
    n443,
    n1182
  );


  xor
  g1350
  (
    n1241,
    n647,
    n366,
    n499,
    n722
  );


  nand
  g1351
  (
    n1213,
    n633,
    n657,
    n1179,
    n526
  );


  and
  g1352
  (
    n1422,
    n607,
    n343,
    n1133,
    n1112
  );


  nor
  g1353
  (
    n1633,
    n521,
    n682,
    n719,
    n1142
  );


  xor
  g1354
  (
    n1409,
    n1113,
    n699,
    n519,
    n1135
  );


  or
  g1355
  (
    n1559,
    n681,
    n1160,
    n386,
    n675
  );


  nand
  g1356
  (
    n1306,
    n1180,
    n552,
    n555,
    n611
  );


  xnor
  g1357
  (
    KeyWire_0_42,
    n680,
    n586,
    n515,
    n1128
  );


  nor
  g1358
  (
    n1545,
    n613,
    n501,
    n410,
    n1123
  );


  nor
  g1359
  (
    n1519,
    n544,
    n1100,
    n683,
    n1111
  );


  nand
  g1360
  (
    n1357,
    n1159,
    n1091,
    n681,
    n1101
  );


  and
  g1361
  (
    n1391,
    n503,
    n691,
    n606,
    n444
  );


  or
  g1362
  (
    n1300,
    n572,
    n702,
    n1187,
    n696
  );


  and
  g1363
  (
    n1525,
    n503,
    n341,
    n408,
    n620
  );


  nor
  g1364
  (
    n1382,
    n672,
    n440,
    n325,
    n517
  );


  and
  g1365
  (
    n1556,
    n585,
    n712,
    n403,
    n679
  );


  and
  g1366
  (
    KeyWire_0_40,
    n446,
    n558,
    n429,
    n509
  );


  and
  g1367
  (
    n1428,
    n1113,
    n552,
    n563,
    n1178
  );


  xor
  g1368
  (
    n1312,
    n517,
    n1149,
    n726,
    n382
  );


  or
  g1369
  (
    n1480,
    n536,
    n502,
    n587,
    n692
  );


  or
  g1370
  (
    n1372,
    n498,
    n454,
    n631,
    n485
  );


  nor
  g1371
  (
    n1370,
    n576,
    n557,
    n1192,
    n483
  );


  nor
  g1372
  (
    n1583,
    n603,
    n1109,
    n375,
    n395
  );


  xnor
  g1373
  (
    n1605,
    n622,
    n514,
    n577,
    n509
  );


  nor
  g1374
  (
    n1564,
    n594,
    n1172,
    n388,
    n610
  );


  or
  g1375
  (
    n1454,
    n477,
    n436,
    n358,
    n313
  );


  nand
  g1376
  (
    n1601,
    n579,
    n534,
    n591,
    n326
  );


  or
  g1377
  (
    n1451,
    n676,
    n725,
    n698,
    n1171
  );


  xnor
  g1378
  (
    n1282,
    n1164,
    n1116,
    n550,
    n1083
  );


  nand
  g1379
  (
    n1563,
    n526,
    n1142,
    n461,
    n690
  );


  and
  g1380
  (
    n1259,
    n709,
    n1132,
    n642,
    n1109
  );


  and
  g1381
  (
    n1641,
    n523,
    n667,
    n532,
    n322
  );


  xnor
  g1382
  (
    n1629,
    n614,
    n614,
    n674,
    n667
  );


  xor
  g1383
  (
    n1219,
    n618,
    n398,
    n586,
    n1134
  );


  and
  g1384
  (
    n1458,
    n1179,
    n713,
    n516,
    n501
  );


  and
  g1385
  (
    n1510,
    n1178,
    n701,
    n407,
    n706
  );


  xor
  g1386
  (
    n1578,
    n1084,
    n494,
    n1175,
    n448
  );


  xor
  g1387
  (
    KeyWire_0_57,
    n309,
    n402,
    n657,
    n694
  );


  or
  g1388
  (
    n1355,
    n1162,
    n581,
    n631,
    n522
  );


  nand
  g1389
  (
    n1279,
    n718,
    n402,
    n492,
    n627
  );


  nor
  g1390
  (
    n1269,
    n1143,
    n334,
    n1162,
    n655
  );


  nor
  g1391
  (
    n1602,
    n589,
    n647,
    n1030,
    n1089
  );


  nand
  g1392
  (
    n1587,
    n1133,
    n1173,
    n415,
    n424
  );


  nor
  g1393
  (
    n1474,
    n480,
    n1169,
    n420,
    n510
  );


  nand
  g1394
  (
    n1477,
    n315,
    n453,
    n687,
    n1096
  );


  and
  g1395
  (
    n1570,
    n324,
    n719,
    n619,
    n1089
  );


  xnor
  g1396
  (
    n1345,
    n1133,
    n307,
    n672,
    n717
  );


  xor
  g1397
  (
    n1296,
    n371,
    n413,
    n563,
    n504
  );


  nand
  g1398
  (
    n1638,
    n1128,
    n583,
    n593,
    n529
  );


  or
  g1399
  (
    n1619,
    n508,
    n474,
    n1098,
    n436
  );


  or
  g1400
  (
    n1371,
    n704,
    n556,
    n1104,
    n690
  );


  or
  g1401
  (
    n1273,
    n721,
    n390,
    n1138,
    n704
  );


  nand
  g1402
  (
    n1227,
    n1109,
    n612,
    n720,
    n609
  );


  xor
  g1403
  (
    n1496,
    n569,
    n1121,
    n689,
    n638
  );


  xor
  g1404
  (
    KeyWire_0_59,
    n445,
    n725,
    n1161,
    n1090
  );


  nand
  g1405
  (
    n1437,
    n664,
    n1191,
    n593,
    n588
  );


  xor
  g1406
  (
    n1365,
    n505,
    n584,
    n354,
    n600
  );


  or
  g1407
  (
    n1509,
    n477,
    n345,
    n1184,
    n421
  );


  nand
  g1408
  (
    n1214,
    n539,
    n705,
    n1168,
    n1167
  );


  xnor
  g1409
  (
    n1336,
    n411,
    n486,
    n582,
    n641
  );


  xnor
  g1410
  (
    n1565,
    n553,
    n682,
    n545,
    n631
  );


  nor
  g1411
  (
    n1254,
    n709,
    n356,
    n704,
    n1170
  );


  and
  g1412
  (
    n1414,
    n1167,
    n1138,
    n1122,
    n464
  );


  and
  g1413
  (
    n1569,
    n1130,
    n352,
    n1108,
    n667
  );


  or
  g1414
  (
    n1290,
    n1117,
    n619,
    n573,
    n604
  );


  and
  g1415
  (
    n1276,
    n615,
    n1125,
    n503,
    n1178
  );


  xor
  g1416
  (
    n1212,
    n373,
    n1100,
    n626,
    n1114
  );


  nor
  g1417
  (
    n1518,
    n701,
    n426,
    n573,
    n466
  );


  xor
  g1418
  (
    n1625,
    n613,
    n727,
    n549,
    n1157
  );


  nand
  g1419
  (
    n1211,
    n716,
    n1154,
    n1172,
    n434
  );


  nand
  g1420
  (
    n1374,
    n427,
    n1084,
    n1131,
    n1141
  );


  or
  g1421
  (
    n1487,
    n469,
    n1091,
    n572,
    n646
  );


  nor
  g1422
  (
    n1637,
    n599,
    n567,
    n536,
    n534
  );


  or
  g1423
  (
    n1255,
    n394,
    n671,
    n540,
    n640
  );


  nand
  g1424
  (
    n1577,
    n607,
    n1177,
    n1149,
    n637
  );


  nand
  g1425
  (
    n1600,
    n625,
    n1085,
    n1084,
    n604
  );


  or
  g1426
  (
    n1358,
    n534,
    n1184,
    n697,
    n633
  );


  or
  g1427
  (
    n1399,
    n570,
    n362,
    n554,
    n1096
  );


  xnor
  g1428
  (
    n1235,
    n1105,
    n571,
    n1140,
    n640
  );


  or
  g1429
  (
    n1457,
    n1082,
    n465,
    n368,
    n345
  );


  or
  g1430
  (
    n1216,
    n406,
    n554,
    n673,
    n1174
  );


  xnor
  g1431
  (
    n1402,
    n1178,
    n711,
    n325,
    n447
  );


  or
  g1432
  (
    n1367,
    n567,
    n317,
    n418,
    n1173
  );


  and
  g1433
  (
    n1532,
    n1159,
    n584,
    n617,
    n1165
  );


  nor
  g1434
  (
    n1589,
    n1165,
    n1170,
    n483,
    n510
  );


  nor
  g1435
  (
    n1251,
    n334,
    n474,
    n494,
    n528
  );


  nor
  g1436
  (
    n1508,
    n383,
    n316,
    n406,
    n1026
  );


  xor
  g1437
  (
    n1202,
    n471,
    n662,
    n559,
    n616
  );


  or
  g1438
  (
    n1197,
    n656,
    n466,
    n1155,
    n693
  );


  or
  g1439
  (
    n1328,
    n425,
    n1141,
    n477,
    n1110
  );


  xor
  g1440
  (
    n1237,
    n389,
    n479,
    n511,
    n421
  );


  nand
  g1441
  (
    n1317,
    n1180,
    n640,
    n509,
    n661
  );


  xor
  g1442
  (
    n1359,
    n409,
    n599,
    n600,
    n656
  );


  or
  g1443
  (
    n1432,
    n726,
    n566,
    n594,
    n475
  );


  nand
  g1444
  (
    n1434,
    n400,
    n1113,
    n329,
    n533
  );


  or
  g1445
  (
    n1271,
    n665,
    n544,
    n641,
    n592
  );


  xor
  g1446
  (
    n1580,
    n699,
    n1130,
    n695,
    n330
  );


  xor
  g1447
  (
    KeyWire_0_47,
    n495,
    n1099,
    n586,
    n1119
  );


  nand
  g1448
  (
    n1481,
    n618,
    n652,
    n1151,
    n467
  );


  and
  g1449
  (
    n1442,
    n1163,
    n458,
    n561,
    n685
  );


  and
  g1450
  (
    n1323,
    n439,
    n591,
    n1082,
    n513
  );


  nor
  g1451
  (
    n1360,
    n1140,
    n714,
    n1190,
    n531
  );


  xor
  g1452
  (
    n1204,
    n676,
    n662,
    n529,
    n665
  );


  nor
  g1453
  (
    KeyWire_0_58,
    n1173,
    n350,
    n518,
    n574
  );


  xnor
  g1454
  (
    n1593,
    n1145,
    n357,
    n1162,
    n511
  );


  nand
  g1455
  (
    n1620,
    n679,
    n1125,
    n604,
    n1180
  );


  xor
  g1456
  (
    n1244,
    n596,
    n392,
    n573,
    n1184
  );


  xnor
  g1457
  (
    n1356,
    n560,
    n490,
    n530,
    n519
  );


  nor
  g1458
  (
    n1243,
    n1089,
    n388,
    n580,
    n710
  );


  xnor
  g1459
  (
    n1567,
    n1153,
    n1093,
    n342,
    n512
  );


  xor
  g1460
  (
    n1198,
    n684,
    n586,
    n653,
    n349
  );


  nand
  g1461
  (
    n1537,
    n479,
    n454,
    n1132,
    n608
  );


  nor
  g1462
  (
    n1310,
    n486,
    n638,
    n484,
    n658
  );


  xnor
  g1463
  (
    n1607,
    n698,
    n1154,
    n527,
    n555
  );


  nand
  g1464
  (
    n1383,
    n416,
    n385,
    n515,
    n376
  );


  nor
  g1465
  (
    n1497,
    n380,
    n600,
    n1155,
    n559
  );


  and
  g1466
  (
    n1568,
    n573,
    n534,
    n1168,
    n487
  );


  nand
  g1467
  (
    n1257,
    n1192,
    n1163,
    n344,
    n587
  );


  xor
  g1468
  (
    n1352,
    n523,
    n547,
    n677,
    n597
  );


  nand
  g1469
  (
    n1343,
    n1124,
    n374,
    n671,
    n1118
  );


  and
  g1470
  (
    n1376,
    n540,
    n1153,
    n1097,
    n1148
  );


  xnor
  g1471
  (
    n1413,
    n711,
    n482,
    n551,
    n544
  );


  nand
  g1472
  (
    n1407,
    n580,
    n724,
    n553,
    n1136
  );


  nand
  g1473
  (
    n1473,
    n568,
    n556,
    n535,
    n1115
  );


  nand
  g1474
  (
    n1299,
    n340,
    n1122,
    n465,
    n537
  );


  xor
  g1475
  (
    n1507,
    n496,
    n500,
    n410,
    n1124
  );


  or
  g1476
  (
    n1298,
    n407,
    n569,
    n1183,
    n638
  );


  xnor
  g1477
  (
    n1307,
    n506,
    n705,
    n548,
    n651
  );


  and
  g1478
  (
    n1588,
    n393,
    n1190,
    n716,
    n515
  );


  and
  g1479
  (
    n1334,
    n428,
    n393,
    n1114,
    n347
  );


  xor
  g1480
  (
    n1632,
    n1092,
    n1117,
    n720,
    n710
  );


  xor
  g1481
  (
    n1396,
    n726,
    n531,
    n571,
    n1165
  );


  and
  g1482
  (
    n1295,
    n629,
    n520,
    n637
  );


  xor
  g1483
  (
    n1246,
    n613,
    n435,
    n1174,
    n526
  );


  nor
  g1484
  (
    n1394,
    n600,
    n1134,
    n714,
    n396
  );


  and
  g1485
  (
    n1450,
    n557,
    n417,
    n318,
    n635
  );


  xnor
  g1486
  (
    n1344,
    n1132,
    n476,
    n563,
    n498
  );


  nand
  g1487
  (
    n1364,
    n521,
    n415,
    n643,
    n648
  );


  nand
  g1488
  (
    n1597,
    n1121,
    n482,
    n1126,
    n673
  );


  and
  g1489
  (
    n1266,
    n655,
    n1185,
    n1103,
    n713
  );


  nand
  g1490
  (
    n1339,
    n571,
    n508,
    n635,
    n524
  );


  nor
  g1491
  (
    n1540,
    n404,
    n438,
    n521,
    n1116
  );


  and
  g1492
  (
    n1410,
    n639,
    n697,
    n538,
    n610
  );


  xor
  g1493
  (
    n1228,
    n1183,
    n378,
    n589,
    n1139
  );


  nand
  g1494
  (
    n1463,
    n1100,
    n619,
    n558,
    n702
  );


  nor
  g1495
  (
    n1392,
    n1158,
    n1158,
    n1111,
    n574
  );


  xor
  g1496
  (
    n1482,
    n518,
    n580,
    n646,
    n1119
  );


  and
  g1497
  (
    n1293,
    n621,
    n1171,
    n498,
    n579
  );


  or
  g1498
  (
    n1550,
    n419,
    n352,
    n1169,
    n570
  );


  or
  g1499
  (
    n1571,
    n504,
    n348,
    n583,
    n1146
  );


  and
  g1500
  (
    n1501,
    n682,
    n424,
    n604,
    n1157
  );


  nand
  g1501
  (
    n1264,
    n616,
    n499,
    n1088,
    n484
  );


  or
  g1502
  (
    n1572,
    n308,
    n441,
    n663,
    n1090
  );


  or
  g1503
  (
    n1616,
    n1108,
    n581,
    n598,
    n330
  );


  or
  g1504
  (
    n1249,
    n683,
    n618,
    n727,
    n368
  );


  xnor
  g1505
  (
    n1552,
    n492,
    n664,
    n725,
    n480
  );


  or
  g1506
  (
    n1513,
    n372,
    n685,
    n728,
    n561
  );


  nand
  g1507
  (
    n1354,
    n449,
    n1186,
    n606,
    n714
  );


  xnor
  g1508
  (
    n1260,
    n575,
    n1150,
    n1187,
    n654
  );


  xor
  g1509
  (
    n1401,
    n565,
    n1177,
    n332,
    n1128
  );


  xnor
  g1510
  (
    n1439,
    n645,
    n689,
    n1143,
    n391
  );


  xnor
  g1511
  (
    n1342,
    n626,
    n615,
    n1142,
    n1143
  );


  nand
  g1512
  (
    n1560,
    n707,
    n513,
    n505,
    n1180
  );


  xnor
  g1513
  (
    n1331,
    n687,
    n1096,
    n1137,
    n524
  );


  and
  g1514
  (
    n1351,
    n455,
    n1100,
    n644,
    n1116
  );


  xnor
  g1515
  (
    n1574,
    n1088,
    n1115,
    n518,
    n492
  );


  nor
  g1516
  (
    n1592,
    n1190,
    n652,
    n603,
    n1173
  );


  xor
  g1517
  (
    n1609,
    n666,
    n706,
    n1105,
    n529
  );


  xnor
  g1518
  (
    n1418,
    n597,
    n1149,
    n642,
    n541
  );


  xor
  g1519
  (
    n1575,
    n310,
    n350,
    n564,
    n1114
  );


  nand
  g1520
  (
    n1272,
    n639,
    n560,
    n1191,
    n645
  );


  xnor
  g1521
  (
    n1452,
    n1102,
    n442,
    n488,
    n1106
  );


  xor
  g1522
  (
    n1250,
    n1174,
    n636,
    n365,
    n533
  );


  xnor
  g1523
  (
    n1438,
    n485,
    n1122,
    n588,
    n314
  );


  xnor
  g1524
  (
    n1614,
    n369,
    n1082,
    n394,
    n353
  );


  or
  g1525
  (
    n1466,
    n595,
    n367,
    n414,
    n312
  );


  nor
  g1526
  (
    n1470,
    n723,
    n441,
    n478,
    n495
  );


  xor
  g1527
  (
    n1335,
    n401,
    n1157,
    n1141,
    n652
  );


  xor
  g1528
  (
    n1210,
    n719,
    n339,
    n697,
    n575
  );


  xnor
  g1529
  (
    n1551,
    n1185,
    n592,
    n1160,
    n1123
  );


  and
  g1530
  (
    n1611,
    n623,
    n1085,
    n1130,
    n423
  );


  or
  g1531
  (
    n1461,
    n622,
    n1027,
    n398,
    n1102
  );


  or
  g1532
  (
    n1635,
    n483,
    n510,
    n653,
    n337
  );


  and
  g1533
  (
    n1416,
    n533,
    n627,
    n560,
    n412
  );


  xnor
  g1534
  (
    n1239,
    n593,
    n342,
    n525,
    n1085
  );


  nor
  g1535
  (
    n1503,
    n521,
    n496,
    n552,
    n1169
  );


  nor
  g1536
  (
    n1218,
    n716,
    n547,
    n550,
    n723
  );


  nor
  g1537
  (
    n1494,
    n423,
    n1134,
    n568,
    n590
  );


  nand
  g1538
  (
    KeyWire_0_53,
    n1190,
    n527,
    n619,
    n703
  );


  or
  g1539
  (
    n1516,
    n366,
    n1098,
    n359,
    n505
  );


  xor
  g1540
  (
    n1425,
    n479,
    n702,
    n491,
    n1087
  );


  nor
  g1541
  (
    n1443,
    n387,
    n1103,
    n630,
    n1095
  );


  xnor
  g1542
  (
    n1304,
    n692,
    n576,
    n518,
    n566
  );


  nor
  g1543
  (
    n1387,
    n403,
    n1129,
    n1090,
    n713
  );


  or
  g1544
  (
    n1581,
    n692,
    n437,
    n726,
    n391
  );


  nor
  g1545
  (
    n1340,
    n1179,
    n592,
    n1120,
    n405
  );


  xnor
  g1546
  (
    n1378,
    n1089,
    n328,
    n689,
    n695
  );


  or
  g1547
  (
    n1327,
    n712,
    n541,
    n605,
    n1153
  );


  xor
  g1548
  (
    n1209,
    n1094,
    n605,
    n532,
    n589
  );


  nor
  g1549
  (
    n1302,
    n506,
    n1191,
    n557,
    n686
  );


  xor
  g1550
  (
    n1398,
    n520,
    n1120,
    n1124,
    n703
  );


  xor
  g1551
  (
    n1486,
    n1106,
    n688,
    n494,
    n1131
  );


  nor
  g1552
  (
    n1406,
    n453,
    n717,
    n628,
    n1091
  );


  or
  g1553
  (
    n1294,
    n505,
    n1144,
    n1181,
    n728
  );


  and
  g1554
  (
    n1201,
    n1107,
    n491,
    n506,
    n1143
  );


  or
  g1555
  (
    n1220,
    n1163,
    n696,
    n621,
    n677
  );


  or
  g1556
  (
    n1502,
    n401,
    n356,
    n1172,
    n354
  );


  nor
  g1557
  (
    n1449,
    n588,
    n570,
    n451,
    n688
  );


  and
  g1558
  (
    n1256,
    n316,
    n519,
    n360,
    n674
  );


  xnor
  g1559
  (
    n1623,
    n632,
    n427,
    n1189,
    n1129
  );


  or
  g1560
  (
    n1460,
    n616,
    n319,
    n719,
    n648
  );


  and
  g1561
  (
    n1318,
    n529,
    n315,
    n691,
    n680
  );


  nand
  g1562
  (
    n1385,
    n699,
    n473,
    n558,
    n470
  );


  and
  g1563
  (
    n1258,
    n677,
    n432,
    n596,
    n497
  );


  or
  g1564
  (
    n1341,
    n575,
    n323,
    n669,
    n1029
  );


  xnor
  g1565
  (
    n1504,
    n476,
    n1123,
    n357,
    n1152
  );


  nand
  g1566
  (
    n1639,
    n577,
    n320,
    n627,
    n473
  );


  xor
  g1567
  (
    n1485,
    n555,
    n601,
    n681,
    n503
  );


  nand
  g1568
  (
    n1403,
    n514,
    n641,
    n569,
    n452
  );


  or
  g1569
  (
    n1534,
    n338,
    n709,
    n1141,
    n1179
  );


  or
  g1570
  (
    n1275,
    n724,
    n572,
    n659,
    n399
  );


  nor
  g1571
  (
    n1640,
    n624,
    n493,
    n1108,
    n663
  );


  nor
  g1572
  (
    n1599,
    n1137,
    n588,
    n500,
    n1117
  );


  nand
  g1573
  (
    n1242,
    n605,
    n1101,
    n722,
    n531
  );


  nor
  g1574
  (
    n1505,
    n660,
    n701,
    n1086,
    n632
  );


  nand
  g1575
  (
    n1288,
    n541,
    n1182,
    n1175,
    n565
  );


  xnor
  g1576
  (
    n1573,
    n651,
    n1159,
    n579,
    n1095
  );


  nand
  g1577
  (
    n1305,
    n1106,
    n542,
    n327,
    n496
  );


  or
  g1578
  (
    n1544,
    n547,
    n543,
    n706,
    n493
  );


  xnor
  g1579
  (
    n1234,
    n724,
    n462,
    n1177,
    n624
  );


  xor
  g1580
  (
    n1322,
    n411,
    n323,
    n1183,
    n384
  );


  xor
  g1581
  (
    n1585,
    n614,
    n1140,
    n700,
    n673
  );


  nand
  g1582
  (
    n1280,
    n399,
    n700,
    n353,
    n696
  );


  or
  g1583
  (
    n1263,
    n1101,
    n668,
    n484,
    n536
  );


  xnor
  g1584
  (
    n1268,
    n426,
    n660,
    n318,
    n702
  );


  xor
  g1585
  (
    n1285,
    n686,
    n1104,
    n307,
    n504
  );


  and
  g1586
  (
    n1553,
    n405,
    n598,
    n1172,
    n1192
  );


  nand
  g1587
  (
    n1315,
    n722,
    n655,
    n1183,
    n715
  );


  and
  g1588
  (
    n1324,
    n364,
    n722,
    n623,
    n1082
  );


  xor
  g1589
  (
    n1337,
    n564,
    n674,
    n638,
    n355
  );


  or
  g1590
  (
    n1362,
    n612,
    n384,
    n317,
    n530
  );


  xnor
  g1591
  (
    n1203,
    n675,
    n1163,
    n1187,
    n1109
  );


  xnor
  g1592
  (
    n1223,
    n341,
    n679,
    n429,
    n563
  );


  or
  g1593
  (
    n1309,
    n1098,
    n1131,
    n602,
    n1159
  );


  nor
  g1594
  (
    n1433,
    n674,
    n516,
    n370,
    n609
  );


  nand
  g1595
  (
    n1393,
    n603,
    n1086,
    n717,
    n542
  );


  or
  g1596
  (
    n1455,
    n507,
    n1167,
    n392,
    n377
  );


  xnor
  g1597
  (
    n1642,
    n729,
    n1194
  );


  nor
  g1598
  (
    n1644,
    n729,
    n730
  );


  nor
  g1599
  (
    n1643,
    n729,
    n1642
  );


  not
  g1600
  (
    n1647,
    n1644
  );


  buf
  g1601
  (
    n1650,
    n730
  );


  buf
  g1602
  (
    n1649,
    n1643
  );


  not
  g1603
  (
    n1651,
    n1644
  );


  buf
  g1604
  (
    n1648,
    n1643
  );


  buf
  g1605
  (
    n1646,
    n1643
  );


  xor
  g1606
  (
    n1645,
    n1643,
    n1644
  );


  not
  g1607
  (
    n1663,
    n731
  );


  buf
  g1608
  (
    n1664,
    n1648
  );


  not
  g1609
  (
    n1660,
    n736
  );


  buf
  g1610
  (
    n1661,
    n738
  );


  and
  g1611
  (
    n1656,
    n734,
    n1649,
    n733,
    n737
  );


  xnor
  g1612
  (
    n1657,
    n737,
    n732,
    n1647
  );


  or
  g1613
  (
    n1652,
    n734,
    n737,
    n1649,
    n1646
  );


  or
  g1614
  (
    n1662,
    n736,
    n738,
    n733,
    n1646
  );


  xor
  g1615
  (
    n1654,
    n734,
    n1648,
    n735,
    n1650
  );


  xnor
  g1616
  (
    n1658,
    n1651,
    n735,
    n1650,
    n737
  );


  nor
  g1617
  (
    n1659,
    n736,
    n1647,
    n732,
    n1645
  );


  xnor
  g1618
  (
    n1655,
    n733,
    n731,
    n1645,
    n735
  );


  or
  g1619
  (
    n1665,
    n735,
    n731,
    n1651
  );


  and
  g1620
  (
    n1653,
    n736,
    n732,
    n734,
    n733
  );


  buf
  g1621
  (
    KeyWire_0_31,
    n738
  );


  buf
  g1622
  (
    n1706,
    n1662
  );


  not
  g1623
  (
    n1695,
    n1656
  );


  buf
  g1624
  (
    n1668,
    n1660
  );


  buf
  g1625
  (
    n1708,
    n1661
  );


  not
  g1626
  (
    n1670,
    n1664
  );


  buf
  g1627
  (
    n1678,
    n950
  );


  buf
  g1628
  (
    n1674,
    n1661
  );


  not
  g1629
  (
    n1721,
    n1655
  );


  buf
  g1630
  (
    n1713,
    n948
  );


  buf
  g1631
  (
    n1675,
    n1661
  );


  not
  g1632
  (
    n1707,
    n949
  );


  buf
  g1633
  (
    n1666,
    n1662
  );


  buf
  g1634
  (
    n1690,
    n1659
  );


  buf
  g1635
  (
    n1683,
    n1665
  );


  buf
  g1636
  (
    KeyWire_0_48,
    n949
  );


  buf
  g1637
  (
    n1720,
    n1652
  );


  buf
  g1638
  (
    n1710,
    n1657
  );


  not
  g1639
  (
    n1703,
    n1663
  );


  not
  g1640
  (
    KeyWire_0_14,
    n1657
  );


  not
  g1641
  (
    n1684,
    n950
  );


  not
  g1642
  (
    n1716,
    n1664
  );


  buf
  g1643
  (
    n1715,
    n1662
  );


  not
  g1644
  (
    n1688,
    n1663
  );


  not
  g1645
  (
    n1687,
    n1658
  );


  not
  g1646
  (
    n1702,
    n1654
  );


  buf
  g1647
  (
    n1700,
    n1659
  );


  buf
  g1648
  (
    n1681,
    n1665
  );


  buf
  g1649
  (
    n1669,
    n1657
  );


  buf
  g1650
  (
    n1712,
    n1656
  );


  buf
  g1651
  (
    n1671,
    n1660
  );


  not
  g1652
  (
    n1667,
    n1659
  );


  buf
  g1653
  (
    n1699,
    n740
  );


  not
  g1654
  (
    n1718,
    n1655
  );


  not
  g1655
  (
    n1697,
    n739
  );


  buf
  g1656
  (
    n1709,
    n1664
  );


  nor
  g1657
  (
    n1701,
    n1658,
    n740
  );


  or
  g1658
  (
    KeyWire_0_19,
    n1663,
    n1654
  );


  and
  g1659
  (
    n1677,
    n948,
    n1655
  );


  nor
  g1660
  (
    n1689,
    n1665,
    n1654
  );


  nand
  g1661
  (
    n1680,
    n1658,
    n1655
  );


  xor
  g1662
  (
    n1694,
    n1665,
    n1658
  );


  or
  g1663
  (
    n1719,
    n1661,
    n947
  );


  nand
  g1664
  (
    KeyWire_0_54,
    n1657,
    n1652
  );


  and
  g1665
  (
    n1711,
    n948,
    n1653
  );


  xor
  g1666
  (
    KeyWire_0_7,
    n947,
    n1659
  );


  nand
  g1667
  (
    n1691,
    n739,
    n1656
  );


  xor
  g1668
  (
    n1714,
    n948,
    n1654
  );


  nand
  g1669
  (
    n1693,
    n1656,
    n949
  );


  nor
  g1670
  (
    n1686,
    n1664,
    n739
  );


  and
  g1671
  (
    n1673,
    n738,
    n1660
  );


  and
  g1672
  (
    n1682,
    n949,
    n1660
  );


  buf
  g1673
  (
    n1672,
    n1653
  );


  and
  g1674
  (
    n1717,
    n1652,
    n1662
  );


  and
  g1675
  (
    n1696,
    n739,
    n1653
  );


  xnor
  g1676
  (
    n1685,
    n1652,
    n1663
  );


  xor
  g1677
  (
    n1869,
    n1505,
    n1353,
    n1430,
    n1370
  );


  or
  g1678
  (
    n1824,
    n1467,
    n1703,
    n1678,
    n1477
  );


  xnor
  g1679
  (
    n1755,
    n1461,
    n1448,
    n1293,
    n1236
  );


  xor
  g1680
  (
    n1866,
    n1711,
    n1315,
    n1460,
    n1701
  );


  xor
  g1681
  (
    n1884,
    n1371,
    n1200,
    n1670,
    n1674
  );


  xnor
  g1682
  (
    n1756,
    n1253,
    n1683,
    n1213,
    n1313
  );


  and
  g1683
  (
    n1753,
    n1226,
    n1451,
    n1294,
    n1385
  );


  and
  g1684
  (
    n1877,
    n1346,
    n1690,
    n1519,
    n1286
  );


  and
  g1685
  (
    n1848,
    n1458,
    n1716,
    n1366,
    n1692
  );


  nand
  g1686
  (
    n1921,
    n1247,
    n1686,
    n1237,
    n1254
  );


  xor
  g1687
  (
    n1777,
    n1506,
    n1429,
    n1680,
    n1426
  );


  or
  g1688
  (
    n1727,
    n1509,
    n1515,
    n1490,
    n1326
  );


  or
  g1689
  (
    n1782,
    n1271,
    n1523,
    n1485
  );


  xnor
  g1690
  (
    n1734,
    n1470,
    n1217,
    n1503,
    n1348
  );


  nand
  g1691
  (
    n1752,
    n1239,
    n1702,
    n1697,
    n1400
  );


  xor
  g1692
  (
    n1807,
    n1333,
    n1517,
    n1298,
    n1205
  );


  and
  g1693
  (
    n1793,
    n1673,
    n1198,
    n1700,
    n1669
  );


  nor
  g1694
  (
    n1934,
    n1404,
    n1295,
    n1264,
    n1402
  );


  and
  g1695
  (
    n1754,
    n1203,
    n1479,
    n1687,
    n1484
  );


  nor
  g1696
  (
    n1938,
    n1272,
    n1335,
    n1443,
    n1332
  );


  xnor
  g1697
  (
    n1894,
    n1718,
    n1256,
    n1462,
    n1678
  );


  nand
  g1698
  (
    n1862,
    n1691,
    n1447,
    n1411,
    n1522
  );


  nand
  g1699
  (
    n1937,
    n1299,
    n1680,
    n1387,
    n1310
  );


  nand
  g1700
  (
    n1745,
    n1427,
    n1475,
    n1412,
    n1311
  );


  xnor
  g1701
  (
    n1853,
    n1423,
    n1481,
    n1671,
    n1716
  );


  nor
  g1702
  (
    n1916,
    n1255,
    n1710,
    n1712,
    n1407
  );


  nor
  g1703
  (
    n1943,
    n1418,
    n1291,
    n1357,
    n1227
  );


  or
  g1704
  (
    n1933,
    n1344,
    n1715,
    n1201,
    n1666
  );


  or
  g1705
  (
    n1942,
    n1452,
    n1509,
    n1683,
    n1669
  );


  nand
  g1706
  (
    n1809,
    n1472,
    n1365,
    n1478,
    n1720
  );


  nand
  g1707
  (
    n1749,
    n1273,
    n1238,
    n1359,
    n1484
  );


  xnor
  g1708
  (
    n1819,
    n1339,
    n1717,
    n1489,
    n1214
  );


  or
  g1709
  (
    n1922,
    n1525,
    n1197,
    n1711,
    n1440
  );


  xor
  g1710
  (
    n1902,
    n1324,
    n1392,
    n1415,
    n1224
  );


  or
  g1711
  (
    n1863,
    n1402,
    n1249,
    n1666,
    n1520
  );


  xnor
  g1712
  (
    n1735,
    n1499,
    n1326,
    n1691,
    n1377
  );


  and
  g1713
  (
    n1914,
    n1690,
    n1711,
    n1353,
    n1677
  );


  xor
  g1714
  (
    KeyWire_0_24,
    n1414,
    n1694,
    n1222,
    n1667
  );


  or
  g1715
  (
    n1932,
    n1398,
    n1268,
    n1475,
    n1306
  );


  xnor
  g1716
  (
    n1931,
    n1498,
    n1380,
    n1696,
    n1464
  );


  xnor
  g1717
  (
    n1817,
    n1403,
    n1410,
    n1279,
    n1708
  );


  xor
  g1718
  (
    n1743,
    n1284,
    n1204,
    n1711,
    n1699
  );


  xor
  g1719
  (
    n1887,
    n1294,
    n1252,
    n1208,
    n1695
  );


  xnor
  g1720
  (
    n1876,
    n1396,
    n1720,
    n1684,
    n1457
  );


  nand
  g1721
  (
    n1904,
    n1677,
    n1310,
    n1527,
    n1218
  );


  nor
  g1722
  (
    n1882,
    n1221,
    n1308,
    n1705,
    n1693
  );


  xor
  g1723
  (
    KeyWire_0_23,
    n1416,
    n1707,
    n1283,
    n1299
  );


  or
  g1724
  (
    n1805,
    n1325,
    n1261,
    n1508,
    n1300
  );


  nor
  g1725
  (
    n1913,
    n1694,
    n1721,
    n1376,
    n1290
  );


  nand
  g1726
  (
    KeyWire_0_32,
    n1258,
    n1674,
    n1447,
    n1325
  );


  or
  g1727
  (
    n1796,
    n1221,
    n1675,
    n1211,
    n1695
  );


  or
  g1728
  (
    n1927,
    n1235,
    n1454,
    n1522,
    n1521
  );


  xnor
  g1729
  (
    n1845,
    n1213,
    n1321,
    n1492,
    n1231
  );


  nand
  g1730
  (
    n1764,
    n1705,
    n1700,
    n1514,
    n1273
  );


  nand
  g1731
  (
    n1738,
    n1673,
    n1363,
    n1362,
    n1230
  );


  nand
  g1732
  (
    n1801,
    n1250,
    n1513,
    n1501,
    n1383
  );


  or
  g1733
  (
    n1945,
    n1199,
    n1276,
    n1708,
    n1435
  );


  nand
  g1734
  (
    n1784,
    n1317,
    n1358,
    n1223,
    n1301
  );


  xnor
  g1735
  (
    n1732,
    n1335,
    n1681,
    n1458,
    n1246
  );


  or
  g1736
  (
    n1830,
    n1361,
    n1279,
    n1338,
    n1263
  );


  nor
  g1737
  (
    n1873,
    n1671,
    n1518,
    n1322,
    n1684
  );


  nor
  g1738
  (
    n1911,
    n1449,
    n1212,
    n1375,
    n1333
  );


  nor
  g1739
  (
    n1790,
    n1319,
    n1237,
    n1376,
    n1682
  );


  and
  g1740
  (
    n1729,
    n1697,
    n1667,
    n1291,
    n1719
  );


  xnor
  g1741
  (
    n1818,
    n1685,
    n1349,
    n1476,
    n1448
  );


  xnor
  g1742
  (
    n1840,
    n1429,
    n1394,
    n1362,
    n1316
  );


  nor
  g1743
  (
    n1905,
    n1503,
    n1679,
    n1491,
    n1410
  );


  or
  g1744
  (
    n1821,
    n1331,
    n1255,
    n1283,
    n1232
  );


  or
  g1745
  (
    n1891,
    n1675,
    n1220,
    n1420,
    n1365
  );


  and
  g1746
  (
    n1815,
    n1378,
    n1479,
    n1707,
    n1675
  );


  nor
  g1747
  (
    n1847,
    n1334,
    n1343,
    n1232,
    n1488
  );


  and
  g1748
  (
    n1772,
    n1701,
    n1305,
    n1312,
    n1244
  );


  xnor
  g1749
  (
    n1747,
    n1405,
    n1721,
    n1323,
    n1417
  );


  or
  g1750
  (
    n1926,
    n1713,
    n1369,
    n1425,
    n1201
  );


  nor
  g1751
  (
    n1810,
    n1225,
    n1524,
    n1323,
    n1709
  );


  xnor
  g1752
  (
    n1901,
    n1674,
    n1408,
    n1340,
    n1409
  );


  nand
  g1753
  (
    n1737,
    n1216,
    n1496,
    n1408,
    n1694
  );


  nor
  g1754
  (
    n1800,
    n1680,
    n1462,
    n1206,
    n1241
  );


  nand
  g1755
  (
    n1778,
    n1205,
    n1337,
    n1468,
    n1307
  );


  or
  g1756
  (
    n1892,
    n1530,
    n1682,
    n1498,
    n1710
  );


  and
  g1757
  (
    n1920,
    n1501,
    n1206,
    n1330,
    n1267
  );


  xor
  g1758
  (
    n1751,
    n1262,
    n1349,
    n1413,
    n1712
  );


  xor
  g1759
  (
    n1872,
    n1710,
    n1435,
    n1293,
    n1217
  );


  nand
  g1760
  (
    n1896,
    n1225,
    n1202,
    n1395,
    n1425
  );


  nor
  g1761
  (
    n1730,
    n1352,
    n1691,
    n1233,
    n1274
  );


  nand
  g1762
  (
    n1803,
    n1668,
    n1342,
    n1382,
    n1302
  );


  or
  g1763
  (
    n1785,
    n1690,
    n1396,
    n1679,
    n1714
  );


  xnor
  g1764
  (
    n1919,
    n1504,
    n1336,
    n1392,
    n1407
  );


  or
  g1765
  (
    n1762,
    n1451,
    n1719,
    n1687,
    n1266
  );


  xnor
  g1766
  (
    n1893,
    n1687,
    n1383,
    n1247,
    n1228
  );


  nand
  g1767
  (
    n1774,
    n1494,
    n1379,
    n1249,
    n1469
  );


  nand
  g1768
  (
    n1795,
    n1271,
    n1346,
    n1388,
    n1463
  );


  xor
  g1769
  (
    n1910,
    n1420,
    n1292,
    n1252,
    n1257
  );


  xor
  g1770
  (
    n1741,
    n1482,
    n1713,
    n1441,
    n1275
  );


  nand
  g1771
  (
    n1832,
    n1384,
    n1197,
    n1678,
    n1214
  );


  xor
  g1772
  (
    n1844,
    n1690,
    n1318,
    n1263,
    n1708
  );


  nand
  g1773
  (
    n1890,
    n1430,
    n1385,
    n1389,
    n1443
  );


  xor
  g1774
  (
    n1728,
    n1477,
    n1324,
    n1703,
    n1391
  );


  nor
  g1775
  (
    n1874,
    n1715,
    n1320,
    n1210,
    n1282
  );


  nand
  g1776
  (
    n1804,
    n1703,
    n1287,
    n1675,
    n1270
  );


  or
  g1777
  (
    n1771,
    n1388,
    n1697,
    n1288,
    n1670
  );


  xnor
  g1778
  (
    n1744,
    n1504,
    n1269,
    n1245,
    n1207
  );


  or
  g1779
  (
    n1767,
    n1523,
    n1281,
    n1461,
    n1386
  );


  xnor
  g1780
  (
    n1842,
    n1517,
    n1219,
    n1666,
    n1489
  );


  or
  g1781
  (
    n1806,
    n1234,
    n1195,
    n1478,
    n1483
  );


  xnor
  g1782
  (
    KeyWire_0_4,
    n1681,
    n1238,
    n1227,
    n1280
  );


  or
  g1783
  (
    n1835,
    n1713,
    n1423,
    n1696,
    n1413
  );


  nand
  g1784
  (
    n1731,
    n1712,
    n1487,
    n1695,
    n1672
  );


  nor
  g1785
  (
    KeyWire_0_45,
    n1222,
    n1709,
    n1700,
    n1267
  );


  and
  g1786
  (
    n1859,
    n1719,
    n1511,
    n1455,
    n1260
  );


  nand
  g1787
  (
    n1822,
    n1715,
    n1199,
    n1309,
    n1520
  );


  nand
  g1788
  (
    n1812,
    n1240,
    n1328,
    n1386,
    n1695
  );


  and
  g1789
  (
    n1739,
    n1356,
    n1209,
    n1387,
    n1304
  );


  or
  g1790
  (
    n1829,
    n1702,
    n1720,
    n1196,
    n1474
  );


  or
  g1791
  (
    n1907,
    n1524,
    n1360,
    n1699,
    n1331
  );


  or
  g1792
  (
    n1870,
    n1516,
    n1529,
    n1671,
    n1287
  );


  and
  g1793
  (
    n1799,
    n1688,
    n1668,
    n1431,
    n1313
  );


  or
  g1794
  (
    n1879,
    n1345,
    n1709,
    n1433,
    n1401
  );


  and
  g1795
  (
    n1928,
    n1704,
    n1216,
    n1717,
    n1518
  );


  nor
  g1796
  (
    n1871,
    n1218,
    n1681,
    n1483
  );


  nor
  g1797
  (
    n1758,
    n1466,
    n1277,
    n1317,
    n1521
  );


  nor
  g1798
  (
    n1776,
    n1364,
    n1278,
    n1228,
    n1511
  );


  and
  g1799
  (
    n1827,
    n1231,
    n1482,
    n1262,
    n1699
  );


  xor
  g1800
  (
    n1912,
    n1394,
    n1463,
    n1683,
    n1328
  );


  or
  g1801
  (
    n1820,
    n1209,
    n1716,
    n1366,
    n1693
  );


  xnor
  g1802
  (
    n1779,
    n1347,
    n1710,
    n1230,
    n1411
  );


  or
  g1803
  (
    n1857,
    n1258,
    n1241,
    n1330,
    n1676
  );


  and
  g1804
  (
    n1823,
    n1371,
    n1688,
    n1424,
    n1373
  );


  or
  g1805
  (
    n1723,
    n1373,
    n1672,
    n1685,
    n1698
  );


  or
  g1806
  (
    n1944,
    n1459,
    n1309,
    n1400,
    n1372
  );


  xnor
  g1807
  (
    n1722,
    n1297,
    n1264,
    n1680,
    n1502
  );


  and
  g1808
  (
    n1761,
    n1314,
    n1714,
    n1246,
    n1704
  );


  and
  g1809
  (
    n1833,
    n1686,
    n1245,
    n1421,
    n1490
  );


  xnor
  g1810
  (
    KeyWire_0_29,
    n1314,
    n1256,
    n1381,
    n1673
  );


  and
  g1811
  (
    n1897,
    n1355,
    n1699,
    n1714,
    n1307
  );


  nand
  g1812
  (
    n1787,
    n1244,
    n1397,
    n1459,
    n1677
  );


  nor
  g1813
  (
    n1881,
    n1514,
    n1696,
    n1669,
    n1480
  );


  or
  g1814
  (
    n1856,
    n1334,
    n1526,
    n1250,
    n1248
  );


  and
  g1815
  (
    n1935,
    n1322,
    n1329,
    n1220,
    n1452
  );


  or
  g1816
  (
    n1808,
    n1525,
    n1370,
    n1679
  );


  or
  g1817
  (
    n1781,
    n1401,
    n1465,
    n1687,
    n1685
  );


  xor
  g1818
  (
    n1865,
    n1327,
    n1670,
    n1254,
    n1442
  );


  and
  g1819
  (
    n1736,
    n1445,
    n1682,
    n1471,
    n1357
  );


  and
  g1820
  (
    n1825,
    n1395,
    n1487,
    n1194,
    n1364
  );


  or
  g1821
  (
    n1861,
    n1686,
    n1721,
    n1708,
    n1409
  );


  or
  g1822
  (
    n1794,
    n1692,
    n1706,
    n1721,
    n1368
  );


  and
  g1823
  (
    n1826,
    n1278,
    n1354,
    n1456,
    n1368
  );


  nand
  g1824
  (
    n1757,
    n1689,
    n1464,
    n1688,
    n1332
  );


  or
  g1825
  (
    n1852,
    n1450,
    n1393,
    n1242,
    n1471
  );


  or
  g1826
  (
    n1918,
    n1265,
    n1692,
    n1374,
    n1486
  );


  nand
  g1827
  (
    n1834,
    n1689,
    n1704,
    n1718,
    n1340
  );


  or
  g1828
  (
    n1929,
    n1426,
    n1693,
    n1207,
    n1422
  );


  or
  g1829
  (
    n1750,
    n1363,
    n1428,
    n1678,
    n1285
  );


  nand
  g1830
  (
    n1791,
    n1688,
    n1236,
    n1285,
    n1269
  );


  or
  g1831
  (
    n1868,
    n1441,
    n1251,
    n1668,
    n1442
  );


  or
  g1832
  (
    n1802,
    n1507,
    n1350,
    n1212,
    n1701
  );


  xnor
  g1833
  (
    n1936,
    n1202,
    n1677,
    n1500,
    n1684
  );


  and
  g1834
  (
    n1792,
    n1434,
    n1399,
    n1277,
    n1203
  );


  nand
  g1835
  (
    n1930,
    n1223,
    n1476,
    n1359,
    n1516
  );


  nand
  g1836
  (
    n1814,
    n1488,
    n1327,
    n1268,
    n1718
  );


  xor
  g1837
  (
    n1813,
    n1397,
    n1280,
    n1347,
    n1248
  );


  nor
  g1838
  (
    n1828,
    n1713,
    n1444,
    n1367,
    n1235
  );


  xnor
  g1839
  (
    n1766,
    n1446,
    n1412,
    n1390,
    n1707
  );


  and
  g1840
  (
    n1850,
    n1515,
    n1261,
    n1449,
    n1434
  );


  xnor
  g1841
  (
    n1726,
    n1684,
    n1527,
    n1281,
    n1378
  );


  xnor
  g1842
  (
    n1775,
    n1303,
    n1705,
    n1706
  );


  xnor
  g1843
  (
    n1760,
    n1682,
    n1224,
    n1703,
    n1436
  );


  nand
  g1844
  (
    n1769,
    n1427,
    n1469,
    n1276,
    n1473
  );


  xnor
  g1845
  (
    n1858,
    n1676,
    n1374,
    n1667,
    n1508
  );


  nor
  g1846
  (
    n1789,
    n1671,
    n1337,
    n1338,
    n1305
  );


  or
  g1847
  (
    n1746,
    n1672,
    n1432,
    n1265,
    n1718
  );


  xnor
  g1848
  (
    n1878,
    n1272,
    n1382,
    n1714,
    n1303
  );


  xor
  g1849
  (
    n1940,
    n1361,
    n1473,
    n1666,
    n1715
  );


  xnor
  g1850
  (
    n1788,
    n1355,
    n1507,
    n1226,
    n1505
  );


  and
  g1851
  (
    n1851,
    n1502,
    n1513,
    n1494,
    n1219
  );


  nor
  g1852
  (
    n1880,
    n1351,
    n1510,
    n1512,
    n1290
  );


  and
  g1853
  (
    n1909,
    n1438,
    n1707,
    n1360,
    n1210
  );


  nor
  g1854
  (
    n1843,
    n1312,
    n1422,
    n1344,
    n1297
  );


  nand
  g1855
  (
    n1816,
    n1686,
    n1369,
    n1416,
    n1234
  );


  and
  g1856
  (
    n1923,
    n1289,
    n1381,
    n1419,
    n1698
  );


  nand
  g1857
  (
    n1875,
    n1345,
    n1233,
    n1251,
    n1295
  );


  and
  g1858
  (
    n1831,
    n1292,
    n1689,
    n1698,
    n1493
  );


  and
  g1859
  (
    n1860,
    n1491,
    n1379,
    n1445,
    n1384
  );


  xnor
  g1860
  (
    n1765,
    n1354,
    n1242,
    n1717,
    n1352
  );


  nor
  g1861
  (
    n1786,
    n1480,
    n1367,
    n1301,
    n1428
  );


  nand
  g1862
  (
    n1724,
    n1495,
    n1404,
    n1437,
    n1351
  );


  nor
  g1863
  (
    n1841,
    n1702,
    n1691,
    n1257,
    n1418
  );


  and
  g1864
  (
    n1759,
    n1296,
    n1393,
    n1302,
    n1284
  );


  and
  g1865
  (
    n1903,
    n1709,
    n1319,
    n1424,
    n1229
  );


  or
  g1866
  (
    n1886,
    n1700,
    n1467,
    n1372,
    n1380
  );


  or
  g1867
  (
    n1838,
    n1415,
    n1685,
    n1497,
    n1229
  );


  xor
  g1868
  (
    n1925,
    n1282,
    n1667,
    n1315,
    n1274
  );


  nor
  g1869
  (
    n1908,
    n1198,
    n1674,
    n1286,
    n1196
  );


  xor
  g1870
  (
    n1895,
    n1453,
    n1243,
    n1239,
    n1676
  );


  or
  g1871
  (
    n1883,
    n1253,
    n1712,
    n1270,
    n1719
  );


  and
  g1872
  (
    n1742,
    n1195,
    n1474,
    n1702,
    n1243
  );


  xor
  g1873
  (
    n1939,
    n1720,
    n1529,
    n1500,
    n1439
  );


  xnor
  g1874
  (
    n1740,
    n1512,
    n1468,
    n1215,
    n1266
  );


  and
  g1875
  (
    n1837,
    n1336,
    n1438,
    n1358,
    n1298
  );


  xnor
  g1876
  (
    n1725,
    n1389,
    n1275,
    n1470,
    n1704
  );


  or
  g1877
  (
    n1768,
    n1453,
    n1436,
    n1676,
    n1454
  );


  or
  g1878
  (
    n1900,
    n1433,
    n1450,
    n1697,
    n1444
  );


  nand
  g1879
  (
    n1888,
    n1701,
    n1446,
    n1432,
    n1495
  );


  and
  g1880
  (
    n1846,
    n1717,
    n1406,
    n1403,
    n1670
  );


  nor
  g1881
  (
    n1811,
    n1304,
    n1350,
    n1716,
    n1672
  );


  and
  g1882
  (
    n1855,
    n1497,
    n1506,
    n1668,
    n1419
  );


  nor
  g1883
  (
    n1889,
    n1320,
    n1405,
    n1316,
    n1492
  );


  or
  g1884
  (
    n1780,
    n1431,
    n1694,
    n1215,
    n1342
  );


  xor
  g1885
  (
    n1899,
    n1705,
    n1200,
    n1706,
    n1692
  );


  xnor
  g1886
  (
    n1915,
    n1375,
    n1204,
    n1414,
    n1499
  );


  nor
  g1887
  (
    n1783,
    n1465,
    n1683,
    n1437,
    n1208
  );


  nor
  g1888
  (
    n1839,
    n1439,
    n1339,
    n1308,
    n1460
  );


  xnor
  g1889
  (
    n1773,
    n1288,
    n1696,
    n1417,
    n1348
  );


  nand
  g1890
  (
    n1770,
    n1456,
    n1457,
    n1289,
    n1698
  );


  and
  g1891
  (
    n1867,
    n1496,
    n1486,
    n1669,
    n1329
  );


  or
  g1892
  (
    n1898,
    n1455,
    n1528,
    n1240,
    n1391
  );


  nor
  g1893
  (
    n1763,
    n1211,
    n1472,
    n1406,
    n1341
  );


  and
  g1894
  (
    n1906,
    n1440,
    n1318,
    n1399,
    n1311
  );


  nor
  g1895
  (
    n1885,
    n1356,
    n1673,
    n1259,
    n1321
  );


  nor
  g1896
  (
    n1941,
    n1300,
    n1466,
    n1306,
    n1526
  );


  or
  g1897
  (
    n1748,
    n1343,
    n1296,
    n1260,
    n1481
  );


  nor
  g1898
  (
    n1849,
    n1519,
    n1341,
    n1259,
    n1377
  );


  xnor
  g1899
  (
    n1797,
    n1390,
    n1528,
    n1493,
    n1421
  );


  or
  g1900
  (
    n1854,
    n1693,
    n1689,
    n1510,
    n1398
  );


  xor
  g1901
  (
    n2077,
    n743,
    n866,
    n1936,
    n1843
  );


  and
  g1902
  (
    n2159,
    n744,
    n895,
    n1544,
    n1883
  );


  nand
  g1903
  (
    KeyWire_0_12,
    n1875,
    n1585,
    n766,
    n922
  );


  xor
  g1904
  (
    n2243,
    n1597,
    n1766,
    n1885,
    n1769
  );


  or
  g1905
  (
    n1974,
    n819,
    n1614,
    n1926,
    n1930
  );


  or
  g1906
  (
    n2078,
    n1820,
    n813,
    n784,
    n1726
  );


  xnor
  g1907
  (
    n2124,
    n1736,
    n892,
    n1551,
    n820
  );


  nor
  g1908
  (
    n1961,
    n791,
    n753,
    n1933,
    n1547
  );


  nor
  g1909
  (
    n2001,
    n1909,
    n808,
    n1908,
    n1934
  );


  nand
  g1910
  (
    n2149,
    n1930,
    n877,
    n1887,
    n774
  );


  nor
  g1911
  (
    n2235,
    n1912,
    n1741,
    n1586,
    n1605
  );


  nand
  g1912
  (
    n2215,
    n853,
    n781,
    n907,
    n1586
  );


  nand
  g1913
  (
    n2041,
    n875,
    n1866,
    n1589,
    n1582
  );


  xnor
  g1914
  (
    n2157,
    n751,
    n910,
    n1913,
    n877
  );


  nor
  g1915
  (
    n2282,
    n1621,
    n794,
    n782,
    n888
  );


  xnor
  g1916
  (
    n2017,
    n1830,
    n741,
    n921,
    n1557
  );


  nor
  g1917
  (
    n2137,
    n812,
    n1850,
    n867,
    n852
  );


  nor
  g1918
  (
    n2161,
    n908,
    n1862,
    n817,
    n1608
  );


  and
  g1919
  (
    n2257,
    n1943,
    n1560,
    n863,
    n1740
  );


  and
  g1920
  (
    n2117,
    n770,
    n1562,
    n846,
    n915
  );


  and
  g1921
  (
    n2092,
    n1878,
    n1901,
    n900,
    n889
  );


  or
  g1922
  (
    n2125,
    n817,
    n1724,
    n1592,
    n783
  );


  xor
  g1923
  (
    n2059,
    n1536,
    n744,
    n899,
    n752
  );


  or
  g1924
  (
    n1975,
    n754,
    n749,
    n862,
    n1542
  );


  nor
  g1925
  (
    n2290,
    n1536,
    n1945,
    n807,
    n848
  );


  nand
  g1926
  (
    n2070,
    n1728,
    n872,
    n800,
    n754
  );


  nor
  g1927
  (
    n1956,
    n920,
    n1753,
    n800,
    n888
  );


  and
  g1928
  (
    n2134,
    n795,
    n769,
    n747,
    n1912
  );


  nand
  g1929
  (
    n1976,
    n823,
    n1895,
    n841,
    n1605
  );


  and
  g1930
  (
    n2160,
    n1577,
    n875,
    n1612,
    n916
  );


  and
  g1931
  (
    n2111,
    n915,
    n824,
    n762,
    n1792
  );


  or
  g1932
  (
    n2042,
    n846,
    n1593,
    n1576,
    n1778
  );


  nand
  g1933
  (
    n2130,
    n864,
    n1794,
    n904,
    n1833
  );


  nor
  g1934
  (
    n2270,
    n1797,
    n756,
    n837,
    n1844
  );


  nor
  g1935
  (
    n2007,
    n844,
    n872,
    n868,
    n1600
  );


  nor
  g1936
  (
    n2062,
    n862,
    n1889,
    n1798,
    n1845
  );


  and
  g1937
  (
    n2028,
    n1740,
    n911,
    n1801,
    n1874
  );


  and
  g1938
  (
    n2139,
    n1903,
    n898,
    n904,
    n1623
  );


  nand
  g1939
  (
    n1977,
    n1825,
    n749,
    n875,
    n870
  );


  and
  g1940
  (
    n1972,
    n1921,
    n1756,
    n1749,
    n1869
  );


  xor
  g1941
  (
    n1953,
    n1839,
    n757,
    n1817,
    n1750
  );


  and
  g1942
  (
    n2067,
    n833,
    n1739,
    n838,
    n879
  );


  xor
  g1943
  (
    n2133,
    n1544,
    n760,
    n1823,
    n878
  );


  nor
  g1944
  (
    n2024,
    n1915,
    n881,
    n772,
    n1790
  );


  nand
  g1945
  (
    n2250,
    n815,
    n1754,
    n823,
    n1766
  );


  and
  g1946
  (
    n1990,
    n883,
    n1942,
    n847,
    n803
  );


  nand
  g1947
  (
    n2231,
    n806,
    n883,
    n775,
    n1613
  );


  or
  g1948
  (
    n2104,
    n787,
    n760,
    n1770,
    n1747
  );


  nand
  g1949
  (
    n2262,
    n881,
    n843,
    n923,
    n1602
  );


  xor
  g1950
  (
    n2255,
    n919,
    n1783,
    n1599,
    n898
  );


  nand
  g1951
  (
    n2198,
    n755,
    n816,
    n799,
    n1920
  );


  xnor
  g1952
  (
    n2277,
    n1816,
    n855,
    n890,
    n869
  );


  nor
  g1953
  (
    n2034,
    n780,
    n772,
    n1537,
    n774
  );


  xor
  g1954
  (
    n1991,
    n1893,
    n1589,
    n837,
    n1842
  );


  xor
  g1955
  (
    n2239,
    n786,
    n741,
    n1848,
    n828
  );


  nor
  g1956
  (
    n2109,
    n1533,
    n856,
    n825,
    n1762
  );


  nand
  g1957
  (
    n2146,
    n751,
    n1836,
    n1577,
    n820
  );


  and
  g1958
  (
    n2002,
    n1920,
    n1615,
    n748,
    n744
  );


  or
  g1959
  (
    n1963,
    n1882,
    n1768,
    n783,
    n873
  );


  or
  g1960
  (
    n2174,
    n1541,
    n835,
    n1889,
    n747
  );


  xor
  g1961
  (
    n2088,
    n1780,
    n884,
    n1558
  );


  and
  g1962
  (
    n2266,
    n822,
    n794,
    n1863,
    n782
  );


  and
  g1963
  (
    n2199,
    n1563,
    n917,
    n1798,
    n1590
  );


  xor
  g1964
  (
    n1964,
    n831,
    n1917,
    n905,
    n906
  );


  or
  g1965
  (
    n2195,
    n1869,
    n769,
    n1781,
    n1550
  );


  nand
  g1966
  (
    n2275,
    n757,
    n1729,
    n853,
    n1880
  );


  or
  g1967
  (
    n2165,
    n1610,
    n1744,
    n1893,
    n1859
  );


  xnor
  g1968
  (
    n2208,
    n778,
    n1545,
    n1738,
    n1799
  );


  or
  g1969
  (
    n2203,
    n913,
    n870,
    n1574,
    n920
  );


  xor
  g1970
  (
    n2144,
    n766,
    n906,
    n1882,
    n851
  );


  xnor
  g1971
  (
    n2248,
    n878,
    n1885,
    n806,
    n748
  );


  nand
  g1972
  (
    n2283,
    n901,
    n1779,
    n858,
    n771
  );


  xor
  g1973
  (
    n2219,
    n1813,
    n1905,
    n1846,
    n1726
  );


  nor
  g1974
  (
    n2022,
    n809,
    n902,
    n1552,
    n1918
  );


  or
  g1975
  (
    n2057,
    n1732,
    n912,
    n1932,
    n914
  );


  or
  g1976
  (
    n1994,
    n1813,
    n814,
    n1823,
    n1572
  );


  nor
  g1977
  (
    n2206,
    n758,
    n747,
    n1853,
    n831
  );


  nand
  g1978
  (
    n1989,
    n1620,
    n1533,
    n833,
    n791
  );


  or
  g1979
  (
    n1960,
    n810,
    n825,
    n771,
    n767
  );


  nor
  g1980
  (
    n2014,
    n758,
    n1617,
    n845,
    n1734
  );


  nand
  g1981
  (
    n2269,
    n740,
    n1750,
    n1561,
    n1731
  );


  or
  g1982
  (
    n1987,
    n1548,
    n755,
    n858,
    n786
  );


  nand
  g1983
  (
    n2260,
    n1864,
    n853,
    n1830,
    n1600
  );


  xor
  g1984
  (
    n2240,
    n900,
    n1617,
    n1723,
    n914
  );


  xor
  g1985
  (
    n2251,
    n804,
    n885,
    n857,
    n746
  );


  nor
  g1986
  (
    n2006,
    n850,
    n1582,
    n788,
    n832
  );


  nand
  g1987
  (
    n2263,
    n1770,
    n1847,
    n797,
    n908
  );


  xor
  g1988
  (
    n2136,
    n792,
    n1795,
    n886,
    n862
  );


  xor
  g1989
  (
    n2214,
    n1767,
    n849,
    n776,
    n1596
  );


  nand
  g1990
  (
    n2020,
    n790,
    n879,
    n893,
    n832
  );


  and
  g1991
  (
    n2032,
    n1923,
    n1916,
    n1572,
    n1551
  );


  xor
  g1992
  (
    KeyWire_0_55,
    n1738,
    n1865,
    n1858,
    n909
  );


  or
  g1993
  (
    n2035,
    n1879,
    n1924,
    n889,
    n1538
  );


  and
  g1994
  (
    n2181,
    n779,
    n1918,
    n836,
    n1751
  );


  and
  g1995
  (
    n2221,
    n784,
    n1532,
    n1744,
    n1768
  );


  xor
  g1996
  (
    n2210,
    n859,
    n1809,
    n811,
    n801
  );


  nor
  g1997
  (
    n2039,
    n1587,
    n1545,
    n761,
    n919
  );


  or
  g1998
  (
    n2220,
    n1769,
    n923,
    n1877,
    n1802
  );


  and
  g1999
  (
    n2018,
    n762,
    n763,
    n798,
    n760
  );


  and
  g2000
  (
    n2000,
    n847,
    n1794,
    n1530,
    n1616
  );


  nor
  g2001
  (
    n1978,
    n840,
    n904,
    n1786,
    n1821
  );


  nor
  g2002
  (
    n2213,
    n810,
    n1896,
    n892,
    n798
  );


  nand
  g2003
  (
    n2202,
    n886,
    n815,
    n1914,
    n1888
  );


  nand
  g2004
  (
    n2033,
    n1575,
    n1917,
    n803,
    n780
  );


  or
  g2005
  (
    n2253,
    n791,
    n797,
    n1759,
    n1902
  );


  or
  g2006
  (
    n2147,
    n805,
    n920,
    n1729,
    n1868
  );


  nand
  g2007
  (
    n2140,
    n1618,
    n887,
    n1776,
    n1570
  );


  nand
  g2008
  (
    n1970,
    n1598,
    n1611,
    n755,
    n861
  );


  nand
  g2009
  (
    n1997,
    n758,
    n909,
    n776,
    n767
  );


  or
  g2010
  (
    n2279,
    n918,
    n1807,
    n783,
    n830
  );


  xor
  g2011
  (
    n2172,
    n841,
    n911,
    n1585,
    n1827
  );


  nor
  g2012
  (
    n2040,
    n924,
    n1584,
    n776,
    n1751
  );


  xor
  g2013
  (
    n2212,
    n808,
    n1833,
    n822,
    n1540
  );


  xor
  g2014
  (
    n2112,
    n1815,
    n1852,
    n850,
    n801
  );


  and
  g2015
  (
    n1955,
    n1847,
    n1787,
    n852,
    n779
  );


  nor
  g2016
  (
    n2191,
    n759,
    n1797,
    n830,
    n1782
  );


  xor
  g2017
  (
    n1966,
    n797,
    n833,
    n754,
    n1940
  );


  nand
  g2018
  (
    n2064,
    n1932,
    n917,
    n773,
    n841
  );


  xnor
  g2019
  (
    n2110,
    n1836,
    n824,
    n1607,
    n1808
  );


  nand
  g2020
  (
    n2065,
    n835,
    n1939,
    n762,
    n1725
  );


  or
  g2021
  (
    n2265,
    n892,
    n824,
    n760,
    n786
  );


  nand
  g2022
  (
    n2060,
    n802,
    n857,
    n1848,
    n1878
  );


  xor
  g2023
  (
    n2115,
    n1810,
    n761,
    n874,
    n1743
  );


  xor
  g2024
  (
    n2089,
    n918,
    n1565,
    n1929,
    n1619
  );


  nor
  g2025
  (
    n1951,
    n1834,
    n912,
    n1831,
    n893
  );


  and
  g2026
  (
    n2222,
    n740,
    n890,
    n822,
    n1552
  );


  and
  g2027
  (
    n2171,
    n1888,
    n1565,
    n859,
    n1887
  );


  or
  g2028
  (
    n2236,
    n1567,
    n865,
    n792,
    n1737
  );


  xnor
  g2029
  (
    n2047,
    n863,
    n1602,
    n1825,
    n1730
  );


  and
  g2030
  (
    n2186,
    n826,
    n773,
    n818,
    n1872
  );


  nor
  g2031
  (
    n2087,
    n795,
    n1614,
    n861,
    n1884
  );


  nand
  g2032
  (
    n2197,
    n770,
    n821,
    n843,
    n757
  );


  nand
  g2033
  (
    n2167,
    n1616,
    n1627,
    n801,
    n887
  );


  nor
  g2034
  (
    n2106,
    n1580,
    n1904,
    n818,
    n855
  );


  and
  g2035
  (
    n1949,
    n832,
    n777,
    n834,
    n752
  );


  xor
  g2036
  (
    n2114,
    n771,
    n767,
    n1790,
    n754
  );


  and
  g2037
  (
    n2247,
    n1553,
    n1782,
    n766,
    n1804
  );


  xnor
  g2038
  (
    n2019,
    n1838,
    n751,
    n898,
    n883
  );


  xor
  g2039
  (
    n2141,
    n822,
    n889,
    n1784,
    n1774
  );


  nor
  g2040
  (
    n2154,
    n1815,
    n1806,
    n1743,
    n1626
  );


  and
  g2041
  (
    n2216,
    n769,
    n842,
    n1849,
    n1880
  );


  xnor
  g2042
  (
    n2101,
    n1858,
    n749,
    n829,
    n899
  );


  or
  g2043
  (
    n1995,
    n823,
    n849,
    n782,
    n799
  );


  xnor
  g2044
  (
    n1983,
    n804,
    n1931,
    n1570,
    n1554
  );


  nand
  g2045
  (
    n2152,
    n1856,
    n845,
    n1754,
    n813
  );


  nor
  g2046
  (
    n2090,
    n905,
    n1891,
    n781,
    n1560
  );


  nand
  g2047
  (
    n1959,
    n874,
    n1745,
    n1550,
    n1876
  );


  xor
  g2048
  (
    n2038,
    n859,
    n1890,
    n1580,
    n1826
  );


  xnor
  g2049
  (
    n2280,
    n787,
    n781,
    n819,
    n1911
  );


  nand
  g2050
  (
    n2268,
    n916,
    n911,
    n838,
    n819
  );


  xnor
  g2051
  (
    n2234,
    n1817,
    n795,
    n877,
    n1566
  );


  or
  g2052
  (
    n1986,
    n1573,
    n814,
    n857,
    n750
  );


  and
  g2053
  (
    n2063,
    n833,
    n1837,
    n887,
    n879
  );


  nor
  g2054
  (
    n2244,
    n1569,
    n1827,
    n1757,
    n877
  );


  nor
  g2055
  (
    n2192,
    n775,
    n1892,
    n747,
    n869
  );


  xnor
  g2056
  (
    n2180,
    n913,
    n1855,
    n921,
    n860
  );


  nand
  g2057
  (
    n2122,
    n852,
    n897,
    n1819,
    n888
  );


  and
  g2058
  (
    n2272,
    n1832,
    n869,
    n1741,
    n1591
  );


  and
  g2059
  (
    n2100,
    n815,
    n826,
    n1787,
    n775
  );


  nand
  g2060
  (
    n2037,
    n840,
    n1844,
    n880,
    n895
  );


  nor
  g2061
  (
    n2026,
    n1622,
    n1764,
    n867,
    n756
  );


  xnor
  g2062
  (
    n1980,
    n874,
    n1875,
    n1546,
    n1922
  );


  and
  g2063
  (
    n2223,
    n1615,
    n1800,
    n922,
    n1891
  );


  or
  g2064
  (
    n2278,
    n882,
    n758,
    n1724,
    n893
  );


  and
  g2065
  (
    n2211,
    n1543,
    n1538,
    n1804,
    n882
  );


  or
  g2066
  (
    n2098,
    n1780,
    n886,
    n1599,
    n1596
  );


  xnor
  g2067
  (
    n2209,
    n821,
    n742,
    n830,
    n1877
  );


  nand
  g2068
  (
    n2031,
    n798,
    n839,
    n1543,
    n1742
  );


  xnor
  g2069
  (
    n2258,
    n1808,
    n766,
    n1755,
    n897
  );


  nor
  g2070
  (
    n1993,
    n1776,
    n1913,
    n768,
    n894
  );


  or
  g2071
  (
    KeyWire_0_21,
    n1775,
    n787,
    n1559,
    n1537
  );


  nand
  g2072
  (
    n2185,
    n894,
    n1857,
    n844,
    n1826
  );


  and
  g2073
  (
    n2103,
    n801,
    n780,
    n1862,
    n1564
  );


  nand
  g2074
  (
    n2113,
    n1777,
    n891,
    n1748,
    n903
  );


  nand
  g2075
  (
    n2175,
    n1608,
    n1828,
    n905,
    n844
  );


  xor
  g2076
  (
    n2121,
    n896,
    n880,
    n838,
    n1627
  );


  nand
  g2077
  (
    n2230,
    n742,
    n880,
    n1837,
    n834
  );


  and
  g2078
  (
    KeyWire_0_13,
    n1802,
    n764,
    n809,
    n897
  );


  and
  g2079
  (
    n2027,
    n1843,
    n1890,
    n1898,
    n815
  );


  and
  g2080
  (
    n2120,
    n1789,
    n834,
    n788,
    n1900
  );


  nor
  g2081
  (
    n1984,
    n1871,
    n1783,
    n746,
    n1779
  );


  nand
  g2082
  (
    n1988,
    n789,
    n1730,
    n1903,
    n851
  );


  nand
  g2083
  (
    n1992,
    n867,
    n799,
    n1884,
    n1806
  );


  xnor
  g2084
  (
    n2158,
    n780,
    n768,
    n827,
    n1597
  );


  nor
  g2085
  (
    n2075,
    n1535,
    n890,
    n1727,
    n1777
  );


  nor
  g2086
  (
    KeyWire_0_51,
    n835,
    n868,
    n809,
    n1811
  );


  and
  g2087
  (
    n2123,
    n828,
    n914,
    n1910,
    n1938
  );


  xnor
  g2088
  (
    n2178,
    n1935,
    n800,
    n861,
    n864
  );


  nand
  g2089
  (
    n2030,
    n764,
    n1540,
    n1534,
    n1816
  );


  xor
  g2090
  (
    n2094,
    n804,
    n813,
    n884,
    n881
  );


  nand
  g2091
  (
    n2205,
    n844,
    n871,
    n1886,
    n916
  );


  nor
  g2092
  (
    n2054,
    n790,
    n1814,
    n1619,
    n828
  );


  nor
  g2093
  (
    n1948,
    n1745,
    n1943,
    n1941,
    n854
  );


  nand
  g2094
  (
    n2058,
    n753,
    n773,
    n1598,
    n891
  );


  xnor
  g2095
  (
    n2238,
    n1581,
    n785,
    n778,
    n869
  );


  and
  g2096
  (
    n2008,
    n856,
    n899,
    n1865,
    n765
  );


  xor
  g2097
  (
    n1952,
    n1872,
    n882,
    n746,
    n890
  );


  or
  g2098
  (
    n2189,
    n806,
    n853,
    n860,
    n907
  );


  xnor
  g2099
  (
    n2015,
    n745,
    n854,
    n866,
    n1611
  );


  or
  g2100
  (
    n2029,
    n1557,
    n1934,
    n1625,
    n1841
  );


  and
  g2101
  (
    n2095,
    n1732,
    n1840,
    n1773
  );


  nor
  g2102
  (
    n1998,
    n1805,
    n1924,
    n1907,
    n1739
  );


  xnor
  g2103
  (
    n1958,
    n894,
    n746,
    n817,
    n1603
  );


  or
  g2104
  (
    n1996,
    n1854,
    n793,
    n1612,
    n1556
  );


  or
  g2105
  (
    n2153,
    n842,
    n1906,
    n892,
    n912
  );


  nand
  g2106
  (
    n2048,
    n871,
    n763,
    n897,
    n789
  );


  xnor
  g2107
  (
    n2036,
    n1727,
    n881,
    n870,
    n834
  );


  nand
  g2108
  (
    n2273,
    n891,
    n1756,
    n1748,
    n1735
  );


  xor
  g2109
  (
    n2150,
    n827,
    n1881,
    n787,
    n814
  );


  and
  g2110
  (
    n2091,
    n1548,
    n1927,
    n850,
    n808
  );


  and
  g2111
  (
    n2143,
    n868,
    n768,
    n1623,
    n788
  );


  or
  g2112
  (
    n2256,
    n1831,
    n761,
    n785,
    n860
  );


  or
  g2113
  (
    n2188,
    n1764,
    n1860,
    n1583,
    n866
  );


  nor
  g2114
  (
    n2267,
    n1935,
    n1604,
    n774,
    n1921
  );


  or
  g2115
  (
    n2055,
    n755,
    n1838,
    n902,
    n1938
  );


  or
  g2116
  (
    n2142,
    n1583,
    n1563,
    n782,
    n1807
  );


  and
  g2117
  (
    n2050,
    n1576,
    n1723,
    n820,
    n793
  );


  xor
  g2118
  (
    n2162,
    n846,
    n916,
    n854,
    n796
  );


  xor
  g2119
  (
    n2168,
    n880,
    n829,
    n868,
    n792
  );


  nand
  g2120
  (
    n2099,
    n1531,
    n784,
    n1933,
    n878
  );


  xor
  g2121
  (
    n2176,
    n829,
    n896,
    n1594,
    n1892
  );


  xor
  g2122
  (
    n1947,
    n808,
    n1579,
    n1899,
    n763
  );


  nand
  g2123
  (
    n2288,
    n1568,
    n839,
    n770,
    n818
  );


  nand
  g2124
  (
    n1968,
    n1812,
    n745,
    n895,
    n807
  );


  nor
  g2125
  (
    n1950,
    n1568,
    n1795,
    n1812,
    n792
  );


  and
  g2126
  (
    n1973,
    n804,
    n875,
    n873,
    n866
  );


  or
  g2127
  (
    n2184,
    n1799,
    n810,
    n913,
    n1822
  );


  nor
  g2128
  (
    n2228,
    n1791,
    n1604,
    n1542,
    n1603
  );


  xnor
  g2129
  (
    n2045,
    n1532,
    n789,
    n921
  );


  nor
  g2130
  (
    n2066,
    n858,
    n816,
    n1626,
    n843
  );


  or
  g2131
  (
    n2164,
    n812,
    n796,
    n1575,
    n745
  );


  or
  g2132
  (
    n2190,
    n863,
    n1855,
    n748,
    n864
  );


  nor
  g2133
  (
    n2148,
    n1607,
    n888,
    n785,
    n903
  );


  or
  g2134
  (
    n2177,
    n1925,
    n1854,
    n1909,
    n1868
  );


  nor
  g2135
  (
    n2227,
    n914,
    n777,
    n1555,
    n825
  );


  xnor
  g2136
  (
    n1971,
    n1852,
    n743,
    n1584,
    n1722
  );


  or
  g2137
  (
    n2056,
    n950,
    n1870,
    n1796,
    n1820
  );


  or
  g2138
  (
    n2271,
    n1883,
    n906,
    n1939,
    n1749
  );


  and
  g2139
  (
    n2052,
    n744,
    n1851,
    n745,
    n1845
  );


  and
  g2140
  (
    n2009,
    n759,
    n803,
    n1613,
    n1767
  );


  and
  g2141
  (
    n1967,
    n827,
    n1898,
    n922,
    n899
  );


  and
  g2142
  (
    n2131,
    n774,
    n1905,
    n839,
    n764
  );


  or
  g2143
  (
    n2108,
    n1937,
    n873,
    n903,
    n752
  );


  xnor
  g2144
  (
    n2082,
    n765,
    n847,
    n1900,
    n887
  );


  or
  g2145
  (
    n2201,
    n1765,
    n922,
    n865,
    n1574
  );


  nand
  g2146
  (
    n2252,
    n885,
    n797,
    n1809,
    n828
  );


  nand
  g2147
  (
    n1979,
    n1904,
    n786,
    n803,
    n1871
  );


  xnor
  g2148
  (
    n2207,
    n920,
    n1908,
    n847,
    n1587
  );


  nor
  g2149
  (
    n2072,
    n1906,
    n865,
    n1914,
    n902
  );


  nand
  g2150
  (
    n2170,
    n1731,
    n1910,
    n1879,
    n743
  );


  xnor
  g2151
  (
    n2119,
    n849,
    n912,
    n1911,
    n840
  );


  xnor
  g2152
  (
    n2237,
    n873,
    n1829,
    n1774,
    n1772
  );


  and
  g2153
  (
    n2053,
    n1942,
    n1788,
    n1725,
    n1571
  );


  xnor
  g2154
  (
    n1999,
    n891,
    n1566,
    n818,
    n1927
  );


  or
  g2155
  (
    n2232,
    n783,
    n1592,
    n852,
    n743
  );


  xor
  g2156
  (
    n2285,
    n759,
    n902,
    n1894,
    n1558
  );


  or
  g2157
  (
    n2126,
    n751,
    n1819,
    n805,
    n1553
  );


  xnor
  g2158
  (
    KeyWire_0_52,
    n1606,
    n841,
    n769,
    n1864
  );


  and
  g2159
  (
    n2138,
    n1781,
    n848,
    n753,
    n872
  );


  nand
  g2160
  (
    n2196,
    n790,
    n900,
    n796,
    n845
  );


  xnor
  g2161
  (
    n2274,
    n1853,
    n832,
    n1734,
    n1578
  );


  nor
  g2162
  (
    n2127,
    n768,
    n842,
    n1928,
    n1922
  );


  or
  g2163
  (
    n2097,
    n1610,
    n772,
    n809,
    n1896
  );


  xor
  g2164
  (
    n2093,
    n1945,
    n827,
    n1840,
    n1867
  );


  nand
  g2165
  (
    n2051,
    n1841,
    n1801,
    n1578,
    n1554
  );


  xnor
  g2166
  (
    n2151,
    n855,
    n856,
    n846,
    n1941
  );


  nor
  g2167
  (
    n2261,
    n923,
    n896,
    n838,
    n876
  );


  and
  g2168
  (
    n2204,
    n826,
    n773,
    n1539,
    n1549
  );


  nor
  g2169
  (
    n2069,
    n850,
    n1534,
    n884,
    n793
  );


  nand
  g2170
  (
    n2128,
    n756,
    n811,
    n918,
    n1863
  );


  nand
  g2171
  (
    n2074,
    n1539,
    n1728,
    n1785,
    n1561
  );


  xor
  g2172
  (
    n2102,
    n872,
    n816,
    n1755,
    n1894
  );


  and
  g2173
  (
    n1946,
    n876,
    n1609,
    n1861,
    n1873
  );


  xor
  g2174
  (
    n2179,
    n917,
    n807,
    n860,
    n1936
  );


  or
  g2175
  (
    n2135,
    n795,
    n1834,
    n1793,
    n779
  );


  xor
  g2176
  (
    n2013,
    n910,
    n859,
    n921,
    n1842
  );


  nor
  g2177
  (
    n1985,
    n1556,
    n1733,
    n1788,
    n830
  );


  xor
  g2178
  (
    n2118,
    n805,
    n910,
    n1818,
    n915
  );


  nor
  g2179
  (
    n2046,
    n790,
    n905,
    n1784,
    n1861
  );


  nor
  g2180
  (
    n2200,
    n1822,
    n1549,
    n1796,
    n1928
  );


  nor
  g2181
  (
    n2011,
    n919,
    n1588,
    n867,
    n901
  );


  nand
  g2182
  (
    n2281,
    n1814,
    n1874,
    n1899,
    n1897
  );


  and
  g2183
  (
    n1962,
    n1569,
    n1824,
    n864,
    n1907
  );


  and
  g2184
  (
    n2049,
    n855,
    n840,
    n1886,
    n919
  );


  xor
  g2185
  (
    n2025,
    n767,
    n904,
    n1546,
    n907
  );


  nor
  g2186
  (
    n1957,
    n741,
    n896,
    n885,
    n1803
  );


  xnor
  g2187
  (
    KeyWire_0_16,
    n1791,
    n1916,
    n1860,
    n759
  );


  or
  g2188
  (
    n2079,
    n862,
    n842,
    n806,
    n765
  );


  or
  g2189
  (
    n2083,
    n826,
    n1763,
    n820,
    n1606
  );


  nor
  g2190
  (
    n2218,
    n1919,
    n1562,
    n794,
    n908
  );


  and
  g2191
  (
    n2012,
    n1761,
    n1573,
    n1747,
    n1785
  );


  xor
  g2192
  (
    n2068,
    n1759,
    n1805,
    n1594,
    n849
  );


  and
  g2193
  (
    n2194,
    n742,
    n781,
    n1940,
    n1601
  );


  or
  g2194
  (
    n2016,
    n788,
    n913,
    n810,
    n1824
  );


  xnor
  g2195
  (
    n2245,
    n791,
    n777,
    n1620,
    n1775
  );


  and
  g2196
  (
    n2129,
    n814,
    n771,
    n1800,
    n1593
  );


  nand
  g2197
  (
    n2073,
    n1762,
    n753,
    n908,
    n909
  );


  and
  g2198
  (
    n2187,
    n1625,
    n1609,
    n879,
    n1761
  );


  or
  g2199
  (
    n2156,
    n1870,
    n1763,
    n1867,
    n807
  );


  and
  g2200
  (
    n2193,
    n1579,
    n1624,
    n901,
    n1595
  );


  and
  g2201
  (
    n2010,
    n1902,
    n1931,
    n798,
    n898
  );


  nor
  g2202
  (
    n2076,
    n848,
    n817,
    n1590,
    n1859
  );


  nand
  g2203
  (
    n2086,
    n915,
    n750,
    n851,
    n1835
  );


  xor
  g2204
  (
    n2224,
    n845,
    n1628,
    n856,
    n799
  );


  nor
  g2205
  (
    n2105,
    n1771,
    n1722,
    n876,
    n835
  );


  xor
  g2206
  (
    n2155,
    n883,
    n1772,
    n813,
    n1757
  );


  nand
  g2207
  (
    n1954,
    n750,
    n1588,
    n1765,
    n901
  );


  nor
  g2208
  (
    n2287,
    n1601,
    n1559,
    n874,
    n821
  );


  xnor
  g2209
  (
    n2084,
    n1535,
    n836,
    n851,
    n1915
  );


  or
  g2210
  (
    n1965,
    n1944,
    n894,
    n1778,
    n843
  );


  nand
  g2211
  (
    n2166,
    n750,
    n765,
    n824,
    n1857
  );


  xor
  g2212
  (
    n2173,
    n785,
    n777,
    n1850,
    n906
  );


  and
  g2213
  (
    n2116,
    n778,
    n1846,
    n1752,
    n857
  );


  and
  g2214
  (
    n2043,
    n865,
    n1866,
    n1829,
    n1839
  );


  xor
  g2215
  (
    n2217,
    n1786,
    n1789,
    n742,
    n831
  );


  xnor
  g2216
  (
    n2021,
    n1760,
    n882,
    n1737,
    n900
  );


  and
  g2217
  (
    n2145,
    n1925,
    n1923,
    n1771,
    n819
  );


  xor
  g2218
  (
    n2254,
    n1929,
    n1746,
    n1881,
    n870
  );


  xor
  g2219
  (
    n2276,
    n917,
    n909,
    n1876,
    n1733
  );


  or
  g2220
  (
    n2226,
    n761,
    n871,
    n764,
    n1618
  );


  nand
  g2221
  (
    n2061,
    n1555,
    n1792,
    n839,
    n889
  );


  xnor
  g2222
  (
    n2163,
    n1818,
    n794,
    n907,
    n836
  );


  nand
  g2223
  (
    n2225,
    n812,
    n816,
    n903,
    n1811
  );


  xnor
  g2224
  (
    n2259,
    n779,
    n885,
    n770,
    n1581
  );


  and
  g2225
  (
    n2183,
    n772,
    n811,
    n749,
    n1897
  );


  xor
  g2226
  (
    n2246,
    n836,
    n1531,
    n1919,
    n1926
  );


  or
  g2227
  (
    n2085,
    n776,
    n1567,
    n831,
    n1803
  );


  and
  g2228
  (
    n1969,
    n878,
    n821,
    n1828,
    n1760
  );


  nor
  g2229
  (
    n2242,
    n811,
    n858,
    n1752,
    n741
  );


  xor
  g2230
  (
    n2289,
    n911,
    n748,
    n1746,
    n886
  );


  nor
  g2231
  (
    n2241,
    n1541,
    n800,
    n1735,
    n1753
  );


  nor
  g2232
  (
    n2286,
    n1742,
    n1851,
    n793,
    n1564
  );


  nand
  g2233
  (
    n2107,
    n1571,
    n895,
    n1622,
    n829
  );


  xor
  g2234
  (
    n2080,
    n756,
    n802,
    n876,
    n1849
  );


  or
  g2235
  (
    n2249,
    n805,
    n1835,
    n812,
    n752
  );


  xor
  g2236
  (
    n2229,
    n923,
    n837,
    n861,
    n784
  );


  nor
  g2237
  (
    n2284,
    n837,
    n796,
    n1901,
    n918
  );


  xnor
  g2238
  (
    n2003,
    n1595,
    n1758,
    n757,
    n1621
  );


  nor
  g2239
  (
    n2169,
    n1810,
    n1736,
    n825,
    n762
  );


  and
  g2240
  (
    n2132,
    n823,
    n775,
    n863,
    n1937
  );


  xor
  g2241
  (
    n2044,
    n778,
    n854,
    n1873,
    n802
  );


  and
  g2242
  (
    n2081,
    n1832,
    n1758,
    n763,
    n1856
  );


  xnor
  g2243
  (
    n2096,
    n910,
    n1591,
    n1944,
    n848
  );


  xor
  g2244
  (
    n2182,
    n1547,
    n1895,
    n871,
    n1821
  );


  nand
  g2245
  (
    n2233,
    n1793,
    n802,
    n893,
    n1624
  );


  xor
  g2246
  (
    n2307,
    n2094,
    n1956,
    n2081,
    n2175
  );


  nor
  g2247
  (
    n2301,
    n2034,
    n1951,
    n2189,
    n2155
  );


  nor
  g2248
  (
    n2379,
    n2236,
    n1985,
    n2017,
    n2158
  );


  nor
  g2249
  (
    n2341,
    n1996,
    n2254,
    n2154,
    n2073
  );


  or
  g2250
  (
    n2387,
    n1990,
    n2184,
    n2009,
    n2064
  );


  nor
  g2251
  (
    n2365,
    n2083,
    n1983,
    n2260,
    n2008
  );


  xor
  g2252
  (
    n2380,
    n1984,
    n2010,
    n2071,
    n2230
  );


  nor
  g2253
  (
    n2393,
    n2139,
    n2178,
    n1975,
    n2179
  );


  nor
  g2254
  (
    n2423,
    n2176,
    n2046,
    n1962,
    n2134
  );


  or
  g2255
  (
    n2319,
    n1949,
    n2164,
    n2225,
    n2018
  );


  nor
  g2256
  (
    n2364,
    n2002,
    n2028,
    n2070,
    n2029
  );


  nand
  g2257
  (
    n2315,
    n2152,
    n2115,
    n2058,
    n1982
  );


  nand
  g2258
  (
    n2360,
    n2077,
    n2204,
    n2145,
    n1961
  );


  xor
  g2259
  (
    n2349,
    n1993,
    n1982,
    n1963,
    n2197
  );


  nand
  g2260
  (
    n2442,
    n2257,
    n2109,
    n2019,
    n2006
  );


  nor
  g2261
  (
    n2425,
    n2160,
    n2198,
    n2255,
    n2171
  );


  xor
  g2262
  (
    n2424,
    n1967,
    n1979,
    n2126,
    n2233
  );


  nand
  g2263
  (
    n2297,
    n2234,
    n2224,
    n2129,
    n2112
  );


  xor
  g2264
  (
    n2299,
    n1952,
    n2111,
    n2050,
    n2216
  );


  xor
  g2265
  (
    n2416,
    n1966,
    n2227,
    n2027,
    n2246
  );


  and
  g2266
  (
    n2399,
    n2269,
    n2059,
    n2214,
    n2154
  );


  xnor
  g2267
  (
    n2342,
    n2200,
    n1965,
    n1983,
    n2078
  );


  xor
  g2268
  (
    n2436,
    n1999,
    n2016,
    n2048,
    n1948
  );


  xor
  g2269
  (
    n2439,
    n2190,
    n2036,
    n1997,
    n2197
  );


  or
  g2270
  (
    n2396,
    n2148,
    n2003,
    n2121,
    n2267
  );


  and
  g2271
  (
    n2420,
    n2006,
    n2260,
    n2156,
    n1970
  );


  nor
  g2272
  (
    n2303,
    n2001,
    n2052,
    n2069,
    n2034
  );


  xor
  g2273
  (
    n2384,
    n2259,
    n2139,
    n2090,
    n2255
  );


  nand
  g2274
  (
    n2441,
    n2016,
    n2040,
    n1989,
    n2194
  );


  or
  g2275
  (
    n2382,
    n2012,
    n2207,
    n2246,
    n2212
  );


  nor
  g2276
  (
    n2337,
    n2211,
    n1964,
    n2262,
    n2159
  );


  nand
  g2277
  (
    n2421,
    n2076,
    n2052,
    n2110,
    n1995
  );


  xnor
  g2278
  (
    n2359,
    n2053,
    n2241,
    n2103,
    n2151
  );


  xor
  g2279
  (
    n2386,
    n2089,
    n2126,
    n2230,
    n2263
  );


  nand
  g2280
  (
    n2374,
    n2263,
    n2147,
    n2184,
    n2210
  );


  xnor
  g2281
  (
    n2409,
    n2042,
    n2183,
    n2082,
    n1976
  );


  nand
  g2282
  (
    n2317,
    n2026,
    n2108,
    n2058,
    n2014
  );


  nand
  g2283
  (
    n2357,
    n2086,
    n2025,
    n1977,
    n2217
  );


  xor
  g2284
  (
    n2348,
    n2186,
    n2047,
    n1947,
    n2232
  );


  nor
  g2285
  (
    n2391,
    n2161,
    n2000,
    n2075,
    n2209
  );


  xnor
  g2286
  (
    n2309,
    n1969,
    n2131,
    n2024,
    n2037
  );


  xnor
  g2287
  (
    n2346,
    n2007,
    n2211,
    n2118,
    n2251
  );


  xor
  g2288
  (
    n2328,
    n2187,
    n2178,
    n2203,
    n2256
  );


  nor
  g2289
  (
    n2339,
    n2202,
    n2103,
    n1999,
    n2113
  );


  xor
  g2290
  (
    n2397,
    n2258,
    n1985,
    n2125,
    n2001
  );


  nand
  g2291
  (
    n2295,
    n2169,
    n2079,
    n2193,
    n1972
  );


  and
  g2292
  (
    n2310,
    n1960,
    n2195,
    n2250,
    n2168
  );


  xnor
  g2293
  (
    n2318,
    n2023,
    n2152,
    n2074,
    n2142
  );


  nand
  g2294
  (
    n2389,
    n2020,
    n2060,
    n2043,
    n2192
  );


  and
  g2295
  (
    n2340,
    n2065,
    n2241,
    n2170,
    n1965
  );


  nor
  g2296
  (
    n2408,
    n2240,
    n2079,
    n2203,
    n2251
  );


  or
  g2297
  (
    n2437,
    n2244,
    n2173,
    n2132,
    n1991
  );


  or
  g2298
  (
    n2324,
    n2123,
    n2008,
    n2149,
    n2143
  );


  nor
  g2299
  (
    n2358,
    n2031,
    n2088,
    n2141,
    n2242
  );


  or
  g2300
  (
    n2417,
    n1992,
    n2061,
    n1980,
    n2073
  );


  xnor
  g2301
  (
    n2450,
    n2035,
    n1946,
    n2122,
    n2096
  );


  and
  g2302
  (
    n2445,
    n1958,
    n2084,
    n2082,
    n2261
  );


  nor
  g2303
  (
    n2291,
    n2237,
    n2117,
    n1949,
    n2156
  );


  or
  g2304
  (
    n2313,
    n2031,
    n2224,
    n1956,
    n1957
  );


  or
  g2305
  (
    n2347,
    n2049,
    n2261,
    n2015,
    n1959
  );


  and
  g2306
  (
    n2452,
    n2011,
    n2166,
    n1970,
    n2124
  );


  and
  g2307
  (
    n2363,
    n2225,
    n2022,
    n1973,
    n1977
  );


  xnor
  g2308
  (
    n2395,
    n2028,
    n2032,
    n2071,
    n2080
  );


  or
  g2309
  (
    n2333,
    n2039,
    n2041,
    n2004,
    n2248
  );


  nor
  g2310
  (
    n2376,
    n2259,
    n2022,
    n2137,
    n2056
  );


  xor
  g2311
  (
    n2311,
    n2145,
    n2165,
    n2213,
    n2134
  );


  xor
  g2312
  (
    n2398,
    n2219,
    n2209,
    n2256,
    n2228
  );


  and
  g2313
  (
    n2426,
    n2097,
    n2170,
    n2137,
    n2038
  );


  xnor
  g2314
  (
    n2418,
    n2242,
    n2207,
    n1987,
    n2039
  );


  xnor
  g2315
  (
    n2413,
    n2101,
    n2267,
    n2102,
    n2062
  );


  and
  g2316
  (
    n2381,
    n2151,
    n2176,
    n2217,
    n2102
  );


  and
  g2317
  (
    n2373,
    n2243,
    n1974,
    n1990,
    n2168
  );


  xnor
  g2318
  (
    n2448,
    n2252,
    n2253,
    n2005,
    n2074
  );


  xnor
  g2319
  (
    n2296,
    n2220,
    n2061,
    n2188,
    n2021
  );


  xor
  g2320
  (
    n2435,
    n1946,
    n2192,
    n2144,
    n2147
  );


  and
  g2321
  (
    n2407,
    n2113,
    n2063,
    n2269,
    n2081
  );


  nand
  g2322
  (
    n2321,
    n1963,
    n1979,
    n2215,
    n2221
  );


  nor
  g2323
  (
    n2371,
    n2012,
    n2153,
    n2140,
    n1998
  );


  and
  g2324
  (
    n2343,
    n2245,
    n2062,
    n1976,
    n2116
  );


  nand
  g2325
  (
    n2306,
    n2084,
    n2050,
    n2185,
    n1988
  );


  or
  g2326
  (
    n2332,
    n2229,
    n2040,
    n2112,
    n2171
  );


  nor
  g2327
  (
    n2304,
    n2085,
    n2138,
    n2066,
    n1989
  );


  and
  g2328
  (
    n2327,
    n2086,
    n2208,
    n2244,
    n2093
  );


  nand
  g2329
  (
    n2316,
    n2146,
    n2108,
    n2070,
    n2055
  );


  xnor
  g2330
  (
    n2350,
    n2106,
    n1968,
    n2268,
    n1957
  );


  or
  g2331
  (
    n2404,
    n2198,
    n2033,
    n2193,
    n2010
  );


  nor
  g2332
  (
    n2427,
    n1958,
    n2100,
    n2181,
    n1967
  );


  and
  g2333
  (
    n2394,
    n1948,
    n2130,
    n2098,
    n2090
  );


  xor
  g2334
  (
    n2366,
    n2142,
    n2257,
    n2076,
    n2120
  );


  xor
  g2335
  (
    n2434,
    n2119,
    n2000,
    n2166,
    n2191
  );


  and
  g2336
  (
    n2432,
    n2132,
    n2054,
    n2239,
    n2165
  );


  xnor
  g2337
  (
    KeyWire_0_44,
    n1955,
    n2115,
    n2180,
    n2107
  );


  xor
  g2338
  (
    n2429,
    n2240,
    n2023,
    n2232,
    n2049
  );


  nand
  g2339
  (
    n2403,
    n2199,
    n2186,
    n2128,
    n2140
  );


  and
  g2340
  (
    n2338,
    n2179,
    n2053,
    n2215,
    n2045
  );


  xnor
  g2341
  (
    n2402,
    n2177,
    n2136,
    n2247,
    n1997
  );


  nand
  g2342
  (
    n2353,
    n2092,
    n2222,
    n2221,
    n2105
  );


  and
  g2343
  (
    n2430,
    n2169,
    n2119,
    n2109,
    n2057
  );


  xnor
  g2344
  (
    n2300,
    n2174,
    n2167,
    n2072,
    n2021
  );


  nor
  g2345
  (
    n2362,
    n2048,
    n2149,
    n2249,
    n2030
  );


  xor
  g2346
  (
    n2370,
    n2219,
    n1984,
    n1978,
    n1952
  );


  and
  g2347
  (
    n2344,
    n2264,
    n1998,
    n1954,
    n2127
  );


  and
  g2348
  (
    n2361,
    n2226,
    n2044,
    n2206,
    n2135
  );


  xnor
  g2349
  (
    n2329,
    n2223,
    n2265,
    n2172,
    n2235
  );


  nor
  g2350
  (
    n2411,
    n2133,
    n2067,
    n2174,
    n2041
  );


  nand
  g2351
  (
    n2314,
    n2208,
    n2004,
    n2005,
    n2007
  );


  and
  g2352
  (
    n2447,
    n1951,
    n2087,
    n2243,
    n1955
  );


  xor
  g2353
  (
    n2449,
    n2032,
    n1994,
    n2066,
    n2051
  );


  nor
  g2354
  (
    n2400,
    n2124,
    n2180,
    n1971,
    n2143
  );


  xor
  g2355
  (
    n2330,
    n2069,
    n2185,
    n2253,
    n2254
  );


  and
  g2356
  (
    n2312,
    n1974,
    n2104,
    n2116,
    n2059
  );


  or
  g2357
  (
    n2444,
    n1973,
    n2068,
    n2250,
    n1960
  );


  nand
  g2358
  (
    n2438,
    n2196,
    n2128,
    n1950,
    n2056
  );


  nand
  g2359
  (
    n2331,
    n2064,
    n2033,
    n2155,
    n2196
  );


  nand
  g2360
  (
    n2345,
    n2172,
    n2054,
    n2017,
    n2099
  );


  nand
  g2361
  (
    n2415,
    n2191,
    n1972,
    n2089,
    n2194
  );


  and
  g2362
  (
    n2336,
    n1966,
    n2121,
    n2038,
    n2092
  );


  and
  g2363
  (
    n2355,
    n1978,
    n2051,
    n2200,
    n2248
  );


  and
  g2364
  (
    n2428,
    n2160,
    n2262,
    n1975,
    n2015
  );


  xnor
  g2365
  (
    n2368,
    n2047,
    n2019,
    n2105,
    n2159
  );


  and
  g2366
  (
    n2405,
    n2231,
    n1962,
    n2029,
    n1953
  );


  nor
  g2367
  (
    n2372,
    n1947,
    n2236,
    n2216,
    n2043
  );


  nand
  g2368
  (
    n2326,
    n2104,
    n2150,
    n1991,
    n2144
  );


  and
  g2369
  (
    n2422,
    n2229,
    n2205,
    n2201,
    n2037
  );


  nor
  g2370
  (
    n2378,
    n1953,
    n2264,
    n2163,
    n2093
  );


  nand
  g2371
  (
    n2302,
    n2057,
    n2183,
    n2018,
    n2095
  );


  or
  g2372
  (
    n2305,
    n1954,
    n2003,
    n2223,
    n2222
  );


  xor
  g2373
  (
    n2375,
    n2233,
    n2227,
    n2158,
    n2096
  );


  nand
  g2374
  (
    n2352,
    n2148,
    n2114,
    n2098,
    n2266
  );


  or
  g2375
  (
    n2412,
    n2212,
    n2122,
    n2065,
    n2060
  );


  xnor
  g2376
  (
    n2351,
    n2157,
    n2234,
    n1986,
    n1988
  );


  nor
  g2377
  (
    n2385,
    n2107,
    n2091,
    n2228,
    n2100
  );


  or
  g2378
  (
    n2410,
    n2177,
    n2097,
    n2009,
    n2175
  );


  nand
  g2379
  (
    n2388,
    n2011,
    n2077,
    n2235,
    n2123
  );


  and
  g2380
  (
    n2356,
    n2120,
    n2091,
    n2106,
    n2266
  );


  and
  g2381
  (
    n2451,
    n2036,
    n1992,
    n2020,
    n2075
  );


  nand
  g2382
  (
    n2390,
    n2117,
    n2182,
    n1959,
    n2094
  );


  nand
  g2383
  (
    n2325,
    n2201,
    n2173,
    n2249,
    n2218
  );


  xnor
  g2384
  (
    n2446,
    n2099,
    n2162,
    n2042,
    n1995
  );


  nor
  g2385
  (
    n2320,
    n2252,
    n2210,
    n2068,
    n1987
  );


  nand
  g2386
  (
    n2406,
    n2202,
    n2214,
    n2161,
    n2181
  );


  and
  g2387
  (
    n2414,
    n2055,
    n1950,
    n2182,
    n2220
  );


  xnor
  g2388
  (
    n2322,
    n1981,
    n2125,
    n2027,
    n2014
  );


  xnor
  g2389
  (
    n2431,
    n2111,
    n2044,
    n2085,
    n2226
  );


  and
  g2390
  (
    n2308,
    n1994,
    n2231,
    n2204,
    n1986
  );


  nor
  g2391
  (
    n2367,
    n2218,
    n2135,
    n2045,
    n2153
  );


  nand
  g2392
  (
    n2443,
    n2035,
    n2187,
    n2206,
    n2088
  );


  nor
  g2393
  (
    n2392,
    n2188,
    n2080,
    n2245,
    n2129
  );


  xnor
  g2394
  (
    n2440,
    n2025,
    n2026,
    n1969,
    n2114
  );


  and
  g2395
  (
    n2292,
    n1964,
    n1971,
    n2133,
    n2213
  );


  and
  g2396
  (
    n2323,
    n2013,
    n2127,
    n2237,
    n2072
  );


  and
  g2397
  (
    n2369,
    n2238,
    n2195,
    n1996,
    n2118
  );


  and
  g2398
  (
    n2377,
    n1961,
    n2002,
    n2138,
    n2205
  );


  xor
  g2399
  (
    n2298,
    n2164,
    n2078,
    n2162,
    n2046
  );


  xnor
  g2400
  (
    n2433,
    n2268,
    n2136,
    n2146,
    n2238
  );


  xnor
  g2401
  (
    n2383,
    n2101,
    n2199,
    n2258,
    n1993
  );


  nor
  g2402
  (
    n2294,
    n2150,
    n1980,
    n2190,
    n2013
  );


  and
  g2403
  (
    n2354,
    n2130,
    n2095,
    n2131,
    n2265
  );


  and
  g2404
  (
    n2419,
    n2083,
    n2087,
    n2067,
    n2239
  );


  xor
  g2405
  (
    n2334,
    n2247,
    n2189,
    n2157,
    n2167
  );


  xnor
  g2406
  (
    n2335,
    n2163,
    n2110,
    n1981,
    n2063
  );


  xnor
  g2407
  (
    n2401,
    n2024,
    n1968,
    n2030,
    n2141
  );


  xnor
  g2408
  (
    n2457,
    n2294,
    n2303,
    n2302,
    n2293
  );


  and
  g2409
  (
    n2454,
    n2304,
    n2299,
    n2291,
    n2307
  );


  nor
  g2410
  (
    n2455,
    n2295,
    n2309,
    n2298,
    n2310
  );


  nor
  g2411
  (
    n2453,
    n2297,
    n2305,
    n2300,
    n2296
  );


  xnor
  g2412
  (
    n2456,
    n2306,
    n2292,
    n2301,
    n2308
  );


  not
  g2413
  (
    n2458,
    n2457
  );


  buf
  g2414
  (
    n2461,
    n2455
  );


  not
  g2415
  (
    n2460,
    n2454
  );


  not
  g2416
  (
    n2459,
    n2456
  );


  buf
  g2417
  (
    n2462,
    n2458
  );


  not
  g2418
  (
    n2463,
    n2458
  );


  buf
  g2419
  (
    n2464,
    n2463
  );


  not
  g2420
  (
    n2466,
    n1030
  );


  xor
  g2421
  (
    n2467,
    n2463,
    n2270,
    n1031,
    n2311
  );


  nand
  g2422
  (
    n2465,
    n1030,
    n2270,
    n2462
  );


  xor
  g2423
  (
    n2470,
    n2317,
    n2314,
    n2465
  );


  nor
  g2424
  (
    n2469,
    n2315,
    n2316,
    n2318
  );


  xor
  g2425
  (
    n2468,
    n2312,
    n2464,
    n2313
  );


  nand
  g2426
  (
    n2478,
    n2319,
    n2339,
    n2345,
    n2468
  );


  nor
  g2427
  (
    n2477,
    n2341,
    n2468,
    n2338
  );


  and
  g2428
  (
    n2474,
    n2334,
    n2324,
    n2469
  );


  nor
  g2429
  (
    n2473,
    n2331,
    n2470,
    n2335,
    n2329
  );


  or
  g2430
  (
    n2472,
    n2470,
    n2320,
    n2343,
    n2322
  );


  xor
  g2431
  (
    n2476,
    n2340,
    n2337,
    n2469,
    n2328
  );


  xor
  g2432
  (
    n2479,
    n2327,
    n2325,
    n2333,
    n2336
  );


  or
  g2433
  (
    n2475,
    n2326,
    n2344,
    n2321,
    n2342
  );


  xor
  g2434
  (
    KeyWire_0_46,
    n2470,
    n2323,
    n2330,
    n2332
  );


  nand
  g2435
  (
    n2484,
    n2358,
    n2346,
    n2357,
    n2474
  );


  or
  g2436
  (
    n2480,
    n2352,
    n2359,
    n2356,
    n2350
  );


  or
  g2437
  (
    n2482,
    n2354,
    n2472,
    n2473,
    n2360
  );


  or
  g2438
  (
    n2481,
    n2347,
    n2348,
    n2475,
    n2349
  );


  nor
  g2439
  (
    n2483,
    n2351,
    n2471,
    n2355,
    n2353
  );


  nand
  g2440
  (
    n2486,
    n2364,
    n2372,
    n2369,
    n2363
  );


  nand
  g2441
  (
    n2488,
    n2365,
    n2484,
    n2361,
    n2362
  );


  nor
  g2442
  (
    n2485,
    n2481,
    n2366,
    n2371,
    n2368
  );


  xor
  g2443
  (
    n2487,
    n2367,
    n2483,
    n2482,
    n2370
  );


  xor
  g2444
  (
    n2500,
    n1633,
    n2458,
    n2459,
    n2486
  );


  nand
  g2445
  (
    n2499,
    n2467,
    n2488,
    n2485,
    n2460
  );


  nand
  g2446
  (
    n2493,
    n2373,
    n2461,
    n2459
  );


  nor
  g2447
  (
    n2490,
    n1631,
    n2486,
    n2487
  );


  or
  g2448
  (
    n2489,
    n2458,
    n1640,
    n2460,
    n1628
  );


  xnor
  g2449
  (
    n2491,
    n1634,
    n2485,
    n2486,
    n1639
  );


  xor
  g2450
  (
    n2497,
    n1634,
    n2485,
    n2461
  );


  xor
  g2451
  (
    n2503,
    n1641,
    n2461,
    n2465,
    n1637
  );


  or
  g2452
  (
    n2504,
    n2487,
    n2488,
    n1638,
    n2466
  );


  xnor
  g2453
  (
    n2501,
    n2466,
    n2485,
    n1630,
    n1629
  );


  nand
  g2454
  (
    n2502,
    n1640,
    n1636,
    n1630,
    n1641
  );


  nand
  g2455
  (
    n2498,
    n2487,
    n2488,
    n1632,
    n1031
  );


  and
  g2456
  (
    n2494,
    n2460,
    n1631,
    n1638,
    n2374
  );


  xor
  g2457
  (
    n2496,
    n2460,
    n2487,
    n1636,
    n1639
  );


  xnor
  g2458
  (
    n2495,
    n2488,
    n1635,
    n1633,
    n2459
  );


  xnor
  g2459
  (
    n2492,
    n1632,
    n1635,
    n1629,
    n1637
  );


  and
  g2460
  (
    n2517,
    n2496,
    n2500,
    n1003,
    n2377
  );


  or
  g2461
  (
    n2508,
    n2499,
    n2497,
    n2491,
    n2496
  );


  nor
  g2462
  (
    n2516,
    n2495,
    n2381,
    n2501,
    n950
  );


  and
  g2463
  (
    n2511,
    n2498,
    n2492,
    n2490,
    n2495
  );


  xnor
  g2464
  (
    n2510,
    n2491,
    n2504,
    n2500
  );


  nand
  g2465
  (
    n2506,
    n2494,
    n2378,
    n2492,
    n2376
  );


  xor
  g2466
  (
    n2512,
    n2382,
    n2498,
    n2500,
    n2467
  );


  xor
  g2467
  (
    n2513,
    n2502,
    n2499,
    n2489,
    n2380
  );


  or
  g2468
  (
    n2519,
    n2500,
    n2497,
    n2501
  );


  and
  g2469
  (
    n2518,
    n2497,
    n2503,
    n2498,
    n2504
  );


  or
  g2470
  (
    n2514,
    n2494,
    n2499,
    n2501
  );


  and
  g2471
  (
    n2507,
    n2490,
    n2502,
    n2504,
    n2493
  );


  nand
  g2472
  (
    n2509,
    n2375,
    n1003,
    n2503
  );


  nor
  g2473
  (
    n2505,
    n2379,
    n2497,
    n2489,
    n2502
  );


  nor
  g2474
  (
    n2515,
    n2502,
    n2503,
    n2498,
    n2493
  );


  nor
  g2475
  (
    n2524,
    n2516,
    n2508,
    n2510,
    n2505
  );


  or
  g2476
  (
    n2521,
    n2513,
    n2515,
    n2506,
    n2517
  );


  nor
  g2477
  (
    n2522,
    n2518,
    n2511,
    n2512,
    n2515
  );


  xnor
  g2478
  (
    n2520,
    n2510,
    n2509,
    n2514,
    n2508
  );


  xnor
  g2479
  (
    n2526,
    n2512,
    n2505,
    n2507,
    n2509
  );


  xor
  g2480
  (
    n2523,
    n2507,
    n2513,
    n2518,
    n2516
  );


  and
  g2481
  (
    n2525,
    n2514,
    n2517,
    n2511,
    n2506
  );


  nand
  g2482
  (
    n2527,
    n2384,
    n2387,
    n2526,
    n2386
  );


  and
  g2483
  (
    n2528,
    n2388,
    n2525,
    n2385,
    n2383
  );


  nor
  g2484
  (
    n2532,
    n2527,
    n2528,
    n1052,
    n2477
  );


  nor
  g2485
  (
    n2534,
    n2519,
    n2527,
    n2478,
    n2391
  );


  nand
  g2486
  (
    n2531,
    n2528,
    n1053,
    n2390
  );


  nand
  g2487
  (
    n2530,
    n2528,
    n1015,
    n2527,
    n2479
  );


  nand
  g2488
  (
    n2533,
    n2527,
    n2528,
    n2389,
    n2479
  );


  xor
  g2489
  (
    n2529,
    n2476,
    n1015,
    n924,
    n1644
  );


  nand
  g2490
  (
    n2536,
    n1031,
    n1052,
    n1051
  );


  and
  g2491
  (
    n2535,
    n1053,
    n924,
    n2519
  );


  nor
  g2492
  (
    n2544,
    n2529,
    n2284,
    n2282,
    n2277
  );


  or
  g2493
  (
    n2537,
    n2536,
    n2286,
    n973,
    n2280
  );


  nor
  g2494
  (
    n2549,
    n2272,
    n2290,
    n2533,
    n2273
  );


  nand
  g2495
  (
    n2543,
    n2286,
    n2283,
    n2287,
    n2532
  );


  xnor
  g2496
  (
    n2552,
    n2394,
    n2281,
    n2397,
    n2534
  );


  or
  g2497
  (
    n2547,
    n2275,
    n2278,
    n2289,
    n2271
  );


  nor
  g2498
  (
    n2538,
    n2279,
    n2288,
    n2393,
    n2532
  );


  xnor
  g2499
  (
    n2539,
    n2281,
    n2276,
    n2535
  );


  xnor
  g2500
  (
    n2551,
    n2279,
    n2277,
    n973,
    n2534
  );


  or
  g2501
  (
    n2540,
    n2282,
    n2536,
    n2392,
    n2531
  );


  xor
  g2502
  (
    n2548,
    n2290,
    n2274,
    n2272,
    n2531
  );


  or
  g2503
  (
    n2546,
    n2284,
    n2396,
    n2280,
    n2530
  );


  nor
  g2504
  (
    n2542,
    n2289,
    n2288,
    n2395,
    n2287
  );


  nand
  g2505
  (
    n2541,
    n2285,
    n2529,
    n2273,
    n2274
  );


  nor
  g2506
  (
    n2545,
    n2285,
    n2271,
    n2275,
    n2278
  );


  nor
  g2507
  (
    n2550,
    n2530,
    n2533,
    n2283,
    n2535
  );


  xor
  g2508
  (
    n2576,
    n2446,
    n2540,
    n2544,
    n2452
  );


  xnor
  g2509
  (
    n2562,
    n2551,
    n2428,
    n2430,
    n2548
  );


  and
  g2510
  (
    n2573,
    n2418,
    n2444,
    n2542,
    n2420
  );


  xor
  g2511
  (
    n2559,
    n2539,
    n2404,
    n2552,
    n2448
  );


  and
  g2512
  (
    n2564,
    n2405,
    n2542,
    n2440,
    n2452
  );


  xor
  g2513
  (
    n2565,
    n2444,
    n2436,
    n2417,
    n2410
  );


  xnor
  g2514
  (
    n2556,
    n2451,
    n2412,
    n2422,
    n2450
  );


  xnor
  g2515
  (
    n2572,
    n2449,
    n2428,
    n2437,
    n2540
  );


  nor
  g2516
  (
    n2577,
    n2547,
    n2543,
    n2439,
    n2415
  );


  and
  g2517
  (
    n2580,
    n2401,
    n2430,
    n2431,
    n2451
  );


  nand
  g2518
  (
    n2583,
    n2445,
    n2550,
    n2426,
    n2425
  );


  or
  g2519
  (
    n2568,
    n2441,
    n2538,
    n2424,
    n2413
  );


  xnor
  g2520
  (
    n2579,
    n2450,
    n2408,
    n2411,
    n2399
  );


  and
  g2521
  (
    n2563,
    n2543,
    n2435,
    n2551,
    n2446
  );


  nor
  g2522
  (
    n2558,
    n2549,
    n2443,
    n2437,
    n2422
  );


  xnor
  g2523
  (
    n2554,
    n2416,
    n2546,
    n2442,
    n2420
  );


  and
  g2524
  (
    n2578,
    n2429,
    n2545,
    n2447,
    n2441
  );


  xnor
  g2525
  (
    n2553,
    n2439,
    n2541,
    n2539,
    n2424
  );


  or
  g2526
  (
    n2574,
    n2414,
    n2415,
    n2541,
    n2421
  );


  or
  g2527
  (
    n2582,
    n2445,
    n2426,
    n2416,
    n2425
  );


  and
  g2528
  (
    n2571,
    n2547,
    n2545,
    n2438,
    n2419
  );


  xor
  g2529
  (
    n2584,
    n2537,
    n2447,
    n2433,
    n2436
  );


  nand
  g2530
  (
    n2561,
    n2449,
    n2412,
    n2423,
    n2442
  );


  xnor
  g2531
  (
    n2581,
    n2548,
    n2431,
    n2413,
    n2427
  );


  nor
  g2532
  (
    n2566,
    n2421,
    n2432,
    n2418,
    n2414
  );


  xor
  g2533
  (
    n2567,
    n2538,
    n2409,
    n2448,
    n2433
  );


  nor
  g2534
  (
    n2560,
    n2423,
    n2427,
    n2440,
    n2398
  );


  xnor
  g2535
  (
    n2575,
    n2403,
    n2406,
    n2550,
    n2435
  );


  and
  g2536
  (
    n2557,
    n2419,
    n2549,
    n2546,
    n2417
  );


  xnor
  g2537
  (
    n2570,
    n2432,
    n2438,
    n2402,
    n2434
  );


  xnor
  g2538
  (
    n2569,
    n2434,
    n2544,
    n2552,
    n2537
  );


  and
  g2539
  (
    n2555,
    n2429,
    n2400,
    n2407,
    n2443
  );


  xnor
  KeyGate_0_0
  (
    n1143,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n824,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    KeyNOTWire_0_2,
    keyIn_0_2,
    KeyWire_0_2
  );


  not
  KeyNOTGate_0_2
  (
    n782,
    KeyNOTWire_0_2
  );


  xor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n399,
    KeyNOTWire_0_3
  );


  xor
  KeyGate_0_4
  (
    n1798,
    keyIn_0_4,
    KeyWire_0_4
  );


  xnor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n1419,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n1348,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n1692,
    keyIn_0_7,
    KeyWire_0_7
  );


  xor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n128,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n572,
    keyIn_0_9,
    KeyWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n799,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1008,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    KeyNOTWire_0_12,
    keyIn_0_12,
    KeyWire_0_12
  );


  not
  KeyNOTGate_0_12
  (
    n2071,
    KeyNOTWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n1982,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    KeyNOTWire_0_14,
    keyIn_0_14,
    KeyWire_0_14
  );


  not
  KeyNOTGate_0_14
  (
    n1679,
    KeyNOTWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n1010,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n2264,
    keyIn_0_16,
    KeyWire_0_16
  );


  xor
  KeyGate_0_17
  (
    n392,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    KeyNOTWire_0_18,
    keyIn_0_18,
    KeyWire_0_18
  );


  not
  KeyNOTGate_0_18
  (
    n768,
    KeyNOTWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n1676,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n805,
    keyIn_0_20,
    KeyWire_0_20
  );


  xnor
  KeyGate_0_21
  (
    KeyNOTWire_0_21,
    keyIn_0_21,
    KeyWire_0_21
  );


  not
  KeyNOTGate_0_21
  (
    n1981,
    KeyNOTWire_0_21
  );


  xnor
  KeyGate_0_22
  (
    n422,
    keyIn_0_22,
    KeyWire_0_22
  );


  xor
  KeyGate_0_23
  (
    KeyNOTWire_0_23,
    keyIn_0_23,
    KeyWire_0_23
  );


  not
  KeyNOTGate_0_23
  (
    n1733,
    KeyNOTWire_0_23
  );


  xor
  KeyGate_0_24
  (
    n1924,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    KeyNOTWire_0_25,
    keyIn_0_25,
    KeyWire_0_25
  );


  not
  KeyNOTGate_0_25
  (
    n610,
    KeyNOTWire_0_25
  );


  xor
  KeyGate_0_26
  (
    KeyNOTWire_0_26,
    keyIn_0_26,
    KeyWire_0_26
  );


  not
  KeyNOTGate_0_26
  (
    n63,
    KeyNOTWire_0_26
  );


  xor
  KeyGate_0_27
  (
    KeyNOTWire_0_27,
    keyIn_0_27,
    KeyWire_0_27
  );


  not
  KeyNOTGate_0_27
  (
    n1004,
    KeyNOTWire_0_27
  );


  xnor
  KeyGate_0_28
  (
    n1147,
    keyIn_0_28,
    KeyWire_0_28
  );


  xor
  KeyGate_0_29
  (
    KeyNOTWire_0_29,
    keyIn_0_29,
    KeyWire_0_29
  );


  not
  KeyNOTGate_0_29
  (
    n1864,
    KeyNOTWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    KeyNOTWire_0_30,
    keyIn_0_30,
    KeyWire_0_30
  );


  not
  KeyNOTGate_0_30
  (
    n738,
    KeyNOTWire_0_30
  );


  xor
  KeyGate_0_31
  (
    KeyNOTWire_0_31,
    keyIn_0_31,
    KeyWire_0_31
  );


  not
  KeyNOTGate_0_31
  (
    n1705,
    KeyNOTWire_0_31
  );


  xor
  KeyGate_0_32
  (
    n1917,
    keyIn_0_32,
    KeyWire_0_32
  );


  xnor
  KeyGate_0_33
  (
    KeyNOTWire_0_33,
    keyIn_0_33,
    KeyWire_0_33
  );


  not
  KeyNOTGate_0_33
  (
    n1247,
    KeyNOTWire_0_33
  );


  xor
  KeyGate_0_34
  (
    n59,
    keyIn_0_34,
    KeyWire_0_34
  );


  xnor
  KeyGate_0_35
  (
    n1091,
    keyIn_0_35,
    KeyWire_0_35
  );


  xor
  KeyGate_0_36
  (
    n1554,
    keyIn_0_36,
    KeyWire_0_36
  );


  xor
  KeyGate_0_37
  (
    n207,
    keyIn_0_37,
    KeyWire_0_37
  );


  xor
  KeyGate_0_38
  (
    KeyNOTWire_0_38,
    keyIn_0_38,
    KeyWire_0_38
  );


  not
  KeyNOTGate_0_38
  (
    n1115,
    KeyNOTWire_0_38
  );


  xor
  KeyGate_0_39
  (
    n70,
    keyIn_0_39,
    KeyWire_0_39
  );


  xnor
  KeyGate_0_40
  (
    n1301,
    keyIn_0_40,
    KeyWire_0_40
  );


  xor
  KeyGate_0_41
  (
    n375,
    keyIn_0_41,
    KeyWire_0_41
  );


  xor
  KeyGate_0_42
  (
    KeyNOTWire_0_42,
    keyIn_0_42,
    KeyWire_0_42
  );


  not
  KeyNOTGate_0_42
  (
    n1445,
    KeyNOTWire_0_42
  );


  xnor
  KeyGate_0_43
  (
    n1100,
    keyIn_0_43,
    KeyWire_0_43
  );


  xnor
  KeyGate_0_44
  (
    KeyNOTWire_0_44,
    keyIn_0_44,
    KeyWire_0_44
  );


  not
  KeyNOTGate_0_44
  (
    n2293,
    KeyNOTWire_0_44
  );


  xnor
  KeyGate_0_45
  (
    n1836,
    keyIn_0_45,
    KeyWire_0_45
  );


  xnor
  KeyGate_0_46
  (
    KeyNOTWire_0_46,
    keyIn_0_46,
    KeyWire_0_46
  );


  not
  KeyNOTGate_0_46
  (
    n2471,
    KeyNOTWire_0_46
  );


  xnor
  KeyGate_0_47
  (
    KeyNOTWire_0_47,
    keyIn_0_47,
    KeyWire_0_47
  );


  not
  KeyNOTGate_0_47
  (
    n1539,
    KeyNOTWire_0_47
  );


  xor
  KeyGate_0_48
  (
    KeyNOTWire_0_48,
    keyIn_0_48,
    KeyWire_0_48
  );


  not
  KeyNOTGate_0_48
  (
    n1704,
    KeyNOTWire_0_48
  );


  xnor
  KeyGate_0_49
  (
    n1613,
    keyIn_0_49,
    KeyWire_0_49
  );


  xor
  KeyGate_0_50
  (
    KeyNOTWire_0_50,
    keyIn_0_50,
    KeyWire_0_50
  );


  not
  KeyNOTGate_0_50
  (
    n723,
    KeyNOTWire_0_50
  );


  xnor
  KeyGate_0_51
  (
    n2004,
    keyIn_0_51,
    KeyWire_0_51
  );


  xnor
  KeyGate_0_52
  (
    KeyNOTWire_0_52,
    keyIn_0_52,
    KeyWire_0_52
  );


  not
  KeyNOTGate_0_52
  (
    n2005,
    KeyNOTWire_0_52
  );


  xor
  KeyGate_0_53
  (
    KeyNOTWire_0_53,
    keyIn_0_53,
    KeyWire_0_53
  );


  not
  KeyNOTGate_0_53
  (
    n1465,
    KeyNOTWire_0_53
  );


  xor
  KeyGate_0_54
  (
    n1698,
    keyIn_0_54,
    KeyWire_0_54
  );


  xnor
  KeyGate_0_55
  (
    n2023,
    keyIn_0_55,
    KeyWire_0_55
  );


  xnor
  KeyGate_0_56
  (
    KeyNOTWire_0_56,
    keyIn_0_56,
    KeyWire_0_56
  );


  not
  KeyNOTGate_0_56
  (
    n1542,
    KeyNOTWire_0_56
  );


  xor
  KeyGate_0_57
  (
    n1584,
    keyIn_0_57,
    KeyWire_0_57
  );


  xnor
  KeyGate_0_58
  (
    KeyNOTWire_0_58,
    keyIn_0_58,
    KeyWire_0_58
  );


  not
  KeyNOTGate_0_58
  (
    n1397,
    KeyNOTWire_0_58
  );


  xnor
  KeyGate_0_59
  (
    KeyNOTWire_0_59,
    keyIn_0_59,
    KeyWire_0_59
  );


  not
  KeyNOTGate_0_59
  (
    n1608,
    KeyNOTWire_0_59
  );


  xnor
  KeyGate_0_60
  (
    KeyNOTWire_0_60,
    keyIn_0_60,
    KeyWire_0_60
  );


  not
  KeyNOTGate_0_60
  (
    n975,
    KeyNOTWire_0_60
  );


  xor
  KeyGate_0_61
  (
    KeyNOTWire_0_61,
    keyIn_0_61,
    KeyWire_0_61
  );


  not
  KeyNOTGate_0_61
  (
    n499,
    KeyNOTWire_0_61
  );


  xor
  KeyGate_0_62
  (
    n964,
    keyIn_0_62,
    KeyWire_0_62
  );


  xor
  KeyGate_0_63
  (
    n840,
    keyIn_0_63,
    KeyWire_0_63
  );


endmodule

