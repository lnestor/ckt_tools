

module Stat_392_937
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n399,
  n403,
  n395,
  n396,
  n408,
  n397,
  n414,
  n405,
  n410,
  n398,
  n411,
  n413,
  n407,
  n400,
  n393,
  n409,
  n402,
  n415,
  n404,
  n401,
  n394,
  n412,
  n406
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n399;output n403;output n395;output n396;output n408;output n397;output n414;output n405;output n410;output n398;output n411;output n413;output n407;output n400;output n393;output n409;output n402;output n415;output n404;output n401;output n394;output n412;output n406;
  wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire KeyWire_0_0;wire KeyNOTWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyNOTWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyNOTWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyNOTWire_0_15;

  not
  g0
  (
    n24,
    n1
  );


  not
  g1
  (
    n37,
    n4
  );


  not
  g2
  (
    n29,
    n2
  );


  not
  g3
  (
    n33,
    n2
  );


  buf
  g4
  (
    n25,
    n1
  );


  not
  g5
  (
    n30,
    n1
  );


  not
  g6
  (
    n36,
    n3
  );


  not
  g7
  (
    n26,
    n3
  );


  not
  g8
  (
    n32,
    n2
  );


  buf
  g9
  (
    n35,
    n4
  );


  buf
  g10
  (
    n34,
    n1
  );


  buf
  g11
  (
    n31,
    n3
  );


  buf
  g12
  (
    n27,
    n2
  );


  not
  g13
  (
    n28,
    n3
  );


  not
  g14
  (
    n50,
    n24
  );


  buf
  g15
  (
    n41,
    n29
  );


  buf
  g16
  (
    n59,
    n28
  );


  buf
  g17
  (
    n55,
    n27
  );


  buf
  g18
  (
    n42,
    n26
  );


  buf
  g19
  (
    n43,
    n25
  );


  buf
  g20
  (
    n48,
    n26
  );


  not
  g21
  (
    n58,
    n24
  );


  buf
  g22
  (
    n52,
    n29
  );


  buf
  g23
  (
    n57,
    n27
  );


  buf
  g24
  (
    n39,
    n24
  );


  buf
  g25
  (
    n46,
    n27
  );


  not
  g26
  (
    n44,
    n25
  );


  buf
  g27
  (
    n40,
    n24
  );


  buf
  g28
  (
    n45,
    n30
  );


  not
  g29
  (
    n38,
    n27
  );


  not
  g30
  (
    n53,
    n26
  );


  buf
  g31
  (
    n60,
    n25
  );


  buf
  g32
  (
    n56,
    n28
  );


  buf
  g33
  (
    n51,
    n29
  );


  not
  g34
  (
    n54,
    n26
  );


  not
  g35
  (
    n47,
    n28
  );


  buf
  g36
  (
    n61,
    n28
  );


  not
  g37
  (
    n62,
    n25
  );


  not
  g38
  (
    n49,
    n29
  );


  not
  g39
  (
    n75,
    n39
  );


  buf
  g40
  (
    n68,
    n45
  );


  not
  g41
  (
    n83,
    n40
  );


  not
  g42
  (
    n78,
    n41
  );


  buf
  g43
  (
    n73,
    n42
  );


  buf
  g44
  (
    n79,
    n46
  );


  buf
  g45
  (
    n66,
    n39
  );


  buf
  g46
  (
    n65,
    n38
  );


  not
  g47
  (
    n80,
    n42
  );


  buf
  g48
  (
    n76,
    n48
  );


  not
  g49
  (
    n64,
    n47
  );


  not
  g50
  (
    n71,
    n46
  );


  buf
  g51
  (
    KeyWire_0_9,
    n45
  );


  not
  g52
  (
    n69,
    n43
  );


  not
  g53
  (
    n72,
    n43
  );


  buf
  g54
  (
    n70,
    n41
  );


  not
  g55
  (
    n82,
    n47
  );


  buf
  g56
  (
    n67,
    n44
  );


  buf
  g57
  (
    n74,
    n44
  );


  buf
  g58
  (
    n81,
    n48
  );


  not
  g59
  (
    n63,
    n40
  );


  buf
  g60
  (
    n105,
    n71
  );


  buf
  g61
  (
    n136,
    n63
  );


  not
  g62
  (
    n107,
    n70
  );


  buf
  g63
  (
    n93,
    n65
  );


  buf
  g64
  (
    KeyWire_0_8,
    n63
  );


  buf
  g65
  (
    n114,
    n75
  );


  not
  g66
  (
    n87,
    n76
  );


  buf
  g67
  (
    n96,
    n69
  );


  not
  g68
  (
    n89,
    n68
  );


  not
  g69
  (
    n110,
    n68
  );


  not
  g70
  (
    KeyWire_0_7,
    n71
  );


  not
  g71
  (
    n104,
    n74
  );


  not
  g72
  (
    n102,
    n64
  );


  not
  g73
  (
    n113,
    n65
  );


  buf
  g74
  (
    n116,
    n73
  );


  buf
  g75
  (
    n126,
    n66
  );


  not
  g76
  (
    n106,
    n67
  );


  not
  g77
  (
    n88,
    n70
  );


  buf
  g78
  (
    n123,
    n75
  );


  buf
  g79
  (
    n86,
    n70
  );


  buf
  g80
  (
    n98,
    n69
  );


  buf
  g81
  (
    n109,
    n74
  );


  not
  g82
  (
    n131,
    n69
  );


  buf
  g83
  (
    KeyWire_0_3,
    n66
  );


  not
  g84
  (
    n135,
    n75
  );


  not
  g85
  (
    n118,
    n63
  );


  not
  g86
  (
    n108,
    n72
  );


  buf
  g87
  (
    n115,
    n72
  );


  not
  g88
  (
    n85,
    n74
  );


  buf
  g89
  (
    n99,
    n74
  );


  not
  g90
  (
    n133,
    n64
  );


  not
  g91
  (
    n117,
    n63
  );


  not
  g92
  (
    n125,
    n76
  );


  not
  g93
  (
    n132,
    n72
  );


  buf
  g94
  (
    n122,
    n69
  );


  buf
  g95
  (
    n95,
    n72
  );


  not
  g96
  (
    n134,
    n73
  );


  buf
  g97
  (
    n121,
    n75
  );


  buf
  g98
  (
    n97,
    n67
  );


  not
  g99
  (
    n101,
    n70
  );


  not
  g100
  (
    n90,
    n71
  );


  buf
  g101
  (
    n103,
    n67
  );


  buf
  g102
  (
    n130,
    n76
  );


  not
  g103
  (
    n111,
    n68
  );


  buf
  g104
  (
    n139,
    n65
  );


  buf
  g105
  (
    n129,
    n67
  );


  not
  g106
  (
    n127,
    n73
  );


  not
  g107
  (
    n120,
    n71
  );


  buf
  g108
  (
    n84,
    n68
  );


  not
  g109
  (
    n92,
    n73
  );


  buf
  g110
  (
    n119,
    n66
  );


  not
  g111
  (
    n112,
    n66
  );


  not
  g112
  (
    n94,
    n76
  );


  not
  g113
  (
    n100,
    n65
  );


  not
  g114
  (
    n138,
    n64
  );


  buf
  g115
  (
    n124,
    n64
  );


  not
  g116
  (
    n199,
    n116
  );


  not
  g117
  (
    n183,
    n96
  );


  not
  g118
  (
    n181,
    n111
  );


  not
  g119
  (
    n155,
    n22
  );


  not
  g120
  (
    n141,
    n84
  );


  buf
  g121
  (
    n158,
    n125
  );


  buf
  g122
  (
    n178,
    n86
  );


  not
  g123
  (
    n184,
    n101
  );


  not
  g124
  (
    KeyWire_0_11,
    n5
  );


  not
  g125
  (
    n145,
    n112
  );


  not
  g126
  (
    n186,
    n100
  );


  buf
  g127
  (
    n177,
    n118
  );


  not
  g128
  (
    n148,
    n90
  );


  not
  g129
  (
    n195,
    n115
  );


  and
  g130
  (
    n176,
    n95,
    n112,
    n11,
    n86
  );


  nor
  g131
  (
    n206,
    n120,
    n22,
    n121,
    n92
  );


  nor
  g132
  (
    n157,
    n110,
    n116,
    n106,
    n92
  );


  xnor
  g133
  (
    n191,
    n84,
    n14,
    n113,
    n115
  );


  nor
  g134
  (
    n179,
    n85,
    n113,
    n104,
    n110
  );


  nor
  g135
  (
    n156,
    n12,
    n120,
    n18,
    n104
  );


  nor
  g136
  (
    n162,
    n115,
    n10,
    n12,
    n101
  );


  nand
  g137
  (
    n147,
    n119,
    n93,
    n90,
    n100
  );


  nand
  g138
  (
    n182,
    n102,
    n21,
    n119,
    n118
  );


  xnor
  g139
  (
    n154,
    n125,
    n114,
    n5,
    n97
  );


  xor
  g140
  (
    n149,
    n15,
    n113,
    n122,
    n21
  );


  nand
  g141
  (
    n205,
    n10,
    n12,
    n7,
    n95
  );


  xnor
  g142
  (
    KeyWire_0_5,
    n87,
    n10,
    n19,
    n14
  );


  xnor
  g143
  (
    n172,
    n98,
    n86,
    n18,
    n95
  );


  xnor
  g144
  (
    n152,
    n85,
    n102,
    n98,
    n124
  );


  or
  g145
  (
    n194,
    n93,
    n20,
    n13,
    n89
  );


  xnor
  g146
  (
    n207,
    n5,
    n94,
    n95,
    n86
  );


  nand
  g147
  (
    n203,
    n123,
    n14,
    n104,
    n119
  );


  xor
  g148
  (
    n165,
    n11,
    n122,
    n124,
    n109
  );


  xor
  g149
  (
    n200,
    n8,
    n104,
    n22,
    n93
  );


  nor
  g150
  (
    n174,
    n90,
    n119,
    n109,
    n107
  );


  nor
  g151
  (
    n167,
    n121,
    n85,
    n108,
    n4
  );


  xor
  g152
  (
    n202,
    n106,
    n102,
    n96,
    n89
  );


  or
  g153
  (
    n185,
    n6,
    n17,
    n124,
    n111
  );


  xnor
  g154
  (
    n159,
    n114,
    n102,
    n92,
    n108
  );


  or
  g155
  (
    n196,
    n121,
    n84,
    n93,
    n17
  );


  nor
  g156
  (
    n198,
    n21,
    n18,
    n94,
    n88
  );


  xor
  g157
  (
    KeyWire_0_13,
    n117,
    n112,
    n6,
    n22
  );


  nand
  g158
  (
    n146,
    n8,
    n88,
    n106,
    n107
  );


  nor
  g159
  (
    n144,
    n105,
    n96,
    n111,
    n13
  );


  xnor
  g160
  (
    n201,
    n88,
    n15,
    n87,
    n97
  );


  xor
  g161
  (
    n175,
    n113,
    n120,
    n122,
    n16
  );


  nand
  g162
  (
    n142,
    n108,
    n8,
    n7,
    n18
  );


  xnor
  g163
  (
    n153,
    n111,
    n94,
    n96,
    n91
  );


  and
  g164
  (
    n190,
    n13,
    n7,
    n100,
    n9
  );


  nor
  g165
  (
    n150,
    n84,
    n109,
    n6,
    n100
  );


  xnor
  g166
  (
    n197,
    n91,
    n5,
    n121,
    n17
  );


  and
  g167
  (
    n192,
    n123,
    n99,
    n98,
    n21
  );


  or
  g168
  (
    n168,
    n124,
    n15,
    n103,
    n90
  );


  nor
  g169
  (
    n204,
    n8,
    n108,
    n16,
    n103
  );


  and
  g170
  (
    n143,
    n15,
    n20,
    n13,
    n114
  );


  nand
  g171
  (
    n160,
    n20,
    n94,
    n19,
    n120
  );


  nand
  g172
  (
    n193,
    n91,
    n11,
    n110,
    n17
  );


  xor
  g173
  (
    n208,
    n122,
    n16,
    n106,
    n9
  );


  xnor
  g174
  (
    n189,
    n107,
    n97,
    n12,
    n89
  );


  nor
  g175
  (
    n166,
    n101,
    n99,
    n23,
    n16
  );


  or
  g176
  (
    n171,
    n117,
    n9,
    n116,
    n92
  );


  or
  g177
  (
    n161,
    n114,
    n123,
    n101,
    n105
  );


  and
  g178
  (
    n151,
    n19,
    n118,
    n105,
    n112
  );


  and
  g179
  (
    n163,
    n103,
    n118,
    n9,
    n14
  );


  nand
  g180
  (
    n209,
    n117,
    n116,
    n19,
    n87
  );


  xnor
  g181
  (
    n187,
    n110,
    n88,
    n91,
    n87
  );


  nor
  g182
  (
    n180,
    n10,
    n89,
    n7,
    n6
  );


  xnor
  g183
  (
    n170,
    n109,
    n23,
    n115,
    n117
  );


  or
  g184
  (
    n188,
    n11,
    n103,
    n99,
    n20
  );


  nor
  g185
  (
    n140,
    n98,
    n85,
    n97,
    n107
  );


  xor
  g186
  (
    n164,
    n105,
    n123,
    n4,
    n99
  );


  buf
  g187
  (
    n259,
    n162
  );


  not
  g188
  (
    n223,
    n158
  );


  buf
  g189
  (
    n219,
    n156
  );


  not
  g190
  (
    n231,
    n153
  );


  not
  g191
  (
    n220,
    n166
  );


  not
  g192
  (
    n255,
    n153
  );


  not
  g193
  (
    n243,
    n164
  );


  buf
  g194
  (
    n237,
    n156
  );


  not
  g195
  (
    n236,
    n165
  );


  not
  g196
  (
    n214,
    n151
  );


  not
  g197
  (
    n215,
    n163
  );


  not
  g198
  (
    n252,
    n144
  );


  buf
  g199
  (
    n249,
    n171
  );


  buf
  g200
  (
    n253,
    n174
  );


  buf
  g201
  (
    n212,
    n167
  );


  not
  g202
  (
    n230,
    n168
  );


  buf
  g203
  (
    KeyWire_0_2,
    n150
  );


  buf
  g204
  (
    n216,
    n172
  );


  buf
  g205
  (
    n261,
    n157
  );


  not
  g206
  (
    n222,
    n162
  );


  buf
  g207
  (
    n227,
    n152
  );


  not
  g208
  (
    n257,
    n164
  );


  not
  g209
  (
    KeyWire_0_12,
    n155
  );


  buf
  g210
  (
    n260,
    n166
  );


  buf
  g211
  (
    n244,
    n170
  );


  buf
  g212
  (
    n213,
    n168
  );


  buf
  g213
  (
    n238,
    n165
  );


  buf
  g214
  (
    n258,
    n163
  );


  not
  g215
  (
    n226,
    n167
  );


  not
  g216
  (
    n228,
    n150
  );


  not
  g217
  (
    n248,
    n157
  );


  not
  g218
  (
    n232,
    n161
  );


  buf
  g219
  (
    n239,
    n148
  );


  buf
  g220
  (
    n240,
    n155
  );


  buf
  g221
  (
    n224,
    n149
  );


  buf
  g222
  (
    n221,
    n154
  );


  buf
  g223
  (
    n241,
    n175
  );


  buf
  g224
  (
    n229,
    n151
  );


  not
  g225
  (
    n235,
    n175
  );


  not
  g226
  (
    n211,
    n170
  );


  buf
  g227
  (
    n246,
    n176
  );


  buf
  g228
  (
    n254,
    n141
  );


  buf
  g229
  (
    n217,
    n158
  );


  buf
  g230
  (
    n262,
    n143
  );


  buf
  g231
  (
    n247,
    n172
  );


  not
  g232
  (
    KeyWire_0_15,
    n173
  );


  not
  g233
  (
    n245,
    n146
  );


  buf
  g234
  (
    n242,
    n173
  );


  xnor
  g235
  (
    n233,
    n174,
    n159,
    n169,
    n161
  );


  xor
  g236
  (
    n218,
    n160,
    n149,
    n159,
    n169
  );


  and
  g237
  (
    n250,
    n160,
    n154,
    n147,
    n142
  );


  nor
  g238
  (
    n234,
    n145,
    n152,
    n140,
    n171
  );


  or
  g239
  (
    n315,
    n208,
    n202,
    n225,
    n199
  );


  nand
  g240
  (
    n299,
    n229,
    n227,
    n197,
    n177
  );


  and
  g241
  (
    n331,
    n204,
    n201,
    n254,
    n229
  );


  or
  g242
  (
    n302,
    n204,
    n240,
    n202,
    n255
  );


  nand
  g243
  (
    n274,
    n207,
    n260,
    n252,
    n190
  );


  nand
  g244
  (
    n319,
    n218,
    n230,
    n236,
    n256
  );


  nor
  g245
  (
    n291,
    n183,
    n241,
    n255,
    n246
  );


  nor
  g246
  (
    n306,
    n199,
    n215,
    n252,
    n253
  );


  xor
  g247
  (
    n280,
    n194,
    n206,
    n259,
    n180
  );


  or
  g248
  (
    n344,
    n33,
    n182,
    n200,
    n219
  );


  and
  g249
  (
    n263,
    n228,
    n185,
    n243,
    n180
  );


  nand
  g250
  (
    n296,
    n254,
    n254,
    n49,
    n196
  );


  or
  g251
  (
    n316,
    n225,
    n258,
    n213,
    n256
  );


  nor
  g252
  (
    n339,
    n203,
    n58,
    n222,
    n259
  );


  xor
  g253
  (
    n286,
    n235,
    n217,
    n176,
    n224
  );


  nand
  g254
  (
    n295,
    n230,
    n233,
    n262,
    n208
  );


  xor
  g255
  (
    n334,
    n223,
    n216,
    n183,
    n227
  );


  xnor
  g256
  (
    n325,
    n209,
    n210,
    n187,
    n217
  );


  or
  g257
  (
    n345,
    n247,
    n205,
    n34,
    n202
  );


  or
  g258
  (
    n271,
    n236,
    n52,
    n228,
    n50
  );


  nand
  g259
  (
    n355,
    n238,
    n185,
    n226,
    n178
  );


  xor
  g260
  (
    n288,
    n232,
    n57,
    n33,
    n240
  );


  nand
  g261
  (
    n273,
    n213,
    n216,
    n234,
    n30
  );


  nor
  g262
  (
    n303,
    n245,
    n178,
    n181,
    n220
  );


  nor
  g263
  (
    n323,
    n230,
    n195,
    n248,
    n228
  );


  nor
  g264
  (
    n298,
    n62,
    n246,
    n60,
    n204
  );


  xor
  g265
  (
    n264,
    n203,
    n221,
    n248,
    n179
  );


  xnor
  g266
  (
    n292,
    n196,
    n198,
    n257,
    n237
  );


  and
  g267
  (
    n324,
    n257,
    n195,
    n53,
    n238
  );


  xnor
  g268
  (
    n279,
    n211,
    n198,
    n53,
    n260
  );


  and
  g269
  (
    n352,
    n190,
    n198,
    n33,
    n32
  );


  xor
  g270
  (
    n276,
    n249,
    n258,
    n219,
    n177
  );


  xnor
  g271
  (
    n275,
    n251,
    n258,
    n32,
    n252
  );


  nand
  g272
  (
    n332,
    n193,
    n210,
    n239,
    n214
  );


  and
  g273
  (
    n343,
    n237,
    n193,
    n52,
    n31
  );


  xnor
  g274
  (
    n349,
    n199,
    n214,
    n207,
    n210
  );


  and
  g275
  (
    n267,
    n184,
    n259,
    n215,
    n261
  );


  nor
  g276
  (
    n317,
    n197,
    n30,
    n227,
    n242
  );


  or
  g277
  (
    KeyWire_0_0,
    n250,
    n222,
    n229,
    n232
  );


  xnor
  g278
  (
    n328,
    n59,
    n235,
    n221,
    n191
  );


  nor
  g279
  (
    n351,
    n187,
    n215,
    n186,
    n238
  );


  nand
  g280
  (
    n341,
    n54,
    n250,
    n242,
    n193
  );


  and
  g281
  (
    n300,
    n225,
    n247,
    n233,
    n198
  );


  and
  g282
  (
    n333,
    n219,
    n251,
    n246,
    n248
  );


  nand
  g283
  (
    n304,
    n245,
    n243,
    n261,
    n31
  );


  nor
  g284
  (
    n294,
    n182,
    n34,
    n197,
    n212
  );


  or
  g285
  (
    n322,
    n234,
    n236,
    n190,
    n215
  );


  nor
  g286
  (
    n283,
    n253,
    n35,
    n61,
    n216
  );


  or
  g287
  (
    n270,
    n184,
    n209,
    n260,
    n186
  );


  or
  g288
  (
    n312,
    n192,
    n234,
    n194,
    n23
  );


  nand
  g289
  (
    n301,
    n235,
    n207,
    n241,
    n210
  );


  xnor
  g290
  (
    n313,
    n254,
    n194,
    n196,
    n244
  );


  xor
  g291
  (
    KeyWire_0_6,
    n245,
    n230,
    n229,
    n255
  );


  xor
  g292
  (
    n284,
    n239,
    n214,
    n244,
    n192
  );


  and
  g293
  (
    n268,
    n257,
    n208,
    n255,
    n233
  );


  or
  g294
  (
    n307,
    n189,
    n189,
    n219,
    n221
  );


  nand
  g295
  (
    n277,
    n61,
    n227,
    n197,
    n261
  );


  xnor
  g296
  (
    n290,
    n231,
    n200,
    n220,
    n30
  );


  xnor
  g297
  (
    n348,
    n221,
    n202,
    n231,
    n56
  );


  xnor
  g298
  (
    n272,
    n32,
    n31,
    n238,
    n239
  );


  and
  g299
  (
    n326,
    n54,
    n223,
    n182,
    n257
  );


  nor
  g300
  (
    n356,
    n192,
    n256,
    n232,
    n199
  );


  nand
  g301
  (
    n338,
    n188,
    n249,
    n204,
    n245
  );


  nand
  g302
  (
    n309,
    n212,
    n201,
    n49,
    n250
  );


  xor
  g303
  (
    n269,
    n50,
    n212,
    n183,
    n251
  );


  xnor
  g304
  (
    n327,
    n185,
    n187,
    n188,
    n205
  );


  or
  g305
  (
    n311,
    n253,
    n222,
    n191,
    n205
  );


  and
  g306
  (
    n285,
    n218,
    n225,
    n224,
    n188
  );


  or
  g307
  (
    n308,
    n195,
    n243,
    n59,
    n248
  );


  and
  g308
  (
    n310,
    n240,
    n247,
    n193,
    n218
  );


  and
  g309
  (
    n337,
    n251,
    n182,
    n207,
    n208
  );


  nand
  g310
  (
    n318,
    n241,
    n226,
    n234,
    n224
  );


  and
  g311
  (
    n346,
    n31,
    n55,
    n214,
    n216
  );


  nor
  g312
  (
    n314,
    n223,
    n190,
    n256,
    n262
  );


  nand
  g313
  (
    n329,
    n247,
    n51,
    n60,
    n261
  );


  or
  g314
  (
    n297,
    n184,
    n262,
    n236,
    n200
  );


  xor
  g315
  (
    n320,
    n258,
    n181,
    n253,
    n239
  );


  and
  g316
  (
    KeyWire_0_10,
    n246,
    n189,
    n58,
    n213
  );


  xor
  g317
  (
    n350,
    n185,
    n220,
    n206,
    n188
  );


  xnor
  g318
  (
    n335,
    n206,
    n241,
    n209,
    n203
  );


  and
  g319
  (
    n357,
    n194,
    n212,
    n237,
    n235
  );


  nor
  g320
  (
    KeyWire_0_14,
    n183,
    n217,
    n213
  );


  xnor
  g321
  (
    n266,
    n203,
    n243,
    n201,
    n244
  );


  and
  g322
  (
    n293,
    n262,
    n226,
    n55,
    n231
  );


  nor
  g323
  (
    n358,
    n201,
    n249,
    n244,
    n224
  );


  nor
  g324
  (
    n282,
    n191,
    n220,
    n249,
    n184
  );


  xnor
  g325
  (
    n336,
    n192,
    n260,
    n237,
    n196
  );


  xor
  g326
  (
    n265,
    n242,
    n223,
    n179,
    n189
  );


  nor
  g327
  (
    n281,
    n259,
    n205,
    n51,
    n186
  );


  and
  g328
  (
    n330,
    n57,
    n56,
    n250,
    n195
  );


  nor
  g329
  (
    n340,
    n187,
    n206,
    n232,
    n222
  );


  and
  g330
  (
    n321,
    n209,
    n211,
    n33,
    n34
  );


  and
  g331
  (
    n354,
    n228,
    n181,
    n218,
    n32
  );


  or
  g332
  (
    n287,
    n252,
    n200,
    n233,
    n23
  );


  xor
  g333
  (
    n305,
    n242,
    n186,
    n191,
    n240
  );


  nand
  g334
  (
    n289,
    n181,
    n231,
    n34,
    n226
  );


  nor
  g335
  (
    n380,
    n355,
    n340,
    n290,
    n62
  );


  nand
  g336
  (
    n373,
    n281,
    n83,
    n351,
    n36
  );


  or
  g337
  (
    n364,
    n343,
    n319,
    n317,
    n35
  );


  nor
  g338
  (
    n377,
    n273,
    n282,
    n287,
    n35
  );


  xor
  g339
  (
    n367,
    n350,
    n323,
    n306,
    n81
  );


  xor
  g340
  (
    n387,
    n325,
    n302,
    n283,
    n295
  );


  nand
  g341
  (
    n362,
    n298,
    n313,
    n336,
    n288
  );


  xnor
  g342
  (
    n389,
    n324,
    n307,
    n81,
    n82
  );


  or
  g343
  (
    n375,
    n80,
    n83,
    n267,
    n345
  );


  nor
  g344
  (
    n392,
    n321,
    n37,
    n286,
    n263
  );


  xnor
  g345
  (
    n388,
    n80,
    n320,
    n266,
    n277
  );


  nand
  g346
  (
    n383,
    n356,
    n301,
    n357,
    n82
  );


  xor
  g347
  (
    n363,
    n352,
    n304,
    n312,
    n293
  );


  nor
  g348
  (
    n365,
    n272,
    n36,
    n309,
    n78
  );


  xor
  g349
  (
    n374,
    n82,
    n81,
    n303,
    n326
  );


  and
  g350
  (
    n390,
    n308,
    n331,
    n83,
    n285
  );


  xnor
  g351
  (
    n384,
    n289,
    n344,
    n314,
    n341
  );


  nor
  g352
  (
    n391,
    n280,
    n354,
    n318,
    n347
  );


  and
  g353
  (
    n376,
    n316,
    n268,
    n78,
    n264
  );


  or
  g354
  (
    n368,
    n77,
    n333,
    n353,
    n327
  );


  and
  g355
  (
    n359,
    n346,
    n77,
    n274,
    n35
  );


  xor
  g356
  (
    n360,
    n37,
    n339,
    n292,
    n80
  );


  nand
  g357
  (
    n382,
    n335,
    n279,
    n77,
    n278
  );


  nand
  g358
  (
    n371,
    n83,
    n322,
    n358,
    n79
  );


  nand
  g359
  (
    n370,
    n79,
    n37,
    n299,
    n82
  );


  xnor
  g360
  (
    n372,
    n300,
    n276,
    n37,
    n275
  );


  or
  g361
  (
    n385,
    n349,
    n310,
    n315,
    n338
  );


  xor
  g362
  (
    n379,
    n328,
    n305,
    n79,
    n78
  );


  and
  g363
  (
    n381,
    n296,
    n79,
    n311,
    n80
  );


  nand
  g364
  (
    n369,
    n297,
    n36,
    n77,
    n348
  );


  nor
  g365
  (
    n366,
    n337,
    n294,
    n270,
    n265
  );


  or
  g366
  (
    KeyWire_0_4,
    n269,
    n291,
    n81,
    n334
  );


  or
  g367
  (
    n386,
    n332,
    n78,
    n36,
    n271
  );


  and
  g368
  (
    n378,
    n342,
    n330,
    n284,
    n329
  );


  and
  g369
  (
    n411,
    n129,
    n132,
    n374
  );


  nor
  g370
  (
    n399,
    n377,
    n133,
    n130,
    n135
  );


  xnor
  g371
  (
    n415,
    n371,
    n130,
    n135,
    n139
  );


  or
  g372
  (
    n397,
    n128,
    n131,
    n137
  );


  nor
  g373
  (
    n414,
    n135,
    n375,
    n360,
    n385
  );


  or
  g374
  (
    n405,
    n128,
    n128,
    n138,
    n129
  );


  xnor
  g375
  (
    n398,
    n132,
    n362,
    n134,
    n126
  );


  nor
  g376
  (
    KeyWire_0_1,
    n384,
    n380,
    n369,
    n129
  );


  nand
  g377
  (
    n401,
    n364,
    n390,
    n135,
    n139
  );


  nand
  g378
  (
    n407,
    n359,
    n368,
    n125,
    n131
  );


  nand
  g379
  (
    n400,
    n125,
    n373,
    n131,
    n138
  );


  or
  g380
  (
    n394,
    n379,
    n386,
    n365,
    n367
  );


  xor
  g381
  (
    n413,
    n134,
    n137,
    n361,
    n139
  );


  xnor
  g382
  (
    n403,
    n127,
    n370,
    n388,
    n392
  );


  or
  g383
  (
    n406,
    n139,
    n126,
    n382,
    n137
  );


  nor
  g384
  (
    n409,
    n391,
    n133,
    n387,
    n372
  );


  xnor
  g385
  (
    n410,
    n126,
    n127,
    n133,
    n130
  );


  xnor
  g386
  (
    n395,
    n136,
    n378,
    n130,
    n138
  );


  xor
  g387
  (
    n412,
    n389,
    n134,
    n127
  );


  and
  g388
  (
    n393,
    n366,
    n128,
    n127,
    n136
  );


  nand
  g389
  (
    n402,
    n126,
    n133,
    n137,
    n138
  );


  xor
  g390
  (
    n404,
    n383,
    n132,
    n363,
    n136
  );


  xor
  g391
  (
    n396,
    n376,
    n129,
    n381,
    n136
  );


  xor
  KeyGate_0_0
  (
    KeyNOTWire_0_0,
    keyIn_0_0,
    KeyWire_0_0
  );


  not
  KeyNOTGate_0_0
  (
    n353,
    KeyNOTWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n408,
    keyIn_0_1,
    KeyWire_0_1
  );


  xnor
  KeyGate_0_2
  (
    n225,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    KeyNOTWire_0_3,
    keyIn_0_3,
    KeyWire_0_3
  );


  not
  KeyNOTGate_0_3
  (
    n128,
    KeyNOTWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n361,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    KeyNOTWire_0_5,
    keyIn_0_5,
    KeyWire_0_5
  );


  not
  KeyNOTGate_0_5
  (
    n173,
    KeyNOTWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n342,
    keyIn_0_6,
    KeyWire_0_6
  );


  xor
  KeyGate_0_7
  (
    n137,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n91,
    KeyNOTWire_0_8
  );


  xor
  KeyGate_0_9
  (
    n77,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n278,
    KeyNOTWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n210,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n256,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n169,
    KeyNOTWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n347,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    KeyNOTWire_0_15,
    keyIn_0_15,
    KeyWire_0_15
  );


  not
  KeyNOTGate_0_15
  (
    n251,
    KeyNOTWire_0_15
  );


endmodule


