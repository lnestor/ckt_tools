

module Stat_3000_326
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n22,
  n23,
  n24,
  n25,
  n26,
  n27,
  n28,
  n29,
  n30,
  n31,
  n32,
  n2795,
  n2851,
  n2849,
  n2847,
  n2848,
  n2852,
  n2846,
  n2844,
  n2845,
  n3028,
  n3013,
  n3029,
  n3019,
  n3011,
  n3015,
  n3022,
  n3032,
  n3023,
  n3026,
  n3010,
  n3031,
  n3012,
  n3014,
  n3021,
  n3024,
  n3017,
  n3018,
  n3025,
  n3020,
  n3016,
  n3030,
  n3027
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input n22;input n23;input n24;input n25;input n26;input n27;input n28;input n29;input n30;input n31;input n32;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;
  output n2795;output n2851;output n2849;output n2847;output n2848;output n2852;output n2846;output n2844;output n2845;output n3028;output n3013;output n3029;output n3019;output n3011;output n3015;output n3022;output n3032;output n3023;output n3026;output n3010;output n3031;output n3012;output n3014;output n3021;output n3024;output n3017;output n3018;output n3025;output n3020;output n3016;output n3030;output n3027;
  wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1763;wire n1764;wire n1765;wire n1766;wire n1767;wire n1768;wire n1769;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1829;wire n1830;wire n1831;wire n1832;wire n1833;wire n1834;wire n1835;wire n1836;wire n1837;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1861;wire n1862;wire n1863;wire n1864;wire n1865;wire n1866;wire n1867;wire n1868;wire n1869;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire n1878;wire n1879;wire n1880;wire n1881;wire n1882;wire n1883;wire n1884;wire n1885;wire n1886;wire n1887;wire n1888;wire n1889;wire n1890;wire n1891;wire n1892;wire n1893;wire n1894;wire n1895;wire n1896;wire n1897;wire n1898;wire n1899;wire n1900;wire n1901;wire n1902;wire n1903;wire n1904;wire n1905;wire n1906;wire n1907;wire n1908;wire n1909;wire n1910;wire n1911;wire n1912;wire n1913;wire n1914;wire n1915;wire n1916;wire n1917;wire n1918;wire n1919;wire n1920;wire n1921;wire n1922;wire n1923;wire n1924;wire n1925;wire n1926;wire n1927;wire n1928;wire n1929;wire n1930;wire n1931;wire n1932;wire n1933;wire n1934;wire n1935;wire n1936;wire n1937;wire n1938;wire n1939;wire n1940;wire n1941;wire n1942;wire n1943;wire n1944;wire n1945;wire n1946;wire n1947;wire n1948;wire n1949;wire n1950;wire n1951;wire n1952;wire n1953;wire n1954;wire n1955;wire n1956;wire n1957;wire n1958;wire n1959;wire n1960;wire n1961;wire n1962;wire n1963;wire n1964;wire n1965;wire n1966;wire n1967;wire n1968;wire n1969;wire n1970;wire n1971;wire n1972;wire n1973;wire n1974;wire n1975;wire n1976;wire n1977;wire n1978;wire n1979;wire n1980;wire n1981;wire n1982;wire n1983;wire n1984;wire n1985;wire n1986;wire n1987;wire n1988;wire n1989;wire n1990;wire n1991;wire n1992;wire n1993;wire n1994;wire n1995;wire n1996;wire n1997;wire n1998;wire n1999;wire n2000;wire n2001;wire n2002;wire n2003;wire n2004;wire n2005;wire n2006;wire n2007;wire n2008;wire n2009;wire n2010;wire n2011;wire n2012;wire n2013;wire n2014;wire n2015;wire n2016;wire n2017;wire n2018;wire n2019;wire n2020;wire n2021;wire n2022;wire n2023;wire n2024;wire n2025;wire n2026;wire n2027;wire n2028;wire n2029;wire n2030;wire n2031;wire n2032;wire n2033;wire n2034;wire n2035;wire n2036;wire n2037;wire n2038;wire n2039;wire n2040;wire n2041;wire n2042;wire n2043;wire n2044;wire n2045;wire n2046;wire n2047;wire n2048;wire n2049;wire n2050;wire n2051;wire n2052;wire n2053;wire n2054;wire n2055;wire n2056;wire n2057;wire n2058;wire n2059;wire n2060;wire n2061;wire n2062;wire n2063;wire n2064;wire n2065;wire n2066;wire n2067;wire n2068;wire n2069;wire n2070;wire n2071;wire n2072;wire n2073;wire n2074;wire n2075;wire n2076;wire n2077;wire n2078;wire n2079;wire n2080;wire n2081;wire n2082;wire n2083;wire n2084;wire n2085;wire n2086;wire n2087;wire n2088;wire n2089;wire n2090;wire n2091;wire n2092;wire n2093;wire n2094;wire n2095;wire n2096;wire n2097;wire n2098;wire n2099;wire n2100;wire n2101;wire n2102;wire n2103;wire n2104;wire n2105;wire n2106;wire n2107;wire n2108;wire n2109;wire n2110;wire n2111;wire n2112;wire n2113;wire n2114;wire n2115;wire n2116;wire n2117;wire n2118;wire n2119;wire n2120;wire n2121;wire n2122;wire n2123;wire n2124;wire n2125;wire n2126;wire n2127;wire n2128;wire n2129;wire n2130;wire n2131;wire n2132;wire n2133;wire n2134;wire n2135;wire n2136;wire n2137;wire n2138;wire n2139;wire n2140;wire n2141;wire n2142;wire n2143;wire n2144;wire n2145;wire n2146;wire n2147;wire n2148;wire n2149;wire n2150;wire n2151;wire n2152;wire n2153;wire n2154;wire n2155;wire n2156;wire n2157;wire n2158;wire n2159;wire n2160;wire n2161;wire n2162;wire n2163;wire n2164;wire n2165;wire n2166;wire n2167;wire n2168;wire n2169;wire n2170;wire n2171;wire n2172;wire n2173;wire n2174;wire n2175;wire n2176;wire n2177;wire n2178;wire n2179;wire n2180;wire n2181;wire n2182;wire n2183;wire n2184;wire n2185;wire n2186;wire n2187;wire n2188;wire n2189;wire n2190;wire n2191;wire n2192;wire n2193;wire n2194;wire n2195;wire n2196;wire n2197;wire n2198;wire n2199;wire n2200;wire n2201;wire n2202;wire n2203;wire n2204;wire n2205;wire n2206;wire n2207;wire n2208;wire n2209;wire n2210;wire n2211;wire n2212;wire n2213;wire n2214;wire n2215;wire n2216;wire n2217;wire n2218;wire n2219;wire n2220;wire n2221;wire n2222;wire n2223;wire n2224;wire n2225;wire n2226;wire n2227;wire n2228;wire n2229;wire n2230;wire n2231;wire n2232;wire n2233;wire n2234;wire n2235;wire n2236;wire n2237;wire n2238;wire n2239;wire n2240;wire n2241;wire n2242;wire n2243;wire n2244;wire n2245;wire n2246;wire n2247;wire n2248;wire n2249;wire n2250;wire n2251;wire n2252;wire n2253;wire n2254;wire n2255;wire n2256;wire n2257;wire n2258;wire n2259;wire n2260;wire n2261;wire n2262;wire n2263;wire n2264;wire n2265;wire n2266;wire n2267;wire n2268;wire n2269;wire n2270;wire n2271;wire n2272;wire n2273;wire n2274;wire n2275;wire n2276;wire n2277;wire n2278;wire n2279;wire n2280;wire n2281;wire n2282;wire n2283;wire n2284;wire n2285;wire n2286;wire n2287;wire n2288;wire n2289;wire n2290;wire n2291;wire n2292;wire n2293;wire n2294;wire n2295;wire n2296;wire n2297;wire n2298;wire n2299;wire n2300;wire n2301;wire n2302;wire n2303;wire n2304;wire n2305;wire n2306;wire n2307;wire n2308;wire n2309;wire n2310;wire n2311;wire n2312;wire n2313;wire n2314;wire n2315;wire n2316;wire n2317;wire n2318;wire n2319;wire n2320;wire n2321;wire n2322;wire n2323;wire n2324;wire n2325;wire n2326;wire n2327;wire n2328;wire n2329;wire n2330;wire n2331;wire n2332;wire n2333;wire n2334;wire n2335;wire n2336;wire n2337;wire n2338;wire n2339;wire n2340;wire n2341;wire n2342;wire n2343;wire n2344;wire n2345;wire n2346;wire n2347;wire n2348;wire n2349;wire n2350;wire n2351;wire n2352;wire n2353;wire n2354;wire n2355;wire n2356;wire n2357;wire n2358;wire n2359;wire n2360;wire n2361;wire n2362;wire n2363;wire n2364;wire n2365;wire n2366;wire n2367;wire n2368;wire n2369;wire n2370;wire n2371;wire n2372;wire n2373;wire n2374;wire n2375;wire n2376;wire n2377;wire n2378;wire n2379;wire n2380;wire n2381;wire n2382;wire n2383;wire n2384;wire n2385;wire n2386;wire n2387;wire n2388;wire n2389;wire n2390;wire n2391;wire n2392;wire n2393;wire n2394;wire n2395;wire n2396;wire n2397;wire n2398;wire n2399;wire n2400;wire n2401;wire n2402;wire n2403;wire n2404;wire n2405;wire n2406;wire n2407;wire n2408;wire n2409;wire n2410;wire n2411;wire n2412;wire n2413;wire n2414;wire n2415;wire n2416;wire n2417;wire n2418;wire n2419;wire n2420;wire n2421;wire n2422;wire n2423;wire n2424;wire n2425;wire n2426;wire n2427;wire n2428;wire n2429;wire n2430;wire n2431;wire n2432;wire n2433;wire n2434;wire n2435;wire n2436;wire n2437;wire n2438;wire n2439;wire n2440;wire n2441;wire n2442;wire n2443;wire n2444;wire n2445;wire n2446;wire n2447;wire n2448;wire n2449;wire n2450;wire n2451;wire n2452;wire n2453;wire n2454;wire n2455;wire n2456;wire n2457;wire n2458;wire n2459;wire n2460;wire n2461;wire n2462;wire n2463;wire n2464;wire n2465;wire n2466;wire n2467;wire n2468;wire n2469;wire n2470;wire n2471;wire n2472;wire n2473;wire n2474;wire n2475;wire n2476;wire n2477;wire n2478;wire n2479;wire n2480;wire n2481;wire n2482;wire n2483;wire n2484;wire n2485;wire n2486;wire n2487;wire n2488;wire n2489;wire n2490;wire n2491;wire n2492;wire n2493;wire n2494;wire n2495;wire n2496;wire n2497;wire n2498;wire n2499;wire n2500;wire n2501;wire n2502;wire n2503;wire n2504;wire n2505;wire n2506;wire n2507;wire n2508;wire n2509;wire n2510;wire n2511;wire n2512;wire n2513;wire n2514;wire n2515;wire n2516;wire n2517;wire n2518;wire n2519;wire n2520;wire n2521;wire n2522;wire n2523;wire n2524;wire n2525;wire n2526;wire n2527;wire n2528;wire n2529;wire n2530;wire n2531;wire n2532;wire n2533;wire n2534;wire n2535;wire n2536;wire n2537;wire n2538;wire n2539;wire n2540;wire n2541;wire n2542;wire n2543;wire n2544;wire n2545;wire n2546;wire n2547;wire n2548;wire n2549;wire n2550;wire n2551;wire n2552;wire n2553;wire n2554;wire n2555;wire n2556;wire n2557;wire n2558;wire n2559;wire n2560;wire n2561;wire n2562;wire n2563;wire n2564;wire n2565;wire n2566;wire n2567;wire n2568;wire n2569;wire n2570;wire n2571;wire n2572;wire n2573;wire n2574;wire n2575;wire n2576;wire n2577;wire n2578;wire n2579;wire n2580;wire n2581;wire n2582;wire n2583;wire n2584;wire n2585;wire n2586;wire n2587;wire n2588;wire n2589;wire n2590;wire n2591;wire n2592;wire n2593;wire n2594;wire n2595;wire n2596;wire n2597;wire n2598;wire n2599;wire n2600;wire n2601;wire n2602;wire n2603;wire n2604;wire n2605;wire n2606;wire n2607;wire n2608;wire n2609;wire n2610;wire n2611;wire n2612;wire n2613;wire n2614;wire n2615;wire n2616;wire n2617;wire n2618;wire n2619;wire n2620;wire n2621;wire n2622;wire n2623;wire n2624;wire n2625;wire n2626;wire n2627;wire n2628;wire n2629;wire n2630;wire n2631;wire n2632;wire n2633;wire n2634;wire n2635;wire n2636;wire n2637;wire n2638;wire n2639;wire n2640;wire n2641;wire n2642;wire n2643;wire n2644;wire n2645;wire n2646;wire n2647;wire n2648;wire n2649;wire n2650;wire n2651;wire n2652;wire n2653;wire n2654;wire n2655;wire n2656;wire n2657;wire n2658;wire n2659;wire n2660;wire n2661;wire n2662;wire n2663;wire n2664;wire n2665;wire n2666;wire n2667;wire n2668;wire n2669;wire n2670;wire n2671;wire n2672;wire n2673;wire n2674;wire n2675;wire n2676;wire n2677;wire n2678;wire n2679;wire n2680;wire n2681;wire n2682;wire n2683;wire n2684;wire n2685;wire n2686;wire n2687;wire n2688;wire n2689;wire n2690;wire n2691;wire n2692;wire n2693;wire n2694;wire n2695;wire n2696;wire n2697;wire n2698;wire n2699;wire n2700;wire n2701;wire n2702;wire n2703;wire n2704;wire n2705;wire n2706;wire n2707;wire n2708;wire n2709;wire n2710;wire n2711;wire n2712;wire n2713;wire n2714;wire n2715;wire n2716;wire n2717;wire n2718;wire n2719;wire n2720;wire n2721;wire n2722;wire n2723;wire n2724;wire n2725;wire n2726;wire n2727;wire n2728;wire n2729;wire n2730;wire n2731;wire n2732;wire n2733;wire n2734;wire n2735;wire n2736;wire n2737;wire n2738;wire n2739;wire n2740;wire n2741;wire n2742;wire n2743;wire n2744;wire n2745;wire n2746;wire n2747;wire n2748;wire n2749;wire n2750;wire n2751;wire n2752;wire n2753;wire n2754;wire n2755;wire n2756;wire n2757;wire n2758;wire n2759;wire n2760;wire n2761;wire n2762;wire n2763;wire n2764;wire n2765;wire n2766;wire n2767;wire n2768;wire n2769;wire n2770;wire n2771;wire n2772;wire n2773;wire n2774;wire n2775;wire n2776;wire n2777;wire n2778;wire n2779;wire n2780;wire n2781;wire n2782;wire n2783;wire n2784;wire n2785;wire n2786;wire n2787;wire n2788;wire n2789;wire n2790;wire n2791;wire n2792;wire n2793;wire n2794;wire n2796;wire n2797;wire n2798;wire n2799;wire n2800;wire n2801;wire n2802;wire n2803;wire n2804;wire n2805;wire n2806;wire n2807;wire n2808;wire n2809;wire n2810;wire n2811;wire n2812;wire n2813;wire n2814;wire n2815;wire n2816;wire n2817;wire n2818;wire n2819;wire n2820;wire n2821;wire n2822;wire n2823;wire n2824;wire n2825;wire n2826;wire n2827;wire n2828;wire n2829;wire n2830;wire n2831;wire n2832;wire n2833;wire n2834;wire n2835;wire n2836;wire n2837;wire n2838;wire n2839;wire n2840;wire n2841;wire n2842;wire n2843;wire n2850;wire n2853;wire n2854;wire n2855;wire n2856;wire n2857;wire n2858;wire n2859;wire n2860;wire n2861;wire n2862;wire n2863;wire n2864;wire n2865;wire n2866;wire n2867;wire n2868;wire n2869;wire n2870;wire n2871;wire n2872;wire n2873;wire n2874;wire n2875;wire n2876;wire n2877;wire n2878;wire n2879;wire n2880;wire n2881;wire n2882;wire n2883;wire n2884;wire n2885;wire n2886;wire n2887;wire n2888;wire n2889;wire n2890;wire n2891;wire n2892;wire n2893;wire n2894;wire n2895;wire n2896;wire n2897;wire n2898;wire n2899;wire n2900;wire n2901;wire n2902;wire n2903;wire n2904;wire n2905;wire n2906;wire n2907;wire n2908;wire n2909;wire n2910;wire n2911;wire n2912;wire n2913;wire n2914;wire n2915;wire n2916;wire n2917;wire n2918;wire n2919;wire n2920;wire n2921;wire n2922;wire n2923;wire n2924;wire n2925;wire n2926;wire n2927;wire n2928;wire n2929;wire n2930;wire n2931;wire n2932;wire n2933;wire n2934;wire n2935;wire n2936;wire n2937;wire n2938;wire n2939;wire n2940;wire n2941;wire n2942;wire n2943;wire n2944;wire n2945;wire n2946;wire n2947;wire n2948;wire n2949;wire n2950;wire n2951;wire n2952;wire n2953;wire n2954;wire n2955;wire n2956;wire n2957;wire n2958;wire n2959;wire n2960;wire n2961;wire n2962;wire n2963;wire n2964;wire n2965;wire n2966;wire n2967;wire n2968;wire n2969;wire n2970;wire n2971;wire n2972;wire n2973;wire n2974;wire n2975;wire n2976;wire n2977;wire n2978;wire n2979;wire n2980;wire n2981;wire n2982;wire n2983;wire n2984;wire n2985;wire n2986;wire n2987;wire n2988;wire n2989;wire n2990;wire n2991;wire n2992;wire n2993;wire n2994;wire n2995;wire n2996;wire n2997;wire n2998;wire n2999;wire n3000;wire n3001;wire n3002;wire n3003;wire n3004;wire n3005;wire n3006;wire n3007;wire n3008;wire n3009;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyNOTWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyNOTWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyNOTWire_0_7;wire KeyWire_0_8;wire KeyNOTWire_0_8;wire KeyWire_0_9;wire KeyNOTWire_0_9;wire KeyWire_0_10;wire KeyNOTWire_0_10;wire KeyWire_0_11;wire KeyNOTWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyNOTWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;

  not
  g0
  (
    n79,
    n14
  );


  not
  g1
  (
    n156,
    n7
  );


  buf
  g2
  (
    n128,
    n12
  );


  not
  g3
  (
    n78,
    n3
  );


  buf
  g4
  (
    n139,
    n29
  );


  not
  g5
  (
    n53,
    n14
  );


  not
  g6
  (
    n132,
    n3
  );


  not
  g7
  (
    n35,
    n13
  );


  buf
  g8
  (
    n112,
    n5
  );


  not
  g9
  (
    n100,
    n19
  );


  not
  g10
  (
    n37,
    n25
  );


  not
  g11
  (
    n134,
    n22
  );


  buf
  g12
  (
    n107,
    n16
  );


  not
  g13
  (
    n65,
    n25
  );


  buf
  g14
  (
    n38,
    n27
  );


  not
  g15
  (
    n131,
    n24
  );


  not
  g16
  (
    n152,
    n15
  );


  not
  g17
  (
    n146,
    n10
  );


  not
  g18
  (
    n101,
    n10
  );


  buf
  g19
  (
    n59,
    n2
  );


  buf
  g20
  (
    n133,
    n25
  );


  not
  g21
  (
    n158,
    n26
  );


  buf
  g22
  (
    n102,
    n18
  );


  buf
  g23
  (
    n115,
    n29
  );


  not
  g24
  (
    n41,
    n26
  );


  not
  g25
  (
    n89,
    n23
  );


  not
  g26
  (
    n33,
    n28
  );


  buf
  g27
  (
    n140,
    n17
  );


  buf
  g28
  (
    n46,
    n30
  );


  not
  g29
  (
    n138,
    n15
  );


  buf
  g30
  (
    n88,
    n12
  );


  buf
  g31
  (
    n76,
    n15
  );


  buf
  g32
  (
    n135,
    n8
  );


  not
  g33
  (
    n141,
    n29
  );


  buf
  g34
  (
    n99,
    n30
  );


  not
  g35
  (
    n60,
    n9
  );


  buf
  g36
  (
    n98,
    n1
  );


  not
  g37
  (
    n54,
    n4
  );


  not
  g38
  (
    n155,
    n3
  );


  not
  g39
  (
    n147,
    n27
  );


  not
  g40
  (
    n149,
    n11
  );


  buf
  g41
  (
    n103,
    n23
  );


  not
  g42
  (
    n83,
    n26
  );


  buf
  g43
  (
    n67,
    n7
  );


  buf
  g44
  (
    n116,
    n1
  );


  buf
  g45
  (
    n34,
    n5
  );


  buf
  g46
  (
    n143,
    n6
  );


  buf
  g47
  (
    n86,
    n32
  );


  not
  g48
  (
    n127,
    n24
  );


  buf
  g49
  (
    n75,
    n20
  );


  buf
  g50
  (
    n63,
    n8
  );


  buf
  g51
  (
    n137,
    n30
  );


  not
  g52
  (
    n95,
    n5
  );


  buf
  g53
  (
    n104,
    n14
  );


  buf
  g54
  (
    n117,
    n4
  );


  not
  g55
  (
    n50,
    n25
  );


  buf
  g56
  (
    n96,
    n22
  );


  buf
  g57
  (
    n44,
    n12
  );


  not
  g58
  (
    n153,
    n4
  );


  not
  g59
  (
    n70,
    n10
  );


  not
  g60
  (
    n136,
    n9
  );


  buf
  g61
  (
    n81,
    n11
  );


  buf
  g62
  (
    n122,
    n14
  );


  not
  g63
  (
    n119,
    n21
  );


  buf
  g64
  (
    n142,
    n8
  );


  buf
  g65
  (
    n154,
    n28
  );


  buf
  g66
  (
    n123,
    n16
  );


  buf
  g67
  (
    n90,
    n11
  );


  not
  g68
  (
    n121,
    n8
  );


  not
  g69
  (
    n150,
    n19
  );


  buf
  g70
  (
    n159,
    n2
  );


  not
  g71
  (
    n97,
    n29
  );


  buf
  g72
  (
    n42,
    n17
  );


  not
  g73
  (
    n40,
    n21
  );


  not
  g74
  (
    n92,
    n24
  );


  not
  g75
  (
    n120,
    n30
  );


  buf
  g76
  (
    n52,
    n13
  );


  buf
  g77
  (
    n125,
    n22
  );


  not
  g78
  (
    n77,
    n19
  );


  not
  g79
  (
    n49,
    n17
  );


  not
  g80
  (
    n129,
    n13
  );


  buf
  g81
  (
    n57,
    n6
  );


  buf
  g82
  (
    n105,
    n28
  );


  buf
  g83
  (
    n61,
    n31
  );


  buf
  g84
  (
    n47,
    n2
  );


  not
  g85
  (
    n110,
    n20
  );


  not
  g86
  (
    n87,
    n31
  );


  buf
  g87
  (
    n85,
    n21
  );


  not
  g88
  (
    n151,
    n27
  );


  buf
  g89
  (
    n91,
    n1
  );


  not
  g90
  (
    n36,
    n24
  );


  not
  g91
  (
    n157,
    n32
  );


  not
  g92
  (
    n108,
    n9
  );


  buf
  g93
  (
    n145,
    n32
  );


  buf
  g94
  (
    n109,
    n7
  );


  buf
  g95
  (
    n160,
    n18
  );


  not
  g96
  (
    n51,
    n15
  );


  buf
  g97
  (
    n114,
    n5
  );


  not
  g98
  (
    n56,
    n6
  );


  not
  g99
  (
    n72,
    n23
  );


  buf
  g100
  (
    n94,
    n4
  );


  not
  g101
  (
    n71,
    n16
  );


  not
  g102
  (
    n73,
    n16
  );


  not
  g103
  (
    n39,
    n3
  );


  not
  g104
  (
    n66,
    n10
  );


  not
  g105
  (
    n82,
    n27
  );


  not
  g106
  (
    n144,
    n18
  );


  not
  g107
  (
    n58,
    n18
  );


  buf
  g108
  (
    n118,
    n20
  );


  not
  g109
  (
    n48,
    n22
  );


  not
  g110
  (
    n130,
    n28
  );


  not
  g111
  (
    n148,
    n26
  );


  not
  g112
  (
    n45,
    n11
  );


  buf
  g113
  (
    n68,
    n9
  );


  not
  g114
  (
    n80,
    n2
  );


  buf
  g115
  (
    n55,
    n23
  );


  not
  g116
  (
    n69,
    n17
  );


  not
  g117
  (
    n106,
    n20
  );


  not
  g118
  (
    n84,
    n6
  );


  not
  g119
  (
    n43,
    n1
  );


  not
  g120
  (
    n93,
    n31
  );


  buf
  g121
  (
    n124,
    n21
  );


  not
  g122
  (
    n74,
    n13
  );


  buf
  g123
  (
    n62,
    n32
  );


  buf
  g124
  (
    n113,
    n12
  );


  buf
  g125
  (
    n126,
    n19
  );


  buf
  g126
  (
    n111,
    n7
  );


  not
  g127
  (
    n64,
    n31
  );


  not
  g128
  (
    n535,
    n118
  );


  not
  g129
  (
    n589,
    n102
  );


  buf
  g130
  (
    n668,
    n117
  );


  not
  g131
  (
    n405,
    n38
  );


  buf
  g132
  (
    n232,
    n133
  );


  buf
  g133
  (
    n480,
    n55
  );


  buf
  g134
  (
    n427,
    n36
  );


  not
  g135
  (
    n521,
    n128
  );


  buf
  g136
  (
    n340,
    n64
  );


  not
  g137
  (
    n555,
    n70
  );


  not
  g138
  (
    n345,
    n122
  );


  not
  g139
  (
    n550,
    n142
  );


  buf
  g140
  (
    n182,
    n65
  );


  not
  g141
  (
    n625,
    n69
  );


  not
  g142
  (
    n635,
    n119
  );


  not
  g143
  (
    n397,
    n59
  );


  buf
  g144
  (
    n367,
    n93
  );


  not
  g145
  (
    n643,
    n97
  );


  buf
  g146
  (
    n177,
    n150
  );


  not
  g147
  (
    n473,
    n111
  );


  buf
  g148
  (
    n219,
    n152
  );


  not
  g149
  (
    n465,
    n88
  );


  not
  g150
  (
    n167,
    n53
  );


  not
  g151
  (
    n663,
    n81
  );


  not
  g152
  (
    n201,
    n43
  );


  buf
  g153
  (
    n343,
    n98
  );


  buf
  g154
  (
    n446,
    n150
  );


  buf
  g155
  (
    n517,
    n73
  );


  not
  g156
  (
    n544,
    n156
  );


  not
  g157
  (
    n303,
    n94
  );


  not
  g158
  (
    n672,
    n95
  );


  not
  g159
  (
    n531,
    n74
  );


  buf
  g160
  (
    n394,
    n157
  );


  buf
  g161
  (
    n618,
    n129
  );


  buf
  g162
  (
    n518,
    n137
  );


  not
  g163
  (
    n667,
    n58
  );


  not
  g164
  (
    n601,
    n133
  );


  not
  g165
  (
    n671,
    n119
  );


  buf
  g166
  (
    n223,
    n36
  );


  not
  g167
  (
    n417,
    n147
  );


  buf
  g168
  (
    n658,
    n141
  );


  buf
  g169
  (
    n291,
    n106
  );


  not
  g170
  (
    n273,
    n117
  );


  buf
  g171
  (
    n263,
    n90
  );


  buf
  g172
  (
    n504,
    n80
  );


  buf
  g173
  (
    n323,
    n53
  );


  not
  g174
  (
    n324,
    n116
  );


  not
  g175
  (
    n311,
    n101
  );


  not
  g176
  (
    n578,
    n117
  );


  buf
  g177
  (
    n486,
    n145
  );


  buf
  g178
  (
    n224,
    n33
  );


  not
  g179
  (
    n174,
    n115
  );


  buf
  g180
  (
    n363,
    n45
  );


  not
  g181
  (
    n186,
    n157
  );


  not
  g182
  (
    n422,
    n127
  );


  buf
  g183
  (
    n423,
    n97
  );


  buf
  g184
  (
    n470,
    n94
  );


  not
  g185
  (
    KeyWire_0_6,
    n78
  );


  not
  g186
  (
    n431,
    n48
  );


  not
  g187
  (
    n301,
    n120
  );


  buf
  g188
  (
    n294,
    n155
  );


  buf
  g189
  (
    n548,
    n84
  );


  not
  g190
  (
    n295,
    n41
  );


  buf
  g191
  (
    n662,
    n157
  );


  buf
  g192
  (
    n314,
    n138
  );


  not
  g193
  (
    n464,
    n87
  );


  not
  g194
  (
    n241,
    n74
  );


  not
  g195
  (
    n561,
    n132
  );


  buf
  g196
  (
    n488,
    n101
  );


  not
  g197
  (
    n510,
    n99
  );


  not
  g198
  (
    n451,
    n138
  );


  not
  g199
  (
    n288,
    n101
  );


  not
  g200
  (
    n297,
    n109
  );


  buf
  g201
  (
    n636,
    n159
  );


  not
  g202
  (
    n378,
    n39
  );


  buf
  g203
  (
    n437,
    n118
  );


  buf
  g204
  (
    n180,
    n150
  );


  buf
  g205
  (
    n655,
    n46
  );


  buf
  g206
  (
    n306,
    n98
  );


  buf
  g207
  (
    n347,
    n49
  );


  not
  g208
  (
    n577,
    n79
  );


  buf
  g209
  (
    n406,
    n136
  );


  not
  g210
  (
    n381,
    n81
  );


  buf
  g211
  (
    n315,
    n39
  );


  buf
  g212
  (
    n403,
    n124
  );


  not
  g213
  (
    n173,
    n72
  );


  not
  g214
  (
    n598,
    n143
  );


  buf
  g215
  (
    n370,
    n116
  );


  buf
  g216
  (
    n187,
    n81
  );


  not
  g217
  (
    n322,
    n124
  );


  not
  g218
  (
    n163,
    n128
  );


  buf
  g219
  (
    n565,
    n61
  );


  buf
  g220
  (
    n214,
    n49
  );


  not
  g221
  (
    n538,
    n46
  );


  buf
  g222
  (
    n243,
    n108
  );


  buf
  g223
  (
    n244,
    n54
  );


  not
  g224
  (
    n525,
    n50
  );


  not
  g225
  (
    n633,
    n33
  );


  buf
  g226
  (
    n176,
    n50
  );


  not
  g227
  (
    n559,
    n70
  );


  not
  g228
  (
    n246,
    n80
  );


  not
  g229
  (
    n260,
    n134
  );


  not
  g230
  (
    n566,
    n84
  );


  not
  g231
  (
    n429,
    n129
  );


  not
  g232
  (
    n569,
    n124
  );


  not
  g233
  (
    n387,
    n114
  );


  not
  g234
  (
    n179,
    n62
  );


  not
  g235
  (
    n513,
    n118
  );


  buf
  g236
  (
    n557,
    n153
  );


  not
  g237
  (
    n197,
    n112
  );


  not
  g238
  (
    n299,
    n46
  );


  not
  g239
  (
    n638,
    n154
  );


  not
  g240
  (
    n206,
    n69
  );


  not
  g241
  (
    n623,
    n90
  );


  buf
  g242
  (
    n271,
    n156
  );


  not
  g243
  (
    n484,
    n64
  );


  buf
  g244
  (
    n198,
    n143
  );


  not
  g245
  (
    n329,
    n102
  );


  not
  g246
  (
    n629,
    n37
  );


  buf
  g247
  (
    n462,
    n87
  );


  not
  g248
  (
    n424,
    n111
  );


  not
  g249
  (
    n584,
    n41
  );


  buf
  g250
  (
    n419,
    n82
  );


  not
  g251
  (
    n653,
    n71
  );


  buf
  g252
  (
    n659,
    n154
  );


  not
  g253
  (
    n649,
    n104
  );


  buf
  g254
  (
    n547,
    n135
  );


  buf
  g255
  (
    n570,
    n80
  );


  not
  g256
  (
    n384,
    n53
  );


  buf
  g257
  (
    n400,
    n70
  );


  not
  g258
  (
    n185,
    n139
  );


  not
  g259
  (
    n328,
    n92
  );


  not
  g260
  (
    n285,
    n121
  );


  not
  g261
  (
    n238,
    n106
  );


  buf
  g262
  (
    n240,
    n67
  );


  not
  g263
  (
    n287,
    n56
  );


  buf
  g264
  (
    n571,
    n151
  );


  buf
  g265
  (
    n597,
    n128
  );


  buf
  g266
  (
    n228,
    n96
  );


  not
  g267
  (
    n515,
    n87
  );


  not
  g268
  (
    n490,
    n44
  );


  not
  g269
  (
    n316,
    n57
  );


  buf
  g270
  (
    n546,
    n36
  );


  buf
  g271
  (
    n450,
    n94
  );


  buf
  g272
  (
    n594,
    n34
  );


  buf
  g273
  (
    n389,
    n89
  );


  not
  g274
  (
    n614,
    n85
  );


  not
  g275
  (
    n261,
    n107
  );


  buf
  g276
  (
    n596,
    n122
  );


  not
  g277
  (
    n600,
    n130
  );


  buf
  g278
  (
    n567,
    n146
  );


  not
  g279
  (
    n619,
    n146
  );


  not
  g280
  (
    n496,
    n88
  );


  buf
  g281
  (
    n218,
    n55
  );


  not
  g282
  (
    n505,
    n75
  );


  not
  g283
  (
    n642,
    n110
  );


  buf
  g284
  (
    n611,
    n84
  );


  not
  g285
  (
    n242,
    n113
  );


  not
  g286
  (
    n237,
    n63
  );


  not
  g287
  (
    n425,
    n126
  );


  buf
  g288
  (
    n568,
    n42
  );


  buf
  g289
  (
    n617,
    n104
  );


  not
  g290
  (
    n634,
    n132
  );


  not
  g291
  (
    n599,
    n91
  );


  buf
  g292
  (
    n469,
    n133
  );


  buf
  g293
  (
    n249,
    n113
  );


  not
  g294
  (
    n317,
    n140
  );


  buf
  g295
  (
    n660,
    n88
  );


  buf
  g296
  (
    n494,
    n40
  );


  not
  g297
  (
    n447,
    n151
  );


  buf
  g298
  (
    n239,
    n125
  );


  not
  g299
  (
    n284,
    n86
  );


  not
  g300
  (
    n277,
    n71
  );


  not
  g301
  (
    n349,
    n74
  );


  not
  g302
  (
    n575,
    n123
  );


  not
  g303
  (
    n326,
    n131
  );


  not
  g304
  (
    n579,
    n115
  );


  buf
  g305
  (
    n290,
    n48
  );


  buf
  g306
  (
    n292,
    n76
  );


  buf
  g307
  (
    n318,
    n156
  );


  not
  g308
  (
    n580,
    n135
  );


  not
  g309
  (
    n354,
    n82
  );


  buf
  g310
  (
    n353,
    n73
  );


  not
  g311
  (
    n651,
    n68
  );


  not
  g312
  (
    n592,
    n104
  );


  buf
  g313
  (
    n632,
    n78
  );


  not
  g314
  (
    n355,
    n148
  );


  buf
  g315
  (
    n573,
    n100
  );


  not
  g316
  (
    n443,
    n127
  );


  not
  g317
  (
    n361,
    n140
  );


  buf
  g318
  (
    n362,
    n158
  );


  buf
  g319
  (
    n615,
    n48
  );


  buf
  g320
  (
    n171,
    n52
  );


  buf
  g321
  (
    n452,
    n77
  );


  buf
  g322
  (
    n283,
    n67
  );


  not
  g323
  (
    n553,
    n68
  );


  not
  g324
  (
    n460,
    n60
  );


  not
  g325
  (
    n175,
    n63
  );


  buf
  g326
  (
    n613,
    n143
  );


  not
  g327
  (
    n269,
    n33
  );


  not
  g328
  (
    n657,
    n148
  );


  not
  g329
  (
    n491,
    n126
  );


  buf
  g330
  (
    n351,
    n56
  );


  not
  g331
  (
    n274,
    n66
  );


  buf
  g332
  (
    n390,
    n99
  );


  not
  g333
  (
    n170,
    n39
  );


  not
  g334
  (
    n270,
    n140
  );


  not
  g335
  (
    n670,
    n84
  );


  buf
  g336
  (
    n217,
    n103
  );


  buf
  g337
  (
    n254,
    n125
  );


  buf
  g338
  (
    n250,
    n123
  );


  buf
  g339
  (
    n514,
    n47
  );


  not
  g340
  (
    n500,
    n83
  );


  buf
  g341
  (
    n374,
    n74
  );


  not
  g342
  (
    n407,
    n155
  );


  buf
  g343
  (
    n162,
    n44
  );


  buf
  g344
  (
    n280,
    n79
  );


  buf
  g345
  (
    n428,
    n95
  );


  buf
  g346
  (
    n476,
    n116
  );


  buf
  g347
  (
    n524,
    n93
  );


  not
  g348
  (
    n449,
    n132
  );


  buf
  g349
  (
    n563,
    n63
  );


  not
  g350
  (
    n586,
    n58
  );


  buf
  g351
  (
    n554,
    n114
  );


  not
  g352
  (
    n661,
    n44
  );


  buf
  g353
  (
    n439,
    n130
  );


  not
  g354
  (
    n479,
    n88
  );


  not
  g355
  (
    n220,
    n54
  );


  buf
  g356
  (
    n430,
    n117
  );


  not
  g357
  (
    n233,
    n106
  );


  not
  g358
  (
    n607,
    n90
  );


  buf
  g359
  (
    n414,
    n149
  );


  buf
  g360
  (
    n627,
    n158
  );


  not
  g361
  (
    n388,
    n79
  );


  not
  g362
  (
    n421,
    n103
  );


  buf
  g363
  (
    n161,
    n109
  );


  buf
  g364
  (
    n166,
    n147
  );


  not
  g365
  (
    n365,
    n135
  );


  not
  g366
  (
    n172,
    n93
  );


  not
  g367
  (
    n435,
    n51
  );


  not
  g368
  (
    n252,
    n57
  );


  not
  g369
  (
    n485,
    n137
  );


  not
  g370
  (
    n341,
    n152
  );


  buf
  g371
  (
    n641,
    n151
  );


  buf
  g372
  (
    n195,
    n150
  );


  buf
  g373
  (
    n385,
    n40
  );


  not
  g374
  (
    n595,
    n59
  );


  buf
  g375
  (
    n231,
    n85
  );


  not
  g376
  (
    n247,
    n57
  );


  not
  g377
  (
    n475,
    n92
  );


  buf
  g378
  (
    n640,
    n91
  );


  buf
  g379
  (
    n646,
    n136
  );


  not
  g380
  (
    n539,
    n61
  );


  buf
  g381
  (
    n298,
    n37
  );


  buf
  g382
  (
    n213,
    n131
  );


  not
  g383
  (
    n506,
    n33
  );


  buf
  g384
  (
    n256,
    n121
  );


  buf
  g385
  (
    n380,
    n144
  );


  not
  g386
  (
    n621,
    n59
  );


  buf
  g387
  (
    n307,
    n34
  );


  not
  g388
  (
    n321,
    n34
  );


  buf
  g389
  (
    n320,
    n69
  );


  buf
  g390
  (
    n308,
    n81
  );


  buf
  g391
  (
    n281,
    n131
  );


  buf
  g392
  (
    n178,
    n110
  );


  buf
  g393
  (
    n227,
    n76
  );


  not
  g394
  (
    n393,
    n66
  );


  buf
  g395
  (
    n511,
    n132
  );


  not
  g396
  (
    n519,
    n145
  );


  not
  g397
  (
    n536,
    n160
  );


  not
  g398
  (
    n606,
    n110
  );


  buf
  g399
  (
    n296,
    n137
  );


  not
  g400
  (
    n204,
    n144
  );


  not
  g401
  (
    n262,
    n153
  );


  buf
  g402
  (
    n272,
    n42
  );


  buf
  g403
  (
    n327,
    n63
  );


  buf
  g404
  (
    n558,
    n152
  );


  not
  g405
  (
    n352,
    n97
  );


  buf
  g406
  (
    n276,
    n103
  );


  buf
  g407
  (
    n184,
    n138
  );


  buf
  g408
  (
    n540,
    n78
  );


  buf
  g409
  (
    n202,
    n159
  );


  buf
  g410
  (
    n528,
    n38
  );


  buf
  g411
  (
    n442,
    n35
  );


  buf
  g412
  (
    n650,
    n75
  );


  not
  g413
  (
    n501,
    n100
  );


  not
  g414
  (
    n616,
    n135
  );


  buf
  g415
  (
    n583,
    n82
  );


  buf
  g416
  (
    n604,
    n83
  );


  not
  g417
  (
    n537,
    n120
  );


  not
  g418
  (
    n368,
    n157
  );


  not
  g419
  (
    n289,
    n160
  );


  not
  g420
  (
    n523,
    n94
  );


  not
  g421
  (
    n412,
    n129
  );


  not
  g422
  (
    n286,
    n126
  );


  not
  g423
  (
    n235,
    n58
  );


  not
  g424
  (
    n582,
    n79
  );


  not
  g425
  (
    n502,
    n75
  );


  buf
  g426
  (
    n482,
    n136
  );


  not
  g427
  (
    n481,
    n156
  );


  not
  g428
  (
    n564,
    n102
  );


  buf
  g429
  (
    n631,
    n62
  );


  not
  g430
  (
    n265,
    n51
  );


  not
  g431
  (
    n401,
    n78
  );


  not
  g432
  (
    n225,
    n105
  );


  buf
  g433
  (
    n608,
    n95
  );


  not
  g434
  (
    n216,
    n41
  );


  buf
  g435
  (
    n507,
    n77
  );


  not
  g436
  (
    n335,
    n104
  );


  buf
  g437
  (
    n572,
    n52
  );


  buf
  g438
  (
    n612,
    n45
  );


  buf
  g439
  (
    n192,
    n61
  );


  buf
  g440
  (
    n226,
    n72
  );


  not
  g441
  (
    n207,
    n111
  );


  buf
  g442
  (
    n526,
    n34
  );


  not
  g443
  (
    n372,
    n124
  );


  not
  g444
  (
    n603,
    n37
  );


  not
  g445
  (
    n416,
    n42
  );


  not
  g446
  (
    n196,
    n101
  );


  not
  g447
  (
    n512,
    n52
  );


  buf
  g448
  (
    n645,
    n143
  );


  not
  g449
  (
    n312,
    n146
  );


  buf
  g450
  (
    n399,
    n43
  );


  not
  g451
  (
    n533,
    n148
  );


  not
  g452
  (
    n478,
    n116
  );


  buf
  g453
  (
    n477,
    n98
  );


  not
  g454
  (
    n605,
    n144
  );


  buf
  g455
  (
    n319,
    n141
  );


  not
  g456
  (
    n587,
    n115
  );


  buf
  g457
  (
    n602,
    n70
  );


  not
  g458
  (
    n221,
    n91
  );


  buf
  g459
  (
    n333,
    n160
  );


  buf
  g460
  (
    n455,
    n141
  );


  not
  g461
  (
    n356,
    n122
  );


  not
  g462
  (
    n665,
    n151
  );


  buf
  g463
  (
    n453,
    n122
  );


  buf
  g464
  (
    n331,
    n159
  );


  buf
  g465
  (
    n543,
    n58
  );


  buf
  g466
  (
    n245,
    n40
  );


  not
  g467
  (
    n551,
    n103
  );


  buf
  g468
  (
    n279,
    n50
  );


  buf
  g469
  (
    n278,
    n60
  );


  not
  g470
  (
    n357,
    n128
  );


  buf
  g471
  (
    n304,
    n67
  );


  buf
  g472
  (
    n541,
    n83
  );


  buf
  g473
  (
    n325,
    n118
  );


  buf
  g474
  (
    n574,
    n36
  );


  not
  g475
  (
    n209,
    n115
  );


  not
  g476
  (
    n330,
    n54
  );


  buf
  g477
  (
    n499,
    n153
  );


  not
  g478
  (
    n637,
    n55
  );


  not
  g479
  (
    n342,
    n134
  );


  not
  g480
  (
    n253,
    n148
  );


  not
  g481
  (
    n610,
    n57
  );


  not
  g482
  (
    n440,
    n96
  );


  not
  g483
  (
    n652,
    n147
  );


  not
  g484
  (
    n248,
    n97
  );


  buf
  g485
  (
    n386,
    n73
  );


  not
  g486
  (
    n310,
    n52
  );


  buf
  g487
  (
    n444,
    n160
  );


  buf
  g488
  (
    n305,
    n133
  );


  buf
  g489
  (
    n199,
    n73
  );


  not
  g490
  (
    n522,
    n62
  );


  not
  g491
  (
    n268,
    n91
  );


  buf
  g492
  (
    n588,
    n51
  );


  buf
  g493
  (
    n474,
    n43
  );


  buf
  g494
  (
    KeyWire_0_15,
    n144
  );


  buf
  g495
  (
    n593,
    n68
  );


  buf
  g496
  (
    n576,
    n85
  );


  buf
  g497
  (
    n483,
    n92
  );


  not
  g498
  (
    n251,
    n45
  );


  buf
  g499
  (
    n293,
    n140
  );


  not
  g500
  (
    n516,
    n105
  );


  not
  g501
  (
    n164,
    n86
  );


  not
  g502
  (
    n259,
    n112
  );


  not
  g503
  (
    n350,
    n76
  );


  not
  g504
  (
    n339,
    n64
  );


  not
  g505
  (
    n211,
    n45
  );


  not
  g506
  (
    n545,
    n93
  );


  buf
  g507
  (
    n445,
    n89
  );


  not
  g508
  (
    n609,
    n152
  );


  buf
  g509
  (
    n492,
    n39
  );


  not
  g510
  (
    n282,
    n51
  );


  not
  g511
  (
    n420,
    n38
  );


  buf
  g512
  (
    n591,
    n149
  );


  not
  g513
  (
    n337,
    n114
  );


  buf
  g514
  (
    n191,
    n35
  );


  buf
  g515
  (
    n626,
    n108
  );


  not
  g516
  (
    n458,
    n126
  );


  buf
  g517
  (
    n459,
    n158
  );


  buf
  g518
  (
    n257,
    n40
  );


  not
  g519
  (
    n183,
    n90
  );


  buf
  g520
  (
    n471,
    n96
  );


  buf
  g521
  (
    n630,
    n153
  );


  not
  g522
  (
    n426,
    n69
  );


  buf
  g523
  (
    n495,
    n119
  );


  buf
  g524
  (
    n433,
    n119
  );


  buf
  g525
  (
    n467,
    n139
  );


  buf
  g526
  (
    n549,
    n71
  );


  not
  g527
  (
    n472,
    n102
  );


  buf
  g528
  (
    n463,
    n123
  );


  not
  g529
  (
    n366,
    n120
  );


  buf
  g530
  (
    n382,
    n46
  );


  not
  g531
  (
    n654,
    n100
  );


  buf
  g532
  (
    n411,
    n92
  );


  buf
  g533
  (
    n520,
    n155
  );


  buf
  g534
  (
    n418,
    n61
  );


  buf
  g535
  (
    n267,
    n65
  );


  not
  g536
  (
    n364,
    n38
  );


  not
  g537
  (
    n181,
    n47
  );


  buf
  g538
  (
    n255,
    n130
  );


  not
  g539
  (
    n530,
    n139
  );


  buf
  g540
  (
    n360,
    n66
  );


  not
  g541
  (
    n487,
    n142
  );


  buf
  g542
  (
    n348,
    n77
  );


  not
  g543
  (
    n620,
    n158
  );


  buf
  g544
  (
    n664,
    n127
  );


  buf
  g545
  (
    n336,
    n109
  );


  not
  g546
  (
    n234,
    n83
  );


  buf
  g547
  (
    n377,
    n65
  );


  buf
  g548
  (
    KeyWire_0_7,
    n89
  );


  not
  g549
  (
    n169,
    n67
  );


  buf
  g550
  (
    n466,
    n134
  );


  not
  g551
  (
    n300,
    n138
  );


  not
  g552
  (
    KeyWire_0_0,
    n65
  );


  buf
  g553
  (
    n205,
    n60
  );


  buf
  g554
  (
    n552,
    n145
  );


  not
  g555
  (
    n168,
    n134
  );


  buf
  g556
  (
    n562,
    n49
  );


  buf
  g557
  (
    n628,
    n121
  );


  not
  g558
  (
    n236,
    n123
  );


  not
  g559
  (
    n489,
    n112
  );


  buf
  g560
  (
    n373,
    n131
  );


  buf
  g561
  (
    n408,
    n48
  );


  buf
  g562
  (
    n188,
    n76
  );


  not
  g563
  (
    n436,
    n106
  );


  not
  g564
  (
    n509,
    n130
  );


  buf
  g565
  (
    n529,
    n59
  );


  not
  g566
  (
    n590,
    n154
  );


  buf
  g567
  (
    n194,
    n86
  );


  not
  g568
  (
    n379,
    n56
  );


  buf
  g569
  (
    n457,
    n86
  );


  not
  g570
  (
    n493,
    n121
  );


  not
  g571
  (
    n338,
    n42
  );


  not
  g572
  (
    n454,
    n54
  );


  not
  g573
  (
    n193,
    n56
  );


  buf
  g574
  (
    n229,
    n105
  );


  not
  g575
  (
    n275,
    n82
  );


  buf
  g576
  (
    n391,
    n55
  );


  buf
  g577
  (
    n448,
    n125
  );


  buf
  g578
  (
    n332,
    n68
  );


  not
  g579
  (
    n415,
    n113
  );


  not
  g580
  (
    n190,
    n96
  );


  not
  g581
  (
    n556,
    n62
  );


  not
  g582
  (
    n375,
    n107
  );


  not
  g583
  (
    n302,
    n109
  );


  not
  g584
  (
    n508,
    n154
  );


  not
  g585
  (
    n497,
    n146
  );


  not
  g586
  (
    n230,
    n35
  );


  not
  g587
  (
    n434,
    n142
  );


  buf
  g588
  (
    n534,
    n149
  );


  not
  g589
  (
    n648,
    n136
  );


  not
  g590
  (
    n438,
    n99
  );


  not
  g591
  (
    n581,
    n141
  );


  buf
  g592
  (
    n503,
    n127
  );


  buf
  g593
  (
    n165,
    n107
  );


  buf
  g594
  (
    n369,
    n72
  );


  not
  g595
  (
    n441,
    n50
  );


  not
  g596
  (
    n542,
    n105
  );


  not
  g597
  (
    n266,
    n64
  );


  buf
  g598
  (
    n585,
    n47
  );


  buf
  g599
  (
    n264,
    n155
  );


  not
  g600
  (
    n200,
    n49
  );


  not
  g601
  (
    n258,
    n66
  );


  buf
  g602
  (
    n371,
    n98
  );


  not
  g603
  (
    n413,
    n99
  );


  not
  g604
  (
    n395,
    n147
  );


  buf
  g605
  (
    KeyWire_0_4,
    n72
  );


  not
  g606
  (
    n532,
    n41
  );


  buf
  g607
  (
    n644,
    n53
  );


  not
  g608
  (
    n309,
    n149
  );


  buf
  g609
  (
    n189,
    n95
  );


  buf
  g610
  (
    n432,
    n35
  );


  buf
  g611
  (
    n222,
    n43
  );


  buf
  g612
  (
    n210,
    n108
  );


  buf
  g613
  (
    n456,
    n114
  );


  not
  g614
  (
    n622,
    n44
  );


  not
  g615
  (
    n461,
    n111
  );


  buf
  g616
  (
    n468,
    n110
  );


  not
  g617
  (
    n313,
    n112
  );


  buf
  g618
  (
    n402,
    n85
  );


  not
  g619
  (
    n203,
    n159
  );


  buf
  g620
  (
    n359,
    n120
  );


  buf
  g621
  (
    n212,
    n100
  );


  not
  g622
  (
    n404,
    n137
  );


  not
  g623
  (
    n409,
    n71
  );


  buf
  g624
  (
    n208,
    n129
  );


  not
  g625
  (
    n215,
    n108
  );


  not
  g626
  (
    n656,
    n87
  );


  buf
  g627
  (
    n398,
    n77
  );


  buf
  g628
  (
    n647,
    n47
  );


  not
  g629
  (
    n346,
    n75
  );


  buf
  g630
  (
    n392,
    n89
  );


  not
  g631
  (
    n376,
    n80
  );


  not
  g632
  (
    n383,
    n142
  );


  buf
  g633
  (
    n666,
    n145
  );


  not
  g634
  (
    n344,
    n113
  );


  buf
  g635
  (
    n396,
    n125
  );


  not
  g636
  (
    n624,
    n107
  );


  not
  g637
  (
    KeyWire_0_10,
    n37
  );


  buf
  g638
  (
    n639,
    n139
  );


  not
  g639
  (
    n358,
    n60
  );


  not
  g640
  (
    n1258,
    n478
  );


  buf
  g641
  (
    n814,
    n231
  );


  not
  g642
  (
    n827,
    n445
  );


  not
  g643
  (
    n1145,
    n512
  );


  buf
  g644
  (
    n1452,
    n545
  );


  not
  g645
  (
    n1058,
    n404
  );


  buf
  g646
  (
    n1035,
    n325
  );


  not
  g647
  (
    n1338,
    n605
  );


  buf
  g648
  (
    n843,
    n450
  );


  not
  g649
  (
    n683,
    n210
  );


  not
  g650
  (
    n1050,
    n221
  );


  not
  g651
  (
    n1027,
    n491
  );


  buf
  g652
  (
    n1417,
    n650
  );


  not
  g653
  (
    n988,
    n267
  );


  not
  g654
  (
    n1101,
    n175
  );


  buf
  g655
  (
    n1365,
    n561
  );


  not
  g656
  (
    n1360,
    n645
  );


  not
  g657
  (
    n719,
    n419
  );


  not
  g658
  (
    n833,
    n291
  );


  not
  g659
  (
    n1203,
    n369
  );


  buf
  g660
  (
    n1356,
    n632
  );


  buf
  g661
  (
    n942,
    n495
  );


  buf
  g662
  (
    n1292,
    n331
  );


  buf
  g663
  (
    n806,
    n583
  );


  not
  g664
  (
    n1275,
    n550
  );


  buf
  g665
  (
    n849,
    n205
  );


  not
  g666
  (
    n1507,
    n261
  );


  buf
  g667
  (
    n766,
    n255
  );


  buf
  g668
  (
    KeyWire_0_13,
    n453
  );


  not
  g669
  (
    n983,
    n561
  );


  not
  g670
  (
    n1157,
    n372
  );


  buf
  g671
  (
    n899,
    n259
  );


  buf
  g672
  (
    n673,
    n283
  );


  buf
  g673
  (
    n1331,
    n339
  );


  not
  g674
  (
    n1450,
    n379
  );


  not
  g675
  (
    n1500,
    n292
  );


  buf
  g676
  (
    n742,
    n441
  );


  not
  g677
  (
    n1502,
    n547
  );


  buf
  g678
  (
    n1361,
    n268
  );


  not
  g679
  (
    n1043,
    n349
  );


  not
  g680
  (
    n1174,
    n496
  );


  not
  g681
  (
    n868,
    n234
  );


  not
  g682
  (
    n1152,
    n287
  );


  buf
  g683
  (
    n1374,
    n287
  );


  buf
  g684
  (
    n1086,
    n585
  );


  not
  g685
  (
    n1148,
    n405
  );


  buf
  g686
  (
    n1337,
    n525
  );


  not
  g687
  (
    n1104,
    n445
  );


  not
  g688
  (
    n961,
    n336
  );


  not
  g689
  (
    n944,
    n660
  );


  buf
  g690
  (
    n1391,
    n427
  );


  not
  g691
  (
    n1256,
    n199
  );


  not
  g692
  (
    n998,
    n406
  );


  buf
  g693
  (
    n694,
    n329
  );


  not
  g694
  (
    n720,
    n219
  );


  buf
  g695
  (
    n863,
    n338
  );


  not
  g696
  (
    n1363,
    n596
  );


  buf
  g697
  (
    n970,
    n394
  );


  not
  g698
  (
    n1321,
    n337
  );


  not
  g699
  (
    n731,
    n617
  );


  not
  g700
  (
    n1129,
    n383
  );


  not
  g701
  (
    n1436,
    n473
  );


  buf
  g702
  (
    n1113,
    n623
  );


  not
  g703
  (
    n1271,
    n339
  );


  buf
  g704
  (
    n1103,
    n620
  );


  buf
  g705
  (
    n1080,
    n538
  );


  buf
  g706
  (
    n1210,
    n290
  );


  buf
  g707
  (
    n1497,
    n659
  );


  buf
  g708
  (
    n755,
    n492
  );


  not
  g709
  (
    n1056,
    n255
  );


  not
  g710
  (
    n1480,
    n347
  );


  not
  g711
  (
    n1230,
    n524
  );


  buf
  g712
  (
    n1441,
    n665
  );


  buf
  g713
  (
    n1471,
    n243
  );


  not
  g714
  (
    n1438,
    n637
  );


  buf
  g715
  (
    n1389,
    n283
  );


  buf
  g716
  (
    n1161,
    n489
  );


  buf
  g717
  (
    n1309,
    n161
  );


  not
  g718
  (
    n1039,
    n640
  );


  not
  g719
  (
    n839,
    n369
  );


  buf
  g720
  (
    n947,
    n500
  );


  buf
  g721
  (
    n1037,
    n513
  );


  not
  g722
  (
    n1310,
    n417
  );


  buf
  g723
  (
    n1238,
    n395
  );


  not
  g724
  (
    n1327,
    n452
  );


  buf
  g725
  (
    n823,
    n225
  );


  buf
  g726
  (
    n1151,
    n433
  );


  not
  g727
  (
    n697,
    n437
  );


  buf
  g728
  (
    n785,
    n444
  );


  buf
  g729
  (
    n767,
    n461
  );


  not
  g730
  (
    n1070,
    n206
  );


  not
  g731
  (
    n920,
    n365
  );


  buf
  g732
  (
    n1162,
    n457
  );


  buf
  g733
  (
    n735,
    n341
  );


  buf
  g734
  (
    n1493,
    n402
  );


  buf
  g735
  (
    n1375,
    n385
  );


  buf
  g736
  (
    n1137,
    n627
  );


  buf
  g737
  (
    n780,
    n576
  );


  buf
  g738
  (
    n1269,
    n446
  );


  buf
  g739
  (
    n1277,
    n394
  );


  buf
  g740
  (
    n1454,
    n385
  );


  not
  g741
  (
    n1078,
    n531
  );


  buf
  g742
  (
    n993,
    n499
  );


  not
  g743
  (
    n852,
    n388
  );


  not
  g744
  (
    n812,
    n653
  );


  buf
  g745
  (
    n759,
    n434
  );


  buf
  g746
  (
    n1366,
    n212
  );


  not
  g747
  (
    n792,
    n252
  );


  buf
  g748
  (
    n1018,
    n536
  );


  buf
  g749
  (
    n1233,
    n628
  );


  not
  g750
  (
    n1353,
    n551
  );


  buf
  g751
  (
    n705,
    n197
  );


  buf
  g752
  (
    n957,
    n463
  );


  not
  g753
  (
    n674,
    n273
  );


  buf
  g754
  (
    n1390,
    n290
  );


  buf
  g755
  (
    n917,
    n323
  );


  buf
  g756
  (
    n1227,
    n332
  );


  buf
  g757
  (
    n765,
    n455
  );


  not
  g758
  (
    n739,
    n479
  );


  not
  g759
  (
    n1064,
    n218
  );


  not
  g760
  (
    n1220,
    n270
  );


  not
  g761
  (
    n885,
    n401
  );


  not
  g762
  (
    n1147,
    n648
  );


  buf
  g763
  (
    n1300,
    n511
  );


  buf
  g764
  (
    n994,
    n638
  );


  buf
  g765
  (
    n1046,
    n202
  );


  buf
  g766
  (
    n1117,
    n529
  );


  not
  g767
  (
    n699,
    n399
  );


  buf
  g768
  (
    n1213,
    n652
  );


  buf
  g769
  (
    n700,
    n244
  );


  not
  g770
  (
    n1424,
    n334
  );


  buf
  g771
  (
    n1205,
    n407
  );


  not
  g772
  (
    n1279,
    n546
  );


  buf
  g773
  (
    n1307,
    n578
  );


  not
  g774
  (
    n1301,
    n646
  );


  not
  g775
  (
    n789,
    n447
  );


  not
  g776
  (
    n1163,
    n534
  );


  not
  g777
  (
    n1000,
    n481
  );


  buf
  g778
  (
    n1431,
    n271
  );


  not
  g779
  (
    n1120,
    n585
  );


  not
  g780
  (
    n1044,
    n548
  );


  buf
  g781
  (
    n1215,
    n333
  );


  not
  g782
  (
    n1042,
    n280
  );


  buf
  g783
  (
    n986,
    n162
  );


  buf
  g784
  (
    n702,
    n667
  );


  buf
  g785
  (
    n684,
    n484
  );


  not
  g786
  (
    n955,
    n618
  );


  buf
  g787
  (
    n1426,
    n549
  );


  buf
  g788
  (
    n1180,
    n566
  );


  not
  g789
  (
    n1176,
    n608
  );


  buf
  g790
  (
    n1135,
    n253
  );


  not
  g791
  (
    n1296,
    n271
  );


  buf
  g792
  (
    n741,
    n224
  );


  buf
  g793
  (
    n1351,
    n371
  );


  buf
  g794
  (
    n1150,
    n528
  );


  not
  g795
  (
    n838,
    n396
  );


  buf
  g796
  (
    n1340,
    n164
  );


  buf
  g797
  (
    n1249,
    n555
  );


  buf
  g798
  (
    n1383,
    n293
  );


  buf
  g799
  (
    n1112,
    n318
  );


  not
  g800
  (
    n747,
    n288
  );


  buf
  g801
  (
    n732,
    n231
  );


  buf
  g802
  (
    n1384,
    n600
  );


  not
  g803
  (
    n1019,
    n439
  );


  buf
  g804
  (
    n875,
    n254
  );


  not
  g805
  (
    n1494,
    n174
  );


  buf
  g806
  (
    n1052,
    n595
  );


  not
  g807
  (
    n835,
    n588
  );


  not
  g808
  (
    n908,
    n276
  );


  not
  g809
  (
    n882,
    n381
  );


  not
  g810
  (
    n810,
    n561
  );


  buf
  g811
  (
    n748,
    n529
  );


  not
  g812
  (
    n1287,
    n233
  );


  not
  g813
  (
    n1388,
    n481
  );


  not
  g814
  (
    n1167,
    n568
  );


  not
  g815
  (
    n1010,
    n303
  );


  buf
  g816
  (
    n1187,
    n462
  );


  buf
  g817
  (
    n876,
    n652
  );


  buf
  g818
  (
    n715,
    n470
  );


  buf
  g819
  (
    n1025,
    n547
  );


  buf
  g820
  (
    n1297,
    n611
  );


  buf
  g821
  (
    n1482,
    n359
  );


  not
  g822
  (
    n924,
    n640
  );


  buf
  g823
  (
    n1322,
    n609
  );


  not
  g824
  (
    n695,
    n194
  );


  not
  g825
  (
    n1293,
    n304
  );


  not
  g826
  (
    n1057,
    n587
  );


  buf
  g827
  (
    n1405,
    n650
  );


  buf
  g828
  (
    n680,
    n308
  );


  buf
  g829
  (
    n1226,
    n559
  );


  not
  g830
  (
    n853,
    n618
  );


  not
  g831
  (
    n902,
    n469
  );


  not
  g832
  (
    n919,
    n507
  );


  not
  g833
  (
    n1055,
    n634
  );


  buf
  g834
  (
    n1362,
    n344
  );


  buf
  g835
  (
    n1212,
    n439
  );


  not
  g836
  (
    n678,
    n667
  );


  buf
  g837
  (
    n1122,
    n344
  );


  not
  g838
  (
    n1067,
    n615
  );


  buf
  g839
  (
    n1175,
    n622
  );


  not
  g840
  (
    n1065,
    n181
  );


  buf
  g841
  (
    n786,
    n279
  );


  not
  g842
  (
    n963,
    n575
  );


  buf
  g843
  (
    n1001,
    n173
  );


  buf
  g844
  (
    n1208,
    n374
  );


  not
  g845
  (
    n973,
    n347
  );


  not
  g846
  (
    n841,
    n353
  );


  buf
  g847
  (
    n1252,
    n209
  );


  buf
  g848
  (
    n1154,
    n392
  );


  not
  g849
  (
    n1221,
    n312
  );


  buf
  g850
  (
    n1105,
    n654
  );


  buf
  g851
  (
    n991,
    n272
  );


  not
  g852
  (
    n1246,
    n447
  );


  buf
  g853
  (
    n758,
    n251
  );


  not
  g854
  (
    n817,
    n487
  );


  buf
  g855
  (
    n984,
    n382
  );


  not
  g856
  (
    n1047,
    n330
  );


  buf
  g857
  (
    n1443,
    n434
  );


  not
  g858
  (
    n1425,
    n427
  );


  buf
  g859
  (
    n1341,
    n625
  );


  not
  g860
  (
    n1315,
    n630
  );


  buf
  g861
  (
    n1165,
    n599
  );


  not
  g862
  (
    n779,
    n512
  );


  buf
  g863
  (
    n907,
    n167
  );


  not
  g864
  (
    n768,
    n392
  );


  buf
  g865
  (
    n721,
    n360
  );


  buf
  g866
  (
    n1091,
    n614
  );


  not
  g867
  (
    n826,
    n316
  );


  buf
  g868
  (
    n749,
    n327
  );


  buf
  g869
  (
    n1476,
    n586
  );


  buf
  g870
  (
    n1392,
    n383
  );


  not
  g871
  (
    n709,
    n162
  );


  not
  g872
  (
    n1160,
    n437
  );


  buf
  g873
  (
    n774,
    n559
  );


  buf
  g874
  (
    n1229,
    n324
  );


  not
  g875
  (
    n858,
    n445
  );


  not
  g876
  (
    n1179,
    n384
  );


  not
  g877
  (
    n1059,
    n357
  );


  buf
  g878
  (
    n1207,
    n375
  );


  not
  g879
  (
    n1231,
    n602
  );


  buf
  g880
  (
    n1396,
    n534
  );


  buf
  g881
  (
    n1209,
    n304
  );


  buf
  g882
  (
    n855,
    n325
  );


  not
  g883
  (
    n888,
    n517
  );


  buf
  g884
  (
    n712,
    n503
  );


  not
  g885
  (
    n738,
    n311
  );


  not
  g886
  (
    n750,
    n570
  );


  buf
  g887
  (
    n681,
    n580
  );


  buf
  g888
  (
    n1168,
    n410
  );


  not
  g889
  (
    n1280,
    n255
  );


  buf
  g890
  (
    n1026,
    n307
  );


  buf
  g891
  (
    n1469,
    n186
  );


  not
  g892
  (
    n1114,
    n471
  );


  not
  g893
  (
    n972,
    n583
  );


  buf
  g894
  (
    n1393,
    n400
  );


  buf
  g895
  (
    n1263,
    n190
  );


  buf
  g896
  (
    n936,
    n573
  );


  buf
  g897
  (
    n1232,
    n560
  );


  not
  g898
  (
    n1447,
    n170
  );


  buf
  g899
  (
    n1036,
    n641
  );


  buf
  g900
  (
    n1029,
    n564
  );


  not
  g901
  (
    n1326,
    n374
  );


  buf
  g902
  (
    n939,
    n398
  );


  not
  g903
  (
    n808,
    n390
  );


  not
  g904
  (
    n1041,
    n569
  );


  not
  g905
  (
    n1017,
    n587
  );


  not
  g906
  (
    n1126,
    n174
  );


  buf
  g907
  (
    n743,
    n243
  );


  buf
  g908
  (
    n704,
    n237
  );


  not
  g909
  (
    n1236,
    n359
  );


  not
  g910
  (
    n1475,
    n666
  );


  buf
  g911
  (
    n718,
    n373
  );


  not
  g912
  (
    n1185,
    n322
  );


  not
  g913
  (
    n1247,
    n448
  );


  buf
  g914
  (
    n1347,
    n460
  );


  buf
  g915
  (
    n914,
    n221
  );


  buf
  g916
  (
    n772,
    n542
  );


  buf
  g917
  (
    n1143,
    n467
  );


  not
  g918
  (
    n1380,
    n474
  );


  not
  g919
  (
    n787,
    n331
  );


  not
  g920
  (
    n1456,
    n240
  );


  not
  g921
  (
    n1149,
    n357
  );


  not
  g922
  (
    n815,
    n368
  );


  buf
  g923
  (
    n846,
    n162
  );


  not
  g924
  (
    n1022,
    n424
  );


  buf
  g925
  (
    n964,
    n533
  );


  not
  g926
  (
    n1011,
    n443
  );


  not
  g927
  (
    n1407,
    n475
  );


  buf
  g928
  (
    n1082,
    n265
  );


  buf
  g929
  (
    n1427,
    n459
  );


  not
  g930
  (
    n906,
    n316
  );


  not
  g931
  (
    n1499,
    n314
  );


  buf
  g932
  (
    n1422,
    n473
  );


  not
  g933
  (
    n679,
    n347
  );


  buf
  g934
  (
    n1262,
    n312
  );


  not
  g935
  (
    n800,
    n192
  );


  not
  g936
  (
    n1298,
    n392
  );


  buf
  g937
  (
    n745,
    n656
  );


  not
  g938
  (
    n860,
    n371
  );


  not
  g939
  (
    n1352,
    n532
  );


  not
  g940
  (
    n845,
    n375
  );


  not
  g941
  (
    n698,
    n473
  );


  not
  g942
  (
    n1478,
    n178
  );


  not
  g943
  (
    n816,
    n205
  );


  buf
  g944
  (
    n706,
    n587
  );


  not
  g945
  (
    n1075,
    n203
  );


  buf
  g946
  (
    n1420,
    n541
  );


  buf
  g947
  (
    n791,
    n583
  );


  buf
  g948
  (
    n1344,
    n205
  );


  not
  g949
  (
    n935,
    n456
  );


  not
  g950
  (
    n883,
    n572
  );


  not
  g951
  (
    n1295,
    n548
  );


  not
  g952
  (
    n938,
    n336
  );


  not
  g953
  (
    n1140,
    n550
  );


  buf
  g954
  (
    n761,
    n490
  );


  not
  g955
  (
    n1198,
    n644
  );


  buf
  g956
  (
    n1194,
    n334
  );


  not
  g957
  (
    n1468,
    n282
  );


  not
  g958
  (
    n744,
    n663
  );


  buf
  g959
  (
    n728,
    n353
  );


  buf
  g960
  (
    n1239,
    n643
  );


  not
  g961
  (
    n891,
    n414
  );


  not
  g962
  (
    n1429,
    n186
  );


  buf
  g963
  (
    n825,
    n457
  );


  buf
  g964
  (
    n1357,
    n562
  );


  not
  g965
  (
    n811,
    n161
  );


  buf
  g966
  (
    n754,
    n609
  );


  buf
  g967
  (
    n689,
    n370
  );


  buf
  g968
  (
    n982,
    n486
  );


  buf
  g969
  (
    n1021,
    n515
  );


  not
  g970
  (
    n934,
    n594
  );


  buf
  g971
  (
    n1173,
    n372
  );


  not
  g972
  (
    n836,
    n208
  );


  buf
  g973
  (
    n1444,
    n572
  );


  buf
  g974
  (
    n1432,
    n477
  );


  not
  g975
  (
    n820,
    n275
  );


  not
  g976
  (
    n1354,
    n357
  );


  buf
  g977
  (
    n1459,
    n171
  );


  not
  g978
  (
    n1118,
    n642
  );


  buf
  g979
  (
    n1281,
    n546
  );


  not
  g980
  (
    n1138,
    n415
  );


  not
  g981
  (
    n1483,
    n302
  );


  buf
  g982
  (
    n1192,
    n593
  );


  buf
  g983
  (
    n1462,
    n352
  );


  not
  g984
  (
    n873,
    n442
  );


  not
  g985
  (
    n1381,
    n479
  );


  buf
  g986
  (
    n1433,
    n218
  );


  buf
  g987
  (
    n903,
    n269
  );


  not
  g988
  (
    n1061,
    n453
  );


  not
  g989
  (
    n824,
    n657
  );


  not
  g990
  (
    n1242,
    n240
  );


  buf
  g991
  (
    n1474,
    n331
  );


  buf
  g992
  (
    n777,
    n588
  );


  buf
  g993
  (
    n1100,
    n364
  );


  buf
  g994
  (
    n1186,
    n632
  );


  not
  g995
  (
    n1385,
    n378
  );


  not
  g996
  (
    n848,
    n373
  );


  not
  g997
  (
    n1153,
    n527
  );


  buf
  g998
  (
    n1189,
    n277
  );


  buf
  g999
  (
    n1339,
    n220
  );


  not
  g1000
  (
    n1094,
    n266
  );


  buf
  g1001
  (
    n1428,
    n383
  );


  not
  g1002
  (
    n1504,
    n616
  );


  buf
  g1003
  (
    n740,
    n581
  );


  buf
  g1004
  (
    n1378,
    n557
  );


  buf
  g1005
  (
    n1166,
    n554
  );


  not
  g1006
  (
    n716,
    n195
  );


  not
  g1007
  (
    n1072,
    n182
  );


  buf
  g1008
  (
    n954,
    n358
  );


  buf
  g1009
  (
    n1283,
    n397
  );


  not
  g1010
  (
    n985,
    n166
  );


  buf
  g1011
  (
    n949,
    n415
  );


  not
  g1012
  (
    n974,
    n421
  );


  not
  g1013
  (
    n1486,
    n322
  );


  not
  g1014
  (
    n752,
    n164
  );


  buf
  g1015
  (
    n830,
    n230
  );


  buf
  g1016
  (
    n1409,
    n609
  );


  not
  g1017
  (
    n1254,
    n550
  );


  buf
  g1018
  (
    n918,
    n207
  );


  not
  g1019
  (
    n1219,
    n578
  );


  not
  g1020
  (
    n737,
    n178
  );


  not
  g1021
  (
    n893,
    n417
  );


  not
  g1022
  (
    n867,
    n465
  );


  not
  g1023
  (
    n1084,
    n451
  );


  buf
  g1024
  (
    n948,
    n592
  );


  buf
  g1025
  (
    n776,
    n468
  );


  not
  g1026
  (
    n898,
    n501
  );


  not
  g1027
  (
    n685,
    n170
  );


  not
  g1028
  (
    n797,
    n398
  );


  buf
  g1029
  (
    KeyWire_0_3,
    n275
  );


  not
  g1030
  (
    n1463,
    n205
  );


  buf
  g1031
  (
    n805,
    n667
  );


  not
  g1032
  (
    n701,
    n260
  );


  buf
  g1033
  (
    n1003,
    n446
  );


  buf
  g1034
  (
    n724,
    n465
  );


  not
  g1035
  (
    n1446,
    n635
  );


  not
  g1036
  (
    n1481,
    n413
  );


  not
  g1037
  (
    n1121,
    n281
  );


  buf
  g1038
  (
    n1127,
    n415
  );


  not
  g1039
  (
    n1144,
    n621
  );


  buf
  g1040
  (
    n1107,
    n189
  );


  buf
  g1041
  (
    n1235,
    n268
  );


  not
  g1042
  (
    n925,
    n539
  );


  not
  g1043
  (
    n1131,
    n277
  );


  not
  g1044
  (
    n1068,
    n369
  );


  buf
  g1045
  (
    n1373,
    n167
  );


  buf
  g1046
  (
    n859,
    n466
  );


  buf
  g1047
  (
    n1023,
    n390
  );


  not
  g1048
  (
    n892,
    n240
  );


  not
  g1049
  (
    n1421,
    n294
  );


  buf
  g1050
  (
    n995,
    n389
  );


  not
  g1051
  (
    n967,
    n299
  );


  not
  g1052
  (
    n1330,
    n656
  );


  not
  g1053
  (
    n1156,
    n505
  );


  not
  g1054
  (
    n1132,
    n539
  );


  not
  g1055
  (
    n1098,
    n492
  );


  buf
  g1056
  (
    n912,
    n559
  );


  not
  g1057
  (
    n1303,
    n225
  );


  not
  g1058
  (
    n951,
    n443
  );


  not
  g1059
  (
    n1045,
    n651
  );


  buf
  g1060
  (
    n1024,
    n503
  );


  not
  g1061
  (
    n1332,
    n560
  );


  not
  g1062
  (
    n1183,
    n169
  );


  buf
  g1063
  (
    n1170,
    n454
  );


  not
  g1064
  (
    n760,
    n201
  );


  not
  g1065
  (
    n1009,
    n639
  );


  buf
  g1066
  (
    n794,
    n325
  );


  not
  g1067
  (
    n1290,
    n201
  );


  buf
  g1068
  (
    n1218,
    n298
  );


  buf
  g1069
  (
    n1503,
    n329
  );


  not
  g1070
  (
    n1485,
    n440
  );


  buf
  g1071
  (
    n677,
    n364
  );


  buf
  g1072
  (
    n1460,
    n621
  );


  nand
  g1073
  (
    n1284,
    n636,
    n435,
    n414
  );


  nor
  g1074
  (
    n1190,
    n362,
    n309,
    n454,
    n443
  );


  xnor
  g1075
  (
    n793,
    n170,
    n613,
    n387,
    n350
  );


  and
  g1076
  (
    n1191,
    n489,
    n450,
    n522,
    n521
  );


  xnor
  g1077
  (
    n889,
    n464,
    n626,
    n319,
    n188
  );


  or
  g1078
  (
    n1299,
    n622,
    n236,
    n191,
    n586
  );


  and
  g1079
  (
    n1419,
    n624,
    n584,
    n668,
    n249
  );


  xnor
  g1080
  (
    n1085,
    n337,
    n472,
    n354,
    n247
  );


  xor
  g1081
  (
    n1164,
    n252,
    n259,
    n214,
    n264
  );


  xnor
  g1082
  (
    n1336,
    n352,
    n547,
    n476,
    n274
  );


  nand
  g1083
  (
    n1395,
    n366,
    n603,
    n236,
    n488
  );


  xor
  g1084
  (
    n1069,
    n628,
    n590,
    n658,
    n198
  );


  xnor
  g1085
  (
    n1193,
    n646,
    n597,
    n352,
    n395
  );


  xor
  g1086
  (
    n1223,
    n410,
    n173,
    n240,
    n197
  );


  and
  g1087
  (
    n992,
    n567,
    n214,
    n425,
    n422
  );


  or
  g1088
  (
    n1142,
    n558,
    n643,
    n320,
    n210
  );


  or
  g1089
  (
    n987,
    n193,
    n444,
    n657,
    n474
  );


  xor
  g1090
  (
    n1030,
    n461,
    n477,
    n371,
    n408
  );


  or
  g1091
  (
    n1423,
    n656,
    n507,
    n635,
    n280
  );


  and
  g1092
  (
    n770,
    n481,
    n501,
    n242,
    n267
  );


  xor
  g1093
  (
    n1081,
    n295,
    n250,
    n591,
    n289
  );


  xnor
  g1094
  (
    n1076,
    n236,
    n644,
    n228,
    n478
  );


  nor
  g1095
  (
    n1372,
    n460,
    n166,
    n580,
    n604
  );


  nand
  g1096
  (
    n746,
    n615,
    n203,
    n247,
    n351
  );


  or
  g1097
  (
    n676,
    n227,
    n444,
    n200,
    n516
  );


  nor
  g1098
  (
    n926,
    n215,
    n647,
    n237,
    n313
  );


  xor
  g1099
  (
    n822,
    n355,
    n568,
    n420,
    n647
  );


  and
  g1100
  (
    n691,
    n165,
    n310,
    n461,
    n426
  );


  and
  g1101
  (
    n900,
    n270,
    n597,
    n176,
    n576
  );


  xnor
  g1102
  (
    n751,
    n182,
    n176,
    n376,
    n556
  );


  xnor
  g1103
  (
    n1286,
    n477,
    n621,
    n179,
    n324
  );


  nor
  g1104
  (
    n968,
    n346,
    n662,
    n500,
    n344
  );


  xor
  g1105
  (
    n1466,
    n560,
    n253,
    n607,
    n565
  );


  xnor
  g1106
  (
    n921,
    n660,
    n234,
    n239,
    n590
  );


  nand
  g1107
  (
    n763,
    n601,
    n451,
    n308,
    n176
  );


  xor
  g1108
  (
    n871,
    n173,
    n612,
    n638,
    n366
  );


  xor
  g1109
  (
    n1416,
    n620,
    n499,
    n585,
    n459
  );


  xor
  g1110
  (
    n1370,
    n632,
    n436,
    n595,
    n520
  );


  nor
  g1111
  (
    n764,
    n319,
    n374,
    n432,
    n533
  );


  or
  g1112
  (
    n1334,
    n393,
    n342,
    n429,
    n565
  );


  xnor
  g1113
  (
    n1412,
    n603,
    n573,
    n196,
    n661
  );


  nor
  g1114
  (
    n1034,
    n379,
    n335,
    n564,
    n579
  );


  nand
  g1115
  (
    n1439,
    n511,
    n191,
    n406,
    n289
  );


  xnor
  g1116
  (
    n953,
    n600,
    n370,
    n326,
    n272
  );


  nand
  g1117
  (
    n922,
    n613,
    n268,
    n216,
    n403
  );


  xnor
  g1118
  (
    n1066,
    n652,
    n551,
    n246,
    n290
  );


  and
  g1119
  (
    n801,
    n395,
    n624,
    n317,
    n350
  );


  nor
  g1120
  (
    n1400,
    n269,
    n239,
    n424,
    n563
  );


  nand
  g1121
  (
    n976,
    n530,
    n578,
    n362,
    n466
  );


  or
  g1122
  (
    n1367,
    n296,
    n214,
    n642,
    n588
  );


  or
  g1123
  (
    n1033,
    n551,
    n540,
    n310,
    n669
  );


  or
  g1124
  (
    n733,
    n518,
    n423,
    n422,
    n354
  );


  nor
  g1125
  (
    n1377,
    n552,
    n280,
    n582,
    n666
  );


  nand
  g1126
  (
    n1028,
    n643,
    n291,
    n248,
    n196
  );


  or
  g1127
  (
    n1477,
    n178,
    n616,
    n318,
    n448
  );


  xor
  g1128
  (
    n933,
    n519,
    n495,
    n597,
    n631
  );


  xor
  g1129
  (
    n1241,
    n423,
    n340,
    n663,
    n360
  );


  xnor
  g1130
  (
    n971,
    n568,
    n312,
    n319,
    n424
  );


  or
  g1131
  (
    n1244,
    n489,
    n512,
    n166,
    n235
  );


  xor
  g1132
  (
    n707,
    n229,
    n361,
    n348,
    n534
  );


  or
  g1133
  (
    n865,
    n418,
    n589,
    n574,
    n606
  );


  nand
  g1134
  (
    n1272,
    n543,
    n194,
    n417,
    n482
  );


  and
  g1135
  (
    n1312,
    n320,
    n293,
    n572,
    n297
  );


  or
  g1136
  (
    n1285,
    n658,
    n671,
    n432,
    n553
  );


  nand
  g1137
  (
    n1401,
    n486,
    n567,
    n670,
    n519
  );


  xnor
  g1138
  (
    n1211,
    n289,
    n377,
    n161,
    n548
  );


  xnor
  g1139
  (
    n1448,
    n295,
    n663,
    n397,
    n399
  );


  xnor
  g1140
  (
    n1333,
    n600,
    n645,
    n630,
    n522
  );


  xor
  g1141
  (
    n1197,
    n330,
    n654,
    n498,
    n670
  );


  or
  g1142
  (
    n874,
    n592,
    n484,
    n413,
    n215
  );


  xnor
  g1143
  (
    n1004,
    n313,
    n419,
    n181,
    n454
  );


  xnor
  g1144
  (
    n864,
    n663,
    n432,
    n549,
    n248
  );


  and
  g1145
  (
    n1267,
    n429,
    n405,
    n502,
    n529
  );


  or
  g1146
  (
    n1006,
    n238,
    n169,
    n245,
    n520
  );


  or
  g1147
  (
    n1199,
    n472,
    n515,
    n475,
    n259
  );


  nor
  g1148
  (
    n753,
    n262,
    n429,
    n415,
    n540
  );


  nor
  g1149
  (
    n1371,
    n204,
    n400,
    n370,
    n441
  );


  xor
  g1150
  (
    n1491,
    n209,
    n248,
    n657,
    n520
  );


  nand
  g1151
  (
    n840,
    n589,
    n549,
    n229,
    n224
  );


  xor
  g1152
  (
    n890,
    n384,
    n202,
    n490,
    n190
  );


  nor
  g1153
  (
    n1288,
    n496,
    n506,
    n460,
    n202
  );


  nor
  g1154
  (
    n905,
    n566,
    n260,
    n531,
    n340
  );


  and
  g1155
  (
    n975,
    n311,
    n624,
    n264,
    n332
  );


  nand
  g1156
  (
    n1146,
    n342,
    n275,
    n211,
    n607
  );


  or
  g1157
  (
    n717,
    n419,
    n268,
    n422,
    n359
  );


  nor
  g1158
  (
    n1250,
    n626,
    n263,
    n245,
    n484
  );


  xor
  g1159
  (
    n941,
    n343,
    n253,
    n518,
    n347
  );


  nor
  g1160
  (
    n775,
    n335,
    n385,
    n326,
    n423
  );


  or
  g1161
  (
    n913,
    n585,
    n556,
    n507,
    n617
  );


  nor
  g1162
  (
    n710,
    n525,
    n467,
    n648,
    n486
  );


  xnor
  g1163
  (
    n1111,
    n317,
    n403,
    n409,
    n372
  );


  nor
  g1164
  (
    n1413,
    n452,
    n541,
    n393,
    n599
  );


  nor
  g1165
  (
    n1414,
    n623,
    n499,
    n433,
    n409
  );


  or
  g1166
  (
    n1228,
    n632,
    n622,
    n529,
    n671
  );


  nor
  g1167
  (
    n757,
    n553,
    n655,
    n476,
    n361
  );


  xor
  g1168
  (
    n1455,
    n474,
    n317,
    n333,
    n219
  );


  nor
  g1169
  (
    n929,
    n671,
    n531,
    n418,
    n298
  );


  and
  g1170
  (
    n877,
    n265,
    n523,
    n567,
    n370
  );


  xnor
  g1171
  (
    n1324,
    n247,
    n289,
    n266,
    n349
  );


  or
  g1172
  (
    n959,
    n314,
    n265,
    n609,
    n408
  );


  xnor
  g1173
  (
    n818,
    n224,
    n231,
    n601,
    n275
  );


  nand
  g1174
  (
    n1014,
    n493,
    n582,
    n418,
    n398
  );


  or
  g1175
  (
    n1355,
    n188,
    n273,
    n469,
    n217
  );


  or
  g1176
  (
    n819,
    n281,
    n343,
    n497,
    n437
  );


  and
  g1177
  (
    n1268,
    n285,
    n526,
    n546,
    n619
  );


  xnor
  g1178
  (
    n1479,
    n235,
    n296,
    n532,
    n604
  );


  nand
  g1179
  (
    n688,
    n180,
    n253,
    n367,
    n207
  );


  and
  g1180
  (
    n1158,
    n386,
    n468,
    n218,
    n436
  );


  or
  g1181
  (
    n729,
    n525,
    n554,
    n244,
    n301
  );


  nor
  g1182
  (
    n1225,
    n274,
    n525,
    n391,
    n228
  );


  nand
  g1183
  (
    n1093,
    n396,
    n426,
    n168,
    n323
  );


  nand
  g1184
  (
    n1079,
    n340,
    n335,
    n619,
    n202
  );


  nor
  g1185
  (
    n1265,
    n571,
    n563,
    n490,
    n171
  );


  nor
  g1186
  (
    n1434,
    n350,
    n542,
    n497,
    n603
  );


  nand
  g1187
  (
    n862,
    n636,
    n499,
    n296,
    n556
  );


  and
  g1188
  (
    n1253,
    n280,
    n418,
    n363,
    n500
  );


  nor
  g1189
  (
    n1133,
    n553,
    n263,
    n589,
    n483
  );


  xor
  g1190
  (
    n1005,
    n646,
    n260,
    n168,
    n391
  );


  nor
  g1191
  (
    n847,
    n604,
    n295,
    n197,
    n230
  );


  nor
  g1192
  (
    n1032,
    n644,
    n577,
    n626,
    n634
  );


  xnor
  g1193
  (
    n931,
    n637,
    n401,
    n501,
    n478
  );


  and
  g1194
  (
    n894,
    n434,
    n261,
    n643,
    n516
  );


  xor
  g1195
  (
    n1294,
    n171,
    n654,
    n574,
    n208
  );


  nand
  g1196
  (
    n1451,
    n433,
    n465,
    n666,
    n668
  );


  xnor
  g1197
  (
    n1002,
    n226,
    n232,
    n270,
    n352
  );


  nand
  g1198
  (
    n1106,
    n425,
    n396,
    n558,
    n575
  );


  xnor
  g1199
  (
    n781,
    n591,
    n287,
    n286,
    n225
  );


  and
  g1200
  (
    n1016,
    n579,
    n378,
    n664,
    n368
  );


  nor
  g1201
  (
    n1467,
    n476,
    n254,
    n642,
    n488
  );


  nand
  g1202
  (
    n1410,
    n256,
    n510,
    n327,
    n192
  );


  xnor
  g1203
  (
    n1089,
    n570,
    n180,
    n328,
    n318
  );


  or
  g1204
  (
    n1109,
    n406,
    n391,
    n411,
    n185
  );


  xnor
  g1205
  (
    KeyWire_0_8,
    n670,
    n605,
    n367,
    n305
  );


  or
  g1206
  (
    n1449,
    n274,
    n408,
    n610,
    n222
  );


  nor
  g1207
  (
    n1496,
    n217,
    n310,
    n446,
    n548
  );


  xnor
  g1208
  (
    n1264,
    n428,
    n188,
    n577,
    n492
  );


  nor
  g1209
  (
    n714,
    n653,
    n668,
    n321,
    n483
  );


  and
  g1210
  (
    n1345,
    n324,
    n250,
    n436,
    n484
  );


  and
  g1211
  (
    n1087,
    n463,
    n569,
    n650,
    n574
  );


  nor
  g1212
  (
    n1484,
    n590,
    n539,
    n315,
    n487
  );


  xnor
  g1213
  (
    n997,
    n466,
    n380,
    n333,
    n204
  );


  nand
  g1214
  (
    n1077,
    n477,
    n523,
    n322,
    n619
  );


  nor
  g1215
  (
    n1430,
    n371,
    n276,
    n624,
    n301
  );


  and
  g1216
  (
    n1134,
    n365,
    n633,
    n599,
    n187
  );


  xnor
  g1217
  (
    n981,
    n326,
    n239,
    n432,
    n640
  );


  and
  g1218
  (
    n1335,
    n508,
    n665,
    n266,
    n331
  );


  or
  g1219
  (
    n958,
    n342,
    n649,
    n526,
    n430
  );


  and
  g1220
  (
    n1125,
    n211,
    n263,
    n290,
    n498
  );


  or
  g1221
  (
    n1397,
    n425,
    n301,
    n598,
    n497
  );


  nor
  g1222
  (
    n1308,
    n206,
    n229,
    n457,
    n203
  );


  or
  g1223
  (
    n1495,
    n353,
    n210,
    n319,
    n555
  );


  or
  g1224
  (
    n1240,
    n442,
    n221,
    n264,
    n321
  );


  nor
  g1225
  (
    n960,
    n388,
    n416,
    n501,
    n288
  );


  xnor
  g1226
  (
    n945,
    n185,
    n412,
    n644,
    n479
  );


  nand
  g1227
  (
    n1155,
    n660,
    n430,
    n657,
    n261
  );


  xnor
  g1228
  (
    n769,
    n504,
    n629,
    n637,
    n428
  );


  or
  g1229
  (
    n952,
    n345,
    n318,
    n276,
    n164
  );


  nor
  g1230
  (
    n978,
    n239,
    n316,
    n181,
    n299
  );


  nor
  g1231
  (
    n807,
    n485,
    n554,
    n236,
    n203
  );


  xnor
  g1232
  (
    n965,
    n332,
    n615,
    n271,
    n307
  );


  nor
  g1233
  (
    n910,
    n193,
    n630,
    n402,
    n258
  );


  and
  g1234
  (
    n1435,
    n172,
    n390,
    n183,
    n366
  );


  xnor
  g1235
  (
    n1234,
    n379,
    n330,
    n668,
    n412
  );


  nand
  g1236
  (
    n886,
    n645,
    n343,
    n337,
    n630
  );


  xor
  g1237
  (
    n1399,
    n506,
    n517,
    n629,
    n528
  );


  and
  g1238
  (
    n930,
    n256,
    n468,
    n452,
    n329
  );


  xor
  g1239
  (
    n809,
    n592,
    n444,
    n175,
    n220
  );


  nor
  g1240
  (
    n1403,
    n198,
    n505,
    n669,
    n222
  );


  and
  g1241
  (
    n795,
    n243,
    n633,
    n358,
    n216
  );


  and
  g1242
  (
    n722,
    n613,
    n338,
    n620,
    n393
  );


  nand
  g1243
  (
    n1110,
    n530,
    n175,
    n320,
    n358
  );


  or
  g1244
  (
    n996,
    n356,
    n242,
    n269,
    n616
  );


  and
  g1245
  (
    n1130,
    n601,
    n552,
    n544,
    n438
  );


  nor
  g1246
  (
    n1049,
    n281,
    n216,
    n495,
    n508
  );


  nor
  g1247
  (
    n943,
    n469,
    n262,
    n344,
    n633
  );


  or
  g1248
  (
    n1102,
    n232,
    n163,
    n323,
    n297
  );


  nor
  g1249
  (
    n1508,
    n488,
    n310,
    n469,
    n356
  );


  nor
  g1250
  (
    n813,
    n506,
    n384,
    n521,
    n233
  );


  nor
  g1251
  (
    n1096,
    n547,
    n380,
    n278,
    n315
  );


  xnor
  g1252
  (
    n804,
    n387,
    n384,
    n465,
    n558
  );


  xor
  g1253
  (
    n1054,
    n421,
    n378,
    n576,
    n475
  );


  xor
  g1254
  (
    n1139,
    n590,
    n305,
    n177,
    n169
  );


  nor
  g1255
  (
    n782,
    n187,
    n503,
    n658,
    n563
  );


  nand
  g1256
  (
    n725,
    n300,
    n231,
    n245,
    n409
  );


  nand
  g1257
  (
    n870,
    n509,
    n233,
    n213,
    n262
  );


  nand
  g1258
  (
    n1411,
    n315,
    n494,
    n564,
    n601
  );


  or
  g1259
  (
    n1342,
    n392,
    n391,
    n594,
    n449
  );


  or
  g1260
  (
    n1171,
    n382,
    n587,
    n459,
    n583
  );


  and
  g1261
  (
    n1099,
    n261,
    n662,
    n652,
    n185
  );


  nand
  g1262
  (
    n1473,
    n179,
    n172,
    n214,
    n500
  );


  and
  g1263
  (
    n854,
    n440,
    n213,
    n513,
    n273
  );


  and
  g1264
  (
    n682,
    n610,
    n165,
    n438,
    n625
  );


  xnor
  g1265
  (
    n1060,
    n616,
    n379,
    n452,
    n311
  );


  or
  g1266
  (
    n1464,
    n651,
    n662,
    n397,
    n196
  );


  xor
  g1267
  (
    n896,
    n284,
    n278,
    n440,
    n387
  );


  or
  g1268
  (
    n1368,
    n180,
    n191,
    n578,
    n199
  );


  xnor
  g1269
  (
    n884,
    n387,
    n343,
    n232,
    n224
  );


  xor
  g1270
  (
    n784,
    n505,
    n190,
    n478,
    n535
  );


  xnor
  g1271
  (
    n756,
    n435,
    n241,
    n278,
    n345
  );


  xnor
  g1272
  (
    n1038,
    n439,
    n480,
    n430,
    n365
  );


  nand
  g1273
  (
    n844,
    n226,
    n639,
    n586,
    n169
  );


  xnor
  g1274
  (
    n1040,
    n456,
    n413,
    n322,
    n213
  );


  xor
  g1275
  (
    n1348,
    n634,
    n222,
    n244,
    n192
  );


  and
  g1276
  (
    n1313,
    n260,
    n365,
    n522,
    n412
  );


  nor
  g1277
  (
    n1195,
    n286,
    n411,
    n279,
    n472
  );


  and
  g1278
  (
    n1159,
    n303,
    n451,
    n533,
    n332
  );


  nor
  g1279
  (
    n1311,
    n555,
    n542,
    n431,
    n374
  );


  and
  g1280
  (
    n1095,
    n284,
    n491,
    n250,
    n530
  );


  nand
  g1281
  (
    n1248,
    n504,
    n607,
    n502,
    n641
  );


  xnor
  g1282
  (
    n1008,
    n651,
    n431,
    n217,
    n582
  );


  nor
  g1283
  (
    n1188,
    n238,
    n610,
    n177,
    n633
  );


  nor
  g1284
  (
    n904,
    n195,
    n438,
    n615,
    n443
  );


  nor
  g1285
  (
    n1498,
    n262,
    n316,
    n659,
    n638
  );


  nand
  g1286
  (
    n1051,
    n398,
    n481,
    n403,
    n266
  );


  nor
  g1287
  (
    n675,
    n385,
    n498,
    n216,
    n237
  );


  nand
  g1288
  (
    n1063,
    n305,
    n537,
    n220,
    n649
  );


  and
  g1289
  (
    n1453,
    n251,
    n345,
    n623,
    n254
  );


  and
  g1290
  (
    n1305,
    n167,
    n467,
    n494,
    n197
  );


  or
  g1291
  (
    n1346,
    n185,
    n564,
    n493,
    n669
  );


  nand
  g1292
  (
    n1222,
    n300,
    n404,
    n346,
    n228
  );


  nor
  g1293
  (
    n895,
    n509,
    n581,
    n470,
    n209
  );


  nand
  g1294
  (
    n1136,
    n445,
    n300,
    n227,
    n426
  );


  or
  g1295
  (
    n1359,
    n346,
    n219,
    n388,
    n504
  );


  nand
  g1296
  (
    n962,
    n603,
    n222,
    n607,
    n406
  );


  nand
  g1297
  (
    n1440,
    n251,
    n641,
    n250,
    n163
  );


  xor
  g1298
  (
    n1470,
    n372,
    n636,
    n561,
    n409
  );


  or
  g1299
  (
    n1274,
    n272,
    n282,
    n389,
    n402
  );


  nor
  g1300
  (
    n950,
    n512,
    n524,
    n453,
    n296
  );


  xor
  g1301
  (
    n969,
    n360,
    n584,
    n242,
    n453
  );


  nand
  g1302
  (
    n1369,
    n233,
    n212,
    n270,
    n170
  );


  xnor
  g1303
  (
    n897,
    n246,
    n416,
    n625,
    n671
  );


  xor
  g1304
  (
    n1116,
    n552,
    n514,
    n364,
    n612
  );


  xor
  g1305
  (
    n911,
    n249,
    n183,
    n229,
    n464
  );


  nand
  g1306
  (
    n937,
    n381,
    n517,
    n246,
    n284
  );


  nand
  g1307
  (
    n1323,
    n368,
    n577,
    n287,
    n613
  );


  or
  g1308
  (
    n1224,
    n614,
    n248,
    n466,
    n598
  );


  nand
  g1309
  (
    n693,
    n235,
    n327,
    n199,
    n187
  );


  and
  g1310
  (
    n1490,
    n346,
    n241,
    n605,
    n376
  );


  xnor
  g1311
  (
    n1097,
    n189,
    n541,
    n382,
    n208
  );


  and
  g1312
  (
    n856,
    n566,
    n628,
    n355,
    n505
  );


  or
  g1313
  (
    n932,
    n184,
    n336,
    n665,
    n593
  );


  xor
  g1314
  (
    n1214,
    n467,
    n227,
    n520,
    n182
  );


  xnor
  g1315
  (
    n1270,
    n226,
    n184,
    n621,
    n302
  );


  or
  g1316
  (
    n790,
    n569,
    n362,
    n441,
    n538
  );


  nand
  g1317
  (
    n1506,
    n618,
    n637,
    n446,
    n416
  );


  xnor
  g1318
  (
    n1115,
    n408,
    n494,
    n244,
    n277
  );


  nand
  g1319
  (
    n1257,
    n430,
    n354,
    n434,
    n475
  );


  and
  g1320
  (
    n1387,
    n200,
    n543,
    n523,
    n653
  );


  nand
  g1321
  (
    n1251,
    n461,
    n437,
    n173,
    n305
  );


  and
  g1322
  (
    n762,
    n227,
    n519,
    n271,
    n373
  );


  or
  g1323
  (
    n940,
    n256,
    n394,
    n407,
    n183
  );


  and
  g1324
  (
    n1181,
    n464,
    n458,
    n510,
    n165
  );


  xor
  g1325
  (
    n723,
    n225,
    n423,
    n532,
    n463
  );


  xor
  g1326
  (
    n1172,
    n350,
    n457,
    n329,
    n531
  );


  and
  g1327
  (
    n1329,
    n462,
    n297,
    n215,
    n513
  );


  xor
  g1328
  (
    n829,
    n618,
    n560,
    n455,
    n502
  );


  xor
  g1329
  (
    n999,
    n596,
    n363,
    n255,
    n375
  );


  nand
  g1330
  (
    n857,
    n518,
    n472,
    n441,
    n295
  );


  nand
  g1331
  (
    n1505,
    n195,
    n521,
    n336,
    n308
  );


  xor
  g1332
  (
    n1364,
    n491,
    n402,
    n312,
    n545
  );


  xor
  g1333
  (
    n1048,
    n631,
    n544,
    n653,
    n264
  );


  nand
  g1334
  (
    n1415,
    n661,
    n629,
    n258,
    n655
  );


  nor
  g1335
  (
    n834,
    n639,
    n544,
    n664,
    n162
  );


  or
  g1336
  (
    n1457,
    n186,
    n306,
    n167,
    n381
  );


  xor
  g1337
  (
    n837,
    n369,
    n237,
    n509,
    n462
  );


  and
  g1338
  (
    n1406,
    n608,
    n470,
    n599,
    n297
  );


  or
  g1339
  (
    n1261,
    n306,
    n364,
    n219,
    n659
  );


  xnor
  g1340
  (
    n842,
    n342,
    n442,
    n377,
    n474
  );


  and
  g1341
  (
    n1465,
    n456,
    n355,
    n642,
    n299
  );


  nor
  g1342
  (
    n1108,
    n184,
    n304,
    n582,
    n635
  );


  or
  g1343
  (
    n887,
    n636,
    n620,
    n591,
    n598
  );


  xnor
  g1344
  (
    n832,
    n381,
    n605,
    n314,
    n519
  );


  nand
  g1345
  (
    n1343,
    n285,
    n424,
    n427,
    n334
  );


  xnor
  g1346
  (
    n1349,
    n597,
    n375,
    n614,
    n192
  );


  or
  g1347
  (
    n1398,
    n458,
    n435,
    n320,
    n401
  );


  and
  g1348
  (
    n1074,
    n257,
    n399,
    n625,
    n258
  );


  nand
  g1349
  (
    n726,
    n405,
    n328,
    n313,
    n507
  );


  nor
  g1350
  (
    n869,
    n277,
    n186,
    n356,
    n514
  );


  xnor
  g1351
  (
    n1289,
    n602,
    n389,
    n517,
    n670
  );


  xnor
  g1352
  (
    n1204,
    n604,
    n194,
    n535,
    n557
  );


  nor
  g1353
  (
    n708,
    n341,
    n400,
    n367,
    n450
  );


  xnor
  g1354
  (
    n783,
    n303,
    n188,
    n496,
    n411
  );


  xnor
  g1355
  (
    n989,
    n390,
    n168,
    n660,
    n163
  );


  xor
  g1356
  (
    n928,
    n284,
    n204,
    n508,
    n213
  );


  and
  g1357
  (
    n1169,
    n172,
    n614,
    n235,
    n460
  );


  nand
  g1358
  (
    n851,
    n536,
    n627,
    n527,
    n514
  );


  nand
  g1359
  (
    n1200,
    n362,
    n538,
    n285,
    n395
  );


  xnor
  g1360
  (
    n1314,
    n401,
    n556,
    n639,
    n574
  );


  nor
  g1361
  (
    n1012,
    n459,
    n349,
    n377,
    n476
  );


  xnor
  g1362
  (
    n1053,
    n448,
    n348,
    n666,
    n195
  );


  and
  g1363
  (
    n927,
    n575,
    n489,
    n610,
    n246
  );


  or
  g1364
  (
    n909,
    n655,
    n537,
    n389,
    n321
  );


  nand
  g1365
  (
    n1201,
    n557,
    n515,
    n497,
    n382
  );


  xnor
  g1366
  (
    n1237,
    n513,
    n521,
    n338,
    n317
  );


  or
  g1367
  (
    n1325,
    n581,
    n487,
    n361,
    n183
  );


  nand
  g1368
  (
    n1217,
    n363,
    n351,
    n646,
    n611
  );


  or
  g1369
  (
    n866,
    n542,
    n311,
    n177,
    n492
  );


  and
  g1370
  (
    n1282,
    n228,
    n241,
    n598,
    n544
  );


  xnor
  g1371
  (
    n1092,
    n470,
    n210,
    n626,
    n282
  );


  or
  g1372
  (
    n1320,
    n417,
    n166,
    n291,
    n580
  );


  nand
  g1373
  (
    n703,
    n339,
    n665,
    n485
  );


  xnor
  g1374
  (
    n977,
    n217,
    n493,
    n568,
    n640
  );


  xor
  g1375
  (
    n1123,
    n286,
    n458,
    n577,
    n480
  );


  nand
  g1376
  (
    n1073,
    n309,
    n234,
    n537,
    n571
  );


  nand
  g1377
  (
    n956,
    n532,
    n193,
    n198,
    n540
  );


  xnor
  g1378
  (
    n771,
    n274,
    n360,
    n498,
    n405
  );


  xor
  g1379
  (
    n1291,
    n428,
    n524,
    n579,
    n288
  );


  and
  g1380
  (
    n1488,
    n412,
    n543,
    n523,
    n440
  );


  xor
  g1381
  (
    n1083,
    n410,
    n341,
    n283,
    n535
  );


  or
  g1382
  (
    n879,
    n206,
    n608,
    n309,
    n656
  );


  and
  g1383
  (
    n711,
    n165,
    n627,
    n485,
    n267
  );


  and
  g1384
  (
    n1243,
    n543,
    n238,
    n661,
    n562
  );


  nand
  g1385
  (
    n1316,
    n491,
    n308,
    n482,
    n638
  );


  nor
  g1386
  (
    n881,
    n429,
    n552,
    n258,
    n545
  );


  nor
  g1387
  (
    n734,
    n530,
    n483,
    n161,
    n535
  );


  xnor
  g1388
  (
    n1273,
    n662,
    n664,
    n201,
    n283
  );


  or
  g1389
  (
    n1458,
    n508,
    n407,
    n172,
    n303
  );


  nor
  g1390
  (
    n687,
    n580,
    n553,
    n403,
    n292
  );


  xor
  g1391
  (
    n946,
    n480,
    n510,
    n182,
    n357
  );


  nand
  g1392
  (
    n1501,
    n345,
    n573,
    n293,
    n177
  );


  or
  g1393
  (
    n713,
    n174,
    n528,
    n506,
    n249
  );


  xor
  g1394
  (
    n1119,
    n200,
    n292,
    n302,
    n327
  );


  and
  g1395
  (
    n1182,
    n307,
    n526,
    n591,
    n294
  );


  nor
  g1396
  (
    n880,
    n571,
    n651,
    n249,
    n448
  );


  xor
  g1397
  (
    n979,
    n176,
    n394,
    n230,
    n355
  );


  and
  g1398
  (
    n1442,
    n397,
    n340,
    n259,
    n252
  );


  xor
  g1399
  (
    n1318,
    n339,
    n584,
    n218,
    n629
  );


  xor
  g1400
  (
    n915,
    n439,
    n273,
    n359,
    n606
  );


  xor
  g1401
  (
    n923,
    n539,
    n647,
    n257,
    n534
  );


  nor
  g1402
  (
    n690,
    n488,
    n279,
    n526,
    n163
  );


  nand
  g1403
  (
    n1071,
    n404,
    n562,
    n455,
    n314
  );


  nand
  g1404
  (
    n1386,
    n537,
    n404,
    n363,
    n431
  );


  and
  g1405
  (
    n1245,
    n455,
    n358,
    n278,
    n223
  );


  xnor
  g1406
  (
    n1379,
    n495,
    n458,
    n376,
    n285
  );


  or
  g1407
  (
    n1472,
    n414,
    n326,
    n212,
    n449
  );


  xor
  g1408
  (
    n1141,
    n276,
    n450,
    n425,
    n242
  );


  or
  g1409
  (
    n916,
    n223,
    n269,
    n596,
    n575
  );


  xor
  g1410
  (
    n831,
    n600,
    n649,
    n428,
    n399
  );


  xor
  g1411
  (
    n990,
    n565,
    n641,
    n386,
    n514
  );


  nand
  g1412
  (
    n1255,
    n486,
    n584,
    n581,
    n545
  );


  xnor
  g1413
  (
    n1015,
    n279,
    n635,
    n516,
    n386
  );


  xnor
  g1414
  (
    n1177,
    n281,
    n356,
    n551,
    n215
  );


  xor
  g1415
  (
    n980,
    n420,
    n348,
    n380,
    n411
  );


  xor
  g1416
  (
    n1437,
    n571,
    n496,
    n267,
    n407
  );


  xnor
  g1417
  (
    n1178,
    n627,
    n421,
    n315,
    n306
  );


  nor
  g1418
  (
    n861,
    n617,
    n612,
    n309,
    n566
  );


  nand
  g1419
  (
    n778,
    n245,
    n299,
    n234,
    n546
  );


  and
  g1420
  (
    n1445,
    n232,
    n378,
    n257,
    n464
  );


  nor
  g1421
  (
    n1376,
    n540,
    n324,
    n572,
    n265
  );


  nand
  g1422
  (
    n1013,
    n661,
    n252,
    n628,
    n473
  );


  and
  g1423
  (
    n1007,
    n482,
    n669,
    n386,
    n282
  );


  xnor
  g1424
  (
    n966,
    n321,
    n528,
    n414,
    n212
  );


  and
  g1425
  (
    n1124,
    n456,
    n471,
    n479,
    n426
  );


  xor
  g1426
  (
    n1317,
    n490,
    n550,
    n200,
    n655
  );


  xor
  g1427
  (
    n1304,
    n549,
    n612,
    n462,
    n193
  );


  xnor
  g1428
  (
    n788,
    n419,
    n622,
    n361,
    n323
  );


  nor
  g1429
  (
    n1276,
    n421,
    n288,
    n380,
    n338
  );


  nand
  g1430
  (
    n1088,
    n293,
    n223,
    n595,
    n206
  );


  or
  g1431
  (
    n798,
    n483,
    n334,
    n383,
    n207
  );


  nand
  g1432
  (
    n1306,
    n608,
    n468,
    n353,
    n377
  );


  nand
  g1433
  (
    n1266,
    n178,
    n570,
    n648,
    n208
  );


  and
  g1434
  (
    n1302,
    n611,
    n368,
    n241,
    n511
  );


  or
  g1435
  (
    n1031,
    n187,
    n204,
    n431,
    n207
  );


  and
  g1436
  (
    n773,
    n494,
    n602,
    n420,
    n196
  );


  nor
  g1437
  (
    n1402,
    n595,
    n373,
    n194,
    n198
  );


  or
  g1438
  (
    n1184,
    n191,
    n301,
    n589,
    n588
  );


  xnor
  g1439
  (
    n1492,
    n422,
    n410,
    n650,
    n179
  );


  nand
  g1440
  (
    n1206,
    n554,
    n328,
    n438,
    n658
  );


  or
  g1441
  (
    n696,
    n337,
    n451,
    n223,
    n263
  );


  xnor
  g1442
  (
    n1408,
    n487,
    n168,
    n557,
    n654
  );


  xnor
  g1443
  (
    n692,
    n645,
    n503,
    n536,
    n509
  );


  xnor
  g1444
  (
    n901,
    n522,
    n349,
    n593,
    n209
  );


  nand
  g1445
  (
    n1382,
    n366,
    n471,
    n541,
    n563
  );


  xnor
  g1446
  (
    n1196,
    n524,
    n201,
    n667,
    n251
  );


  nor
  g1447
  (
    n1350,
    n436,
    n602,
    n619,
    n307
  );


  or
  g1448
  (
    n850,
    n576,
    n504,
    n648,
    n376
  );


  nor
  g1449
  (
    n730,
    n647,
    n294,
    n555,
    n211
  );


  xor
  g1450
  (
    n1259,
    n175,
    n396,
    n515,
    n180
  );


  xnor
  g1451
  (
    n1487,
    n341,
    n659,
    n330,
    n335
  );


  nand
  g1452
  (
    n799,
    n272,
    n562,
    n413,
    n493
  );


  nand
  g1453
  (
    n686,
    n634,
    n435,
    n300,
    n221
  );


  nand
  g1454
  (
    n1489,
    n570,
    n433,
    n291,
    n292
  );


  nor
  g1455
  (
    n796,
    n594,
    n400,
    n333,
    n325
  );


  or
  g1456
  (
    n1216,
    n516,
    n211,
    n511,
    n164
  );


  or
  g1457
  (
    n736,
    n306,
    n567,
    n447,
    n569
  );


  xnor
  g1458
  (
    n1418,
    n592,
    n631,
    n573,
    n181
  );


  nor
  g1459
  (
    n1090,
    n388,
    n596,
    n427,
    n199
  );


  nor
  g1460
  (
    n1394,
    n447,
    n294,
    n631,
    n238
  );


  xor
  g1461
  (
    n803,
    n579,
    n510,
    n538,
    n533
  );


  nor
  g1462
  (
    n828,
    n393,
    n179,
    n559,
    n606
  );


  xor
  g1463
  (
    n1020,
    n454,
    n649,
    n593,
    n354
  );


  nor
  g1464
  (
    n1319,
    n254,
    n304,
    n328,
    n586
  );


  and
  g1465
  (
    n1358,
    n527,
    n480,
    n351,
    n286
  );


  xnor
  g1466
  (
    n1404,
    n226,
    n184,
    n536,
    n565
  );


  or
  g1467
  (
    n1202,
    n243,
    n527,
    n256,
    n247
  );


  nand
  g1468
  (
    n1260,
    n623,
    n298,
    n313,
    n189
  );


  and
  g1469
  (
    n878,
    n611,
    n518,
    n171,
    n302
  );


  nor
  g1470
  (
    n1328,
    n351,
    n189,
    n594,
    n230
  );


  xnor
  g1471
  (
    n821,
    n617,
    n348,
    n471,
    n190
  );


  and
  g1472
  (
    n1062,
    n416,
    n257,
    n420,
    n367
  );


  nand
  g1473
  (
    n1128,
    n664,
    n449,
    n606
  );


  nor
  g1474
  (
    n1278,
    n174,
    n220,
    n442,
    n482
  );


  xnor
  g1475
  (
    n872,
    n502,
    n463,
    n558,
    n298
  );


  xor
  g1476
  (
    n1567,
    n1288,
    n784,
    n1270,
    n971
  );


  or
  g1477
  (
    n1692,
    n921,
    n1383,
    n919,
    n1394
  );


  or
  g1478
  (
    n1716,
    n1320,
    n1019,
    n689,
    n697
  );


  xnor
  g1479
  (
    n1611,
    n814,
    n942,
    n868,
    n764
  );


  nand
  g1480
  (
    n1657,
    n1252,
    n1022,
    n840,
    n759
  );


  or
  g1481
  (
    n1694,
    n1494,
    n1221,
    n748,
    n928
  );


  nand
  g1482
  (
    n1690,
    n1009,
    n1406,
    n1445,
    n1005
  );


  nor
  g1483
  (
    n1645,
    n1124,
    n904,
    n1430,
    n973
  );


  xnor
  g1484
  (
    n1672,
    n1021,
    n968,
    n685,
    n1246
  );


  nand
  g1485
  (
    n1678,
    n1032,
    n747,
    n714,
    n986
  );


  or
  g1486
  (
    n1558,
    n1327,
    n873,
    n1219,
    n930
  );


  nor
  g1487
  (
    n1531,
    n1467,
    n982,
    n954,
    n1042
  );


  or
  g1488
  (
    n1658,
    n831,
    n1287,
    n789,
    n1249
  );


  and
  g1489
  (
    n1516,
    n965,
    n1055,
    n1163,
    n679
  );


  xor
  g1490
  (
    n1615,
    n1261,
    n1492,
    n1217,
    n737
  );


  and
  g1491
  (
    n1579,
    n754,
    n755,
    n843,
    n1096
  );


  xor
  g1492
  (
    n1613,
    n1197,
    n1420,
    n774,
    n966
  );


  nor
  g1493
  (
    n1556,
    n1179,
    n1316,
    n884,
    n981
  );


  and
  g1494
  (
    n1619,
    n1384,
    n1385,
    n1321,
    n984
  );


  xor
  g1495
  (
    n1641,
    n802,
    n1356,
    n993,
    n1285
  );


  nor
  g1496
  (
    n1626,
    n687,
    n1284,
    n1489,
    n864
  );


  nand
  g1497
  (
    n1515,
    n1426,
    n1110,
    n866,
    n1157
  );


  or
  g1498
  (
    n1527,
    n1235,
    n1460,
    n1162,
    n943
  );


  xor
  g1499
  (
    n1532,
    n1264,
    n1132,
    n811,
    n886
  );


  or
  g1500
  (
    n1595,
    n1154,
    n1414,
    n1410,
    n1324
  );


  and
  g1501
  (
    n1715,
    n1073,
    n1029,
    n1388,
    n901
  );


  xor
  g1502
  (
    n1517,
    n1160,
    n1381,
    n1033,
    n703
  );


  nand
  g1503
  (
    n1636,
    n1234,
    n1375,
    n847,
    n959
  );


  xnor
  g1504
  (
    n1679,
    n997,
    n1496,
    n1165,
    n990
  );


  or
  g1505
  (
    n1589,
    n1215,
    n941,
    n1178,
    n974
  );


  nand
  g1506
  (
    n1696,
    n1501,
    n1499,
    n918,
    n807
  );


  and
  g1507
  (
    n1709,
    n785,
    n1277,
    n1440,
    n760
  );


  or
  g1508
  (
    n1540,
    n900,
    n936,
    n1167,
    n684
  );


  or
  g1509
  (
    n1536,
    n1276,
    n1501,
    n1408,
    n1074
  );


  or
  g1510
  (
    n1684,
    n793,
    n1002,
    n1101,
    n1245
  );


  nand
  g1511
  (
    n1622,
    n882,
    n1115,
    n1172,
    n1208
  );


  xor
  g1512
  (
    n1616,
    n1044,
    n1407,
    n960,
    n1150
  );


  nor
  g1513
  (
    n1566,
    n1393,
    n850,
    n826,
    n915
  );


  and
  g1514
  (
    n1618,
    n1243,
    n1098,
    n751,
    n835
  );


  or
  g1515
  (
    n1583,
    n875,
    n1299,
    n1065,
    n989
  );


  xor
  g1516
  (
    n1648,
    n768,
    n1006,
    n1199,
    n828
  );


  nor
  g1517
  (
    n1565,
    n979,
    n792,
    n682,
    n795
  );


  nand
  g1518
  (
    n1581,
    n842,
    n1118,
    n1143,
    n1242
  );


  xor
  g1519
  (
    n1548,
    n1409,
    n934,
    n1402,
    n1418
  );


  xnor
  g1520
  (
    n1545,
    n1224,
    n1386,
    n1265,
    n1366
  );


  nor
  g1521
  (
    n1651,
    n1419,
    n818,
    n1416,
    n681
  );


  nand
  g1522
  (
    n1599,
    n863,
    n1020,
    n1175,
    n956
  );


  xor
  g1523
  (
    n1713,
    n1293,
    n1308,
    n1369,
    n937
  );


  or
  g1524
  (
    n1546,
    n1377,
    n1348,
    n719,
    n933
  );


  or
  g1525
  (
    n1659,
    n721,
    n991,
    n1100,
    n1198
  );


  nand
  g1526
  (
    n1711,
    n1345,
    n694,
    n765,
    n1269
  );


  xor
  g1527
  (
    n1642,
    n1423,
    n1341,
    n1183,
    n1099
  );


  or
  g1528
  (
    n1551,
    n1278,
    n1194,
    n1336,
    n976
  );


  and
  g1529
  (
    n1597,
    n995,
    n1403,
    n844,
    n1257
  );


  nor
  g1530
  (
    n1509,
    n822,
    n674,
    n683,
    n762
  );


  or
  g1531
  (
    n1529,
    n1010,
    n962,
    n806,
    n1184
  );


  nor
  g1532
  (
    n1701,
    n810,
    n1429,
    n1425,
    n961
  );


  nand
  g1533
  (
    n1568,
    n1411,
    n895,
    n829,
    n1023
  );


  xnor
  g1534
  (
    n1654,
    n1181,
    n1361,
    n848,
    n1247
  );


  xor
  g1535
  (
    n1510,
    n996,
    n1240,
    n1030,
    n841
  );


  xor
  g1536
  (
    n1526,
    n1059,
    n1086,
    n756,
    n1189
  );


  or
  g1537
  (
    n1530,
    n927,
    n1213,
    n1084,
    n1093
  );


  xnor
  g1538
  (
    n1564,
    n1202,
    n1012,
    n1380,
    n838
  );


  or
  g1539
  (
    n1535,
    n1041,
    n914,
    n770,
    n1360
  );


  or
  g1540
  (
    n1680,
    n1130,
    n923,
    n1045,
    n1289
  );


  nor
  g1541
  (
    n1649,
    n947,
    n820,
    n913,
    n1335
  );


  xor
  g1542
  (
    n1561,
    n897,
    n1347,
    n1436,
    n1103
  );


  xnor
  g1543
  (
    n1699,
    n704,
    n733,
    n776,
    n1122
  );


  or
  g1544
  (
    n1643,
    n1333,
    n790,
    n1034,
    n1260
  );


  nand
  g1545
  (
    n1698,
    n1142,
    n1129,
    n1050,
    n1151
  );


  or
  g1546
  (
    n1646,
    n780,
    n1112,
    n1200,
    n1368
  );


  nand
  g1547
  (
    n1668,
    n722,
    n1295,
    n1433,
    n805
  );


  and
  g1548
  (
    n1537,
    n1483,
    n769,
    n1001,
    n1185
  );


  nor
  g1549
  (
    n1604,
    n1363,
    n1229,
    n720,
    n808
  );


  nand
  g1550
  (
    n1630,
    n1051,
    n912,
    n1227,
    n1049
  );


  xor
  g1551
  (
    n1519,
    n1382,
    n839,
    n1232,
    n1353
  );


  nand
  g1552
  (
    n1596,
    n783,
    n1095,
    n909,
    n1451
  );


  or
  g1553
  (
    n1640,
    n1474,
    n1271,
    n1392,
    n1313
  );


  nand
  g1554
  (
    n1559,
    n1486,
    n1091,
    n1447,
    n696
  );


  xor
  g1555
  (
    n1600,
    n1127,
    n1067,
    n753,
    n1241
  );


  and
  g1556
  (
    n1691,
    n1139,
    n1135,
    n1456,
    n861
  );


  or
  g1557
  (
    n1573,
    n1155,
    n1236,
    n824,
    n1343
  );


  and
  g1558
  (
    n1562,
    n1226,
    n1144,
    n920,
    n778
  );


  nor
  g1559
  (
    n1703,
    n1253,
    n876,
    n1087,
    n1290
  );


  and
  g1560
  (
    n1670,
    n732,
    n1203,
    n1294,
    n1117
  );


  nor
  g1561
  (
    n1514,
    n1092,
    n1003,
    n1319,
    n975
  );


  nor
  g1562
  (
    n1550,
    n711,
    n1334,
    n1475,
    n1216
  );


  nor
  g1563
  (
    n1598,
    n1116,
    n1431,
    n1318,
    n728
  );


  nor
  g1564
  (
    n1666,
    n1309,
    n924,
    n1088,
    n1070
  );


  nand
  g1565
  (
    n1702,
    n1370,
    n899,
    n1259,
    n1036
  );


  xor
  g1566
  (
    n1712,
    n1491,
    n1105,
    n1066,
    n1441
  );


  or
  g1567
  (
    n1655,
    n834,
    n1106,
    n929,
    n750
  );


  xnor
  g1568
  (
    n1588,
    n1444,
    n1013,
    n825,
    n1238
  );


  nor
  g1569
  (
    n1534,
    n1109,
    n1297,
    n977,
    n1428
  );


  and
  g1570
  (
    n1586,
    n1258,
    n1282,
    n1137,
    n1323
  );


  xor
  g1571
  (
    n1625,
    n1193,
    n1108,
    n857,
    n891
  );


  xnor
  g1572
  (
    n1542,
    n856,
    n1164,
    n1374,
    n1176
  );


  xnor
  g1573
  (
    n1523,
    n1471,
    n763,
    n1169,
    n1090
  );


  xor
  g1574
  (
    n1681,
    n731,
    n1272,
    n1121,
    n893
  );


  or
  g1575
  (
    n1677,
    n1082,
    n1302,
    n987,
    n1040
  );


  and
  g1576
  (
    n1632,
    n1396,
    n1104,
    n745,
    n1046
  );


  xnor
  g1577
  (
    n1620,
    n678,
    n1330,
    n1404,
    n902
  );


  and
  g1578
  (
    n1639,
    n816,
    n1391,
    n1018,
    n1296
  );


  xor
  g1579
  (
    n1660,
    n1493,
    n761,
    n1415,
    n1220
  );


  nand
  g1580
  (
    n1673,
    n1079,
    n1329,
    n837,
    n1379
  );


  nand
  g1581
  (
    KeyWire_0_1,
    n707,
    n1254,
    n1482,
    n879
  );


  nand
  g1582
  (
    n1555,
    n1083,
    n1071,
    n1057,
    n1301
  );


  and
  g1583
  (
    n1675,
    n1286,
    n1291,
    n1281,
    n1028
  );


  or
  g1584
  (
    n1631,
    n1180,
    n1283,
    n948,
    n992
  );


  nor
  g1585
  (
    n1671,
    n827,
    n1187,
    n782,
    n906
  );


  nor
  g1586
  (
    n1528,
    n1279,
    n691,
    n1113,
    n926
  );


  xor
  g1587
  (
    n1682,
    n1039,
    n967,
    n777,
    n740
  );


  xor
  g1588
  (
    n1656,
    n1463,
    n1325,
    n1468,
    n862
  );


  nand
  g1589
  (
    n1635,
    n1047,
    n1089,
    n1478,
    n729
  );


  nand
  g1590
  (
    n1584,
    n1459,
    n1417,
    n1053,
    n889
  );


  xnor
  g1591
  (
    n1617,
    n1263,
    n985,
    n1058,
    n686
  );


  xnor
  g1592
  (
    n1544,
    n1500,
    n855,
    n1223,
    n1307
  );


  xnor
  g1593
  (
    n1661,
    n677,
    n758,
    n1367,
    n1111
  );


  nand
  g1594
  (
    n1521,
    n980,
    n1170,
    n1437,
    n724
  );


  or
  g1595
  (
    n1689,
    n1008,
    n970,
    n903,
    n1310
  );


  xor
  g1596
  (
    n1563,
    n885,
    n1351,
    n1357,
    n713
  );


  or
  g1597
  (
    n1601,
    n1401,
    n712,
    n949,
    n1472
  );


  xor
  g1598
  (
    n1614,
    n1371,
    n1097,
    n766,
    n1068
  );


  xnor
  g1599
  (
    n1663,
    n821,
    n860,
    n1488,
    n1056
  );


  xor
  g1600
  (
    n1697,
    n922,
    n1275,
    n925,
    n1114
  );


  nand
  g1601
  (
    n1533,
    n1233,
    n1063,
    n775,
    n950
  );


  xnor
  g1602
  (
    n1578,
    n1485,
    n1487,
    n972,
    n1432
  );


  and
  g1603
  (
    n1553,
    n1182,
    n1075,
    n1495,
    n953
  );


  or
  g1604
  (
    n1638,
    n788,
    n1077,
    n705,
    n951
  );


  nand
  g1605
  (
    n1522,
    n1438,
    n892,
    n1457,
    n1126
  );


  or
  g1606
  (
    n1554,
    n695,
    n1133,
    n1349,
    n852
  );


  xnor
  g1607
  (
    n1539,
    n1048,
    n1465,
    n1214,
    n699
  );


  nand
  g1608
  (
    n1714,
    n858,
    n1128,
    n801,
    n794
  );


  nor
  g1609
  (
    n1585,
    n1119,
    n1473,
    n692,
    n871
  );


  xor
  g1610
  (
    n1577,
    n1365,
    n1266,
    n1443,
    n1145
  );


  nand
  g1611
  (
    n1688,
    n716,
    n1267,
    n1340,
    n817
  );


  or
  g1612
  (
    n1549,
    n1421,
    n1346,
    n738,
    n1156
  );


  or
  g1613
  (
    n1628,
    n1054,
    n1204,
    n883,
    n1205
  );


  or
  g1614
  (
    n1710,
    n1373,
    n1458,
    n1314,
    n1354
  );


  or
  g1615
  (
    n1524,
    n1424,
    n787,
    n1031,
    n1102
  );


  or
  g1616
  (
    n1706,
    n1141,
    n823,
    n877,
    n1280
  );


  and
  g1617
  (
    n1647,
    n888,
    n932,
    n1362,
    n796
  );


  nor
  g1618
  (
    n1602,
    n1484,
    n1338,
    n1399,
    n1120
  );


  xnor
  g1619
  (
    n1612,
    n1490,
    n978,
    n1298,
    n894
  );


  and
  g1620
  (
    n1541,
    n1094,
    n1435,
    n815,
    n1397
  );


  nor
  g1621
  (
    n1592,
    n1427,
    n1081,
    n1177,
    n1337
  );


  nor
  g1622
  (
    n1574,
    n700,
    n742,
    n1251,
    n994
  );


  or
  g1623
  (
    n1609,
    n1376,
    n1140,
    n1107,
    n1387
  );


  or
  g1624
  (
    n1571,
    n786,
    n1211,
    n1466,
    n800
  );


  xnor
  g1625
  (
    n1605,
    n708,
    n741,
    n846,
    n791
  );


  xnor
  g1626
  (
    n1610,
    n917,
    n1480,
    n1372,
    n1007
  );


  nor
  g1627
  (
    n1685,
    n767,
    n1123,
    n1125,
    n969
  );


  nor
  g1628
  (
    n1569,
    n1452,
    n819,
    n1210,
    n1025
  );


  nand
  g1629
  (
    n1704,
    n905,
    n1331,
    n1461,
    n1476
  );


  xor
  g1630
  (
    KeyWire_0_2,
    n1317,
    n725,
    n809,
    n749
  );


  nor
  g1631
  (
    n1525,
    n1000,
    n1448,
    n1153,
    n1359
  );


  xnor
  g1632
  (
    n1518,
    n735,
    n1477,
    n1136,
    n1218
  );


  nor
  g1633
  (
    n1603,
    n726,
    n1188,
    n1501,
    n908
  );


  xor
  g1634
  (
    n1538,
    n715,
    n1171,
    n867,
    n1131
  );


  or
  g1635
  (
    n1644,
    n693,
    n675,
    n1239,
    n1352
  );


  nor
  g1636
  (
    n1572,
    n1434,
    n803,
    n1231,
    n1152
  );


  nor
  g1637
  (
    n1634,
    n1225,
    n1061,
    n1332,
    n1052
  );


  xor
  g1638
  (
    n1637,
    n870,
    n710,
    n958,
    n1207
  );


  xor
  g1639
  (
    n1520,
    n1389,
    n881,
    n832,
    n1481
  );


  nand
  g1640
  (
    n1683,
    n1305,
    n880,
    n952,
    n1442
  );


  or
  g1641
  (
    n1607,
    n718,
    n890,
    n836,
    n1147
  );


  nor
  g1642
  (
    n1513,
    n773,
    n1148,
    n1405,
    n723
  );


  xnor
  g1643
  (
    n1627,
    n1292,
    n944,
    n946,
    n1268
  );


  nor
  g1644
  (
    n1608,
    n701,
    n1395,
    n676,
    n939
  );


  xor
  g1645
  (
    n1590,
    n1026,
    n1038,
    n1439,
    n911
  );


  nor
  g1646
  (
    n1674,
    n673,
    n887,
    n845,
    n1390
  );


  and
  g1647
  (
    n1593,
    n1174,
    n813,
    n688,
    n1422
  );


  nand
  g1648
  (
    n1543,
    n1024,
    n771,
    n757,
    n898
  );


  xnor
  g1649
  (
    n1580,
    n1138,
    n833,
    n1322,
    n963
  );


  xnor
  g1650
  (
    n1695,
    n799,
    n1355,
    n709,
    n907
  );


  nand
  g1651
  (
    n1669,
    n746,
    n1446,
    n1454,
    n853
  );


  nor
  g1652
  (
    n1591,
    n916,
    n935,
    n854,
    n999
  );


  and
  g1653
  (
    n1606,
    n1015,
    n706,
    n1350,
    n1469
  );


  and
  g1654
  (
    n1633,
    n1146,
    n1035,
    n1158,
    n896
  );


  nand
  g1655
  (
    n1512,
    n730,
    n910,
    n1168,
    n957
  );


  and
  g1656
  (
    n1557,
    n1072,
    n1449,
    n938,
    n1470
  );


  or
  g1657
  (
    n1629,
    n1064,
    n1237,
    n964,
    n1255
  );


  or
  g1658
  (
    n1650,
    n1250,
    n931,
    n1501,
    n998
  );


  xor
  g1659
  (
    n1687,
    n1016,
    n1195,
    n812,
    n851
  );


  nor
  g1660
  (
    n1667,
    n798,
    n1230,
    n945,
    n1378
  );


  nor
  g1661
  (
    n1570,
    n1027,
    n772,
    n1413,
    n878
  );


  or
  g1662
  (
    n1552,
    n869,
    n797,
    n1306,
    n1339
  );


  or
  g1663
  (
    n1686,
    n1190,
    n874,
    n1244,
    n1479
  );


  nand
  g1664
  (
    n1560,
    n1300,
    n1069,
    n1166,
    n1398
  );


  xor
  g1665
  (
    n1665,
    n1315,
    n988,
    n1186,
    n1206
  );


  or
  g1666
  (
    n1653,
    n1060,
    n1159,
    n1273,
    n1173
  );


  xor
  g1667
  (
    n1582,
    n1209,
    n1326,
    n1080,
    n1192
  );


  nand
  g1668
  (
    n1676,
    n1222,
    n1196,
    n1364,
    n698
  );


  xor
  g1669
  (
    n1575,
    n1274,
    n1212,
    n1149,
    n680
  );


  nor
  g1670
  (
    n1700,
    n1256,
    n849,
    n804,
    n752
  );


  xnor
  g1671
  (
    n1576,
    n1076,
    n830,
    n1085,
    n1455
  );


  or
  g1672
  (
    n1511,
    n734,
    n744,
    n955,
    n736
  );


  or
  g1673
  (
    n1693,
    n1134,
    n1248,
    n1342,
    n690
  );


  and
  g1674
  (
    n1662,
    n1228,
    n1017,
    n1004,
    n865
  );


  or
  g1675
  (
    n1624,
    n1453,
    n1043,
    n702,
    n1450
  );


  nand
  g1676
  (
    n1621,
    n940,
    n1344,
    n872,
    n739
  );


  nand
  g1677
  (
    n1587,
    n1078,
    n1191,
    n717,
    n1262
  );


  xnor
  g1678
  (
    n1708,
    n983,
    n727,
    n1497,
    n781
  );


  and
  g1679
  (
    n1652,
    n743,
    n1412,
    n1311,
    n1011
  );


  nor
  g1680
  (
    n1707,
    n1037,
    n1201,
    n1303,
    n1328
  );


  or
  g1681
  (
    n1705,
    n1462,
    n859,
    n1062,
    n1161
  );


  and
  g1682
  (
    n1594,
    n1312,
    n1014,
    n1304,
    n1400
  );


  xor
  g1683
  (
    n1623,
    n1498,
    n779,
    n1464,
    n1358
  );


  not
  g1684
  (
    n1944,
    n1546
  );


  not
  g1685
  (
    n1792,
    n1528
  );


  buf
  g1686
  (
    n2045,
    n1510
  );


  buf
  g1687
  (
    n1896,
    n1629
  );


  buf
  g1688
  (
    n2029,
    n1517
  );


  not
  g1689
  (
    n1753,
    n1671
  );


  not
  g1690
  (
    n1804,
    n1626
  );


  not
  g1691
  (
    n1966,
    n1528
  );


  not
  g1692
  (
    n1921,
    n1632
  );


  buf
  g1693
  (
    n2211,
    n1515
  );


  buf
  g1694
  (
    n1904,
    n1642
  );


  not
  g1695
  (
    n2102,
    n1538
  );


  buf
  g1696
  (
    n2153,
    n1557
  );


  buf
  g1697
  (
    n1809,
    n1533
  );


  buf
  g1698
  (
    n1721,
    n1649
  );


  not
  g1699
  (
    KeyWire_0_12,
    n1556
  );


  not
  g1700
  (
    n1852,
    n1606
  );


  not
  g1701
  (
    n2196,
    n1645
  );


  not
  g1702
  (
    n1913,
    n1543
  );


  not
  g1703
  (
    n2210,
    n1553
  );


  not
  g1704
  (
    n1854,
    n1671
  );


  not
  g1705
  (
    n1801,
    n1522
  );


  not
  g1706
  (
    n2048,
    n1607
  );


  not
  g1707
  (
    n2152,
    n1582
  );


  buf
  g1708
  (
    n1786,
    n1620
  );


  not
  g1709
  (
    n2138,
    n1587
  );


  buf
  g1710
  (
    n1848,
    n1662
  );


  buf
  g1711
  (
    n1937,
    n1614
  );


  not
  g1712
  (
    n2109,
    n1607
  );


  not
  g1713
  (
    n1898,
    n1510
  );


  buf
  g1714
  (
    n2177,
    n1571
  );


  not
  g1715
  (
    n2189,
    n1624
  );


  buf
  g1716
  (
    n1778,
    n1532
  );


  not
  g1717
  (
    n2022,
    n1558
  );


  buf
  g1718
  (
    n2169,
    n1611
  );


  not
  g1719
  (
    n2005,
    n1576
  );


  buf
  g1720
  (
    n2155,
    n1647
  );


  buf
  g1721
  (
    n1925,
    n1515
  );


  buf
  g1722
  (
    n1763,
    n1639
  );


  not
  g1723
  (
    n2150,
    n1645
  );


  buf
  g1724
  (
    n1872,
    n1637
  );


  buf
  g1725
  (
    n1874,
    n1595
  );


  not
  g1726
  (
    n1783,
    n1644
  );


  buf
  g1727
  (
    n1779,
    n1670
  );


  not
  g1728
  (
    n1907,
    n1515
  );


  buf
  g1729
  (
    n1719,
    n1541
  );


  buf
  g1730
  (
    n2052,
    n1551
  );


  buf
  g1731
  (
    n2069,
    n1538
  );


  buf
  g1732
  (
    n1948,
    n1638
  );


  buf
  g1733
  (
    n2062,
    n1579
  );


  buf
  g1734
  (
    n1892,
    n1611
  );


  not
  g1735
  (
    n1916,
    n1548
  );


  not
  g1736
  (
    n1806,
    n1670
  );


  not
  g1737
  (
    n1875,
    n1617
  );


  not
  g1738
  (
    n2188,
    n1654
  );


  buf
  g1739
  (
    n1825,
    n1565
  );


  not
  g1740
  (
    n1762,
    n1615
  );


  not
  g1741
  (
    n2122,
    n1646
  );


  not
  g1742
  (
    n1794,
    n1525
  );


  buf
  g1743
  (
    n1782,
    n1580
  );


  not
  g1744
  (
    n2010,
    n1621
  );


  not
  g1745
  (
    n1994,
    n1548
  );


  buf
  g1746
  (
    n1769,
    n1550
  );


  not
  g1747
  (
    n2175,
    n1509
  );


  not
  g1748
  (
    n2217,
    n1604
  );


  buf
  g1749
  (
    n2146,
    n1661
  );


  buf
  g1750
  (
    n1850,
    n1623
  );


  buf
  g1751
  (
    n1957,
    n1657
  );


  buf
  g1752
  (
    n1985,
    n1659
  );


  not
  g1753
  (
    n2149,
    n1633
  );


  not
  g1754
  (
    n2162,
    n1539
  );


  buf
  g1755
  (
    n1968,
    n1530
  );


  not
  g1756
  (
    n2186,
    n1554
  );


  buf
  g1757
  (
    n1755,
    n1669
  );


  buf
  g1758
  (
    n1929,
    n1650
  );


  buf
  g1759
  (
    n1918,
    n1558
  );


  buf
  g1760
  (
    n2070,
    n1562
  );


  buf
  g1761
  (
    n2118,
    n1528
  );


  not
  g1762
  (
    n1775,
    n1520
  );


  buf
  g1763
  (
    n2013,
    n1572
  );


  not
  g1764
  (
    n1747,
    n1600
  );


  not
  g1765
  (
    n1839,
    n1667
  );


  buf
  g1766
  (
    n1866,
    n1565
  );


  buf
  g1767
  (
    n1784,
    n1592
  );


  not
  g1768
  (
    n2044,
    n1540
  );


  not
  g1769
  (
    n1882,
    n1650
  );


  not
  g1770
  (
    n1869,
    n1650
  );


  not
  g1771
  (
    n2023,
    n1616
  );


  not
  g1772
  (
    n2043,
    n1577
  );


  not
  g1773
  (
    n1761,
    n1558
  );


  not
  g1774
  (
    n2063,
    n1587
  );


  buf
  g1775
  (
    n1733,
    n1660
  );


  buf
  g1776
  (
    n1973,
    n1596
  );


  buf
  g1777
  (
    n2220,
    n1556
  );


  not
  g1778
  (
    n1991,
    n1663
  );


  buf
  g1779
  (
    n2132,
    n1540
  );


  buf
  g1780
  (
    n1876,
    n1557
  );


  not
  g1781
  (
    n1780,
    n1570
  );


  not
  g1782
  (
    n1902,
    n1545
  );


  not
  g1783
  (
    n1971,
    n1614
  );


  not
  g1784
  (
    n2086,
    n1624
  );


  buf
  g1785
  (
    n1956,
    n1597
  );


  buf
  g1786
  (
    n2130,
    n1530
  );


  buf
  g1787
  (
    n1964,
    n1608
  );


  buf
  g1788
  (
    n1886,
    n1572
  );


  not
  g1789
  (
    KeyWire_0_11,
    n1531
  );


  not
  g1790
  (
    n2190,
    n1589
  );


  buf
  g1791
  (
    n2215,
    n1636
  );


  buf
  g1792
  (
    n1742,
    n1580
  );


  not
  g1793
  (
    n1770,
    n1548
  );


  not
  g1794
  (
    n2075,
    n1642
  );


  buf
  g1795
  (
    n2124,
    n1622
  );


  not
  g1796
  (
    n2147,
    n1534
  );


  not
  g1797
  (
    n1877,
    n1610
  );


  not
  g1798
  (
    n1795,
    n1610
  );


  buf
  g1799
  (
    n2142,
    n1596
  );


  not
  g1800
  (
    n2046,
    n1569
  );


  not
  g1801
  (
    n1920,
    n1628
  );


  not
  g1802
  (
    n1952,
    n1565
  );


  buf
  g1803
  (
    n1989,
    n1645
  );


  not
  g1804
  (
    n1807,
    n1601
  );


  not
  g1805
  (
    n2145,
    n1589
  );


  not
  g1806
  (
    n1776,
    n1613
  );


  buf
  g1807
  (
    n2207,
    n1520
  );


  not
  g1808
  (
    n1894,
    n1595
  );


  not
  g1809
  (
    n2158,
    n1654
  );


  not
  g1810
  (
    n2135,
    n1586
  );


  buf
  g1811
  (
    n2038,
    n1590
  );


  not
  g1812
  (
    n2055,
    n1630
  );


  not
  g1813
  (
    n2097,
    n1559
  );


  buf
  g1814
  (
    n1828,
    n1627
  );


  not
  g1815
  (
    n1914,
    n1536
  );


  not
  g1816
  (
    n1924,
    n1627
  );


  buf
  g1817
  (
    n1734,
    n1568
  );


  buf
  g1818
  (
    n2057,
    n1624
  );


  buf
  g1819
  (
    n1889,
    n1613
  );


  not
  g1820
  (
    n1865,
    n1557
  );


  not
  g1821
  (
    n2164,
    n1672
  );


  buf
  g1822
  (
    n1931,
    n1527
  );


  buf
  g1823
  (
    n2068,
    n1535
  );


  buf
  g1824
  (
    n2119,
    n1583
  );


  buf
  g1825
  (
    n1815,
    n1598
  );


  not
  g1826
  (
    n1899,
    n1588
  );


  not
  g1827
  (
    n2095,
    n1575
  );


  buf
  g1828
  (
    n1908,
    n1517
  );


  not
  g1829
  (
    n1977,
    n1590
  );


  buf
  g1830
  (
    n2128,
    n1551
  );


  buf
  g1831
  (
    n2017,
    n1656
  );


  not
  g1832
  (
    n2085,
    n1521
  );


  buf
  g1833
  (
    n2194,
    n1603
  );


  buf
  g1834
  (
    n1960,
    n1559
  );


  buf
  g1835
  (
    n2099,
    n1526
  );


  buf
  g1836
  (
    n2157,
    n1552
  );


  buf
  g1837
  (
    n2137,
    n1567
  );


  not
  g1838
  (
    n2131,
    n1661
  );


  not
  g1839
  (
    n2074,
    n1524
  );


  buf
  g1840
  (
    n2006,
    n1664
  );


  not
  g1841
  (
    n2081,
    n1649
  );


  buf
  g1842
  (
    n1810,
    n1663
  );


  buf
  g1843
  (
    n1954,
    n1549
  );


  not
  g1844
  (
    n2178,
    n1541
  );


  buf
  g1845
  (
    n2028,
    n1595
  );


  buf
  g1846
  (
    n2064,
    n1522
  );


  not
  g1847
  (
    n2192,
    n1619
  );


  not
  g1848
  (
    n1917,
    n1578
  );


  buf
  g1849
  (
    n2101,
    n1509
  );


  not
  g1850
  (
    n2144,
    n1665
  );


  not
  g1851
  (
    n2092,
    n1524
  );


  buf
  g1852
  (
    n2042,
    n1642
  );


  not
  g1853
  (
    n1945,
    n1516
  );


  not
  g1854
  (
    n1867,
    n1641
  );


  buf
  g1855
  (
    n1981,
    n1537
  );


  buf
  g1856
  (
    n2143,
    n1661
  );


  buf
  g1857
  (
    n1912,
    n1665
  );


  not
  g1858
  (
    n1791,
    n1564
  );


  not
  g1859
  (
    n2051,
    n1651
  );


  buf
  g1860
  (
    n1789,
    n1544
  );


  buf
  g1861
  (
    n1950,
    n1593
  );


  not
  g1862
  (
    n1717,
    n1543
  );


  buf
  g1863
  (
    n1802,
    n1583
  );


  buf
  g1864
  (
    n1843,
    n1596
  );


  not
  g1865
  (
    n1861,
    n1544
  );


  not
  g1866
  (
    n2203,
    n1600
  );


  buf
  g1867
  (
    n2026,
    n1579
  );


  buf
  g1868
  (
    n1891,
    n1513
  );


  buf
  g1869
  (
    n1765,
    n1541
  );


  not
  g1870
  (
    n1987,
    n1586
  );


  not
  g1871
  (
    n1943,
    n1653
  );


  buf
  g1872
  (
    n1883,
    n1660
  );


  not
  g1873
  (
    n1797,
    n1574
  );


  buf
  g1874
  (
    n1999,
    n1518
  );


  not
  g1875
  (
    n2035,
    n1665
  );


  not
  g1876
  (
    n2030,
    n1613
  );


  not
  g1877
  (
    n1855,
    n1595
  );


  not
  g1878
  (
    n2176,
    n1655
  );


  not
  g1879
  (
    n2111,
    n1603
  );


  buf
  g1880
  (
    n1725,
    n1591
  );


  buf
  g1881
  (
    n1911,
    n1639
  );


  not
  g1882
  (
    n1955,
    n1579
  );


  not
  g1883
  (
    n2066,
    n1659
  );


  buf
  g1884
  (
    n1811,
    n1621
  );


  buf
  g1885
  (
    n2165,
    n1518
  );


  not
  g1886
  (
    n2151,
    n1568
  );


  not
  g1887
  (
    n2139,
    n1632
  );


  buf
  g1888
  (
    n2033,
    n1535
  );


  not
  g1889
  (
    n1774,
    n1569
  );


  not
  g1890
  (
    n2218,
    n1533
  );


  buf
  g1891
  (
    n1893,
    n1605
  );


  not
  g1892
  (
    n2183,
    n1657
  );


  not
  g1893
  (
    n1777,
    n1537
  );


  not
  g1894
  (
    n1736,
    n1615
  );


  buf
  g1895
  (
    n1737,
    n1617
  );


  not
  g1896
  (
    n1895,
    n1616
  );


  not
  g1897
  (
    n2008,
    n1594
  );


  buf
  g1898
  (
    n2123,
    n1659
  );


  buf
  g1899
  (
    n1731,
    n1585
  );


  buf
  g1900
  (
    n1919,
    n1570
  );


  not
  g1901
  (
    n1750,
    n1670
  );


  not
  g1902
  (
    n1746,
    n1566
  );


  buf
  g1903
  (
    n1961,
    n1581
  );


  buf
  g1904
  (
    n1748,
    n1514
  );


  not
  g1905
  (
    n2072,
    n1548
  );


  not
  g1906
  (
    n1724,
    n1586
  );


  not
  g1907
  (
    n1773,
    n1630
  );


  buf
  g1908
  (
    n2133,
    n1523
  );


  not
  g1909
  (
    n1933,
    n1623
  );


  buf
  g1910
  (
    n1788,
    n1614
  );


  not
  g1911
  (
    n2170,
    n1573
  );


  buf
  g1912
  (
    n1967,
    n1644
  );


  not
  g1913
  (
    n1820,
    n1651
  );


  buf
  g1914
  (
    n1941,
    n1668
  );


  buf
  g1915
  (
    n1836,
    n1618
  );


  buf
  g1916
  (
    n1881,
    n1519
  );


  buf
  g1917
  (
    n2012,
    n1628
  );


  buf
  g1918
  (
    n2093,
    n1658
  );


  buf
  g1919
  (
    n1816,
    n1520
  );


  not
  g1920
  (
    n2129,
    n1511
  );


  not
  g1921
  (
    n2173,
    n1574
  );


  buf
  g1922
  (
    n1969,
    n1671
  );


  not
  g1923
  (
    n2019,
    n1509
  );


  buf
  g1924
  (
    n2058,
    n1636
  );


  buf
  g1925
  (
    n2025,
    n1568
  );


  not
  g1926
  (
    n2065,
    n1526
  );


  not
  g1927
  (
    n2113,
    n1531
  );


  not
  g1928
  (
    n2202,
    n1531
  );


  buf
  g1929
  (
    n2121,
    n1665
  );


  buf
  g1930
  (
    n2160,
    n1557
  );


  not
  g1931
  (
    n2180,
    n1617
  );


  buf
  g1932
  (
    n1880,
    n1583
  );


  buf
  g1933
  (
    n1901,
    n1592
  );


  not
  g1934
  (
    n2037,
    n1549
  );


  buf
  g1935
  (
    n1868,
    n1543
  );


  not
  g1936
  (
    n2054,
    n1550
  );


  buf
  g1937
  (
    n1793,
    n1542
  );


  buf
  g1938
  (
    n1909,
    n1542
  );


  buf
  g1939
  (
    n2212,
    n1634
  );


  buf
  g1940
  (
    n2179,
    n1545
  );


  not
  g1941
  (
    n2014,
    n1621
  );


  buf
  g1942
  (
    n2089,
    n1534
  );


  buf
  g1943
  (
    n1982,
    n1577
  );


  buf
  g1944
  (
    n2087,
    n1550
  );


  buf
  g1945
  (
    n1887,
    n1574
  );


  not
  g1946
  (
    n2027,
    n1524
  );


  buf
  g1947
  (
    n1873,
    n1519
  );


  buf
  g1948
  (
    n1740,
    n1646
  );


  buf
  g1949
  (
    n1878,
    n1620
  );


  not
  g1950
  (
    n2040,
    n1668
  );


  buf
  g1951
  (
    n1781,
    n1643
  );


  not
  g1952
  (
    n2071,
    n1620
  );


  not
  g1953
  (
    n1767,
    n1630
  );


  buf
  g1954
  (
    n2205,
    n1576
  );


  not
  g1955
  (
    n1915,
    n1647
  );


  not
  g1956
  (
    n2039,
    n1616
  );


  buf
  g1957
  (
    n1757,
    n1620
  );


  not
  g1958
  (
    n2098,
    n1599
  );


  not
  g1959
  (
    n1939,
    n1594
  );


  buf
  g1960
  (
    n2204,
    n1590
  );


  not
  g1961
  (
    n2168,
    n1660
  );


  buf
  g1962
  (
    n2015,
    n1562
  );


  buf
  g1963
  (
    n1864,
    n1509
  );


  buf
  g1964
  (
    n2004,
    n1597
  );


  buf
  g1965
  (
    n2105,
    n1611
  );


  not
  g1966
  (
    n2009,
    n1601
  );


  buf
  g1967
  (
    n1800,
    n1649
  );


  not
  g1968
  (
    n1818,
    n1654
  );


  not
  g1969
  (
    n2182,
    n1581
  );


  not
  g1970
  (
    n1846,
    n1584
  );


  not
  g1971
  (
    n1817,
    n1564
  );


  buf
  g1972
  (
    n2213,
    n1534
  );


  not
  g1973
  (
    n2020,
    n1658
  );


  buf
  g1974
  (
    n1980,
    n1535
  );


  not
  g1975
  (
    n1728,
    n1541
  );


  buf
  g1976
  (
    n2167,
    n1610
  );


  buf
  g1977
  (
    n2107,
    n1514
  );


  buf
  g1978
  (
    n1845,
    n1652
  );


  not
  g1979
  (
    n2082,
    n1641
  );


  buf
  g1980
  (
    n2115,
    n1550
  );


  buf
  g1981
  (
    n1758,
    n1565
  );


  buf
  g1982
  (
    n1726,
    n1554
  );


  not
  g1983
  (
    n1910,
    n1594
  );


  buf
  g1984
  (
    n1739,
    n1663
  );


  buf
  g1985
  (
    n2104,
    n1561
  );


  not
  g1986
  (
    n1903,
    n1658
  );


  not
  g1987
  (
    n1975,
    n1536
  );


  not
  g1988
  (
    n1935,
    n1570
  );


  not
  g1989
  (
    n1853,
    n1523
  );


  buf
  g1990
  (
    n2011,
    n1544
  );


  buf
  g1991
  (
    n2047,
    n1587
  );


  buf
  g1992
  (
    n2050,
    n1556
  );


  buf
  g1993
  (
    n2067,
    n1577
  );


  not
  g1994
  (
    n1805,
    n1521
  );


  not
  g1995
  (
    n2049,
    n1593
  );


  buf
  g1996
  (
    n1744,
    n1652
  );


  not
  g1997
  (
    n2084,
    n1511
  );


  buf
  g1998
  (
    n1813,
    n1553
  );


  not
  g1999
  (
    n2002,
    n1600
  );


  not
  g2000
  (
    n1841,
    n1523
  );


  not
  g2001
  (
    n1993,
    n1575
  );


  buf
  g2002
  (
    n1722,
    n1536
  );


  not
  g2003
  (
    n2166,
    n1607
  );


  not
  g2004
  (
    n2148,
    n1558
  );


  buf
  g2005
  (
    n1940,
    n1640
  );


  not
  g2006
  (
    n2079,
    n1591
  );


  not
  g2007
  (
    n2078,
    n1606
  );


  not
  g2008
  (
    n2096,
    n1618
  );


  buf
  g2009
  (
    n1738,
    n1629
  );


  buf
  g2010
  (
    n1862,
    n1537
  );


  not
  g2011
  (
    n1796,
    n1669
  );


  not
  g2012
  (
    n1953,
    n1644
  );


  not
  g2013
  (
    n1819,
    n1552
  );


  not
  g2014
  (
    n1847,
    n1610
  );


  buf
  g2015
  (
    n1986,
    n1633
  );


  buf
  g2016
  (
    n1998,
    n1631
  );


  not
  g2017
  (
    n1827,
    n1614
  );


  buf
  g2018
  (
    n1832,
    n1580
  );


  not
  g2019
  (
    n1997,
    n1646
  );


  not
  g2020
  (
    n1934,
    n1651
  );


  not
  g2021
  (
    n1962,
    n1649
  );


  not
  g2022
  (
    n2156,
    n1626
  );


  buf
  g2023
  (
    n1897,
    n1623
  );


  buf
  g2024
  (
    n1718,
    n1622
  );


  buf
  g2025
  (
    n1946,
    n1539
  );


  buf
  g2026
  (
    n2134,
    n1592
  );


  not
  g2027
  (
    n1870,
    n1608
  );


  not
  g2028
  (
    n1942,
    n1533
  );


  buf
  g2029
  (
    n1859,
    n1619
  );


  not
  g2030
  (
    n1983,
    n1534
  );


  buf
  g2031
  (
    n2059,
    n1569
  );


  not
  g2032
  (
    n2120,
    n1609
  );


  buf
  g2033
  (
    n1996,
    n1615
  );


  not
  g2034
  (
    n2161,
    n1582
  );


  buf
  g2035
  (
    n1764,
    n1664
  );


  buf
  g2036
  (
    n2159,
    n1672
  );


  buf
  g2037
  (
    n1808,
    n1535
  );


  not
  g2038
  (
    n1829,
    n1549
  );


  not
  g2039
  (
    n1821,
    n1611
  );


  buf
  g2040
  (
    n2125,
    n1656
  );


  buf
  g2041
  (
    n1745,
    n1582
  );


  not
  g2042
  (
    n2088,
    n1533
  );


  buf
  g2043
  (
    n2191,
    n1596
  );


  buf
  g2044
  (
    n1923,
    n1560
  );


  buf
  g2045
  (
    n2041,
    n1612
  );


  buf
  g2046
  (
    n2198,
    n1635
  );


  not
  g2047
  (
    n2100,
    n1643
  );


  buf
  g2048
  (
    n2208,
    n1601
  );


  buf
  g2049
  (
    n2021,
    n1636
  );


  buf
  g2050
  (
    n1799,
    n1652
  );


  not
  g2051
  (
    n1976,
    n1529
  );


  not
  g2052
  (
    n1972,
    n1563
  );


  not
  g2053
  (
    n1838,
    n1528
  );


  buf
  g2054
  (
    n1790,
    n1571
  );


  not
  g2055
  (
    n1823,
    n1646
  );


  buf
  g2056
  (
    n2083,
    n1601
  );


  not
  g2057
  (
    n1992,
    n1542
  );


  not
  g2058
  (
    n2117,
    n1532
  );


  buf
  g2059
  (
    n1858,
    n1529
  );


  buf
  g2060
  (
    n1970,
    n1667
  );


  not
  g2061
  (
    n1727,
    n1584
  );


  buf
  g2062
  (
    n2174,
    n1512
  );


  buf
  g2063
  (
    n2024,
    n1669
  );


  not
  g2064
  (
    n1749,
    n1608
  );


  buf
  g2065
  (
    n1735,
    n1667
  );


  not
  g2066
  (
    n1768,
    n1571
  );


  buf
  g2067
  (
    n1723,
    n1514
  );


  not
  g2068
  (
    n2108,
    n1625
  );


  not
  g2069
  (
    n1772,
    n1648
  );


  buf
  g2070
  (
    n2080,
    n1564
  );


  buf
  g2071
  (
    n1787,
    n1612
  );


  buf
  g2072
  (
    n1849,
    n1526
  );


  not
  g2073
  (
    n1798,
    n1605
  );


  not
  g2074
  (
    n2181,
    n1647
  );


  buf
  g2075
  (
    n1835,
    n1639
  );


  buf
  g2076
  (
    n2091,
    n1585
  );


  not
  g2077
  (
    n2000,
    n1627
  );


  not
  g2078
  (
    n1759,
    n1621
  );


  not
  g2079
  (
    n1834,
    n1530
  );


  not
  g2080
  (
    n1833,
    n1644
  );


  buf
  g2081
  (
    n1812,
    n1560
  );


  buf
  g2082
  (
    n2034,
    n1524
  );


  buf
  g2083
  (
    n2016,
    n1536
  );


  not
  g2084
  (
    n1990,
    n1584
  );


  buf
  g2085
  (
    n2114,
    n1667
  );


  not
  g2086
  (
    n1760,
    n1510
  );


  not
  g2087
  (
    n1837,
    n1641
  );


  buf
  g2088
  (
    n1885,
    n1618
  );


  buf
  g2089
  (
    n1766,
    n1572
  );


  not
  g2090
  (
    n1932,
    n1616
  );


  not
  g2091
  (
    n1928,
    n1547
  );


  not
  g2092
  (
    n1851,
    n1554
  );


  not
  g2093
  (
    n1732,
    n1522
  );


  not
  g2094
  (
    n2163,
    n1545
  );


  buf
  g2095
  (
    n1922,
    n1561
  );


  buf
  g2096
  (
    n1756,
    n1566
  );


  not
  g2097
  (
    n1754,
    n1578
  );


  buf
  g2098
  (
    n1936,
    n1597
  );


  buf
  g2099
  (
    n1822,
    n1510
  );


  buf
  g2100
  (
    n1771,
    n1546
  );


  buf
  g2101
  (
    n1884,
    n1600
  );


  buf
  g2102
  (
    n1857,
    n1663
  );


  not
  g2103
  (
    n2061,
    n1602
  );


  buf
  g2104
  (
    n2103,
    n1563
  );


  not
  g2105
  (
    n2206,
    n1637
  );


  not
  g2106
  (
    n1720,
    n1638
  );


  not
  g2107
  (
    n2053,
    n1660
  );


  not
  g2108
  (
    n2197,
    n1634
  );


  buf
  g2109
  (
    n2018,
    n1562
  );


  buf
  g2110
  (
    n1803,
    n1546
  );


  not
  g2111
  (
    n1949,
    n1564
  );


  not
  g2112
  (
    n1743,
    n1635
  );


  buf
  g2113
  (
    n2221,
    n1530
  );


  buf
  g2114
  (
    n2184,
    n1647
  );


  buf
  g2115
  (
    n2200,
    n1547
  );


  buf
  g2116
  (
    n2219,
    n1605
  );


  not
  g2117
  (
    n2110,
    n1636
  );


  buf
  g2118
  (
    n2106,
    n1531
  );


  buf
  g2119
  (
    n2126,
    n1594
  );


  not
  g2120
  (
    n2077,
    n1655
  );


  not
  g2121
  (
    n2154,
    n1628
  );


  not
  g2122
  (
    n1963,
    n1598
  );


  not
  g2123
  (
    n1814,
    n1518
  );


  not
  g2124
  (
    n2171,
    n1619
  );


  buf
  g2125
  (
    n1988,
    n1623
  );


  buf
  g2126
  (
    n1951,
    n1527
  );


  not
  g2127
  (
    n1995,
    n1648
  );


  not
  g2128
  (
    n1751,
    n1588
  );


  buf
  g2129
  (
    n2056,
    n1604
  );


  not
  g2130
  (
    n2216,
    n1525
  );


  buf
  g2131
  (
    n2201,
    n1518
  );


  not
  g2132
  (
    n1927,
    n1516
  );


  not
  g2133
  (
    n1890,
    n1670
  );


  not
  g2134
  (
    n1905,
    n1566
  );


  buf
  g2135
  (
    n1984,
    n1593
  );


  not
  g2136
  (
    n1729,
    n1662
  );


  not
  g2137
  (
    n1741,
    n1578
  );


  buf
  g2138
  (
    n2032,
    n1589
  );


  xor
  g2139
  (
    n1938,
    n1554,
    n1598,
    n1573,
    n1542
  );


  xor
  g2140
  (
    n2209,
    n1629,
    n1653,
    n1657,
    n1584
  );


  xnor
  g2141
  (
    n1900,
    n1575,
    n1615,
    n1589,
    n1625
  );


  xnor
  g2142
  (
    n1860,
    n1650,
    n1525,
    n1640,
    n1648
  );


  nor
  g2143
  (
    n1871,
    n1617,
    n1519,
    n1512,
    n1576
  );


  xor
  g2144
  (
    n2172,
    n1515,
    n1597,
    n1604,
    n1632
  );


  nor
  g2145
  (
    n1974,
    n1513,
    n1664,
    n1560,
    n1619
  );


  xnor
  g2146
  (
    n2195,
    n1606,
    n1656,
    n1538,
    n1553
  );


  nor
  g2147
  (
    n2060,
    n1563,
    n1561,
    n1574,
    n1666
  );


  nand
  g2148
  (
    n2199,
    n1624,
    n1532,
    n1592,
    n1512
  );


  nand
  g2149
  (
    n1830,
    n1572,
    n1513,
    n1659,
    n1571
  );


  nand
  g2150
  (
    n1785,
    n1608,
    n1643,
    n1599,
    n1543
  );


  nor
  g2151
  (
    n1888,
    n1630,
    n1552,
    n1587,
    n1629
  );


  xor
  g2152
  (
    n2187,
    n1583,
    n1537,
    n1511,
    n1622
  );


  nand
  g2153
  (
    n1979,
    n1562,
    n1627,
    n1522,
    n1599
  );


  nor
  g2154
  (
    n2214,
    n1567,
    n1545,
    n1516,
    n1529
  );


  or
  g2155
  (
    n2073,
    n1577,
    n1590,
    n1626,
    n1566
  );


  or
  g2156
  (
    n1826,
    n1573,
    n1631,
    n1672,
    n1637
  );


  nor
  g2157
  (
    n2036,
    n1661,
    n1591,
    n1638,
    n1593
  );


  xor
  g2158
  (
    n1930,
    n1652,
    n1523,
    n1602,
    n1585
  );


  xnor
  g2159
  (
    n1842,
    n1613,
    n1559,
    n1546,
    n1580
  );


  xnor
  g2160
  (
    n1879,
    n1511,
    n1612,
    n1521,
    n1634
  );


  nor
  g2161
  (
    n1978,
    n1547,
    n1609,
    n1604,
    n1521
  );


  xor
  g2162
  (
    n1947,
    n1657,
    n1655,
    n1555,
    n1628
  );


  and
  g2163
  (
    n1906,
    n1637,
    n1642,
    n1575,
    n1581
  );


  xor
  g2164
  (
    n2140,
    n1605,
    n1551,
    n1532,
    n1598
  );


  and
  g2165
  (
    n1752,
    n1512,
    n1603,
    n1602,
    n1653
  );


  nor
  g2166
  (
    n2007,
    n1585,
    n1640,
    n1654,
    n1612
  );


  nor
  g2167
  (
    n1863,
    n1549,
    n1603,
    n1607,
    n1519
  );


  nand
  g2168
  (
    n2116,
    n1567,
    n1602,
    n1671,
    n1517
  );


  and
  g2169
  (
    n2193,
    n1561,
    n1578,
    n1666,
    n1540
  );


  xnor
  g2170
  (
    n1831,
    n1544,
    n1622,
    n1539,
    n1570
  );


  xor
  g2171
  (
    n1958,
    n1588,
    n1635,
    n1520,
    n1555
  );


  and
  g2172
  (
    n1856,
    n1631,
    n1579,
    n1666,
    n1555
  );


  nor
  g2173
  (
    n1965,
    n1552,
    n1540,
    n1539,
    n1586
  );


  or
  g2174
  (
    n2031,
    n1517,
    n1633,
    n1513,
    n1569
  );


  nor
  g2175
  (
    n2090,
    n1668,
    n1529,
    n1609
  );


  xnor
  g2176
  (
    n2094,
    n1666,
    n1645,
    n1632,
    n1633
  );


  nand
  g2177
  (
    n2141,
    n1559,
    n1568,
    n1655,
    n1527
  );


  or
  g2178
  (
    n1959,
    n1638,
    n1576,
    n1538,
    n1527
  );


  xnor
  g2179
  (
    n2003,
    n1551,
    n1656,
    n1662,
    n1560
  );


  or
  g2180
  (
    n2127,
    n1669,
    n1640,
    n1582,
    n1631
  );


  nand
  g2181
  (
    n2136,
    n1556,
    n1668,
    n1651,
    n1626
  );


  nand
  g2182
  (
    n2076,
    n1664,
    n1567,
    n1555,
    n1588
  );


  and
  g2183
  (
    n1824,
    n1618,
    n1643,
    n1625,
    n1547
  );


  nand
  g2184
  (
    n1840,
    n1514,
    n1635,
    n1581,
    n1526
  );


  nand
  g2185
  (
    n2112,
    n1599,
    n1653,
    n1563,
    n1639
  );


  nand
  g2186
  (
    n1926,
    n1658,
    n1662,
    n1606,
    n1525
  );


  and
  g2187
  (
    n2001,
    n1648,
    n1573,
    n1634,
    n1625
  );


  nand
  g2188
  (
    n2185,
    n1591,
    n1553,
    n1641,
    n1516
  );


  nor
  g2189
  (
    n2228,
    n1717,
    n1718,
    n1724,
    n1755
  );


  and
  g2190
  (
    n2226,
    n1756,
    n1738,
    n1735,
    n1732
  );


  nand
  g2191
  (
    n2225,
    n1721,
    n1736,
    n1749,
    n1725
  );


  nand
  g2192
  (
    n2224,
    n1727,
    n1731,
    n1743,
    n1747
  );


  and
  g2193
  (
    n2222,
    n1754,
    n1753,
    n1722,
    n1740
  );


  or
  g2194
  (
    n2227,
    n1723,
    n1739,
    n1730,
    n1737
  );


  or
  g2195
  (
    n2223,
    n1741,
    n1750,
    n1734,
    n1742
  );


  nor
  g2196
  (
    n2230,
    n1726,
    n1752,
    n1748,
    n1720
  );


  or
  g2197
  (
    n2229,
    n1733,
    n1751,
    n1746,
    n1729
  );


  nor
  g2198
  (
    n2231,
    n1728,
    n1719,
    n1745,
    n1744
  );


  buf
  g2199
  (
    n2240,
    n1674
  );


  buf
  g2200
  (
    n2236,
    n2224
  );


  not
  g2201
  (
    n2233,
    n1673
  );


  not
  g2202
  (
    n2232,
    n2222
  );


  not
  g2203
  (
    n2235,
    n1674
  );


  not
  g2204
  (
    n2241,
    n1673
  );


  xor
  g2205
  (
    n2239,
    n2229,
    n1672
  );


  xnor
  g2206
  (
    n2237,
    n2228,
    n1674,
    n1675,
    n2223
  );


  nor
  g2207
  (
    n2238,
    n2231,
    n1673,
    n2230,
    n2225
  );


  or
  g2208
  (
    n2234,
    n2226,
    n1673,
    n1674,
    n2227
  );


  not
  g2209
  (
    n2242,
    n2232
  );


  buf
  g2210
  (
    n2243,
    n2242
  );


  buf
  g2211
  (
    n2245,
    n2242
  );


  not
  g2212
  (
    n2244,
    n2242
  );


  not
  g2213
  (
    n2246,
    n2243
  );


  buf
  g2214
  (
    n2247,
    n2243
  );


  xnor
  g2215
  (
    n2248,
    n2246,
    n1675,
    n2247,
    n1757
  );


  buf
  g2216
  (
    n2250,
    n2248
  );


  buf
  g2217
  (
    n2249,
    n2248
  );


  not
  g2218
  (
    n2252,
    n672
  );


  buf
  g2219
  (
    n2254,
    n2249
  );


  buf
  g2220
  (
    n2251,
    n2250
  );


  not
  g2221
  (
    n2256,
    n2249
  );


  nand
  g2222
  (
    n2253,
    n672,
    n2250
  );


  xnor
  g2223
  (
    n2255,
    n2249,
    n672
  );


  buf
  g2224
  (
    n2261,
    n2252
  );


  buf
  g2225
  (
    n2264,
    n2252
  );


  buf
  g2226
  (
    n2262,
    n2253
  );


  buf
  g2227
  (
    n2263,
    n2252
  );


  buf
  g2228
  (
    n2257,
    n2252
  );


  not
  g2229
  (
    n2258,
    n2253
  );


  buf
  g2230
  (
    n2259,
    n2253
  );


  buf
  g2231
  (
    n2260,
    n2251
  );


  or
  g2232
  (
    n2282,
    n1694,
    n1692,
    n1698
  );


  xor
  g2233
  (
    n2291,
    n2261,
    n2257,
    n1691,
    n1689
  );


  or
  g2234
  (
    n2286,
    n1689,
    n1690,
    n2264,
    n1688
  );


  and
  g2235
  (
    n2288,
    n1688,
    n1684,
    n1699,
    n1681
  );


  nand
  g2236
  (
    n2267,
    n1698,
    n1681,
    n1686,
    n1685
  );


  nor
  g2237
  (
    n2275,
    n1683,
    n2258,
    n1677,
    n2264
  );


  nand
  g2238
  (
    n2273,
    n2257,
    n1697,
    n1693
  );


  nand
  g2239
  (
    n2284,
    n2264,
    n2261,
    n1675,
    n1684
  );


  nand
  g2240
  (
    n2290,
    n2264,
    n1683,
    n1678,
    n2259
  );


  or
  g2241
  (
    KeyWire_0_14,
    n1680,
    n1676,
    n1690,
    n1689
  );


  and
  g2242
  (
    n2269,
    n1684,
    n1687,
    n1696,
    n1686
  );


  and
  g2243
  (
    n2268,
    n1677,
    n1677,
    n1683,
    n1692
  );


  or
  g2244
  (
    n2271,
    n1696,
    n1694,
    n1680
  );


  or
  g2245
  (
    n2279,
    n1690,
    n1682,
    n1681
  );


  and
  g2246
  (
    n2266,
    n1685,
    n1691,
    n2259,
    n2261
  );


  nor
  g2247
  (
    n2285,
    n2261,
    n1677,
    n1693,
    n2263
  );


  and
  g2248
  (
    n2270,
    n1694,
    n1699,
    n1678,
    n2260
  );


  and
  g2249
  (
    n2289,
    n2258,
    n2262,
    n1678,
    n1682
  );


  nand
  g2250
  (
    n2277,
    n1698,
    n1675,
    n2260,
    n2262
  );


  or
  g2251
  (
    n2281,
    n1686,
    n1691,
    n1680,
    n1688
  );


  nor
  g2252
  (
    n2292,
    n2262,
    n2257,
    n2259,
    n1685
  );


  xnor
  g2253
  (
    n2272,
    n2263,
    n1696,
    n1682
  );


  nand
  g2254
  (
    n2287,
    n2258,
    n1695,
    n1698,
    n2260
  );


  nor
  g2255
  (
    n2276,
    n1679,
    n1697,
    n1678,
    n1688
  );


  or
  g2256
  (
    n2294,
    n1681,
    n2258,
    n1695,
    n1676
  );


  or
  g2257
  (
    n2265,
    n1697,
    n1676,
    n2260,
    n1679
  );


  xor
  g2258
  (
    n2283,
    n1690,
    n2259,
    n1692,
    n1687
  );


  xor
  g2259
  (
    n2296,
    n1676,
    n1695,
    n1689,
    n1683
  );


  xor
  g2260
  (
    n2280,
    n1686,
    n1695,
    n2257,
    n1679
  );


  xor
  g2261
  (
    n2295,
    n1687,
    n1697,
    n2263,
    n1685
  );


  xor
  g2262
  (
    n2293,
    n2263,
    n1679,
    n1684,
    n1687
  );


  xnor
  g2263
  (
    n2274,
    n1680,
    n1691,
    n1693,
    n2262
  );


  xor
  g2264
  (
    n2339,
    n2039,
    n1983,
    n2052,
    n1788
  );


  nand
  g2265
  (
    n2377,
    n1966,
    n1926,
    n2292,
    n1855
  );


  or
  g2266
  (
    n2405,
    n1815,
    n1795,
    n2296,
    n1980
  );


  nor
  g2267
  (
    n2365,
    n2122,
    n2043,
    n1827,
    n2269
  );


  or
  g2268
  (
    n2375,
    n1823,
    n2295,
    n1916,
    n1816
  );


  xor
  g2269
  (
    n2319,
    n2295,
    n1776,
    n1762,
    n1871
  );


  nor
  g2270
  (
    n2304,
    n2099,
    n2291,
    n2268,
    n1800
  );


  xnor
  g2271
  (
    n2348,
    n1818,
    n1947,
    n2028,
    n2271
  );


  xnor
  g2272
  (
    n2388,
    n2278,
    n1984,
    n2119,
    n2286
  );


  xor
  g2273
  (
    n2333,
    n2116,
    n1918,
    n1797,
    n1920
  );


  xnor
  g2274
  (
    n2310,
    n2287,
    n2097,
    n2295,
    n1985
  );


  xor
  g2275
  (
    n2312,
    n1865,
    n1950,
    n2030,
    n1952
  );


  xnor
  g2276
  (
    n2316,
    n2274,
    n1896,
    n1942,
    n1775
  );


  xnor
  g2277
  (
    n2361,
    n1851,
    n1939,
    n1921,
    n2283
  );


  or
  g2278
  (
    n2307,
    n1771,
    n1845,
    n1919,
    n1883
  );


  or
  g2279
  (
    n2373,
    n2274,
    n2063,
    n1856,
    n1842
  );


  xor
  g2280
  (
    n2351,
    n2291,
    n2280,
    n2272,
    n1994
  );


  or
  g2281
  (
    n2416,
    n1977,
    n2023,
    n1847,
    n2033
  );


  and
  g2282
  (
    n2363,
    n2289,
    n2106,
    n1938,
    n2286
  );


  or
  g2283
  (
    n2409,
    n2029,
    n2268,
    n2289,
    n1969
  );


  xnor
  g2284
  (
    n2354,
    n1773,
    n2056,
    n1999,
    n2267
  );


  nor
  g2285
  (
    n2299,
    n2283,
    n2038,
    n1790,
    n1804
  );


  xor
  g2286
  (
    n2379,
    n2279,
    n1852,
    n1915,
    n1792
  );


  or
  g2287
  (
    n2328,
    n2288,
    n1914,
    n1840,
    n2037
  );


  or
  g2288
  (
    n2367,
    n2083,
    n2089,
    n1898,
    n1875
  );


  or
  g2289
  (
    n2350,
    n1978,
    n2009,
    n2276,
    n2282
  );


  nand
  g2290
  (
    n2343,
    n1854,
    n1911,
    n1820,
    n2064
  );


  nor
  g2291
  (
    n2318,
    n2294,
    n2133,
    n1990,
    n1974
  );


  nand
  g2292
  (
    n2324,
    n2292,
    n2271,
    n1937,
    n1759
  );


  nor
  g2293
  (
    n2335,
    n2005,
    n2281,
    n1981,
    n1798
  );


  and
  g2294
  (
    n2322,
    n2072,
    n1779,
    n1893,
    n1913
  );


  xor
  g2295
  (
    n2399,
    n2098,
    n2012,
    n2110,
    n2032
  );


  xnor
  g2296
  (
    n2353,
    n2013,
    n1940,
    n2277,
    n2014
  );


  or
  g2297
  (
    n2362,
    n1824,
    n2109,
    n2266,
    n2001
  );


  xor
  g2298
  (
    n2391,
    n2287,
    n2290,
    n1806,
    n2024
  );


  nor
  g2299
  (
    n2407,
    n2291,
    n2291,
    n1897,
    n1763
  );


  xor
  g2300
  (
    n2414,
    n2088,
    n2113,
    n2002,
    n2272
  );


  and
  g2301
  (
    n2386,
    n1768,
    n1760,
    n2293,
    n2008
  );


  xnor
  g2302
  (
    n2410,
    n2101,
    n1941,
    n1967,
    n2280
  );


  and
  g2303
  (
    n2344,
    n1876,
    n1794,
    n2267,
    n1995
  );


  nor
  g2304
  (
    n2355,
    n2130,
    n2059,
    n2265,
    n1767
  );


  xor
  g2305
  (
    n2300,
    n2081,
    n2050,
    n1808,
    n1928
  );


  xnor
  g2306
  (
    n2376,
    n2270,
    n1764,
    n1758,
    n1953
  );


  nand
  g2307
  (
    n2389,
    n2288,
    n2276,
    n1902,
    n2015
  );


  nand
  g2308
  (
    n2338,
    n2281,
    n2279,
    n2117,
    n2266
  );


  xor
  g2309
  (
    n2347,
    n1890,
    n1802,
    n2287,
    n2280
  );


  nor
  g2310
  (
    n2323,
    n2271,
    n1943,
    n1819,
    n2069
  );


  and
  g2311
  (
    n2346,
    n2041,
    n2019,
    n1923,
    n2082
  );


  xor
  g2312
  (
    n2420,
    n2276,
    n1812,
    n2270,
    n1961
  );


  and
  g2313
  (
    n2321,
    n2084,
    n2265,
    n2066,
    n1787
  );


  xnor
  g2314
  (
    n2331,
    n2006,
    n2007,
    n1954,
    n2275
  );


  and
  g2315
  (
    n2345,
    n1860,
    n2294,
    n2138,
    n1844
  );


  xor
  g2316
  (
    n2371,
    n2095,
    n2137,
    n1904,
    n1846
  );


  nand
  g2317
  (
    n2359,
    n2049,
    n1833,
    n2270,
    n1796
  );


  nand
  g2318
  (
    n2400,
    n2285,
    n2091,
    n2273,
    n1781
  );


  or
  g2319
  (
    n2390,
    n2070,
    n1877,
    n2057,
    n1936
  );


  nor
  g2320
  (
    n2412,
    n2278,
    n1888,
    n1793,
    n1836
  );


  or
  g2321
  (
    n2413,
    n1987,
    n2136,
    n2078,
    n1958
  );


  xor
  g2322
  (
    n2384,
    n2284,
    n1934,
    n1979,
    n1887
  );


  nand
  g2323
  (
    n2330,
    n1894,
    n2121,
    n1927,
    n2134
  );


  nor
  g2324
  (
    n2422,
    n2293,
    n2273,
    n1814,
    n2286
  );


  xnor
  g2325
  (
    n2325,
    n1777,
    n2280,
    n1869,
    n2103
  );


  nand
  g2326
  (
    n2370,
    n2283,
    n1799,
    n1935,
    n2061
  );


  nand
  g2327
  (
    n2387,
    n2275,
    n2107,
    n2265,
    n2079
  );


  or
  g2328
  (
    n2401,
    n1971,
    n2139,
    n2086,
    n2020
  );


  nand
  g2329
  (
    n2302,
    n2292,
    n2010,
    n1930,
    n2271
  );


  or
  g2330
  (
    n2334,
    n2274,
    n2292,
    n2269,
    n2293
  );


  nand
  g2331
  (
    n2356,
    n1899,
    n2284,
    n1988,
    n1826
  );


  xnor
  g2332
  (
    n2424,
    n1843,
    n2283,
    n1992,
    n2128
  );


  xor
  g2333
  (
    n2349,
    n1908,
    n2075,
    n1925,
    n1948
  );


  and
  g2334
  (
    n2326,
    n2282,
    n1955,
    n2118,
    n1772
  );


  xnor
  g2335
  (
    n2341,
    n2077,
    n1872,
    n1813,
    n1791
  );


  and
  g2336
  (
    n2374,
    n2285,
    n1830,
    n2042,
    n1803
  );


  nand
  g2337
  (
    n2383,
    n2126,
    n1909,
    n1900,
    n2000
  );


  nand
  g2338
  (
    n2411,
    n1864,
    n1874,
    n1986,
    n1828
  );


  xor
  g2339
  (
    n2305,
    n2273,
    n1862,
    n1809,
    n1963
  );


  xor
  g2340
  (
    n2393,
    n2284,
    n2027,
    n2031,
    n1801
  );


  nand
  g2341
  (
    n2368,
    n2140,
    n2093,
    n1848,
    n2273
  );


  nand
  g2342
  (
    n2403,
    n1905,
    n1837,
    n2114,
    n1962
  );


  xor
  g2343
  (
    n2419,
    n2289,
    n1841,
    n2279,
    n2060
  );


  and
  g2344
  (
    n2364,
    n2108,
    n1817,
    n1972,
    n2054
  );


  nor
  g2345
  (
    n2372,
    n2047,
    n1998,
    n2127,
    n2016
  );


  nor
  g2346
  (
    n2317,
    n2018,
    n1959,
    n2275,
    n2293
  );


  nand
  g2347
  (
    n2336,
    n1835,
    n2267,
    n1821,
    n1857
  );


  xor
  g2348
  (
    n2301,
    n1831,
    n2035,
    n1859,
    n1780
  );


  xor
  g2349
  (
    n2415,
    n2034,
    n2294,
    n1880,
    n1861
  );


  nor
  g2350
  (
    n2421,
    n1910,
    n2295,
    n1901,
    n1964
  );


  xnor
  g2351
  (
    n2395,
    n2120,
    n2132,
    n2296,
    n2269
  );


  xnor
  g2352
  (
    n2313,
    n2294,
    n1783,
    n2266,
    n2080
  );


  or
  g2353
  (
    n2298,
    n1957,
    n1944,
    n1976,
    n1770
  );


  or
  g2354
  (
    n2369,
    n2277,
    n1889,
    n2048,
    n2026
  );


  or
  g2355
  (
    n2418,
    n1968,
    n1895,
    n1785,
    n1769
  );


  xor
  g2356
  (
    n2402,
    n2045,
    n2021,
    n1863,
    n1945
  );


  nor
  g2357
  (
    n2337,
    n2051,
    n2011,
    n2281,
    n1886
  );


  nand
  g2358
  (
    n2320,
    n1993,
    n2266,
    n1965,
    n1807
  );


  nor
  g2359
  (
    n2332,
    n2267,
    n2286,
    n2123,
    n1870
  );


  or
  g2360
  (
    n2360,
    n1881,
    n1832,
    n1811,
    n1879
  );


  or
  g2361
  (
    n2417,
    n1932,
    n2272,
    n2289,
    n2071
  );


  nand
  g2362
  (
    n2315,
    n2285,
    n1853,
    n1867,
    n2277
  );


  nand
  g2363
  (
    n2311,
    n1970,
    n2288,
    n1924,
    n2290
  );


  nand
  g2364
  (
    n2342,
    n2102,
    n2268,
    n2124,
    n2277
  );


  xnor
  g2365
  (
    n2394,
    n2025,
    n1849,
    n1933,
    n1761
  );


  and
  g2366
  (
    n2308,
    n2281,
    n2062,
    n1982,
    n2272
  );


  xor
  g2367
  (
    n2340,
    n2265,
    n1912,
    n1786,
    n1951
  );


  nand
  g2368
  (
    n2329,
    n2036,
    n2085,
    n2296,
    n1891
  );


  nand
  g2369
  (
    n2297,
    n1975,
    n1829,
    n2092,
    n2058
  );


  xnor
  g2370
  (
    n2385,
    n1789,
    n1850,
    n1838,
    n1784
  );


  xor
  g2371
  (
    n2352,
    n2090,
    n2296,
    n2003,
    n1929
  );


  xnor
  g2372
  (
    n2381,
    n1782,
    n1878,
    n2278,
    n2104
  );


  nand
  g2373
  (
    n2396,
    n1931,
    n2282,
    n2094,
    n2111
  );


  nand
  g2374
  (
    n2358,
    n2096,
    n2065,
    n2004,
    n1766
  );


  or
  g2375
  (
    n2314,
    n2053,
    n1946,
    n2055,
    n2046
  );


  xnor
  g2376
  (
    n2309,
    n2279,
    n1991,
    n2044,
    n2135
  );


  xor
  g2377
  (
    n2408,
    n2282,
    n2073,
    n2125,
    n2290
  );


  and
  g2378
  (
    n2404,
    n2067,
    n2288,
    n1903,
    n2284
  );


  or
  g2379
  (
    n2380,
    n2076,
    n1774,
    n1825,
    n2040
  );


  xnor
  g2380
  (
    n2306,
    n1892,
    n1810,
    n1997,
    n1765
  );


  nand
  g2381
  (
    n2423,
    n2074,
    n1949,
    n1884,
    n1866
  );


  nand
  g2382
  (
    n2392,
    n2068,
    n1834,
    n1922,
    n1917
  );


  and
  g2383
  (
    n2327,
    n1873,
    n1885,
    n1907,
    n2100
  );


  or
  g2384
  (
    n2357,
    n2131,
    n2105,
    n1805,
    n2290
  );


  xnor
  g2385
  (
    n2398,
    n2270,
    n2275,
    n1858,
    n2017
  );


  nor
  g2386
  (
    n2382,
    n1989,
    n2274,
    n1868,
    n1822
  );


  and
  g2387
  (
    n2397,
    n2287,
    n2087,
    n2276,
    n1882
  );


  xnor
  g2388
  (
    n2303,
    n2129,
    n1906,
    n2115,
    n2268
  );


  nand
  g2389
  (
    n2406,
    n1996,
    n2278,
    n1956,
    n2112
  );


  and
  g2390
  (
    n2366,
    n1778,
    n1973,
    n2141,
    n2285
  );


  nor
  g2391
  (
    n2378,
    n1960,
    n2022,
    n1839,
    n2269
  );


  not
  g2392
  (
    n2527,
    n2345
  );


  buf
  g2393
  (
    n2508,
    n2339
  );


  buf
  g2394
  (
    n2494,
    n2383
  );


  not
  g2395
  (
    n2498,
    n2328
  );


  buf
  g2396
  (
    n2665,
    n2412
  );


  not
  g2397
  (
    n2530,
    n2339
  );


  not
  g2398
  (
    n2426,
    n2323
  );


  buf
  g2399
  (
    n2500,
    n2310
  );


  buf
  g2400
  (
    n2493,
    n2408
  );


  buf
  g2401
  (
    n2455,
    n2387
  );


  not
  g2402
  (
    n2445,
    n2326
  );


  buf
  g2403
  (
    n2489,
    n2381
  );


  buf
  g2404
  (
    n2459,
    n2321
  );


  not
  g2405
  (
    n2521,
    n2348
  );


  buf
  g2406
  (
    n2545,
    n2382
  );


  not
  g2407
  (
    n2594,
    n2344
  );


  not
  g2408
  (
    n2449,
    n2412
  );


  not
  g2409
  (
    n2541,
    n2415
  );


  not
  g2410
  (
    n2681,
    n2320
  );


  buf
  g2411
  (
    n2713,
    n2360
  );


  not
  g2412
  (
    n2518,
    n2394
  );


  buf
  g2413
  (
    n2559,
    n2378
  );


  not
  g2414
  (
    n2507,
    n2333
  );


  buf
  g2415
  (
    n2663,
    n2418
  );


  buf
  g2416
  (
    n2624,
    n2393
  );


  buf
  g2417
  (
    n2714,
    n2352
  );


  buf
  g2418
  (
    n2573,
    n2349
  );


  not
  g2419
  (
    n2536,
    n2332
  );


  not
  g2420
  (
    n2505,
    n2297
  );


  not
  g2421
  (
    n2655,
    n2302
  );


  not
  g2422
  (
    n2506,
    n2335
  );


  not
  g2423
  (
    n2712,
    n2384
  );


  not
  g2424
  (
    n2437,
    n2392
  );


  not
  g2425
  (
    n2672,
    n2367
  );


  buf
  g2426
  (
    n2605,
    n2397
  );


  not
  g2427
  (
    n2699,
    n2349
  );


  not
  g2428
  (
    n2554,
    n2310
  );


  buf
  g2429
  (
    n2474,
    n2317
  );


  not
  g2430
  (
    n2604,
    n2408
  );


  not
  g2431
  (
    n2718,
    n2397
  );


  not
  g2432
  (
    n2581,
    n2314
  );


  not
  g2433
  (
    n2673,
    n1503
  );


  buf
  g2434
  (
    n2570,
    n2323
  );


  buf
  g2435
  (
    n2482,
    n2375
  );


  buf
  g2436
  (
    n2574,
    n2359
  );


  not
  g2437
  (
    n2577,
    n2376
  );


  buf
  g2438
  (
    n2485,
    n2343
  );


  not
  g2439
  (
    n2662,
    n2254
  );


  not
  g2440
  (
    n2674,
    n2302
  );


  buf
  g2441
  (
    n2644,
    n2328
  );


  not
  g2442
  (
    n2647,
    n2417
  );


  buf
  g2443
  (
    n2586,
    n2338
  );


  buf
  g2444
  (
    KeyWire_0_5,
    n2341
  );


  buf
  g2445
  (
    n2684,
    n2346
  );


  buf
  g2446
  (
    n2467,
    n1508
  );


  not
  g2447
  (
    n2560,
    n2412
  );


  buf
  g2448
  (
    n2457,
    n2312
  );


  buf
  g2449
  (
    n2621,
    n2378
  );


  not
  g2450
  (
    n2638,
    n2394
  );


  not
  g2451
  (
    n2522,
    n2255
  );


  not
  g2452
  (
    n2611,
    n2396
  );


  not
  g2453
  (
    n2593,
    n2314
  );


  not
  g2454
  (
    n2595,
    n2351
  );


  buf
  g2455
  (
    n2450,
    n1508
  );


  buf
  g2456
  (
    n2488,
    n2388
  );


  not
  g2457
  (
    n2452,
    n2376
  );


  buf
  g2458
  (
    n2636,
    n2422
  );


  not
  g2459
  (
    n2525,
    n2352
  );


  buf
  g2460
  (
    n2563,
    n2391
  );


  buf
  g2461
  (
    n2720,
    n2256
  );


  not
  g2462
  (
    n2613,
    n2389
  );


  not
  g2463
  (
    n2568,
    n2311
  );


  buf
  g2464
  (
    n2502,
    n2347
  );


  not
  g2465
  (
    n2519,
    n2299
  );


  buf
  g2466
  (
    n2512,
    n2347
  );


  buf
  g2467
  (
    n2590,
    n2316
  );


  buf
  g2468
  (
    n2626,
    n2388
  );


  not
  g2469
  (
    n2645,
    n2404
  );


  not
  g2470
  (
    n2692,
    n2365
  );


  buf
  g2471
  (
    n2615,
    n2355
  );


  not
  g2472
  (
    n2704,
    n2401
  );


  buf
  g2473
  (
    n2616,
    n2376
  );


  not
  g2474
  (
    n2585,
    n1505
  );


  buf
  g2475
  (
    n2583,
    n2300
  );


  buf
  g2476
  (
    n2435,
    n2256
  );


  not
  g2477
  (
    n2669,
    n2301
  );


  not
  g2478
  (
    n2675,
    n2418
  );


  buf
  g2479
  (
    n2619,
    n2335
  );


  buf
  g2480
  (
    n2690,
    n2321
  );


  not
  g2481
  (
    n2433,
    n2388
  );


  not
  g2482
  (
    n2579,
    n1504
  );


  not
  g2483
  (
    n2628,
    n2362
  );


  not
  g2484
  (
    n2698,
    n1504
  );


  buf
  g2485
  (
    n2706,
    n2400
  );


  buf
  g2486
  (
    n2582,
    n2326
  );


  buf
  g2487
  (
    n2456,
    n2402
  );


  not
  g2488
  (
    n2687,
    n2350
  );


  buf
  g2489
  (
    n2442,
    n2337
  );


  buf
  g2490
  (
    n2461,
    n2329
  );


  buf
  g2491
  (
    n2468,
    n2306
  );


  not
  g2492
  (
    n2623,
    n2393
  );


  not
  g2493
  (
    n2553,
    n2298
  );


  buf
  g2494
  (
    n2620,
    n2298
  );


  not
  g2495
  (
    n2438,
    n2326
  );


  not
  g2496
  (
    n2481,
    n2315
  );


  buf
  g2497
  (
    n2492,
    n2420
  );


  buf
  g2498
  (
    n2668,
    n2324
  );


  not
  g2499
  (
    n2632,
    n2380
  );


  buf
  g2500
  (
    n2483,
    n2346
  );


  not
  g2501
  (
    n2682,
    n2341
  );


  not
  g2502
  (
    n2618,
    n2343
  );


  not
  g2503
  (
    n2496,
    n2340
  );


  buf
  g2504
  (
    n2477,
    n2327
  );


  buf
  g2505
  (
    n2576,
    n2358
  );


  buf
  g2506
  (
    n2533,
    n2412
  );


  buf
  g2507
  (
    n2625,
    n2333
  );


  buf
  g2508
  (
    n2454,
    n1506
  );


  not
  g2509
  (
    n2664,
    n2361
  );


  not
  g2510
  (
    n2513,
    n2382
  );


  not
  g2511
  (
    n2501,
    n2411
  );


  buf
  g2512
  (
    n2598,
    n2411
  );


  not
  g2513
  (
    n2658,
    n2372
  );


  not
  g2514
  (
    n2509,
    n2419
  );


  buf
  g2515
  (
    n2650,
    n2390
  );


  buf
  g2516
  (
    n2648,
    n2394
  );


  not
  g2517
  (
    n2564,
    n2384
  );


  buf
  g2518
  (
    n2520,
    n2305
  );


  not
  g2519
  (
    n2640,
    n2302
  );


  not
  g2520
  (
    n2575,
    n2312
  );


  not
  g2521
  (
    n2444,
    n2423
  );


  buf
  g2522
  (
    n2484,
    n2336
  );


  not
  g2523
  (
    n2617,
    n2393
  );


  not
  g2524
  (
    n2490,
    n2300
  );


  buf
  g2525
  (
    n2466,
    n2363
  );


  not
  g2526
  (
    n2567,
    n2314
  );


  not
  g2527
  (
    n2537,
    n2385
  );


  not
  g2528
  (
    n2486,
    n2305
  );


  buf
  g2529
  (
    n2705,
    n2416
  );


  not
  g2530
  (
    n2471,
    n2403
  );


  not
  g2531
  (
    n2546,
    n2421
  );


  buf
  g2532
  (
    n2446,
    n2403
  );


  not
  g2533
  (
    n2523,
    n2322
  );


  buf
  g2534
  (
    n2580,
    n2350
  );


  buf
  g2535
  (
    n2578,
    n2390
  );


  not
  g2536
  (
    n2549,
    n2405
  );


  buf
  g2537
  (
    n2538,
    n2414
  );


  not
  g2538
  (
    n2517,
    n2411
  );


  buf
  g2539
  (
    n2562,
    n2329
  );


  not
  g2540
  (
    n2453,
    n2303
  );


  buf
  g2541
  (
    n2695,
    n2363
  );


  buf
  g2542
  (
    n2431,
    n2336
  );


  not
  g2543
  (
    n2661,
    n2382
  );


  not
  g2544
  (
    n2646,
    n2418
  );


  buf
  g2545
  (
    n2532,
    n2398
  );


  buf
  g2546
  (
    n2693,
    n2395
  );


  not
  g2547
  (
    n2607,
    n2366
  );


  buf
  g2548
  (
    n2529,
    n1502
  );


  buf
  g2549
  (
    n2463,
    n2323
  );


  buf
  g2550
  (
    n2552,
    n2420
  );


  not
  g2551
  (
    n2473,
    n2356
  );


  buf
  g2552
  (
    n2470,
    n1502
  );


  not
  g2553
  (
    n2680,
    n2317
  );


  buf
  g2554
  (
    n2707,
    n2404
  );


  not
  g2555
  (
    n2475,
    n2330
  );


  not
  g2556
  (
    n2547,
    n2364
  );


  buf
  g2557
  (
    n2641,
    n2416
  );


  not
  g2558
  (
    n2543,
    n2362
  );


  not
  g2559
  (
    n2558,
    n2320
  );


  not
  g2560
  (
    n2643,
    n2314
  );


  not
  g2561
  (
    n2469,
    n2342
  );


  buf
  g2562
  (
    n2528,
    n2312
  );


  buf
  g2563
  (
    n2694,
    n2319
  );


  not
  g2564
  (
    n2434,
    n2415
  );


  not
  g2565
  (
    n2688,
    n2318
  );


  buf
  g2566
  (
    n2629,
    n2316
  );


  buf
  g2567
  (
    n2443,
    n2402
  );


  not
  g2568
  (
    n2597,
    n2327
  );


  buf
  g2569
  (
    n2606,
    n2354
  );


  not
  g2570
  (
    n2497,
    n2256
  );


  not
  g2571
  (
    n2596,
    n2419
  );


  not
  g2572
  (
    n2447,
    n2380
  );


  buf
  g2573
  (
    n2569,
    n2389
  );


  not
  g2574
  (
    n2703,
    n2369
  );


  buf
  g2575
  (
    n2656,
    n2381
  );


  not
  g2576
  (
    n2427,
    n2357
  );


  buf
  g2577
  (
    n2696,
    n2406
  );


  buf
  g2578
  (
    n2588,
    n2336
  );


  not
  g2579
  (
    n2551,
    n2421
  );


  not
  g2580
  (
    n2540,
    n2334
  );


  not
  g2581
  (
    n2710,
    n2348
  );


  buf
  g2582
  (
    n2633,
    n2330
  );


  not
  g2583
  (
    n2544,
    n2413
  );


  not
  g2584
  (
    n2685,
    n2410
  );


  buf
  g2585
  (
    n2709,
    n1505
  );


  buf
  g2586
  (
    n2659,
    n2380
  );


  not
  g2587
  (
    n2539,
    n2372
  );


  buf
  g2588
  (
    n2637,
    n2324
  );


  buf
  g2589
  (
    n2670,
    n2395
  );


  buf
  g2590
  (
    n2702,
    n2424
  );


  buf
  g2591
  (
    n2514,
    n2401
  );


  buf
  g2592
  (
    n2614,
    n2377
  );


  not
  g2593
  (
    n2622,
    n2318
  );


  buf
  g2594
  (
    n2430,
    n2356
  );


  buf
  g2595
  (
    n2472,
    n2363
  );


  not
  g2596
  (
    n2511,
    n2308
  );


  not
  g2597
  (
    n2715,
    n2369
  );


  not
  g2598
  (
    n2440,
    n2334
  );


  buf
  g2599
  (
    n2425,
    n2385
  );


  not
  g2600
  (
    n2701,
    n2364
  );


  not
  g2601
  (
    n2534,
    n2365
  );


  buf
  g2602
  (
    n2627,
    n2302
  );


  not
  g2603
  (
    n2535,
    n2297
  );


  buf
  g2604
  (
    n2557,
    n2313
  );


  and
  g2605
  (
    n2678,
    n2403,
    n2377,
    n2313
  );


  xor
  g2606
  (
    n2499,
    n2311,
    n2319,
    n2381
  );


  nor
  g2607
  (
    n2634,
    n2420,
    n2357,
    n2300,
    n2416
  );


  xnor
  g2608
  (
    n2683,
    n2325,
    n2347,
    n2344,
    n2304
  );


  xnor
  g2609
  (
    n2464,
    n2386,
    n2309,
    n2353,
    n2378
  );


  or
  g2610
  (
    n2612,
    n2418,
    n2297,
    n2376,
    n2408
  );


  or
  g2611
  (
    n2439,
    n2306,
    n2385,
    n2389,
    n2395
  );


  nor
  g2612
  (
    n2436,
    n2395,
    n2308,
    n2370,
    n2368
  );


  nor
  g2613
  (
    n2711,
    n2366,
    n2410
  );


  nand
  g2614
  (
    n2491,
    n2407,
    n2407,
    n2423,
    n2409
  );


  nor
  g2615
  (
    n2719,
    n1507,
    n2320,
    n2373,
    n2332
  );


  and
  g2616
  (
    n2515,
    n2254,
    n2399,
    n2337,
    n1503
  );


  and
  g2617
  (
    n2432,
    n2359,
    n2372,
    n2310,
    n2375
  );


  or
  g2618
  (
    n2603,
    n2301,
    n2407,
    n2330,
    n2383
  );


  or
  g2619
  (
    n2441,
    n2332,
    n2371,
    n2315,
    n2421
  );


  xor
  g2620
  (
    n2686,
    n2341,
    n2398,
    n2301,
    n2399
  );


  xnor
  g2621
  (
    n2708,
    n2385,
    n1502,
    n2403,
    n1505
  );


  nand
  g2622
  (
    n2465,
    n2400,
    n2340,
    n2417,
    n2392
  );


  and
  g2623
  (
    n2479,
    n2371,
    n2374,
    n2399,
    n2386
  );


  or
  g2624
  (
    n2524,
    n2367,
    n2378,
    n2255,
    n2400
  );


  and
  g2625
  (
    n2550,
    n2142,
    n2253,
    n2391,
    n2336
  );


  xnor
  g2626
  (
    n2462,
    n2357,
    n2419,
    n2342,
    n2364
  );


  xnor
  g2627
  (
    n2561,
    n2415,
    n2345,
    n2323,
    n2331
  );


  and
  g2628
  (
    n2571,
    n2309,
    n2320,
    n1506,
    n2359
  );


  xor
  g2629
  (
    n2600,
    n2319,
    n2326,
    n2308,
    n2399
  );


  and
  g2630
  (
    n2448,
    n2372,
    n2304,
    n2353,
    n2406
  );


  xnor
  g2631
  (
    n2587,
    n2255,
    n2306,
    n2368,
    n2310
  );


  nand
  g2632
  (
    n2602,
    n2369,
    n2350,
    n2361
  );


  xor
  g2633
  (
    n2654,
    n2329,
    n2417,
    n2343,
    n2375
  );


  nor
  g2634
  (
    n2555,
    n2363,
    n2312,
    n2332,
    n2360
  );


  nand
  g2635
  (
    n2503,
    n2409,
    n2392,
    n2313,
    n2357
  );


  nand
  g2636
  (
    n2689,
    n2321,
    n2351,
    n2393,
    n2411
  );


  nor
  g2637
  (
    n2548,
    n2345,
    n2379,
    n2331,
    n2382
  );


  or
  g2638
  (
    n2608,
    n2406,
    n2307,
    n2322,
    n2301
  );


  xnor
  g2639
  (
    n2510,
    n2358,
    n2422,
    n2416,
    n1504
  );


  nor
  g2640
  (
    n2631,
    n2396,
    n2366,
    n2303,
    n2368
  );


  xor
  g2641
  (
    n2610,
    n2340,
    n2414,
    n2355,
    n2324
  );


  xor
  g2642
  (
    n2657,
    n2354,
    n2318,
    n2351,
    n2315
  );


  nor
  g2643
  (
    n2565,
    n2344,
    n2254,
    n2405,
    n2328
  );


  xnor
  g2644
  (
    n2639,
    n2390,
    n2408,
    n2371,
    n2327
  );


  xnor
  g2645
  (
    n2476,
    n2309,
    n2405,
    n2370,
    n2383
  );


  or
  g2646
  (
    n2601,
    n1507,
    n2311,
    n2365,
    n2342
  );


  xnor
  g2647
  (
    n2428,
    n2388,
    n2380,
    n2405,
    n2360
  );


  nor
  g2648
  (
    n2591,
    n2337,
    n2414,
    n1507,
    n2341
  );


  xor
  g2649
  (
    n2531,
    n2338,
    n2305,
    n2375,
    n2401
  );


  xnor
  g2650
  (
    n2677,
    n2356,
    n1506,
    n2392,
    n2360
  );


  xor
  g2651
  (
    n2716,
    n2330,
    n2303,
    n2342,
    n2355
  );


  and
  g2652
  (
    n2667,
    n2402,
    n1503,
    n2413,
    n2325
  );


  xor
  g2653
  (
    n2487,
    n2387,
    n2313,
    n2337,
    n2377
  );


  xnor
  g2654
  (
    n2649,
    n2333,
    n2316,
    n2370
  );


  nor
  g2655
  (
    n2566,
    n2397,
    n2345,
    n2348,
    n2374
  );


  nand
  g2656
  (
    n2429,
    n2354,
    n1506,
    n1508,
    n2346
  );


  xnor
  g2657
  (
    n2666,
    n2394,
    n2398,
    n2304,
    n2355
  );


  and
  g2658
  (
    n2495,
    n2352,
    n1508,
    n2373,
    n2300
  );


  xnor
  g2659
  (
    n2589,
    n2391,
    n2379,
    n2422,
    n2297
  );


  and
  g2660
  (
    n2584,
    n2404,
    n2339,
    n2304,
    n2358
  );


  nand
  g2661
  (
    n2679,
    n2340,
    n2349,
    n2322,
    n2367
  );


  xor
  g2662
  (
    n2691,
    n2386,
    n2384,
    n2362,
    n2254
  );


  nor
  g2663
  (
    n2721,
    n2298,
    n2423,
    n2420,
    n2389
  );


  and
  g2664
  (
    n2451,
    n2325,
    n2373,
    n2374,
    n1503
  );


  or
  g2665
  (
    n2526,
    n2401,
    n2346,
    n2383,
    n2379
  );


  and
  g2666
  (
    n2599,
    n2356,
    n2410,
    n2307,
    n2413
  );


  xor
  g2667
  (
    n2642,
    n2307,
    n2347,
    n2417,
    n2335
  );


  and
  g2668
  (
    n2516,
    n2339,
    n2325,
    n2379,
    n2329
  );


  and
  g2669
  (
    n2609,
    n2331,
    n2374,
    n2387,
    n2359
  );


  xnor
  g2670
  (
    n2542,
    n2390,
    n2377,
    n2338,
    n2384
  );


  or
  g2671
  (
    n2652,
    n2371,
    n2365,
    n2321,
    n2353
  );


  xor
  g2672
  (
    n2630,
    n2308,
    n2143,
    n1505,
    n2299
  );


  nand
  g2673
  (
    n2722,
    n2414,
    n2409,
    n2349,
    n2331
  );


  xor
  g2674
  (
    n2653,
    n2317,
    n1502,
    n2335,
    n2387
  );


  nand
  g2675
  (
    n2592,
    n2299,
    n2402,
    n2397,
    n2327
  );


  or
  g2676
  (
    n2717,
    n2409,
    n2299,
    n2381,
    n2311
  );


  xor
  g2677
  (
    n2660,
    n2309,
    n2413,
    n2364,
    n2343
  );


  xnor
  g2678
  (
    n2635,
    n2298,
    n2386,
    n2353,
    n2368
  );


  xor
  g2679
  (
    n2460,
    n2423,
    n2358,
    n2367,
    n2361
  );


  xnor
  g2680
  (
    n2572,
    n2407,
    n2306,
    n1504,
    n2324
  );


  or
  g2681
  (
    n2480,
    n2352,
    n2370,
    n2255,
    n2369
  );


  nand
  g2682
  (
    n2478,
    n2334,
    n2317,
    n2391,
    n2354
  );


  nand
  g2683
  (
    n2504,
    n2348,
    n2415,
    n2328,
    n2421
  );


  nand
  g2684
  (
    n2700,
    n1507,
    n2362,
    n2305,
    n2318
  );


  and
  g2685
  (
    n2697,
    n2334,
    n2333,
    n2422,
    n2398
  );


  and
  g2686
  (
    n2676,
    n2404,
    n2424,
    n2400,
    n2406
  );


  nor
  g2687
  (
    n2651,
    n2315,
    n2351,
    n2373,
    n2322
  );


  xnor
  g2688
  (
    n2556,
    n2303,
    n2344,
    n2419,
    n2396
  );


  xnor
  g2689
  (
    n2458,
    n2307,
    n2396,
    n2338,
    n2361
  );


  nor
  g2690
  (
    n2723,
    n2425,
    n2426
  );


  or
  g2691
  (
    n2724,
    n2144,
    n2723,
    n2146,
    n2145
  );


  and
  g2692
  (
    n2725,
    n2148,
    n2724
  );


  or
  g2693
  (
    n2726,
    n2431,
    n2428,
    n2427,
    n2434
  );


  and
  g2694
  (
    n2727,
    n2430,
    n2429,
    n2436,
    n2432
  );


  nor
  g2695
  (
    n2728,
    n2435,
    n2433,
    n2724,
    n2147
  );


  and
  g2696
  (
    n2730,
    n2446,
    n2728,
    n2453,
    n2441
  );


  or
  g2697
  (
    n2732,
    n2449,
    n2450,
    n2448,
    n2728
  );


  or
  g2698
  (
    n2736,
    n2728,
    n2437,
    n2725,
    n2445
  );


  xor
  g2699
  (
    n2733,
    n2728,
    n2458,
    n2443,
    n2727
  );


  nand
  g2700
  (
    n2729,
    n2456,
    n2452,
    n2454,
    n2439
  );


  nor
  g2701
  (
    n2735,
    n2447,
    n2727,
    n2442,
    n2457
  );


  and
  g2702
  (
    n2734,
    n2438,
    n2451,
    n2459,
    n2455
  );


  nor
  g2703
  (
    n2731,
    n2460,
    n2726,
    n2444,
    n2440
  );


  nand
  g2704
  (
    n2742,
    n1711,
    n1709,
    n2172,
    n1710
  );


  nor
  g2705
  (
    n2751,
    n2179,
    n2152,
    n2151,
    n1702
  );


  xor
  g2706
  (
    n2743,
    n2736,
    n2163,
    n1710,
    n1714
  );


  nor
  g2707
  (
    n2756,
    n2733,
    n2171,
    n2174,
    n1704
  );


  xnor
  g2708
  (
    n2764,
    n2736,
    n2180,
    n1714,
    n2733
  );


  xnor
  g2709
  (
    n2740,
    n1704,
    n2732,
    n1706,
    n1701
  );


  and
  g2710
  (
    n2761,
    n2735,
    n2463,
    n1713,
    n1700
  );


  xor
  g2711
  (
    n2768,
    n1705,
    n2735,
    n2729,
    n1713
  );


  nor
  g2712
  (
    n2745,
    n1703,
    n1711,
    n2730,
    n2176
  );


  or
  g2713
  (
    n2757,
    n2729,
    n1706,
    n2730,
    n2732
  );


  nor
  g2714
  (
    n2766,
    n2165,
    n2162,
    n2736,
    n1707
  );


  and
  g2715
  (
    n2767,
    n1708,
    n1714,
    n2166,
    n2730
  );


  xor
  g2716
  (
    n2759,
    n2731,
    n1699,
    n1708,
    n2178
  );


  nand
  g2717
  (
    n2753,
    n2731,
    n1699,
    n1701,
    n2164
  );


  nor
  g2718
  (
    n2739,
    n2732,
    n1705,
    n1708,
    n2154
  );


  and
  g2719
  (
    n2754,
    n2156,
    n1707,
    n2734,
    n2175
  );


  or
  g2720
  (
    n2752,
    n1704,
    n2177,
    n2169,
    n1708
  );


  xor
  g2721
  (
    n2737,
    n1710,
    n2150,
    n1702,
    n1707
  );


  xor
  g2722
  (
    n2744,
    n1705,
    n1704,
    n2735,
    n1701
  );


  xnor
  g2723
  (
    n2748,
    n1711,
    n1703,
    n2729,
    n2170
  );


  xor
  g2724
  (
    n2763,
    n1710,
    n1706,
    n2161,
    n2462
  );


  xor
  g2725
  (
    n2765,
    n1712,
    n2173,
    n2158,
    n2157
  );


  xor
  g2726
  (
    n2741,
    n1706,
    n2729,
    n2732,
    n2734
  );


  and
  g2727
  (
    n2762,
    n2461,
    n2159,
    n2730,
    n2149
  );


  nand
  g2728
  (
    n2747,
    n2733,
    n1705,
    n2168,
    n1702
  );


  xnor
  g2729
  (
    n2749,
    n1701,
    n1703,
    n1713,
    n2733
  );


  nor
  g2730
  (
    n2750,
    n1712,
    n1712,
    n2736,
    n2160
  );


  xnor
  g2731
  (
    n2746,
    n2731,
    n2734,
    n2735,
    n1702
  );


  nor
  g2732
  (
    n2738,
    n1713,
    n1709,
    n1711,
    n1703
  );


  xor
  g2733
  (
    n2760,
    n2734,
    n1709,
    n1700
  );


  xnor
  g2734
  (
    n2758,
    n1700,
    n2731,
    n1709,
    n2155
  );


  or
  g2735
  (
    n2755,
    n2153,
    n2167,
    n1712,
    n1707
  );


  xnor
  g2736
  (
    n2775,
    n2759,
    n2760,
    n2758,
    n2762
  );


  and
  g2737
  (
    n2779,
    n2182,
    n2757,
    n2746,
    n2737
  );


  and
  g2738
  (
    n2781,
    n2747,
    n2764,
    n2184,
    n2765
  );


  or
  g2739
  (
    n2774,
    n2764,
    n2766,
    n2188,
    n2763
  );


  or
  g2740
  (
    n2780,
    n2754,
    n2192,
    n2185,
    n2767
  );


  and
  g2741
  (
    n2777,
    n2767,
    n2183,
    n2186,
    n2766
  );


  xor
  g2742
  (
    n2773,
    n2764,
    n2767,
    n2187,
    n2766
  );


  and
  g2743
  (
    n2772,
    n2738,
    n2749,
    n2750,
    n2765
  );


  or
  g2744
  (
    n2770,
    n2745,
    n2764,
    n2740,
    n2191
  );


  xnor
  g2745
  (
    n2769,
    n2755,
    n2753,
    n2756,
    n2766
  );


  xnor
  g2746
  (
    n2778,
    n2752,
    n2189,
    n2768,
    n2742
  );


  nor
  g2747
  (
    n2782,
    n2748,
    n2181,
    n2739,
    n2190
  );


  nor
  g2748
  (
    n2771,
    n2767,
    n2751,
    n2741,
    n2765
  );


  xnor
  g2749
  (
    n2776,
    n2765,
    n2743,
    n2761,
    n2744
  );


  buf
  g2750
  (
    n2788,
    n2780
  );


  buf
  g2751
  (
    n2793,
    n2782
  );


  not
  g2752
  (
    n2783,
    n2777
  );


  not
  g2753
  (
    n2795,
    n2780
  );


  not
  g2754
  (
    n2798,
    n2780
  );


  not
  g2755
  (
    n2796,
    n2782
  );


  not
  g2756
  (
    n2803,
    n2776
  );


  buf
  g2757
  (
    n2797,
    n2781
  );


  buf
  g2758
  (
    n2801,
    n2781
  );


  buf
  g2759
  (
    n2789,
    n2779
  );


  not
  g2760
  (
    n2786,
    n2769
  );


  not
  g2761
  (
    n2792,
    n2781
  );


  buf
  g2762
  (
    n2804,
    n2770
  );


  not
  g2763
  (
    n2784,
    n2782
  );


  not
  g2764
  (
    n2787,
    n2780
  );


  not
  g2765
  (
    n2785,
    n2781
  );


  buf
  g2766
  (
    n2805,
    n2773
  );


  buf
  g2767
  (
    n2802,
    n2772
  );


  buf
  g2768
  (
    n2794,
    n2778
  );


  buf
  g2769
  (
    n2791,
    n2782
  );


  buf
  g2770
  (
    n2790,
    n2775
  );


  not
  g2771
  (
    n2799,
    n2774
  );


  xnor
  g2772
  (
    n2800,
    n2771,
    n2256
  );


  not
  g2773
  (
    n2815,
    n2803
  );


  not
  g2774
  (
    n2808,
    n2804
  );


  buf
  g2775
  (
    n2824,
    n2803
  );


  buf
  g2776
  (
    n2835,
    n2805
  );


  buf
  g2777
  (
    n2821,
    n2209
  );


  not
  g2778
  (
    n2813,
    n2798
  );


  not
  g2779
  (
    n2832,
    n2787
  );


  buf
  g2780
  (
    n2819,
    n2783
  );


  not
  g2781
  (
    n2837,
    n2200
  );


  not
  g2782
  (
    n2812,
    n2215
  );


  buf
  g2783
  (
    n2816,
    n2804
  );


  not
  g2784
  (
    n2820,
    n2202
  );


  buf
  g2785
  (
    n2806,
    n2206
  );


  buf
  g2786
  (
    n2810,
    n2207
  );


  buf
  g2787
  (
    n2807,
    n2205
  );


  buf
  g2788
  (
    n2829,
    n2790
  );


  not
  g2789
  (
    n2841,
    n2219
  );


  buf
  g2790
  (
    n2836,
    n2788
  );


  not
  g2791
  (
    n2826,
    n2802
  );


  buf
  g2792
  (
    n2825,
    n2212
  );


  buf
  g2793
  (
    n2822,
    n2793
  );


  not
  g2794
  (
    n2838,
    n2216
  );


  not
  g2795
  (
    n2823,
    n2797
  );


  not
  g2796
  (
    n2842,
    n2799
  );


  not
  g2797
  (
    KeyWire_0_9,
    n2210
  );


  not
  g2798
  (
    n2814,
    n2805
  );


  buf
  g2799
  (
    n2840,
    n2195
  );


  buf
  g2800
  (
    n2843,
    n2804
  );


  xor
  g2801
  (
    n2827,
    n2218,
    n2805
  );


  or
  g2802
  (
    n2834,
    n2800,
    n2203,
    n2789,
    n2794
  );


  xnor
  g2803
  (
    n2817,
    n2193,
    n2803,
    n2791,
    n2211
  );


  nand
  g2804
  (
    n2833,
    n2213,
    n2220,
    n2802,
    n2201
  );


  and
  g2805
  (
    n2818,
    n2217,
    n2802,
    n2784,
    n2804
  );


  nor
  g2806
  (
    n2809,
    n2786,
    n2796,
    n2214,
    n2204
  );


  xor
  g2807
  (
    n2839,
    n2198,
    n2801,
    n2197
  );


  nand
  g2808
  (
    n2828,
    n2792,
    n2802,
    n2199,
    n2208
  );


  nand
  g2809
  (
    n2831,
    n2196,
    n2795,
    n2803,
    n2785
  );


  or
  g2810
  (
    n2811,
    n2805,
    n2801,
    n2194
  );


  nand
  g2811
  (
    n2844,
    n2806,
    n1716,
    n2811,
    n2831
  );


  nor
  g2812
  (
    n2852,
    n1715,
    n2817,
    n2822,
    n2819
  );


  nor
  g2813
  (
    n2848,
    n2826,
    n2827,
    n2816,
    n1716
  );


  nor
  g2814
  (
    n2850,
    n2813,
    n2808,
    n2820,
    n2814
  );


  xor
  g2815
  (
    n2849,
    n2812,
    n2807,
    n2809,
    n1715
  );


  nor
  g2816
  (
    n2847,
    n1715,
    n2832,
    n1716,
    n2824
  );


  nor
  g2817
  (
    n2851,
    n2828,
    n2810,
    n2825,
    n2821
  );


  and
  g2818
  (
    n2846,
    n2815,
    n2818,
    n1716,
    n2823
  );


  xor
  g2819
  (
    n2845,
    n2829,
    n1714,
    n2830,
    n1715
  );


  and
  g2820
  (
    n2853,
    n2221,
    n2852
  );


  nor
  g2821
  (
    n2856,
    n2471,
    n2464,
    n2467,
    n2475
  );


  nand
  g2822
  (
    n2857,
    n2474,
    n2472,
    n2465,
    n2853
  );


  xnor
  g2823
  (
    n2854,
    n2853,
    n2853,
    n2466,
    n2469
  );


  xor
  g2824
  (
    n2855,
    n2470,
    n2473,
    n2853,
    n2468
  );


  or
  g2825
  (
    n2868,
    n2839,
    n2236,
    n2843,
    n2857
  );


  nor
  g2826
  (
    n2867,
    n2842,
    n2238,
    n2840,
    n2854
  );


  xor
  g2827
  (
    n2864,
    n2245,
    n2239,
    n2840,
    n2241
  );


  xor
  g2828
  (
    n2858,
    n2856,
    n2834,
    n2855,
    n2857
  );


  nor
  g2829
  (
    n2861,
    n2243,
    n2841,
    n2835,
    n2245
  );


  and
  g2830
  (
    n2862,
    n2768,
    n2856,
    n2243,
    n2843
  );


  nor
  g2831
  (
    n2870,
    n2244,
    n2245,
    n2854
  );


  nand
  g2832
  (
    n2871,
    n2842,
    n2842,
    n2839,
    n2244
  );


  and
  g2833
  (
    n2869,
    n2234,
    n2856,
    n2857,
    n2840
  );


  and
  g2834
  (
    n2865,
    n2839,
    n2854,
    n2855,
    n2833
  );


  nand
  g2835
  (
    n2866,
    n2244,
    n2768,
    n2838,
    n2237
  );


  xor
  g2836
  (
    n2872,
    n2244,
    n2837,
    n2240,
    n2233
  );


  and
  g2837
  (
    n2873,
    n2856,
    n2841,
    n2768,
    n2235
  );


  and
  g2838
  (
    n2863,
    n2839,
    n2854,
    n2836,
    n2855
  );


  xor
  g2839
  (
    n2859,
    n2855,
    n2841,
    n2857
  );


  nor
  g2840
  (
    n2860,
    n2840,
    n2843,
    n2842
  );


  not
  g2841
  (
    n2877,
    n2869
  );


  buf
  g2842
  (
    n2890,
    n2862
  );


  not
  g2843
  (
    n2897,
    n2865
  );


  not
  g2844
  (
    n2925,
    n2864
  );


  buf
  g2845
  (
    n2884,
    n2868
  );


  buf
  g2846
  (
    n2922,
    n2873
  );


  not
  g2847
  (
    n2904,
    n2872
  );


  buf
  g2848
  (
    n2907,
    n2859
  );


  not
  g2849
  (
    n2893,
    n2863
  );


  buf
  g2850
  (
    n2902,
    n2480
  );


  not
  g2851
  (
    n2892,
    n2859
  );


  not
  g2852
  (
    n2911,
    n2242
  );


  buf
  g2853
  (
    n2886,
    n2873
  );


  not
  g2854
  (
    n2898,
    n2861
  );


  not
  g2855
  (
    n2894,
    n2870
  );


  buf
  g2856
  (
    n2903,
    n2867
  );


  buf
  g2857
  (
    n2908,
    n2867
  );


  not
  g2858
  (
    n2927,
    n2867
  );


  buf
  g2859
  (
    n2914,
    n2863
  );


  not
  g2860
  (
    n2915,
    n2865
  );


  not
  g2861
  (
    n2891,
    n2864
  );


  not
  g2862
  (
    n2887,
    n2869
  );


  buf
  g2863
  (
    n2888,
    n2871
  );


  not
  g2864
  (
    n2923,
    n2866
  );


  not
  g2865
  (
    n2924,
    n2864
  );


  buf
  g2866
  (
    n2918,
    n2868
  );


  buf
  g2867
  (
    n2917,
    n2477
  );


  buf
  g2868
  (
    n2910,
    n2861
  );


  not
  g2869
  (
    n2916,
    n2870
  );


  not
  g2870
  (
    n2921,
    n2865
  );


  not
  g2871
  (
    n2899,
    n2859
  );


  buf
  g2872
  (
    n2913,
    n2872
  );


  buf
  g2873
  (
    n2919,
    n2866
  );


  not
  g2874
  (
    n2909,
    n2872
  );


  buf
  g2875
  (
    n2926,
    n2860
  );


  buf
  g2876
  (
    n2875,
    n2858
  );


  buf
  g2877
  (
    n2880,
    n2872
  );


  buf
  g2878
  (
    n2900,
    n2481
  );


  not
  g2879
  (
    n2882,
    n2870
  );


  buf
  g2880
  (
    n2883,
    n2479
  );


  not
  g2881
  (
    n2905,
    n2866
  );


  buf
  g2882
  (
    n2912,
    n2859
  );


  not
  g2883
  (
    n2885,
    n2864
  );


  not
  g2884
  (
    n2881,
    n2873
  );


  not
  g2885
  (
    n2874,
    n2860
  );


  buf
  g2886
  (
    n2929,
    n2866
  );


  not
  g2887
  (
    n2895,
    n2867
  );


  buf
  g2888
  (
    n2889,
    n2862
  );


  not
  g2889
  (
    n2901,
    n2424
  );


  not
  g2890
  (
    n2878,
    n2869
  );


  nor
  g2891
  (
    n2896,
    n2861,
    n2871,
    n2424,
    n2858
  );


  nor
  g2892
  (
    n2920,
    n2863,
    n2865,
    n2858
  );


  xnor
  g2893
  (
    n2879,
    n2862,
    n2871,
    n2478,
    n2482
  );


  nor
  g2894
  (
    n2876,
    n2868,
    n2870,
    n2862,
    n2476
  );


  or
  g2895
  (
    n2906,
    n2868,
    n2860,
    n2873,
    n2871
  );


  nand
  g2896
  (
    n2928,
    n2860,
    n2863,
    n2861,
    n2869
  );


  xor
  g2897
  (
    n2935,
    n2666,
    n2917,
    n2536,
    n2537
  );


  or
  g2898
  (
    n2980,
    n2497,
    n2628,
    n2664,
    n2541
  );


  xor
  g2899
  (
    n2981,
    n2710,
    n2702,
    n2609,
    n2606
  );


  nand
  g2900
  (
    n2963,
    n2923,
    n2650,
    n2926,
    n2640
  );


  and
  g2901
  (
    n3007,
    n2922,
    n2530,
    n2576,
    n2691
  );


  or
  g2902
  (
    n2991,
    n2910,
    n2543,
    n2544,
    n2717
  );


  nor
  g2903
  (
    n2932,
    n2928,
    n2714,
    n2574,
    n2908
  );


  nor
  g2904
  (
    n2936,
    n2894,
    n2711,
    n2565,
    n2885
  );


  nor
  g2905
  (
    n3006,
    n2644,
    n2923,
    n2491,
    n2903
  );


  xnor
  g2906
  (
    n2942,
    n2487,
    n2629,
    n2922,
    n2483
  );


  or
  g2907
  (
    n2931,
    n2688,
    n2920,
    n2578,
    n2895
  );


  or
  g2908
  (
    n2973,
    n2587,
    n2658,
    n2712,
    n2689
  );


  xnor
  g2909
  (
    n2962,
    n2637,
    n2614,
    n2561,
    n2919
  );


  nor
  g2910
  (
    n2950,
    n2879,
    n2501,
    n2676,
    n2504
  );


  or
  g2911
  (
    n3009,
    n2890,
    n2655,
    n2551,
    n2661
  );


  or
  g2912
  (
    n2979,
    n2569,
    n2534,
    n2613,
    n2566
  );


  xnor
  g2913
  (
    n2995,
    n2602,
    n2696,
    n2485,
    n2620
  );


  or
  g2914
  (
    n2940,
    n2708,
    n2625,
    n2542,
    n2592
  );


  xor
  g2915
  (
    n2941,
    n2900,
    n2580,
    n2627,
    n2589
  );


  nand
  g2916
  (
    n2951,
    n2887,
    n2539,
    n2924,
    n2678
  );


  and
  g2917
  (
    n2983,
    n2904,
    n2921,
    n2646,
    n2682
  );


  nand
  g2918
  (
    n2985,
    n2707,
    n2510,
    n2926,
    n2719
  );


  nor
  g2919
  (
    n2975,
    n2925,
    n2502,
    n2503,
    n2686
  );


  xor
  g2920
  (
    n2961,
    n2700,
    n2924,
    n2633,
    n2572
  );


  nor
  g2921
  (
    n2974,
    n2486,
    n2680,
    n2877,
    n2642
  );


  xnor
  g2922
  (
    n2955,
    n2925,
    n2671,
    n2926,
    n2520
  );


  nand
  g2923
  (
    n2971,
    n2560,
    n2594,
    n2553,
    n2571
  );


  and
  g2924
  (
    n2987,
    n2923,
    n2703,
    n2892,
    n2701
  );


  or
  g2925
  (
    n2957,
    n2662,
    n2876,
    n2564,
    n2590
  );


  xnor
  g2926
  (
    n2947,
    n2493,
    n2922,
    n2718,
    n2660
  );


  nor
  g2927
  (
    n2978,
    n2909,
    n2639,
    n2902,
    n2545
  );


  xor
  g2928
  (
    n2943,
    n2713,
    n2500,
    n2929,
    n2654
  );


  xor
  g2929
  (
    n2964,
    n2923,
    n2618,
    n2684,
    n2605
  );


  and
  g2930
  (
    n2977,
    n2511,
    n2555,
    n2911,
    n2695
  );


  or
  g2931
  (
    n2993,
    n2535,
    n2626,
    n2874,
    n2907
  );


  or
  g2932
  (
    n2956,
    n2704,
    n2657,
    n2693,
    n2600
  );


  nor
  g2933
  (
    n2946,
    n2906,
    n2880,
    n2652,
    n2494
  );


  xnor
  g2934
  (
    n2998,
    n2913,
    n2547,
    n2706,
    n2490
  );


  nand
  g2935
  (
    n2953,
    n2489,
    n2897,
    n2922,
    n2916
  );


  xor
  g2936
  (
    n2930,
    n2531,
    n2929,
    n2518,
    n2601
  );


  xor
  g2937
  (
    n2969,
    n2488,
    n2549,
    n2683,
    n2591
  );


  xor
  g2938
  (
    n2939,
    n2653,
    n2577,
    n2929,
    n2882
  );


  and
  g2939
  (
    n2999,
    n2912,
    n2881,
    n2581,
    n2681
  );


  and
  g2940
  (
    n2954,
    n2550,
    n2675,
    n2603,
    n2679
  );


  nand
  g2941
  (
    n2988,
    n2532,
    n2888,
    n2611,
    n2610
  );


  and
  g2942
  (
    n2986,
    n2599,
    n2925,
    n2616,
    n2573
  );


  xnor
  g2943
  (
    n3001,
    n2673,
    n2538,
    n2694,
    n2516
  );


  xor
  g2944
  (
    n2938,
    n2548,
    n2635,
    n2495,
    n2540
  );


  xnor
  g2945
  (
    n2965,
    n2604,
    n2690,
    n2630,
    n2677
  );


  and
  g2946
  (
    n2972,
    n2685,
    n2927,
    n2558,
    n2659
  );


  or
  g2947
  (
    n2967,
    n2579,
    n2886,
    n2899,
    n2674
  );


  and
  g2948
  (
    n2992,
    n2883,
    n2927,
    n2567,
    n2515
  );


  xnor
  g2949
  (
    n3002,
    n2722,
    n2575,
    n2891,
    n2559
  );


  xor
  g2950
  (
    n3004,
    n2631,
    n2656,
    n2612,
    n2586
  );


  xor
  g2951
  (
    n3008,
    n2529,
    n2632,
    n2557,
    n2492
  );


  nor
  g2952
  (
    n2997,
    n2905,
    n2928,
    n2929,
    n2584
  );


  xnor
  g2953
  (
    n2989,
    n2505,
    n2716,
    n2697,
    n2915
  );


  nor
  g2954
  (
    n2949,
    n2512,
    n2498,
    n2509,
    n2608
  );


  nand
  g2955
  (
    n2945,
    n2526,
    n2552,
    n2617,
    n2667
  );


  xor
  g2956
  (
    n3000,
    n2507,
    n2598,
    n2670,
    n2663
  );


  xnor
  g2957
  (
    n2937,
    n2499,
    n2928,
    n2506,
    n2562
  );


  nor
  g2958
  (
    n2966,
    n2926,
    n2924,
    n2699,
    n2546
  );


  or
  g2959
  (
    n2970,
    n2918,
    n2525,
    n2597,
    n2593
  );


  and
  g2960
  (
    n2990,
    n2568,
    n2508,
    n2641,
    n2636
  );


  nor
  g2961
  (
    n2960,
    n2709,
    n2927,
    n2875,
    n2582
  );


  nand
  g2962
  (
    n2982,
    n2647,
    n2583,
    n2687,
    n2533
  );


  xnor
  g2963
  (
    n2959,
    n2896,
    n2721,
    n2715,
    n2517
  );


  nor
  g2964
  (
    n2994,
    n2901,
    n2924,
    n2698,
    n2893
  );


  or
  g2965
  (
    n2984,
    n2672,
    n2643,
    n2645,
    n2563
  );


  xnor
  g2966
  (
    n2952,
    n2669,
    n2668,
    n2665,
    n2928
  );


  or
  g2967
  (
    n2933,
    n2705,
    n2692,
    n2596,
    n2889
  );


  xnor
  g2968
  (
    n2958,
    n2595,
    n2528,
    n2484,
    n2585
  );


  and
  g2969
  (
    n2996,
    n2624,
    n2914,
    n2884,
    n2927
  );


  nor
  g2970
  (
    n3003,
    n2513,
    n2607,
    n2898,
    n2621
  );


  and
  g2971
  (
    n2948,
    n2878,
    n2514,
    n2556,
    n2588
  );


  and
  g2972
  (
    n2944,
    n2622,
    n2522,
    n2615,
    n2648
  );


  xnor
  g2973
  (
    n2934,
    n2554,
    n2634,
    n2570,
    n2649
  );


  xor
  g2974
  (
    n2976,
    n2651,
    n2521,
    n2524,
    n2623
  );


  xor
  g2975
  (
    n2968,
    n2925,
    n2519,
    n2523,
    n2720
  );


  xor
  g2976
  (
    n3005,
    n2527,
    n2619,
    n2496,
    n2638
  );


  xnor
  g2977
  (
    n3017,
    n3009,
    n2943,
    n2944,
    n2999
  );


  or
  g2978
  (
    n3018,
    n2951,
    n2969,
    n2976,
    n2977
  );


  xnor
  g2979
  (
    n3022,
    n2959,
    n2962,
    n2950,
    n2931
  );


  xor
  g2980
  (
    n3029,
    n2946,
    n3008,
    n2935,
    n3007
  );


  xnor
  g2981
  (
    n3014,
    n3007,
    n2939,
    n2970,
    n2997
  );


  xnor
  g2982
  (
    n3015,
    n2961,
    n2954,
    n3007,
    n2971
  );


  nand
  g2983
  (
    n3024,
    n2998,
    n2934,
    n2981,
    n2960
  );


  xor
  g2984
  (
    n3019,
    n3006,
    n2983,
    n2990,
    n2984
  );


  and
  g2985
  (
    n3025,
    n2973,
    n3007,
    n2938,
    n3009
  );


  xor
  g2986
  (
    n3016,
    n2930,
    n2933,
    n2979,
    n2987
  );


  nor
  g2987
  (
    n3021,
    n2966,
    n2978,
    n2952,
    n2985
  );


  xor
  g2988
  (
    n3030,
    n2975,
    n3002,
    n2936,
    n2982
  );


  nor
  g2989
  (
    n3020,
    n3008,
    n2956,
    n2986,
    n2955
  );


  or
  g2990
  (
    n3027,
    n3009,
    n2953,
    n2949,
    n2941
  );


  and
  g2991
  (
    n3032,
    n2988,
    n3004,
    n2967,
    n3006
  );


  xor
  g2992
  (
    n3013,
    n2937,
    n2940,
    n3008,
    n2948
  );


  and
  g2993
  (
    n3031,
    n2996,
    n3009,
    n2932,
    n2992
  );


  xor
  g2994
  (
    n3012,
    n3006,
    n3006,
    n2965,
    n3000
  );


  and
  g2995
  (
    n3026,
    n2993,
    n2964,
    n2974,
    n2980
  );


  nand
  g2996
  (
    n3028,
    n2989,
    n2995,
    n2991,
    n3008
  );


  and
  g2997
  (
    n3011,
    n2968,
    n2994,
    n2947,
    n3003
  );


  or
  g2998
  (
    n3023,
    n2963,
    n2972,
    n3005,
    n2958
  );


  and
  g2999
  (
    n3010,
    n3001,
    n2945,
    n2957,
    n2942
  );


  xor
  KeyGate_0_0
  (
    n560,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    KeyNOTWire_0_1,
    keyIn_0_1,
    KeyWire_0_1
  );


  not
  KeyNOTGate_0_1
  (
    n1664,
    KeyNOTWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n1547,
    keyIn_0_2,
    KeyWire_0_2
  );


  xnor
  KeyGate_0_3
  (
    n1461,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    KeyNOTWire_0_4,
    keyIn_0_4,
    KeyWire_0_4
  );


  not
  KeyNOTGate_0_4
  (
    n527,
    KeyNOTWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n2671,
    keyIn_0_5,
    KeyWire_0_5
  );


  xor
  KeyGate_0_6
  (
    n410,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    KeyNOTWire_0_7,
    keyIn_0_7,
    KeyWire_0_7
  );


  not
  KeyNOTGate_0_7
  (
    n498,
    KeyNOTWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    KeyNOTWire_0_8,
    keyIn_0_8,
    KeyWire_0_8
  );


  not
  KeyNOTGate_0_8
  (
    n802,
    KeyNOTWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    KeyNOTWire_0_9,
    keyIn_0_9,
    KeyWire_0_9
  );


  not
  KeyNOTGate_0_9
  (
    n2830,
    KeyNOTWire_0_9
  );


  xor
  KeyGate_0_10
  (
    KeyNOTWire_0_10,
    keyIn_0_10,
    KeyWire_0_10
  );


  not
  KeyNOTGate_0_10
  (
    n669,
    KeyNOTWire_0_10
  );


  xnor
  KeyGate_0_11
  (
    KeyNOTWire_0_11,
    keyIn_0_11,
    KeyWire_0_11
  );


  not
  KeyNOTGate_0_11
  (
    n1730,
    KeyNOTWire_0_11
  );


  xnor
  KeyGate_0_12
  (
    n1844,
    keyIn_0_12,
    KeyWire_0_12
  );


  xnor
  KeyGate_0_13
  (
    KeyNOTWire_0_13,
    keyIn_0_13,
    KeyWire_0_13
  );


  not
  KeyNOTGate_0_13
  (
    n727,
    KeyNOTWire_0_13
  );


  xor
  KeyGate_0_14
  (
    n2278,
    keyIn_0_14,
    KeyWire_0_14
  );


  xnor
  KeyGate_0_15
  (
    n334,
    keyIn_0_15,
    KeyWire_0_15
  );


endmodule


