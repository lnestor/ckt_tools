// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_45 written by SynthGen on 2021/04/05 11:08:37
module C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_45 ( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n101, n113, n83, n122, n93, n95, n86, n110,
 n84, n112, n99, n116, n121, n109, n114, n117,
 n120, n107, n106, n111, n118, n102, n128, n124,
 n127, n130, n131, n125, n132, n129, n126, n123);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n101, n113, n83, n122, n93, n95, n86, n110,
 n84, n112, n99, n116, n121, n109, n114, n117,
 n120, n107, n106, n111, n118, n102, n128, n124,
 n127, n130, n131, n125, n132, n129, n126, n123;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n85, n87, n88, n89, n90, n91,
 n92, n94, n96, n97, n98, n100, n103, n104,
 n105, n108, n115, n119;

not  g0 (n47, n2);
buf  g1 (n62, n3);
buf  g2 (n46, n16);
not  g3 (n52, n11);
buf  g4 (n42, n14);
buf  g5 (n61, n25);
buf  g6 (n37, n26);
not  g7 (n35, n29);
not  g8 (n56, n30);
buf  g9 (n58, n24);
buf  g10 (n64, n4);
buf  g11 (n45, n21);
buf  g12 (n33, n6);
buf  g13 (n40, n7);
buf  g14 (n38, n15);
buf  g15 (n63, n32);
not  g16 (n50, n23);
buf  g17 (n57, n9);
not  g18 (n65, n8);
not  g19 (n49, n32);
buf  g20 (n36, n17);
not  g21 (n51, n18);
not  g22 (n59, n20);
not  g23 (n48, n10);
buf  g24 (n66, n31);
buf  g25 (n44, n27);
not  g26 (n55, n1);
buf  g27 (n43, n28);
not  g28 (n41, n19);
buf  g29 (n60, n22);
buf  g30 (n34, n13);
buf  g31 (n53, n12);
buf  g32 (n54, n32);
buf  g33 (n39, n5);
not  g34 (n75, n33);
buf  g35 (n73, n36);
not  g36 (n68, n34);
buf  g37 (n79, n33);
buf  g38 (n80, n36);
buf  g39 (n69, n36);
not  g40 (n70, n36);
not  g41 (n77, n35);
buf  g42 (n67, n34);
not  g43 (n82, n34);
buf  g44 (n71, n35);
not  g45 (n81, n33);
buf  g46 (n72, n35);
not  g47 (n76, n35);
not  g48 (n78, n33);
not  g49 (n74, n34);
xor  g50 (n87, n77, n43, n51, n40);
and  g51 (n120, n71, n39, n41, n72);
or   g52 (n116, n53, n60, n57, n41);
nand g53 (n88, n54, n49, n79, n37);
nor  g54 (n121, n67, n80, n79, n48);
nand g55 (n98, n38, n50, n75, n61);
and  g56 (n100, n52, n45, n43, n73);
xor  g57 (n97, n60, n39, n50);
nor  g58 (n94, n65, n53, n66, n48);
nand g59 (n110, n79, n63, n66, n64);
and  g60 (n111, n59, n49, n41, n42);
nand g61 (n104, n42, n63, n73, n46);
and  g62 (n113, n48, n49, n59, n43);
xnor g63 (n114, n55, n79, n77, n66);
xnor g64 (n119, n40, n73, n52, n74);
nor  g65 (n117, n45, n76, n44);
nand g66 (n84, n37, n72, n77, n46);
nand g67 (n118, n62, n55, n47, n42);
nand g68 (n112, n72, n44, n74, n45);
nor  g69 (n106, n38, n40, n56);
xnor g70 (n90, n56, n75, n45, n78);
or   g71 (n83, n69, n64, n57, n55);
nand g72 (n105, n51, n77, n62, n78);
nand g73 (n86, n38, n51, n61, n75);
and  g74 (n108, n48, n54, n50);
or   g75 (n99, n74, n76, n44, n46);
nand g76 (n93, n61, n57, n59, n80);
xnor g77 (n115, n52, n37, n65, n78);
and  g78 (n92, n60, n65, n70, n63);
xor  g79 (n102, n58, n39, n37, n44);
xnor g80 (n95, n46, n74, n62, n78);
xnor g81 (n101, n54, n54, n64, n76);
and  g82 (n109, n56, n73, n62, n66);
xor  g83 (n85, n49, n61, n51, n75);
xnor g84 (n107, n43, n65, n59, n52);
and  g85 (n96, n58, n53, n57, n68);
nand g86 (n89, n58, n64, n47);
nand g87 (n91, n42, n47, n41, n63);
xor  g88 (n103, n53, n56, n80, n38);
nor  g89 (n122, n72, n58, n60, n55);
buf  g90 (n125, n114);
buf  g91 (n132, n81);
not  g92 (n126, n81);
buf  g93 (n129, n122);
xor  g94 (n130, n119, n110, n105, n106);
or   g95 (n128, n109, n82);
xor  g96 (n123, n81, n116, n107, n108);
and  g97 (n127, n81, n118, n111, n80);
xor  g98 (n124, n115, n113, n32, n121);
xor  g99 (n131, n120, n117, n112, n82);
endmodule
