// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_2000_303 written by SynthGen on 2021/04/05 11:23:41
module Stat_2000_303( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n442, n608, n1990, n2002, n1992, n1987, n1970, n1996,
 n1998, n1973, n1976, n1965, n1995, n1974, n1997, n1999,
 n1989, n1968, n1971, n1985, n2003, n1988, n2001, n1972,
 n1994, n2006, n2007, n2005, n2030, n2031, n2029, n2032);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n442, n608, n1990, n2002, n1992, n1987, n1970, n1996,
 n1998, n1973, n1976, n1965, n1995, n1974, n1997, n1999,
 n1989, n1968, n1971, n1985, n2003, n1988, n2001, n1972,
 n1994, n2006, n2007, n2005, n2030, n2031, n2029, n2032;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n79, n80,
 n81, n82, n83, n84, n85, n86, n87, n88,
 n89, n90, n91, n92, n93, n94, n95, n96,
 n97, n98, n99, n100, n101, n102, n103, n104,
 n105, n106, n107, n108, n109, n110, n111, n112,
 n113, n114, n115, n116, n117, n118, n119, n120,
 n121, n122, n123, n124, n125, n126, n127, n128,
 n129, n130, n131, n132, n133, n134, n135, n136,
 n137, n138, n139, n140, n141, n142, n143, n144,
 n145, n146, n147, n148, n149, n150, n151, n152,
 n153, n154, n155, n156, n157, n158, n159, n160,
 n161, n162, n163, n164, n165, n166, n167, n168,
 n169, n170, n171, n172, n173, n174, n175, n176,
 n177, n178, n179, n180, n181, n182, n183, n184,
 n185, n186, n187, n188, n189, n190, n191, n192,
 n193, n194, n195, n196, n197, n198, n199, n200,
 n201, n202, n203, n204, n205, n206, n207, n208,
 n209, n210, n211, n212, n213, n214, n215, n216,
 n217, n218, n219, n220, n221, n222, n223, n224,
 n225, n226, n227, n228, n229, n230, n231, n232,
 n233, n234, n235, n236, n237, n238, n239, n240,
 n241, n242, n243, n244, n245, n246, n247, n248,
 n249, n250, n251, n252, n253, n254, n255, n256,
 n257, n258, n259, n260, n261, n262, n263, n264,
 n265, n266, n267, n268, n269, n270, n271, n272,
 n273, n274, n275, n276, n277, n278, n279, n280,
 n281, n282, n283, n284, n285, n286, n287, n288,
 n289, n290, n291, n292, n293, n294, n295, n296,
 n297, n298, n299, n300, n301, n302, n303, n304,
 n305, n306, n307, n308, n309, n310, n311, n312,
 n313, n314, n315, n316, n317, n318, n319, n320,
 n321, n322, n323, n324, n325, n326, n327, n328,
 n329, n330, n331, n332, n333, n334, n335, n336,
 n337, n338, n339, n340, n341, n342, n343, n344,
 n345, n346, n347, n348, n349, n350, n351, n352,
 n353, n354, n355, n356, n357, n358, n359, n360,
 n361, n362, n363, n364, n365, n366, n367, n368,
 n369, n370, n371, n372, n373, n374, n375, n376,
 n377, n378, n379, n380, n381, n382, n383, n384,
 n385, n386, n387, n388, n389, n390, n391, n392,
 n393, n394, n395, n396, n397, n398, n399, n400,
 n401, n402, n403, n404, n405, n406, n407, n408,
 n409, n410, n411, n412, n413, n414, n415, n416,
 n417, n418, n419, n420, n421, n422, n423, n424,
 n425, n426, n427, n428, n429, n430, n431, n432,
 n433, n434, n435, n436, n437, n438, n439, n440,
 n441, n443, n444, n445, n446, n447, n448, n449,
 n450, n451, n452, n453, n454, n455, n456, n457,
 n458, n459, n460, n461, n462, n463, n464, n465,
 n466, n467, n468, n469, n470, n471, n472, n473,
 n474, n475, n476, n477, n478, n479, n480, n481,
 n482, n483, n484, n485, n486, n487, n488, n489,
 n490, n491, n492, n493, n494, n495, n496, n497,
 n498, n499, n500, n501, n502, n503, n504, n505,
 n506, n507, n508, n509, n510, n511, n512, n513,
 n514, n515, n516, n517, n518, n519, n520, n521,
 n522, n523, n524, n525, n526, n527, n528, n529,
 n530, n531, n532, n533, n534, n535, n536, n537,
 n538, n539, n540, n541, n542, n543, n544, n545,
 n546, n547, n548, n549, n550, n551, n552, n553,
 n554, n555, n556, n557, n558, n559, n560, n561,
 n562, n563, n564, n565, n566, n567, n568, n569,
 n570, n571, n572, n573, n574, n575, n576, n577,
 n578, n579, n580, n581, n582, n583, n584, n585,
 n586, n587, n588, n589, n590, n591, n592, n593,
 n594, n595, n596, n597, n598, n599, n600, n601,
 n602, n603, n604, n605, n606, n607, n609, n610,
 n611, n612, n613, n614, n615, n616, n617, n618,
 n619, n620, n621, n622, n623, n624, n625, n626,
 n627, n628, n629, n630, n631, n632, n633, n634,
 n635, n636, n637, n638, n639, n640, n641, n642,
 n643, n644, n645, n646, n647, n648, n649, n650,
 n651, n652, n653, n654, n655, n656, n657, n658,
 n659, n660, n661, n662, n663, n664, n665, n666,
 n667, n668, n669, n670, n671, n672, n673, n674,
 n675, n676, n677, n678, n679, n680, n681, n682,
 n683, n684, n685, n686, n687, n688, n689, n690,
 n691, n692, n693, n694, n695, n696, n697, n698,
 n699, n700, n701, n702, n703, n704, n705, n706,
 n707, n708, n709, n710, n711, n712, n713, n714,
 n715, n716, n717, n718, n719, n720, n721, n722,
 n723, n724, n725, n726, n727, n728, n729, n730,
 n731, n732, n733, n734, n735, n736, n737, n738,
 n739, n740, n741, n742, n743, n744, n745, n746,
 n747, n748, n749, n750, n751, n752, n753, n754,
 n755, n756, n757, n758, n759, n760, n761, n762,
 n763, n764, n765, n766, n767, n768, n769, n770,
 n771, n772, n773, n774, n775, n776, n777, n778,
 n779, n780, n781, n782, n783, n784, n785, n786,
 n787, n788, n789, n790, n791, n792, n793, n794,
 n795, n796, n797, n798, n799, n800, n801, n802,
 n803, n804, n805, n806, n807, n808, n809, n810,
 n811, n812, n813, n814, n815, n816, n817, n818,
 n819, n820, n821, n822, n823, n824, n825, n826,
 n827, n828, n829, n830, n831, n832, n833, n834,
 n835, n836, n837, n838, n839, n840, n841, n842,
 n843, n844, n845, n846, n847, n848, n849, n850,
 n851, n852, n853, n854, n855, n856, n857, n858,
 n859, n860, n861, n862, n863, n864, n865, n866,
 n867, n868, n869, n870, n871, n872, n873, n874,
 n875, n876, n877, n878, n879, n880, n881, n882,
 n883, n884, n885, n886, n887, n888, n889, n890,
 n891, n892, n893, n894, n895, n896, n897, n898,
 n899, n900, n901, n902, n903, n904, n905, n906,
 n907, n908, n909, n910, n911, n912, n913, n914,
 n915, n916, n917, n918, n919, n920, n921, n922,
 n923, n924, n925, n926, n927, n928, n929, n930,
 n931, n932, n933, n934, n935, n936, n937, n938,
 n939, n940, n941, n942, n943, n944, n945, n946,
 n947, n948, n949, n950, n951, n952, n953, n954,
 n955, n956, n957, n958, n959, n960, n961, n962,
 n963, n964, n965, n966, n967, n968, n969, n970,
 n971, n972, n973, n974, n975, n976, n977, n978,
 n979, n980, n981, n982, n983, n984, n985, n986,
 n987, n988, n989, n990, n991, n992, n993, n994,
 n995, n996, n997, n998, n999, n1000, n1001, n1002,
 n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
 n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
 n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
 n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
 n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
 n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
 n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
 n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
 n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
 n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
 n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
 n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
 n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
 n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
 n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
 n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
 n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
 n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
 n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
 n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
 n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
 n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
 n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
 n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
 n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
 n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
 n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
 n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
 n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
 n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
 n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
 n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
 n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
 n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
 n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
 n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
 n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
 n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
 n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
 n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
 n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
 n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
 n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
 n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
 n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
 n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
 n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
 n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
 n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
 n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
 n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
 n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
 n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
 n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
 n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
 n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
 n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
 n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
 n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
 n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
 n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
 n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
 n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
 n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
 n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
 n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
 n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
 n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
 n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
 n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
 n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
 n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
 n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
 n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
 n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
 n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
 n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
 n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
 n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
 n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
 n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
 n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
 n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
 n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
 n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
 n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
 n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
 n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
 n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
 n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
 n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
 n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
 n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
 n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
 n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
 n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
 n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
 n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
 n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
 n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
 n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
 n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
 n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
 n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
 n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
 n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
 n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
 n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
 n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
 n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
 n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
 n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
 n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
 n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
 n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
 n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
 n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
 n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946,
 n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
 n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
 n1963, n1964, n1966, n1967, n1969, n1975, n1977, n1978,
 n1979, n1980, n1981, n1982, n1983, n1984, n1986, n1991,
 n1993, n2000, n2004, n2008, n2009, n2010, n2011, n2012,
 n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
 n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028;

not  g0 (n136, n11);
not  g1 (n41, n11);
buf  g2 (n60, n21);
buf  g3 (n96, n7);
not  g4 (n126, n18);
buf  g5 (n44, n7);
buf  g6 (n56, n10);
buf  g7 (n50, n26);
not  g8 (n90, n2);
buf  g9 (n62, n27);
buf  g10 (n103, n10);
not  g11 (n127, n23);
buf  g12 (n77, n4);
not  g13 (n34, n5);
buf  g14 (n63, n8);
not  g15 (n109, n20);
not  g16 (n84, n15);
not  g17 (n137, n13);
buf  g18 (n100, n2);
not  g19 (n133, n22);
not  g20 (n87, n1);
buf  g21 (n33, n21);
not  g22 (n42, n17);
not  g23 (n55, n5);
not  g24 (n97, n25);
buf  g25 (n92, n5);
not  g26 (n106, n9);
not  g27 (n65, n6);
not  g28 (n125, n21);
buf  g29 (n83, n14);
not  g30 (n118, n14);
not  g31 (n135, n2);
buf  g32 (n52, n16);
not  g33 (n112, n26);
buf  g34 (n49, n18);
buf  g35 (n115, n24);
buf  g36 (n73, n9);
buf  g37 (n101, n15);
not  g38 (n57, n6);
not  g39 (n58, n11);
buf  g40 (n107, n5);
buf  g41 (n99, n4);
not  g42 (n70, n12);
not  g43 (n139, n10);
buf  g44 (n82, n1);
not  g45 (n74, n1);
not  g46 (n134, n20);
not  g47 (n132, n7);
not  g48 (n105, n7);
buf  g49 (n102, n16);
buf  g50 (n93, n22);
buf  g51 (n123, n8);
not  g52 (n43, n6);
not  g53 (n98, n27);
buf  g54 (n37, n6);
not  g55 (n48, n24);
buf  g56 (n67, n3);
not  g57 (n45, n16);
buf  g58 (n69, n21);
not  g59 (n85, n4);
buf  g60 (n116, n8);
buf  g61 (n54, n16);
not  g62 (n95, n20);
buf  g63 (n71, n4);
not  g64 (n68, n12);
buf  g65 (n38, n24);
not  g66 (n72, n26);
not  g67 (n88, n10);
buf  g68 (n120, n15);
buf  g69 (n113, n23);
buf  g70 (n75, n13);
buf  g71 (n47, n23);
not  g72 (n91, n27);
buf  g73 (n130, n25);
not  g74 (n138, n1);
not  g75 (n53, n19);
not  g76 (n128, n9);
buf  g77 (n104, n19);
buf  g78 (n80, n13);
not  g79 (n124, n9);
not  g80 (n51, n3);
not  g81 (n89, n22);
not  g82 (n61, n27);
buf  g83 (n121, n13);
buf  g84 (n122, n17);
not  g85 (n40, n14);
not  g86 (n108, n2);
not  g87 (n36, n18);
not  g88 (n114, n11);
not  g89 (n117, n24);
not  g90 (n94, n15);
buf  g91 (n64, n17);
buf  g92 (n111, n17);
buf  g93 (n76, n25);
buf  g94 (n140, n26);
buf  g95 (n129, n12);
buf  g96 (n46, n19);
buf  g97 (n66, n8);
buf  g98 (n131, n18);
buf  g99 (n86, n23);
buf  g100 (n79, n25);
buf  g101 (n78, n3);
buf  g102 (n59, n19);
not  g103 (n39, n20);
not  g104 (n81, n22);
not  g105 (n35, n12);
buf  g106 (n110, n14);
not  g107 (n119, n3);
not  g108 (n177, n87);
xnor g109 (n265, n56, n77);
nor  g110 (n148, n85, n98);
xnor g111 (n253, n45, n88);
and  g112 (n255, n67, n92);
nor  g113 (n164, n37, n64);
nor  g114 (n162, n69, n76);
nand g115 (n232, n65, n40);
nand g116 (n145, n96, n33);
nor  g117 (n243, n86, n73);
xnor g118 (n240, n46, n82);
and  g119 (n270, n78, n88);
nand g120 (n226, n71, n65);
or   g121 (n166, n61, n48);
or   g122 (n173, n79, n47);
and  g123 (n189, n53, n56);
nor  g124 (n249, n62, n64);
xor  g125 (n181, n78, n83);
and  g126 (n225, n51, n71);
xor  g127 (n182, n49, n66);
nand g128 (n196, n56, n88);
xnor g129 (n242, n74, n76);
nor  g130 (n183, n46, n66);
xnor g131 (n223, n55, n89);
xor  g132 (n152, n79, n54);
or   g133 (n208, n48, n71);
xor  g134 (n143, n76, n36);
nor  g135 (n184, n36, n63);
nor  g136 (n150, n75, n50);
xor  g137 (n239, n34, n49);
xnor g138 (n199, n97, n88);
nand g139 (n154, n38, n75);
nor  g140 (n244, n63, n96);
xor  g141 (n172, n73, n74);
nor  g142 (n167, n77, n52);
nand g143 (n187, n43, n58);
xor  g144 (n161, n83, n57);
not  g145 (n227, n42);
or   g146 (n194, n54, n90);
nor  g147 (n262, n33, n81);
or   g148 (n157, n41, n37);
nor  g149 (n178, n85, n36);
and  g150 (n192, n38, n87);
xor  g151 (n160, n84, n92);
or   g152 (n212, n90, n91);
xor  g153 (n169, n71, n79);
and  g154 (n203, n82, n93);
xnor g155 (n258, n64, n97);
xor  g156 (n228, n68, n69);
nor  g157 (n256, n36, n69);
or   g158 (n142, n50, n42);
nor  g159 (n207, n39, n83);
xnor g160 (n146, n66, n51);
xnor g161 (n190, n39, n38);
nand g162 (n245, n84, n87);
or   g163 (n191, n61, n59);
and  g164 (n209, n45, n58);
nand g165 (n264, n34, n54);
and  g166 (n229, n34, n40);
and  g167 (n246, n87, n67);
or   g168 (n260, n58, n89);
nor  g169 (n168, n75, n44);
xnor g170 (n188, n76, n62);
xnor g171 (n214, n44, n56);
and  g172 (n176, n93, n86);
xor  g173 (n269, n59, n81);
or   g174 (n231, n50, n73);
nand g175 (n271, n94, n80);
or   g176 (n211, n62, n83);
xor  g177 (n195, n61, n72);
and  g178 (n216, n47, n99);
nand g179 (n156, n33, n94);
and  g180 (n175, n89, n93);
nor  g181 (n210, n77, n52);
nor  g182 (n248, n90, n60);
or   g183 (n213, n79, n35);
xnor g184 (n247, n53, n69);
xor  g185 (n254, n91, n66);
xnor g186 (n147, n78, n94);
nor  g187 (n219, n95, n55);
nand g188 (n218, n43, n60);
and  g189 (n206, n98, n93);
and  g190 (n221, n98, n99);
nand g191 (n149, n47, n40);
xor  g192 (n220, n68, n70);
nor  g193 (n180, n57, n62);
xor  g194 (n268, n57, n85);
nor  g195 (n165, n41, n44);
nor  g196 (n222, n92, n53);
and  g197 (n174, n80, n84);
nand g198 (n163, n70, n94);
xor  g199 (n198, n74, n70);
or   g200 (n272, n33, n85);
buf  g201 (n201, n48);
nor  g202 (n235, n41, n73);
and  g203 (n186, n96, n44);
or   g204 (n200, n49, n52);
xor  g205 (n202, n60, n43);
xor  g206 (n273, n49, n86);
nand g207 (n153, n96, n84);
xnor g208 (n155, n52, n78);
nand g209 (n144, n82, n45);
xnor g210 (n170, n46, n99);
or   g211 (n251, n42, n46);
and  g212 (n250, n70, n39);
and  g213 (n233, n58, n95);
and  g214 (n158, n41, n54);
nand g215 (n236, n60, n61);
xnor g216 (n237, n51, n91);
nand g217 (n193, n53, n40);
and  g218 (n257, n90, n38);
nor  g219 (n205, n35, n72);
and  g220 (n261, n67, n43);
nor  g221 (n234, n75, n67);
xor  g222 (n171, n50, n97);
xor  g223 (n151, n65, n89);
xor  g224 (n215, n37, n63);
nand g225 (n230, n97, n74);
xor  g226 (n266, n64, n72);
nand g227 (n259, n65, n95);
and  g228 (n224, n59, n47);
and  g229 (n204, n35, n57);
xor  g230 (n252, n37, n86);
xor  g231 (n141, n81, n39);
nor  g232 (n197, n59, n55);
xnor g233 (n238, n80, n55);
xor  g234 (n274, n98, n63);
nand g235 (n263, n45, n72);
and  g236 (n241, n34, n68);
or   g237 (n267, n91, n35);
xnor g238 (n217, n51, n68);
nor  g239 (n179, n95, n92);
xor  g240 (n159, n82, n80);
xor  g241 (n185, n81, n77);
nand g242 (n313, n159, n238, n205, n202);
xor  g243 (n293, n192, n230, n213, n236);
xor  g244 (n346, n170, n193, n167, n228);
or   g245 (n344, n223, n190, n157, n209);
and  g246 (n364, n240, n147, n219, n186);
xor  g247 (n341, n207, n228, n143, n179);
nor  g248 (n279, n177, n231, n199, n232);
or   g249 (n310, n144, n194, n200, n211);
or   g250 (n321, n236, n216, n218, n197);
or   g251 (n315, n196, n146, n177, n167);
nor  g252 (n317, n181, n143, n211, n148);
xor  g253 (n337, n208, n196, n188);
or   g254 (n322, n156, n179, n154, n149);
xor  g255 (n372, n238, n190, n168, n182);
xnor g256 (n365, n215, n205, n145, n159);
or   g257 (n289, n161, n228, n215, n206);
nor  g258 (n299, n163, n156, n180, n220);
nand g259 (n353, n189, n223, n163, n177);
or   g260 (n287, n218, n157, n195, n172);
nor  g261 (n357, n233, n147, n229);
xnor g262 (n366, n235, n158, n191, n148);
and  g263 (n284, n179, n222, n217, n201);
and  g264 (n338, n182, n185, n149, n169);
xnor g265 (n331, n222, n174, n176, n154);
nor  g266 (n318, n189, n143, n192, n157);
nand g267 (n300, n155, n154, n229, n193);
and  g268 (n285, n192, n221, n218, n198);
xor  g269 (n327, n210, n190, n143, n158);
nor  g270 (n294, n155, n182, n153, n187);
or   g271 (n342, n164, n200, n172, n226);
nor  g272 (n340, n181, n183, n175, n194);
nor  g273 (n323, n226, n192, n155, n141);
or   g274 (n339, n175, n226, n239, n223);
nor  g275 (n286, n213, n164, n167, n203);
xor  g276 (n343, n229, n219, n184, n211);
xor  g277 (n311, n180, n225, n202);
and  g278 (n332, n174, n205, n142, n156);
nor  g279 (n280, n145, n232, n151, n236);
and  g280 (n349, n212, n216, n178, n224);
and  g281 (n356, n209, n153, n180, n181);
nor  g282 (n329, n223, n239, n152, n166);
xor  g283 (n374, n186, n239, n204, n146);
nand g284 (n324, n148, n235, n188, n187);
and  g285 (n359, n191, n217, n238, n162);
nor  g286 (n297, n206, n165, n184, n178);
xnor g287 (n291, n215, n176, n166, n237);
or   g288 (n308, n216, n198, n230, n141);
or   g289 (n304, n197, n177, n182, n204);
nand g290 (n369, n199, n199, n204, n184);
xor  g291 (n363, n153, n230, n197, n195);
nand g292 (n358, n201, n175, n199, n168);
xnor g293 (n345, n221, n147, n237);
nand g294 (n367, n174, n186, n170, n222);
nand g295 (n305, n194, n201, n161, n240);
nand g296 (n352, n152, n181, n206, n217);
or   g297 (n334, n166, n171, n205, n173);
xnor g298 (n309, n188, n220, n233, n187);
xnor g299 (n373, n172, n190, n212, n162);
nor  g300 (n288, n234, n148, n217, n150);
or   g301 (n326, n214, n169, n183, n222);
xor  g302 (n348, n164, n237, n240, n226);
and  g303 (n307, n227, n220, n176, n150);
nand g304 (n303, n145, n209, n159, n219);
or   g305 (n278, n146, n147, n200, n171);
xor  g306 (n354, n203, n152, n227, n239);
xnor g307 (n330, n236, n175, n178, n141);
nor  g308 (n290, n146, n227, n185, n233);
nor  g309 (n316, n171, n200, n213, n141);
or   g310 (n301, n232, n184, n151, n193);
and  g311 (n360, n159, n227, n163, n142);
or   g312 (n368, n154, n228, n183, n173);
nand g313 (n296, n149, n225, n238, n233);
nand g314 (n371, n144, n165, n151, n179);
nand g315 (n319, n196, n162, n203, n167);
or   g316 (n347, n224, n170, n153, n160);
nor  g317 (n314, n161, n172, n224, n203);
xor  g318 (n275, n221, n234, n214, n163);
and  g319 (n320, n170, n210, n149, n202);
and  g320 (n282, n150, n144, n186, n232);
xor  g321 (n350, n193, n173, n231, n216);
or   g322 (n298, n191, n207, n208, n152);
or   g323 (n283, n151, n157, n207, n162);
nand g324 (n336, n158, n234, n220, n142);
nand g325 (n295, n144, n218, n178, n188);
nor  g326 (n325, n161, n197, n195, n169);
xnor g327 (n370, n173, n231, n198, n183);
xnor g328 (n302, n180, n168, n145, n165);
and  g329 (n333, n165, n160, n158, n221);
nor  g330 (n281, n240, n219, n214, n230);
nand g331 (n351, n212, n164, n198, n171);
xnor g332 (n362, n209, n195, n231, n185);
xnor g333 (n328, n187, n191, n160, n210);
nand g334 (n292, n189, n208, n234, n210);
nor  g335 (n276, n169, n225, n224, n185);
nor  g336 (n312, n166, n215, n156, n204);
xnor g337 (n355, n189, n235, n211, n225);
xnor g338 (n277, n174, n150, n176, n201);
xor  g339 (n361, n214, n208, n207, n160);
or   g340 (n335, n168, n235, n142, n212);
nor  g341 (n306, n213, n155, n194, n206);
not  g342 (n380, n276);
buf  g343 (n376, n284);
buf  g344 (n377, n299);
buf  g345 (n384, n281);
and  g346 (n382, n278, n279, n297, n292);
and  g347 (n381, n301, n298, n275, n291);
and  g348 (n378, n288, n283, n282, n294);
xnor g349 (n379, n300, n286, n287, n293);
nor  g350 (n383, n289, n302, n277, n295);
nand g351 (n375, n296, n280, n285, n290);
buf  g352 (n405, n250);
not  g353 (n391, n257);
not  g354 (n417, n259);
buf  g355 (n420, n375);
not  g356 (n401, n250);
buf  g357 (n396, n377);
nand g358 (n397, n249, n377);
xor  g359 (n399, n257, n381, n376, n244);
and  g360 (n412, n258, n379, n242, n249);
and  g361 (n407, n244, n251, n250, n247);
nor  g362 (n411, n381, n376, n379, n242);
and  g363 (n385, n260, n378, n382);
xor  g364 (n394, n241, n259, n246, n381);
and  g365 (n421, n380, n303, n261, n262);
xor  g366 (n386, n378, n256, n377, n247);
xor  g367 (n390, n255, n257, n243, n260);
and  g368 (n388, n245, n246, n262, n253);
xor  g369 (n415, n383, n258, n248, n261);
or   g370 (n409, n242, n382, n380, n252);
nand g371 (n403, n251, n246, n253, n254);
nand g372 (n406, n246, n376, n241, n253);
or   g373 (n393, n252, n247, n251, n250);
nand g374 (n400, n241, n260, n245, n379);
nand g375 (n402, n256, n382, n263, n242);
and  g376 (n416, n244, n381, n259, n258);
xor  g377 (n410, n255, n375, n263, n380);
and  g378 (n389, n255, n383, n254, n244);
nor  g379 (n418, n245, n262, n248, n383);
xor  g380 (n413, n243, n254, n251, n259);
and  g381 (n387, n249, n377, n261, n376);
and  g382 (n395, n249, n241, n384, n261);
and  g383 (n414, n243, n254, n256, n248);
nand g384 (n392, n247, n252, n384);
xnor g385 (n419, n380, n383, n260, n248);
xor  g386 (n398, n243, n257, n245, n258);
nand g387 (n408, n375, n253, n256, n379);
xnor g388 (n404, n378, n382, n262, n255);
nor  g389 (n424, n385, n304);
or   g390 (n423, n306, n310, n309, n385);
xor  g391 (n422, n308, n305, n307, n385);
xnor g392 (n426, n266, n265);
or   g393 (n427, n263, n266, n423, n264);
nor  g394 (n425, n422, n266, n423);
nand g395 (n429, n264, n264, n266, n265);
and  g396 (n428, n422, n263, n264, n267);
nand g397 (n436, n333, n320, n317, n313);
nor  g398 (n432, n315, n426, n334, n312);
and  g399 (n430, n325, n332, n425, n427);
and  g400 (n438, n330, n328, n324, n429);
xor  g401 (n437, n340, n327, n429, n336);
or   g402 (n431, n329, n321, n428, n314);
or   g403 (n434, n318, n323, n339, n426);
or   g404 (n439, n322, n428, n425, n335);
xor  g405 (n435, n311, n338, n319, n316);
xnor g406 (n433, n331, n326, n337, n427);
buf  g407 (n440, n432);
buf  g408 (n442, n342);
nor  g409 (n443, n432, n341);
nand g410 (n441, n431, n430);
buf  g411 (n444, n442);
not  g412 (n446, n441);
not  g413 (n445, n443);
nand g414 (n449, n357, n424, n446, n351);
nand g415 (n448, n343, n353, n444);
and  g416 (n457, n352, n363, n346, n362);
nand g417 (n454, n358, n344, n445);
nor  g418 (n452, n362, n355, n358, n444);
xor  g419 (n451, n364, n348, n423, n359);
or   g420 (n450, n357, n356, n424, n446);
xor  g421 (n453, n424, n446, n444, n359);
nor  g422 (n447, n345, n361, n360, n354);
xor  g423 (n455, n347, n363, n445);
nor  g424 (n456, n360, n349, n350, n361);
not  g425 (n464, n451);
not  g426 (n493, n405);
buf  g427 (n478, n456);
buf  g428 (n475, n454);
buf  g429 (n486, n393);
buf  g430 (n487, n397);
not  g431 (n470, n455);
not  g432 (n465, n388);
buf  g433 (n483, n403);
not  g434 (n491, n396);
buf  g435 (n490, n387);
buf  g436 (n474, n390);
buf  g437 (n480, n392);
not  g438 (n462, n399);
not  g439 (n481, n394);
nor  g440 (n479, n451, n447, n403);
nor  g441 (n488, n28, n455, n389, n450);
and  g442 (n468, n395, n405, n449, n404);
and  g443 (n477, n448, n386, n388, n398);
xor  g444 (n469, n388, n457, n402, n404);
or   g445 (n458, n393, n450, n400, n399);
xnor g446 (n461, n386, n454, n389, n447);
or   g447 (n498, n393, n398, n449);
xor  g448 (n459, n453, n401, n393);
xnor g449 (n473, n390, n394, n397, n364);
nand g450 (n495, n391, n449, n453, n387);
or   g451 (n484, n455, n454, n448, n399);
xor  g452 (n471, n395, n396, n385, n392);
xor  g453 (n492, n391, n450, n401, n400);
xor  g454 (n501, n405, n387, n452, n400);
nand g455 (n466, n451, n389, n391, n404);
nand g456 (n476, n386, n395, n448, n405);
and  g457 (n499, n402, n394, n457, n390);
and  g458 (n463, n396, n449, n447, n451);
nor  g459 (n500, n450, n452, n447, n397);
and  g460 (n494, n457, n454, n452, n386);
xor  g461 (n496, n455, n395, n392, n396);
nand g462 (n472, n390, n404, n401, n456);
and  g463 (n482, n388, n448, n365, n402);
xor  g464 (n497, n453, n457, n394, n392);
and  g465 (n489, n453, n456, n403, n406);
or   g466 (n460, n389, n397, n400, n398);
nor  g467 (n485, n456, n403, n402, n399);
xor  g468 (n467, n387, n406, n452, n391);
nor  g469 (n510, n110, n134, n136, n468);
xor  g470 (n559, n476, n136, n488, n114);
xor  g471 (n576, n467, n494, n29, n114);
nand g472 (n505, n469, n463, n135, n484);
xor  g473 (n504, n468, n471, n478, n29);
and  g474 (n519, n130, n129, n466, n125);
nand g475 (n507, n100, n106, n433, n458);
nand g476 (n545, n478, n484, n135, n463);
nand g477 (n551, n471, n115, n113, n111);
xor  g478 (n506, n474, n112, n482, n119);
xor  g479 (n564, n131, n494, n406, n462);
and  g480 (n555, n115, n487, n486, n479);
and  g481 (n521, n458, n111, n117, n480);
or   g482 (n547, n491, n494, n485, n464);
xor  g483 (n580, n439, n474, n461, n477);
nand g484 (n557, n475, n466, n467, n458);
xnor g485 (n556, n116, n108, n480, n106);
nor  g486 (n530, n473, n106, n29, n483);
nor  g487 (n562, n129, n471, n112, n138);
nand g488 (n546, n437, n461, n104, n468);
xnor g489 (n579, n122, n109, n127, n459);
or   g490 (n541, n468, n102, n116, n495);
xnor g491 (n558, n128, n459, n475, n113);
xnor g492 (n554, n137, n129, n133, n484);
nor  g493 (n586, n460, n129, n486, n483);
nor  g494 (n566, n471, n109, n478, n493);
or   g495 (n509, n472, n481, n114, n107);
or   g496 (n532, n459, n488, n120, n110);
xnor g497 (n560, n492, n461, n434, n466);
nand g498 (n582, n117, n28, n496, n121);
and  g499 (n526, n487, n100, n490, n460);
xnor g500 (n525, n109, n490, n120, n123);
and  g501 (n552, n105, n137, n117, n477);
and  g502 (n553, n130, n103, n436, n115);
or   g503 (n534, n492, n118, n100, n137);
nor  g504 (n581, n131, n477, n101, n118);
xnor g505 (n529, n488, n134, n485, n132);
or   g506 (n512, n122, n127, n111, n104);
nor  g507 (n536, n109, n433, n118, n482);
nand g508 (n539, n102, n436, n493, n28);
or   g509 (n520, n465, n496, n481, n108);
xor  g510 (n522, n103, n133, n134, n102);
or   g511 (n550, n118, n267, n497, n481);
or   g512 (n517, n474, n487, n29, n113);
nand g513 (n561, n113, n470, n486, n462);
or   g514 (n538, n136, n492, n481, n127);
nor  g515 (n537, n496, n99, n115, n467);
nand g516 (n578, n110, n476, n121, n131);
nand g517 (n577, n121, n138, n124, n491);
xnor g518 (n514, n125, n124, n470, n112);
and  g519 (n502, n464, n102, n136, n437);
nand g520 (n575, n458, n123, n460, n484);
xor  g521 (n573, n122, n133, n130, n131);
xnor g522 (n503, n438, n128, n488, n473);
or   g523 (n568, n119, n489, n108, n101);
xor  g524 (n535, n107, n493, n494, n476);
xnor g525 (n548, n465, n459, n474, n134);
or   g526 (n565, n110, n135, n107, n130);
or   g527 (n524, n485, n103, n132, n472);
nor  g528 (n515, n126, n487, n467, n116);
nand g529 (n569, n492, n475, n108, n28);
nor  g530 (n584, n497, n101, n434, n138);
xnor g531 (n513, n124, n126, n121, n105);
or   g532 (n585, n125, n101, n462, n119);
and  g533 (n527, n132, n495, n469, n105);
nor  g534 (n528, n482, n463, n133);
nor  g535 (n511, n475, n495, n490, n482);
xor  g536 (n540, n483, n485, n438, n480);
or   g537 (n571, n479, n496, n128, n497);
or   g538 (n533, n476, n103, n267, n132);
nor  g539 (n549, n478, n117, n135, n479);
and  g540 (n508, n490, n105, n472, n435);
and  g541 (n544, n465, n486, n464, n469);
or   g542 (n570, n120, n137, n473, n107);
or   g543 (n523, n470, n483, n104, n480);
xnor g544 (n531, n489, n104, n120, n126);
or   g545 (n574, n124, n493, n464, n491);
nand g546 (n567, n138, n128, n473, n106);
xor  g547 (n518, n125, n462, n116, n489);
or   g548 (n516, n114, n477, n491, n495);
xor  g549 (n583, n470, n123, n466, n461);
nor  g550 (n563, n489, n472, n139, n112);
or   g551 (n572, n123, n435, n479, n122);
and  g552 (n543, n465, n100, n119, n460);
and  g553 (n542, n111, n469, n126, n127);
nor  g554 (n588, n543, n513, n517, n531);
or   g555 (n598, n512, n504, n523, n518);
xnor g556 (n592, n529, n546, n560, n526);
xor  g557 (n590, n539, n541, n552, n506);
or   g558 (n599, n561, n514, n522, n551);
nor  g559 (n591, n532, n559, n511, n528);
xor  g560 (n596, n554, n563, n515, n562);
xnor g561 (n594, n547, n530, n525, n544);
nand g562 (n593, n535, n527, n508, n533);
or   g563 (n602, n545, n542, n502, n555);
nor  g564 (n589, n548, n537, n516, n505);
and  g565 (n597, n507, n553, n524, n556);
nor  g566 (n595, n519, n563, n520, n509);
nand g567 (n601, n521, n550, n503, n557);
nor  g568 (n600, n536, n562, n540, n538);
xor  g569 (n587, n534, n549, n558, n510);
buf  g570 (n603, n365);
nand g571 (n604, n588, n366, n587);
not  g572 (n612, n603);
not  g573 (n608, n603);
not  g574 (n606, n604);
not  g575 (n605, n604);
buf  g576 (n611, n604);
buf  g577 (n610, n603);
buf  g578 (n607, n603);
buf  g579 (n609, n604);
nand g580 (n615, n421, n269, n608, n416);
xnor g581 (n625, n414, n420, n411, n606);
xnor g582 (n639, n420, n408, n610);
xnor g583 (n634, n419, n367, n269, n412);
xnor g584 (n635, n407, n369, n408, n411);
xor  g585 (n627, n499, n418, n610, n417);
and  g586 (n633, n605, n417, n268, n612);
or   g587 (n613, n268, n499, n367, n605);
nor  g588 (n617, n608, n420, n419, n606);
xor  g589 (n640, n416, n416, n500, n608);
and  g590 (n614, n268, n497, n417, n418);
nand g591 (n643, n418, n414, n409, n498);
nand g592 (n631, n370, n407, n609);
nand g593 (n619, n368, n412, n419, n414);
xnor g594 (n618, n607, n415, n410, n421);
nand g595 (n616, n419, n501, n415, n412);
or   g596 (n620, n418, n499, n609, n611);
xnor g597 (n638, n498, n607, n408, n414);
nor  g598 (n623, n612, n268, n609, n611);
xor  g599 (n628, n501, n415, n366, n369);
xnor g600 (n621, n413, n612, n607);
xnor g601 (n637, n610, n409, n412, n370);
xnor g602 (n641, n267, n608, n413, n411);
and  g603 (n636, n415, n408, n416, n611);
xor  g604 (n642, n407, n612, n605, n413);
and  g605 (n630, n421, n407, n370, n410);
nand g606 (n626, n406, n499, n411, n417);
xor  g607 (n632, n368, n409, n606);
or   g608 (n622, n498, n410, n611, n500);
xnor g609 (n629, n413, n409, n410, n500);
nand g610 (n624, n498, n500, n370, n420);
nor  g611 (n644, n613, n564);
not  g612 (n647, n644);
buf  g613 (n648, n644);
buf  g614 (n645, n644);
not  g615 (n646, n644);
or   g616 (n663, n615, n575, n645, n646);
nand g617 (n660, n646, n568, n569, n570);
and  g618 (n650, n572, n421, n614, n621);
nor  g619 (n662, n576, n577, n565);
xnor g620 (n652, n567, n645, n566);
xor  g621 (n655, n647, n647, n580, n575);
and  g622 (n657, n571, n577, n569, n579);
or   g623 (n656, n566, n648, n573);
xnor g624 (n661, n579, n576, n574, n619);
or   g625 (n659, n648, n578, n567, n617);
xor  g626 (n658, n572, n573, n571, n646);
or   g627 (n653, n648, n647, n646, n581);
nand g628 (n651, n580, n574, n578, n620);
nand g629 (n649, n581, n647, n568, n564);
nor  g630 (n654, n618, n570, n645, n616);
buf  g631 (n664, n652);
buf  g632 (n680, n658);
not  g633 (n713, n661);
not  g634 (n671, n661);
buf  g635 (n685, n654);
buf  g636 (n673, n659);
buf  g637 (n710, n649);
buf  g638 (n706, n653);
buf  g639 (n702, n654);
not  g640 (n691, n651);
not  g641 (n701, n663);
not  g642 (n676, n660);
buf  g643 (n716, n649);
not  g644 (n720, n654);
not  g645 (n669, n663);
not  g646 (n718, n650);
buf  g647 (n674, n654);
not  g648 (n703, n652);
not  g649 (n717, n662);
not  g650 (n693, n657);
not  g651 (n712, n649);
not  g652 (n698, n657);
buf  g653 (n686, n655);
not  g654 (n665, n662);
buf  g655 (n677, n650);
not  g656 (n675, n651);
buf  g657 (n672, n656);
not  g658 (n687, n652);
buf  g659 (n709, n659);
not  g660 (n723, n663);
not  g661 (n684, n649);
buf  g662 (n722, n657);
buf  g663 (n695, n659);
buf  g664 (n721, n655);
buf  g665 (n705, n653);
buf  g666 (n689, n652);
not  g667 (n678, n651);
buf  g668 (n697, n653);
not  g669 (n683, n656);
buf  g670 (n719, n655);
not  g671 (n715, n662);
not  g672 (n699, n656);
not  g673 (n681, n653);
not  g674 (n696, n659);
buf  g675 (n714, n661);
not  g676 (n700, n660);
buf  g677 (n707, n660);
not  g678 (n690, n657);
not  g679 (n682, n663);
not  g680 (n668, n660);
buf  g681 (n667, n658);
not  g682 (n666, n651);
not  g683 (n704, n658);
buf  g684 (n708, n650);
not  g685 (n694, n661);
buf  g686 (n670, n662);
not  g687 (n692, n655);
not  g688 (n688, n650);
buf  g689 (n711, n658);
not  g690 (n679, n656);
not  g691 (n724, n669);
buf  g692 (n786, n714);
not  g693 (n765, n698);
not  g694 (n919, n371);
buf  g695 (n735, n372);
not  g696 (n807, n373);
buf  g697 (n817, n682);
buf  g698 (n730, n715);
buf  g699 (n782, n702);
not  g700 (n859, n713);
buf  g701 (n790, n713);
not  g702 (n860, n710);
not  g703 (n749, n677);
buf  g704 (n737, n689);
buf  g705 (n917, n676);
not  g706 (n811, n670);
buf  g707 (n842, n708);
buf  g708 (n814, n673);
buf  g709 (n780, n703);
not  g710 (n747, n697);
buf  g711 (n758, n717);
not  g712 (n836, n678);
buf  g713 (n740, n691);
buf  g714 (n946, n634);
buf  g715 (n886, n696);
buf  g716 (n728, n723);
buf  g717 (n936, n677);
not  g718 (n875, n700);
not  g719 (n962, n675);
not  g720 (n913, n622);
not  g721 (n896, n636);
buf  g722 (n768, n720);
buf  g723 (n871, n667);
not  g724 (n772, n637);
not  g725 (n932, n687);
not  g726 (n947, n679);
not  g727 (n958, n699);
not  g728 (n922, n371);
not  g729 (n907, n679);
not  g730 (n845, n704);
not  g731 (n810, n680);
buf  g732 (n883, n698);
not  g733 (n915, n690);
buf  g734 (n877, n669);
not  g735 (n792, n688);
buf  g736 (n729, n665);
not  g737 (n736, n633);
buf  g738 (n783, n716);
not  g739 (n906, n676);
buf  g740 (n789, n686);
buf  g741 (n956, n721);
buf  g742 (n813, n684);
buf  g743 (n816, n693);
not  g744 (n881, n681);
not  g745 (n808, n624);
not  g746 (n750, n701);
not  g747 (n798, n637);
buf  g748 (n803, n712);
not  g749 (n943, n722);
buf  g750 (n853, n711);
buf  g751 (n929, n706);
buf  g752 (n855, n672);
not  g753 (n933, n688);
not  g754 (n854, n719);
not  g755 (n869, n711);
not  g756 (n914, n704);
buf  g757 (n822, n702);
buf  g758 (n754, n671);
buf  g759 (n741, n718);
not  g760 (n833, n628);
buf  g761 (n752, n707);
buf  g762 (n937, n694);
not  g763 (n820, n683);
buf  g764 (n941, n703);
not  g765 (n910, n722);
not  g766 (n818, n721);
buf  g767 (n872, n664);
buf  g768 (n797, n711);
not  g769 (n951, n686);
buf  g770 (n953, n684);
not  g771 (n903, n691);
buf  g772 (n880, n635);
buf  g773 (n864, n672);
buf  g774 (n934, n664);
not  g775 (n918, n706);
not  g776 (n945, n708);
not  g777 (n759, n632);
not  g778 (n827, n714);
buf  g779 (n891, n706);
buf  g780 (n867, n674);
not  g781 (n844, n668);
not  g782 (n828, n666);
buf  g783 (n756, n709);
buf  g784 (n738, n697);
buf  g785 (n760, n702);
buf  g786 (n847, n688);
not  g787 (n838, n667);
not  g788 (n916, n718);
not  g789 (n744, n680);
not  g790 (n905, n692);
not  g791 (n889, n627);
not  g792 (n858, n699);
buf  g793 (n831, n707);
buf  g794 (n777, n723);
not  g795 (n809, n690);
not  g796 (n748, n373);
buf  g797 (n893, n682);
buf  g798 (n892, n700);
buf  g799 (n961, n714);
buf  g800 (n897, n680);
buf  g801 (n921, n673);
not  g802 (n876, n715);
not  g803 (n767, n372);
not  g804 (n894, n636);
buf  g805 (n887, n669);
buf  g806 (n948, n684);
buf  g807 (n926, n701);
buf  g808 (n931, n692);
not  g809 (n805, n698);
buf  g810 (n726, n710);
not  g811 (n902, n701);
buf  g812 (n954, n678);
not  g813 (n804, n626);
not  g814 (n878, n674);
buf  g815 (n843, n694);
not  g816 (n930, n712);
buf  g817 (n739, n682);
not  g818 (n895, n670);
not  g819 (n944, n700);
buf  g820 (n850, n721);
buf  g821 (n799, n698);
not  g822 (n819, n677);
not  g823 (n841, n687);
not  g824 (n830, n692);
not  g825 (n821, n686);
not  g826 (n837, n722);
not  g827 (n960, n374);
not  g828 (n924, n712);
not  g829 (n778, n675);
buf  g830 (n899, n689);
not  g831 (n800, n715);
buf  g832 (n761, n677);
not  g833 (n794, n711);
not  g834 (n879, n693);
buf  g835 (n862, n681);
buf  g836 (n733, n669);
not  g837 (n755, n716);
not  g838 (n908, n674);
buf  g839 (n766, n694);
buf  g840 (n806, n634);
not  g841 (n776, n671);
not  g842 (n874, n635);
buf  g843 (n762, n371);
not  g844 (n928, n721);
buf  g845 (n882, n708);
buf  g846 (n955, n699);
buf  g847 (n939, n680);
not  g848 (n952, n630);
not  g849 (n863, n720);
buf  g850 (n787, n718);
not  g851 (n823, n670);
not  g852 (n753, n712);
buf  g853 (n791, n705);
buf  g854 (n846, n671);
not  g855 (n912, n690);
buf  g856 (n763, n665);
buf  g857 (n834, n695);
buf  g858 (n774, n701);
not  g859 (n873, n678);
buf  g860 (n795, n697);
buf  g861 (n757, n713);
not  g862 (n745, n679);
not  g863 (n771, n710);
buf  g864 (n963, n630);
not  g865 (n801, n716);
not  g866 (n802, n675);
buf  g867 (n890, n708);
buf  g868 (n796, n691);
buf  g869 (n911, n722);
buf  g870 (n851, n696);
not  g871 (n779, n694);
buf  g872 (n861, n676);
buf  g873 (n781, n705);
buf  g874 (n835, n696);
buf  g875 (n888, n695);
not  g876 (n942, n684);
not  g877 (n923, n666);
not  g878 (n925, n685);
not  g879 (n870, n668);
not  g880 (n865, n665);
buf  g881 (n839, n699);
buf  g882 (n812, n713);
buf  g883 (n950, n679);
buf  g884 (n909, n706);
buf  g885 (n824, n717);
buf  g886 (n770, n631);
not  g887 (n764, n720);
not  g888 (n725, n688);
buf  g889 (n920, n695);
not  g890 (n751, n704);
not  g891 (n832, n692);
xnor g892 (n784, n373, n717);
or   g893 (n826, n674, n683);
or   g894 (n927, n704, n668);
or   g895 (n938, n672, n664);
or   g896 (n940, n690, n629);
nor  g897 (n949, n683, n719);
and  g898 (n769, n681, n685);
or   g899 (n901, n723, n632);
and  g900 (n746, n689, n716);
xnor g901 (n904, n720, n717);
or   g902 (n885, n665, n685);
xnor g903 (n957, n709, n702);
xor  g904 (n900, n373, n686);
nand g905 (n793, n675, n718);
xor  g906 (n732, n714, n673);
nor  g907 (n731, n633, n667);
xnor g908 (n857, n664, n631);
nor  g909 (n856, n672, n673);
or   g910 (n785, n372, n371);
nand g911 (n734, n693, n697);
xnor g912 (n840, n623, n687);
nor  g913 (n849, n374, n696);
nor  g914 (n829, n671, n709);
xnor g915 (n788, n668, n705);
xor  g916 (n825, n707, n695);
xor  g917 (n959, n703, n666);
xor  g918 (n742, n723, n693);
and  g919 (n815, n687, n700);
nor  g920 (n775, n715, n676);
nor  g921 (n727, n710, n678);
xor  g922 (n852, n666, n682);
nor  g923 (n743, n689, n709);
xnor g924 (n884, n670, n691);
and  g925 (n935, n372, n374);
nand g926 (n866, n707, n705);
or   g927 (n773, n625, n683);
xnor g928 (n898, n703, n719);
nor  g929 (n848, n681, n685);
or   g930 (n868, n719, n667);
buf  g931 (n1172, n945);
not  g932 (n1014, n599);
buf  g933 (n1370, n935);
not  g934 (n1528, n272);
buf  g935 (n1614, n866);
not  g936 (n1436, n799);
not  g937 (n1737, n909);
not  g938 (n1306, n760);
not  g939 (n1325, n894);
buf  g940 (n1249, n725);
not  g941 (n1345, n742);
buf  g942 (n1221, n586);
not  g943 (n1755, n862);
not  g944 (n1711, n825);
buf  g945 (n1580, n767);
buf  g946 (n1578, n836);
not  g947 (n1212, n900);
buf  g948 (n1303, n876);
not  g949 (n1242, n934);
not  g950 (n1346, n952);
not  g951 (n1320, n865);
buf  g952 (n1655, n881);
not  g953 (n1584, n867);
buf  g954 (n1270, n844);
buf  g955 (n1289, n942);
buf  g956 (n1665, n585);
buf  g957 (n1656, n782);
not  g958 (n1409, n817);
buf  g959 (n991, n914);
buf  g960 (n1393, n945);
buf  g961 (n1496, n831);
buf  g962 (n1732, n956);
not  g963 (n1471, n733);
not  g964 (n1673, n955);
not  g965 (n1477, n947);
buf  g966 (n1473, n755);
not  g967 (n1426, n799);
buf  g968 (n1093, n851);
not  g969 (n1263, n935);
not  g970 (n1712, n779);
not  g971 (n1326, n926);
buf  g972 (n1161, n851);
not  g973 (n1213, n886);
buf  g974 (n1331, n912);
buf  g975 (n985, n733);
buf  g976 (n1039, n929);
not  g977 (n1020, n940);
not  g978 (n1079, n753);
buf  g979 (n1152, n271);
not  g980 (n1692, n879);
buf  g981 (n1485, n854);
buf  g982 (n1220, n821);
not  g983 (n1650, n642);
not  g984 (n1030, n734);
buf  g985 (n1032, n796);
not  g986 (n1160, n807);
not  g987 (n1304, n826);
buf  g988 (n1599, n798);
not  g989 (n1102, n852);
not  g990 (n1105, n802);
not  g991 (n1691, n816);
buf  g992 (n1222, n828);
buf  g993 (n1744, n913);
not  g994 (n1511, n740);
buf  g995 (n1365, n949);
buf  g996 (n1478, n923);
not  g997 (n1319, n870);
not  g998 (n1150, n927);
buf  g999 (n971, n273);
buf  g1000 (n1410, n953);
not  g1001 (n1038, n783);
buf  g1002 (n1635, n861);
not  g1003 (n1653, n750);
buf  g1004 (n1354, n962);
not  g1005 (n986, n830);
buf  g1006 (n1683, n867);
not  g1007 (n1463, n932);
buf  g1008 (n1620, n961);
buf  g1009 (n1164, n756);
buf  g1010 (n1315, n952);
not  g1011 (n1493, n902);
not  g1012 (n1081, n758);
buf  g1013 (n1028, n833);
buf  g1014 (n1279, n848);
buf  g1015 (n1548, n877);
buf  g1016 (n1392, n851);
not  g1017 (n1417, n943);
buf  g1018 (n1192, n859);
buf  g1019 (n1513, n838);
not  g1020 (n1062, n803);
not  g1021 (n1373, n811);
not  g1022 (n1391, n896);
buf  g1023 (n1372, n845);
not  g1024 (n1272, n910);
buf  g1025 (n1533, n779);
buf  g1026 (n1467, n865);
buf  g1027 (n1281, n950);
not  g1028 (n1660, n931);
not  g1029 (n1701, n894);
not  g1030 (n1215, n803);
buf  g1031 (n1292, n833);
buf  g1032 (n1540, n887);
buf  g1033 (n1512, n812);
buf  g1034 (n1084, n748);
not  g1035 (n1679, n943);
buf  g1036 (n1554, n822);
buf  g1037 (n1006, n945);
not  g1038 (n1336, n858);
buf  g1039 (n1262, n785);
not  g1040 (n1252, n951);
not  g1041 (n1122, n795);
buf  g1042 (n1752, n901);
not  g1043 (n1530, n889);
buf  g1044 (n1033, n843);
buf  g1045 (n1291, n793);
not  g1046 (n1264, n905);
buf  g1047 (n1223, n751);
buf  g1048 (n1570, n743);
buf  g1049 (n1139, n939);
not  g1050 (n1424, n897);
not  g1051 (n1474, n911);
not  g1052 (n1609, n883);
buf  g1053 (n1642, n838);
not  g1054 (n1008, n829);
buf  g1055 (n1562, n878);
not  g1056 (n1425, n807);
not  g1057 (n1438, n952);
buf  g1058 (n1082, n868);
buf  g1059 (n1112, n738);
buf  g1060 (n1608, n932);
buf  g1061 (n1526, n768);
not  g1062 (n994, n743);
not  g1063 (n1042, n791);
buf  g1064 (n1751, n884);
buf  g1065 (n1210, n745);
buf  g1066 (n1064, n954);
buf  g1067 (n1705, n951);
not  g1068 (n1052, n867);
not  g1069 (n1403, n934);
not  g1070 (n1428, n882);
buf  g1071 (n1353, n140);
buf  g1072 (n1416, n819);
not  g1073 (n1063, n881);
not  g1074 (n1509, n783);
buf  g1075 (n1647, n919);
buf  g1076 (n1707, n805);
not  g1077 (n1204, n895);
not  g1078 (n1253, n840);
buf  g1079 (n1747, n931);
not  g1080 (n1132, n769);
not  g1081 (n1120, n790);
not  g1082 (n1230, n863);
buf  g1083 (n1248, n901);
not  g1084 (n1680, n896);
not  g1085 (n1696, n643);
buf  g1086 (n1490, n640);
buf  g1087 (n1114, n727);
not  g1088 (n1521, n787);
buf  g1089 (n1098, n958);
not  g1090 (n1661, n724);
buf  g1091 (n1442, n838);
not  g1092 (n1549, n767);
not  g1093 (n1390, n750);
not  g1094 (n1009, n906);
not  g1095 (n1698, n953);
not  g1096 (n1461, n740);
buf  g1097 (n977, n939);
not  g1098 (n1415, n847);
buf  g1099 (n1268, n934);
buf  g1100 (n1374, n930);
not  g1101 (n1092, n941);
not  g1102 (n1422, n873);
buf  g1103 (n1061, n950);
buf  g1104 (n1563, n831);
not  g1105 (n1706, n835);
buf  g1106 (n1177, n925);
not  g1107 (n1468, n808);
buf  g1108 (n1368, n953);
not  g1109 (n979, n897);
buf  g1110 (n1049, n877);
not  g1111 (n1593, n741);
not  g1112 (n1498, n583);
not  g1113 (n1657, n775);
buf  g1114 (n1420, n591);
buf  g1115 (n1694, n601);
not  g1116 (n1500, n832);
not  g1117 (n1510, n830);
buf  g1118 (n1740, n857);
buf  g1119 (n1545, n871);
buf  g1120 (n1671, n905);
not  g1121 (n1196, n780);
not  g1122 (n1324, n878);
not  g1123 (n1189, n809);
buf  g1124 (n1056, n883);
buf  g1125 (n987, n778);
buf  g1126 (n1095, n777);
not  g1127 (n1273, n954);
not  g1128 (n1481, n790);
not  g1129 (n1700, n885);
buf  g1130 (n1458, n873);
buf  g1131 (n1257, n731);
not  g1132 (n1347, n734);
not  g1133 (n1560, n731);
not  g1134 (n1104, n842);
buf  g1135 (n1143, n886);
buf  g1136 (n1699, n762);
not  g1137 (n1723, n856);
not  g1138 (n1237, n871);
not  g1139 (n1310, n937);
buf  g1140 (n1089, n732);
buf  g1141 (n1394, n915);
buf  g1142 (n1004, n724);
buf  g1143 (n1218, n729);
buf  g1144 (n1234, n820);
buf  g1145 (n1758, n775);
buf  g1146 (n1452, n739);
not  g1147 (n1585, n913);
buf  g1148 (n992, n869);
buf  g1149 (n1497, n739);
buf  g1150 (n1254, n947);
buf  g1151 (n1492, n858);
not  g1152 (n1495, n841);
buf  g1153 (n1440, n749);
not  g1154 (n1746, n936);
buf  g1155 (n1016, n824);
not  g1156 (n1157, n726);
buf  g1157 (n1542, n844);
not  g1158 (n1506, n750);
not  g1159 (n964, n929);
not  g1160 (n1314, n736);
buf  g1161 (n1011, n756);
buf  g1162 (n1553, n765);
not  g1163 (n1516, n760);
buf  g1164 (n1618, n917);
buf  g1165 (n1276, n800);
buf  g1166 (n1571, n866);
buf  g1167 (n1551, n892);
not  g1168 (n1518, n139);
buf  g1169 (n1532, n735);
buf  g1170 (n1734, n856);
not  g1171 (n1280, n947);
buf  g1172 (n1074, n928);
not  g1173 (n1338, n835);
not  g1174 (n1141, n858);
not  g1175 (n1587, n813);
not  g1176 (n1058, n824);
buf  g1177 (n1077, n903);
not  g1178 (n1256, n753);
not  g1179 (n1484, n643);
not  g1180 (n1603, n729);
buf  g1181 (n1115, n847);
buf  g1182 (n1621, n942);
not  g1183 (n1126, n855);
buf  g1184 (n1231, n907);
not  g1185 (n1713, n845);
not  g1186 (n1148, n885);
not  g1187 (n1366, n752);
not  g1188 (n1352, n792);
buf  g1189 (n1630, n731);
not  g1190 (n1298, n846);
buf  g1191 (n1002, n904);
not  g1192 (n1654, n940);
buf  g1193 (n1010, n916);
buf  g1194 (n1146, n798);
not  g1195 (n1174, n954);
buf  g1196 (n1558, n823);
not  g1197 (n1173, n777);
not  g1198 (n1486, n870);
not  g1199 (n1000, n424);
not  g1200 (n1572, n903);
buf  g1201 (n1602, n853);
buf  g1202 (n1382, n735);
not  g1203 (n1536, n792);
buf  g1204 (n1672, n744);
buf  g1205 (n1674, n891);
buf  g1206 (n1638, n898);
buf  g1207 (n1437, n849);
buf  g1208 (n1019, n963);
buf  g1209 (n1730, n919);
not  g1210 (n1524, n934);
not  g1211 (n1592, n914);
buf  g1212 (n1271, n893);
not  g1213 (n1099, n594);
not  g1214 (n1295, n858);
buf  g1215 (n1411, n900);
buf  g1216 (n1034, n780);
buf  g1217 (n1517, n786);
buf  g1218 (n970, n845);
not  g1219 (n1287, n736);
buf  g1220 (n1127, n273);
not  g1221 (n1060, n796);
not  g1222 (n1153, n937);
not  g1223 (n1377, n772);
buf  g1224 (n1219, n589);
not  g1225 (n1693, n828);
buf  g1226 (n1110, n755);
buf  g1227 (n1607, n745);
buf  g1228 (n1329, n931);
not  g1229 (n1227, n879);
not  g1230 (n1434, n961);
not  g1231 (n1397, n139);
buf  g1232 (n1659, n918);
buf  g1233 (n1036, n795);
buf  g1234 (n1318, n923);
not  g1235 (n1119, n945);
not  g1236 (n1332, n829);
not  g1237 (n1266, n811);
buf  g1238 (n1194, n641);
buf  g1239 (n1728, n846);
buf  g1240 (n1349, n940);
not  g1241 (n1547, n790);
not  g1242 (n1670, n807);
not  g1243 (n1235, n802);
not  g1244 (n1616, n962);
buf  g1245 (n1522, n602);
buf  g1246 (n1296, n927);
not  g1247 (n990, n778);
not  g1248 (n1386, n747);
not  g1249 (n1447, n959);
not  g1250 (n1375, n787);
buf  g1251 (n982, n960);
not  g1252 (n1709, n776);
not  g1253 (n1007, n832);
buf  g1254 (n1456, n638);
not  g1255 (n1243, n776);
not  g1256 (n1251, n762);
not  g1257 (n1750, n833);
not  g1258 (n1001, n773);
buf  g1259 (n1406, n958);
buf  g1260 (n1383, n797);
not  g1261 (n1581, n595);
buf  g1262 (n1622, n784);
buf  g1263 (n1340, n840);
not  g1264 (n1688, n911);
buf  g1265 (n1037, n830);
buf  g1266 (n1527, n732);
not  g1267 (n1129, n749);
not  g1268 (n1446, n753);
not  g1269 (n1413, n746);
buf  g1270 (n1283, n868);
buf  g1271 (n1364, n899);
not  g1272 (n1610, n899);
buf  g1273 (n966, n960);
not  g1274 (n1297, n876);
buf  g1275 (n1736, n929);
buf  g1276 (n1258, n764);
buf  g1277 (n1667, n810);
not  g1278 (n1441, n903);
not  g1279 (n1399, n922);
not  g1280 (n1643, n763);
not  g1281 (n1379, n852);
not  g1282 (n1404, n792);
buf  g1283 (n1083, n759);
not  g1284 (n1057, n943);
buf  g1285 (n1429, n761);
not  g1286 (n1175, n766);
not  g1287 (n984, n773);
buf  g1288 (n1309, n582);
not  g1289 (n1151, n785);
not  g1290 (n1641, n772);
buf  g1291 (n1071, n790);
buf  g1292 (n1520, n724);
not  g1293 (n1344, n765);
not  g1294 (n1229, n907);
not  g1295 (n1106, n955);
buf  g1296 (n1305, n956);
not  g1297 (n1717, n837);
buf  g1298 (n1236, n746);
not  g1299 (n1544, n893);
not  g1300 (n1113, n874);
buf  g1301 (n1435, n776);
not  g1302 (n1538, n789);
not  g1303 (n976, n848);
buf  g1304 (n1380, n938);
not  g1305 (n1612, n834);
buf  g1306 (n1443, n813);
buf  g1307 (n1568, n919);
buf  g1308 (n1575, n908);
not  g1309 (n1290, n139);
not  g1310 (n1171, n814);
not  g1311 (n1387, n913);
not  g1312 (n1047, n842);
buf  g1313 (n1162, n850);
buf  g1314 (n1569, n786);
buf  g1315 (n1543, n951);
not  g1316 (n1697, n796);
not  g1317 (n1483, n946);
buf  g1318 (n1250, n942);
not  g1319 (n1480, n743);
buf  g1320 (n1418, n770);
not  g1321 (n1565, n770);
not  g1322 (n1275, n911);
not  g1323 (n1259, n946);
buf  g1324 (n1065, n804);
not  g1325 (n1648, n736);
not  g1326 (n1307, n828);
not  g1327 (n1515, n891);
buf  g1328 (n989, n593);
buf  g1329 (n1742, n887);
not  g1330 (n1464, n874);
buf  g1331 (n1244, n797);
buf  g1332 (n1163, n877);
buf  g1333 (n1133, n791);
not  g1334 (n1024, n794);
buf  g1335 (n1475, n949);
not  g1336 (n1588, n270);
not  g1337 (n1046, n787);
not  g1338 (n1555, n891);
not  g1339 (n1716, n825);
not  g1340 (n1094, n789);
buf  g1341 (n1371, n959);
buf  g1342 (n1460, n862);
buf  g1343 (n1333, n860);
buf  g1344 (n1206, n762);
not  g1345 (n1644, n839);
buf  g1346 (n1482, n961);
buf  g1347 (n1168, n855);
not  g1348 (n1466, n731);
not  g1349 (n1633, n764);
buf  g1350 (n1561, n820);
not  g1351 (n1239, n816);
not  g1352 (n1414, n446);
buf  g1353 (n1240, n823);
not  g1354 (n1187, n937);
buf  g1355 (n1664, n916);
not  g1356 (n1689, n944);
buf  g1357 (n1405, n937);
buf  g1358 (n1255, n847);
buf  g1359 (n1202, n924);
not  g1360 (n1718, n801);
buf  g1361 (n1453, n843);
buf  g1362 (n1041, n768);
buf  g1363 (n1339, n894);
not  g1364 (n1044, n917);
not  g1365 (n1178, n963);
not  g1366 (n1116, n753);
not  g1367 (n1624, n582);
not  g1368 (n1090, n754);
buf  g1369 (n1167, n817);
not  g1370 (n1531, n893);
buf  g1371 (n1499, n933);
buf  g1372 (n1537, n839);
not  g1373 (n1330, n892);
buf  g1374 (n1369, n822);
buf  g1375 (n1327, n830);
buf  g1376 (n1685, n781);
not  g1377 (n1040, n728);
not  g1378 (n1427, n941);
buf  g1379 (n1158, n956);
buf  g1380 (n1743, n922);
not  g1381 (n1704, n801);
buf  g1382 (n1615, n898);
buf  g1383 (n1228, n270);
not  g1384 (n972, n765);
buf  g1385 (n1013, n935);
buf  g1386 (n1015, n866);
buf  g1387 (n1207, n801);
buf  g1388 (n1668, n892);
not  g1389 (n1470, n883);
not  g1390 (n1182, n822);
buf  g1391 (n1634, n770);
not  g1392 (n1702, n792);
buf  g1393 (n1465, n900);
buf  g1394 (n1003, n733);
not  g1395 (n1639, n854);
not  g1396 (n1720, n597);
buf  g1397 (n1640, n863);
buf  g1398 (n1591, n910);
buf  g1399 (n1299, n738);
buf  g1400 (n1505, n737);
buf  g1401 (n1190, n823);
not  g1402 (n1363, n839);
buf  g1403 (n1600, n834);
not  g1404 (n1302, n916);
buf  g1405 (n1606, n882);
buf  g1406 (n1197, n933);
buf  g1407 (n1260, n808);
not  g1408 (n1669, n766);
not  g1409 (n1626, n885);
buf  g1410 (n1051, n948);
buf  g1411 (n1169, n793);
buf  g1412 (n1658, n804);
not  g1413 (n1619, n584);
not  g1414 (n1430, n748);
not  g1415 (n1097, n875);
buf  g1416 (n1376, n272);
not  g1417 (n1636, n896);
buf  g1418 (n1445, n879);
buf  g1419 (n1595, n789);
buf  g1420 (n1574, n748);
not  g1421 (n1385, n771);
buf  g1422 (n1226, n384);
buf  g1423 (n1341, n839);
buf  g1424 (n1494, n939);
buf  g1425 (n999, n772);
not  g1426 (n1101, n794);
not  g1427 (n995, n868);
not  g1428 (n1589, n745);
not  g1429 (n1201, n958);
not  g1430 (n1070, n943);
buf  g1431 (n1193, n793);
not  g1432 (n1165, n746);
not  g1433 (n1423, n917);
not  g1434 (n1209, n909);
buf  g1435 (n1154, n773);
not  g1436 (n1198, n796);
not  g1437 (n1130, n585);
buf  g1438 (n1311, n866);
buf  g1439 (n1225, n761);
buf  g1440 (n1166, n727);
buf  g1441 (n1088, n751);
buf  g1442 (n1159, n940);
buf  g1443 (n1649, n938);
not  g1444 (n1725, n933);
buf  g1445 (n1523, n941);
not  g1446 (n978, n905);
buf  g1447 (n1021, n805);
buf  g1448 (n1611, n861);
buf  g1449 (n1733, n821);
buf  g1450 (n1301, n927);
not  g1451 (n1265, n800);
not  g1452 (n993, n863);
buf  g1453 (n1274, n909);
buf  g1454 (n1053, n829);
not  g1455 (n1432, n758);
not  g1456 (n1738, n819);
buf  g1457 (n1342, n766);
not  g1458 (n1067, n956);
buf  g1459 (n967, n775);
buf  g1460 (n1123, n835);
not  g1461 (n1666, n774);
buf  g1462 (n1459, n788);
not  g1463 (n1337, n880);
not  g1464 (n965, n952);
not  g1465 (n1462, n596);
buf  g1466 (n1586, n841);
not  g1467 (n1048, n764);
buf  g1468 (n1118, n939);
buf  g1469 (n1316, n726);
buf  g1470 (n1613, n781);
not  g1471 (n1245, n782);
buf  g1472 (n1308, n799);
buf  g1473 (n1557, n811);
buf  g1474 (n1055, n271);
buf  g1475 (n1188, n930);
not  g1476 (n1323, n899);
buf  g1477 (n1284, n643);
not  g1478 (n1224, n776);
not  g1479 (n1398, n814);
not  g1480 (n1203, n768);
buf  g1481 (n980, n835);
buf  g1482 (n1722, n846);
buf  g1483 (n1185, n798);
not  g1484 (n1735, n746);
buf  g1485 (n1567, n857);
buf  g1486 (n1170, n895);
not  g1487 (n1328, n907);
buf  g1488 (n1576, n907);
not  g1489 (n1469, n760);
not  g1490 (n1137, n962);
not  g1491 (n1419, n815);
not  g1492 (n1450, n840);
buf  g1493 (n1678, n874);
buf  g1494 (n1507, n890);
not  g1495 (n1519, n925);
buf  g1496 (n1199, n886);
buf  g1497 (n1334, n923);
buf  g1498 (n1031, n906);
not  g1499 (n1078, n826);
not  g1500 (n1147, n806);
not  g1501 (n1401, n957);
buf  g1502 (n1073, n903);
not  g1503 (n1362, n912);
not  g1504 (n1217, n873);
buf  g1505 (n1043, n755);
buf  g1506 (n1686, n735);
not  g1507 (n1682, n958);
buf  g1508 (n1075, n857);
buf  g1509 (n1727, n788);
buf  g1510 (n1457, n271);
not  g1511 (n1195, n725);
buf  g1512 (n983, n782);
buf  g1513 (n1278, n638);
not  g1514 (n1131, n884);
buf  g1515 (n1760, n888);
not  g1516 (n1488, n782);
buf  g1517 (n1508, n946);
buf  g1518 (n1628, n836);
buf  g1519 (n1491, n752);
not  g1520 (n1142, n812);
buf  g1521 (n1068, n774);
not  g1522 (n1233, n908);
buf  g1523 (n1546, n921);
buf  g1524 (n1645, n739);
buf  g1525 (n1756, n639);
not  g1526 (n1294, n810);
buf  g1527 (n1208, n898);
buf  g1528 (n1719, n801);
not  g1529 (n1721, n793);
not  g1530 (n1514, n944);
not  g1531 (n1559, n733);
buf  g1532 (n1487, n814);
not  g1533 (n1214, n744);
buf  g1534 (n1651, n890);
buf  g1535 (n1590, n861);
not  g1536 (n1535, n869);
buf  g1537 (n1502, n768);
not  g1538 (n1069, n741);
buf  g1539 (n1313, n902);
not  g1540 (n1179, n878);
not  g1541 (n1748, n865);
not  g1542 (n1604, n847);
not  g1543 (n1322, n842);
not  g1544 (n975, n912);
not  g1545 (n1005, n820);
buf  g1546 (n1729, n930);
not  g1547 (n1050, n913);
not  g1548 (n1191, n876);
buf  g1549 (n1384, n767);
buf  g1550 (n1121, n849);
not  g1551 (n1541, n947);
not  g1552 (n1180, n850);
not  g1553 (n1138, n846);
buf  g1554 (n1451, n889);
buf  g1555 (n1381, n584);
not  g1556 (n1155, n928);
not  g1557 (n1759, n812);
buf  g1558 (n1583, n730);
not  g1559 (n968, n924);
buf  g1560 (n1646, n883);
buf  g1561 (n1269, n590);
not  g1562 (n1753, n760);
buf  g1563 (n1652, n869);
buf  g1564 (n1277, n732);
not  g1565 (n1087, n951);
buf  g1566 (n1286, n816);
not  g1567 (n1448, n809);
buf  g1568 (n1684, n759);
not  g1569 (n1594, n920);
buf  g1570 (n1109, n642);
buf  g1571 (n1749, n938);
not  g1572 (n1681, n843);
not  g1573 (n1351, n921);
not  g1574 (n973, n586);
buf  g1575 (n1017, n810);
buf  g1576 (n1288, n803);
buf  g1577 (n1731, n900);
not  g1578 (n1388, n898);
not  g1579 (n1378, n936);
buf  g1580 (n1100, n861);
buf  g1581 (n1627, n921);
buf  g1582 (n1757, n725);
buf  g1583 (n1396, n779);
not  g1584 (n1321, n896);
buf  g1585 (n1724, n949);
not  g1586 (n1343, n880);
not  g1587 (n1117, n925);
not  g1588 (n1186, n876);
buf  g1589 (n1504, n742);
not  g1590 (n1282, n859);
not  g1591 (n1476, n734);
buf  g1592 (n1402, n815);
buf  g1593 (n1091, n759);
not  g1594 (n997, n805);
buf  g1595 (n1715, n931);
buf  g1596 (n1356, n916);
not  g1597 (n1745, n882);
not  g1598 (n1472, n919);
buf  g1599 (n1455, n888);
buf  g1600 (n1134, n863);
not  g1601 (n1360, n865);
not  g1602 (n1241, n789);
not  g1603 (n1577, n818);
buf  g1604 (n1348, n875);
buf  g1605 (n1503, n813);
not  g1606 (n1145, n810);
not  g1607 (n1108, n757);
buf  g1608 (n1184, n879);
not  g1609 (n1076, n872);
buf  g1610 (n1022, n836);
buf  g1611 (n1629, n853);
not  g1612 (n1018, n737);
not  g1613 (n1085, n897);
and  g1614 (n1601, n841, n864, n811);
nand g1615 (n1449, n778, n920, n886);
xnor g1616 (n1579, n729, n802, n957);
or   g1617 (n1111, n840, n860, n853);
xor  g1618 (n1663, n780, n751, n809);
nor  g1619 (n1181, n762, n806, n269);
nand g1620 (n1026, n948, n741, n857);
or   g1621 (n1200, n729, n740, n592);
xnor g1622 (n1754, n818, n812, n501);
and  g1623 (n1176, n797, n963, n785);
and  g1624 (n1211, n797, n737, n780);
xor  g1625 (n1066, n926, n915, n869);
and  g1626 (n1444, n754, n953, n769);
nand g1627 (n1261, n821, n800, n927);
and  g1628 (n1625, n908, n855, n904);
xor  g1629 (n1149, n946, n918, n850);
nand g1630 (n1144, n849, n743, n826);
nor  g1631 (n1029, n868, n920, n834);
or   g1632 (n1582, n642, n795, n809);
xnor g1633 (n1439, n852, n909, n806);
xor  g1634 (n1412, n824, n598, n777);
nand g1635 (n1045, n804, n786, n854);
or   g1636 (n1710, n739, n726, n778);
or   g1637 (n1367, n875, n821, n271);
nand g1638 (n1662, n923, n730, n774);
xor  g1639 (n1637, n959, n749, n870);
xor  g1640 (n1489, n901, n758, n836);
xnor g1641 (n1525, n849, n856, n878);
nor  g1642 (n1623, n728, n856, n777);
xor  g1643 (n1361, n906, n851, n727);
xnor g1644 (n1246, n744, n867, n769);
nand g1645 (n1216, n791, n901, n928);
or   g1646 (n1358, n922, n924, n912);
nor  g1647 (n1573, n761, n817, n848);
xor  g1648 (n1598, n825, n882, n870);
xor  g1649 (n1023, n784, n781, n924);
and  g1650 (n1675, n915, n918, n752);
nand g1651 (n1534, n961, n763, n639);
or   g1652 (n1317, n891, n757, n815);
nand g1653 (n1355, n960, n877, n874);
xor  g1654 (n1421, n140, n730, n831);
xnor g1655 (n1035, n771, n841, n270);
nor  g1656 (n1125, n864, n774, n816);
nor  g1657 (n969, n754, n894, n813);
or   g1658 (n1605, n742, n827, n950);
or   g1659 (n981, n765, n837, n962);
nand g1660 (n1300, n764, n751, n860);
or   g1661 (n1726, n758, n959, n795);
nand g1662 (n1359, n833, n756, n842);
nor  g1663 (n1124, n501, n747, n757);
or   g1664 (n1454, n864, n752, n747);
nand g1665 (n1128, n963, n848, n906);
or   g1666 (n1695, n926, n742, n826);
nand g1667 (n1183, n785, n942, n802);
and  g1668 (n1293, n803, n910, n808);
and  g1669 (n1407, n748, n819, n269);
nor  g1670 (n998, n862, n825, n890);
and  g1671 (n1703, n954, n822, n827);
nand g1672 (n1080, n798, n844, n819);
nand g1673 (n1479, n899, n600, n872);
or   g1674 (n1431, n783, n784, n817);
and  g1675 (n1156, n755, n957, n955);
nand g1676 (n1632, n880, n944, n757);
or   g1677 (n1739, n864, n960, n738);
or   g1678 (n1400, n889, n853, n873);
nor  g1679 (n1501, n920, n806, n829);
and  g1680 (n1687, n818, n862, n902);
xnor g1681 (n1617, n881, n941, n827);
nor  g1682 (n1107, n890, n788, n804);
nand g1683 (n1708, n859, n872, n837);
nand g1684 (n1564, n800, n641, n784);
xor  g1685 (n1059, n852, n749, n837);
or   g1686 (n1135, n771, n808, n272);
xor  g1687 (n1232, n730, n726, n740);
nand g1688 (n1136, n914, n832, n875);
nor  g1689 (n1357, n725, n640, n949);
and  g1690 (n1285, n818, n736, n775);
and  g1691 (n1596, n844, n845, n727);
xnor g1692 (n1103, n771, n791, n761);
nand g1693 (n1714, n747, n889, n893);
and  g1694 (n1539, n928, n922, n892);
or   g1695 (n1395, n860, n814, n933);
nor  g1696 (n996, n948, n788, n772);
xnor g1697 (n1205, n834, n904, n807);
and  g1698 (n1072, n885, n735, n884);
nor  g1699 (n1247, n936, n917, n895);
nand g1700 (n1086, n887, n799, n754);
xnor g1701 (n1556, n872, n384, n724);
and  g1702 (n1552, n881, n948, n854);
nor  g1703 (n1350, n728, n859, n783);
nor  g1704 (n1054, n957, n823, n871);
xor  g1705 (n988, n855, n843, n838);
xor  g1706 (n1597, n904, n766, n744);
nor  g1707 (n1025, n759, n767, n779);
or   g1708 (n1027, n932, n888, n918);
xor  g1709 (n1677, n763, n820, n930);
xor  g1710 (n1676, n272, n583, n888);
xnor g1711 (n1012, n769, n815, n935);
and  g1712 (n1335, n737, n925, n832);
and  g1713 (n1408, n728, n770, n944);
nand g1714 (n1433, n773, n850, n955);
or   g1715 (n1631, n750, n929, n887);
xnor g1716 (n1389, n938, n911, n884);
or   g1717 (n1690, n895, n763, n781);
or   g1718 (n1140, n794, n824, n732);
xor  g1719 (n1238, n915, n897, n880);
nor  g1720 (n1312, n932, n921, n871);
nand g1721 (n1529, n905, n910, n827);
or   g1722 (n1566, n741, n805, n914);
xnor g1723 (n1267, n908, n270, n756);
xor  g1724 (n1741, n828, n902, n738);
nand g1725 (n1550, n926, n745, n831);
nand g1726 (n1096, n936, n950, n734);
nand g1727 (n974, n794, n787, n786);
nand g1728 (n1866, n1296, n1584, n1436, n1231);
xnor g1729 (n1874, n1048, n1257, n1386, n1357);
and  g1730 (n1828, n1138, n1235, n1598, n1245);
and  g1731 (n1788, n1538, n1038, n1583, n1555);
nand g1732 (n1887, n1310, n1563, n1327, n1276);
and  g1733 (n1808, n1180, n1335, n1390, n1233);
xor  g1734 (n1765, n1376, n1261, n1447, n1365);
xnor g1735 (n1815, n1501, n1520, n1755, n1504);
and  g1736 (n1837, n1674, n1605, n1179, n1735);
and  g1737 (n1956, n1173, n1422, n1266, n985);
or   g1738 (n1853, n1306, n1575, n1618, n1132);
nor  g1739 (n1813, n1661, n1329, n1711, n1289);
nand g1740 (n1884, n1092, n1258, n1647, n1207);
xor  g1741 (n1958, n1095, n1526, n1644, n991);
or   g1742 (n1782, n1519, n1517, n1359, n1592);
or   g1743 (n1785, n1740, n1637, n1731, n1349);
and  g1744 (n1806, n1251, n1337, n1486, n1604);
and  g1745 (n1886, n1518, n1368, n1712, n1154);
or   g1746 (n1794, n1608, n999, n1225, n1668);
xor  g1747 (n1933, n1030, n1254, n1622, n1283);
and  g1748 (n1950, n1487, n1209, n1750, n1660);
nor  g1749 (n1944, n1081, n1094, n1751, n1698);
xor  g1750 (n1763, n1470, n1722, n1282, n1745);
and  g1751 (n1924, n1279, n1286, n1184, n1114);
xnor g1752 (n1859, n1111, n1272, n1719, n1195);
or   g1753 (n1882, n1280, n1560, n1211, n1333);
nor  g1754 (n1791, n980, n1161, n1688, n1490);
xor  g1755 (n1790, n981, n1435, n1650, n1183);
nand g1756 (n1875, n1489, n1287, n1371, n987);
xor  g1757 (n1830, n1427, n1364, n1221, n1417);
xor  g1758 (n1845, n1193, n1169, n1044, n1640);
or   g1759 (n1904, n1099, n1308, n1194, n31);
xor  g1760 (n1817, n1288, n1240, n993, n1423);
nor  g1761 (n1824, n1260, n1631, n1140, n1402);
nor  g1762 (n1779, n1147, n1186, n1148, n1710);
or   g1763 (n1931, n1293, n1757, n1331, n1119);
nor  g1764 (n1778, n1581, n1013, n32, n1480);
xor  g1765 (n1869, n1466, n1375, n1692, n1336);
xor  g1766 (n1903, n1571, n1174, n1017, n1666);
xor  g1767 (n1955, n1429, n1085, n1050, n1597);
nor  g1768 (n1901, n1524, n1411, n1222, n1426);
or   g1769 (n1927, n1700, n1488, n1314, n1691);
xnor g1770 (n1821, n1029, n1155, n1322, n1468);
nor  g1771 (n1786, n1556, n1086, n1216, n1752);
nand g1772 (n1796, n1239, n986, n1106, n997);
or   g1773 (n1803, n30, n1152, n1215, n1593);
or   g1774 (n1800, n1162, n1016, n1158, n1758);
nor  g1775 (n1776, n1635, n1373, n1671, n1485);
xor  g1776 (n1816, n1479, n1311, n1642, n1213);
and  g1777 (n1825, n1407, n1063, n1075, n1304);
xnor g1778 (n1851, n1709, n1609, n1475, n1274);
nand g1779 (n1841, n1256, n1399, n1277, n1157);
xor  g1780 (n1959, n1118, n1495, n989, n1483);
nand g1781 (n1768, n1549, n1145, n1369, n1476);
xor  g1782 (n1916, n1127, n994, n1393, n1084);
xor  g1783 (n1963, n1238, n1036, n1006, n1060);
or   g1784 (n1784, n1101, n1391, n1658, n1301);
nand g1785 (n1940, n1612, n1267, n1508, n1096);
xnor g1786 (n1829, n1548, n1724, n1250, n1596);
nor  g1787 (n1801, n1345, n1615, n1088, n1482);
xor  g1788 (n1890, n1338, n1024, n1034, n1703);
or   g1789 (n1804, n1143, n1675, n1537, n1190);
xor  g1790 (n1912, n1228, n1116, n1199, n1182);
xor  g1791 (n1952, n1454, n1366, n1634, n1303);
or   g1792 (n1810, n1412, n1129, n1205, n1377);
xnor g1793 (n1879, n1049, n1552, n1672, n1621);
and  g1794 (n1920, n1275, n1643, n1591, n1149);
nand g1795 (n1939, n1577, n1540, n1340, n966);
nand g1796 (n1802, n972, n1684, n1401, n1056);
or   g1797 (n1921, n1108, n1632, n1723, n964);
xor  g1798 (n1792, n971, n1649, n1104, n1421);
xnor g1799 (n1818, n1443, n1565, n1534, n1545);
xnor g1800 (n1907, n1342, n1460, n1410, n1284);
or   g1801 (n1781, n1300, n1396, n1727, n1752);
nor  g1802 (n1949, n1394, n1458, n982, n1522);
xnor g1803 (n1905, n1346, n1478, n1247, n1040);
xor  g1804 (n1926, n31, n1502, n1599, n1290);
nor  g1805 (n1900, n1014, n1619, n1617, n1646);
and  g1806 (n1928, n1586, n1753, n1718, n1419);
xor  g1807 (n1826, n1069, n1414, n1062, n1496);
and  g1808 (n1807, n1015, n1271, n1166, n1601);
xor  g1809 (n1917, n1641, n1744, n1758, n1003);
or   g1810 (n1771, n1620, n1046, n1494, n1319);
nor  g1811 (n1892, n1053, n1384, n30, n1626);
nand g1812 (n1805, n1197, n1507, n1564, n1227);
xor  g1813 (n1895, n1165, n1602, n1613, n1606);
or   g1814 (n1915, n1012, n1756, n1686, n1418);
nand g1815 (n1889, n1332, n1446, n1645, n1202);
xor  g1816 (n1898, n1655, n1362, n1144, n1531);
or   g1817 (n1766, n1754, n1701, n1098, n1582);
xor  g1818 (n1906, n1298, n1743, n1334, n973);
nand g1819 (n1809, n1150, n1570, n1188, n1133);
and  g1820 (n1854, n1058, n1026, n1669, n1192);
nor  g1821 (n1951, n1625, n1051, n1409, n1527);
xnor g1822 (n1902, n1497, n1702, n1455, n975);
nand g1823 (n1919, n1433, n1403, n1268, n1347);
nor  g1824 (n1930, n1474, n1430, n1055, n1262);
xor  g1825 (n1881, n1134, n1413, n1679, n1074);
xor  g1826 (n1774, n1253, n1512, n1082, n1379);
nand g1827 (n1839, n1378, n1153, n1292, n1059);
nand g1828 (n1961, n1243, n1022, n1648, n1208);
xnor g1829 (n1945, n1687, n1543, n1156, n1229);
nand g1830 (n1789, n1083, n1326, n1629, n974);
and  g1831 (n1864, n1318, n1676, n1677, n1071);
nor  g1832 (n1953, n1728, n1370, n1484, n1749);
and  g1833 (n1836, n1350, n1307, n1170, n1664);
nor  g1834 (n1957, n1682, n1442, n1694, n1073);
or   g1835 (n1948, n1547, n1295, n1007, n1313);
nand g1836 (n1764, n1139, n1741, n32, n1043);
xor  g1837 (n1932, n1733, n1544, n1706, n1695);
and  g1838 (n1855, n1027, n1627, n1037, n1492);
or   g1839 (n1850, n1554, n1623, n1562, n1168);
nand g1840 (n1962, n1005, n1693, n1725, n1325);
or   g1841 (n1769, n1230, n1499, n1477, n1690);
nor  g1842 (n1885, n1117, n1103, n1392, n1343);
nor  g1843 (n1812, n1498, n1441, n1328, n1236);
and  g1844 (n1772, n1572, n1210, n1281, n1525);
nor  g1845 (n1822, n1681, n1453, n1039, n1395);
or   g1846 (n1857, n1714, n1491, n1115, n1397);
xor  g1847 (n1835, n1516, n969, n1382, n1737);
xor  g1848 (n1761, n1019, n1273, n1141, n1720);
xor  g1849 (n1783, n1717, n1509, n1330, n1503);
nor  g1850 (n1797, n1579, n1457, n1696, n1107);
nor  g1851 (n1878, n1535, n1473, n1189, n1678);
nor  g1852 (n1844, n1461, n1372, n1406, n1387);
and  g1853 (n1899, n1550, n1360, n1356, n1363);
xnor g1854 (n1873, n1090, n1576, n1532, n1076);
xor  g1855 (n1811, n1341, n1025, n1746, n1351);
nand g1856 (n1888, n1529, n1177, n1175, n1590);
nand g1857 (n1799, n1109, n1546, n1680, n1756);
or   g1858 (n1856, n1699, n1159, n1708, n1748);
xor  g1859 (n1935, n1057, n1573, n1742, n1163);
xnor g1860 (n1954, n1639, n968, n1320, n1408);
xor  g1861 (n1840, n1707, n1381, n1449, n1316);
nand g1862 (n1870, n1067, n30, n1515, n1424);
or   g1863 (n1946, n1469, n31, n1285, n1079);
nor  g1864 (n1923, n1224, n1078, n1726, n1416);
nor  g1865 (n1943, n1070, n978, n1052, n1045);
xnor g1866 (n1929, n1705, n1514, n1234, n1683);
or   g1867 (n1880, n1652, n1252, n1181, n1616);
nor  g1868 (n1838, n1237, n1110, n1588, n976);
xnor g1869 (n1795, n1246, n1054, n1223, n1294);
and  g1870 (n1858, n1673, n1220, n1630, n1715);
xnor g1871 (n1861, n1732, n1611, n1120, n30);
and  g1872 (n1937, n1665, n1729, n1219, n439);
nand g1873 (n1848, n1656, n1511, n32, n1226);
nor  g1874 (n1820, n1077, n1533, n1628, n1578);
nand g1875 (n1787, n1659, n1574, n1481, n1721);
and  g1876 (n1922, n1198, n1380, n1018, n1136);
nand g1877 (n1925, n1551, n1439, n1452, n1603);
and  g1878 (n1918, n1438, n1041, n1204, n1638);
nand g1879 (n1908, n1263, n1259, n1667, n1185);
or   g1880 (n1814, n1353, n1121, n1011, n1035);
nor  g1881 (n1947, n1348, n1172, n1249, n1061);
nand g1882 (n1827, n1309, n1164, n1321, n1305);
nand g1883 (n1767, n1028, n1428, n1214, n1600);
nor  g1884 (n1831, n1142, n1450, n1102, n1066);
or   g1885 (n1798, n1730, n1542, n1355, n1594);
and  g1886 (n1777, n1670, n1033, n1697, n1464);
xnor g1887 (n1942, n1244, n990, n1255, n1171);
xnor g1888 (n1865, n1241, n1462, n1021, n1146);
nor  g1889 (n1909, n1178, n1654, n1009, n1425);
or   g1890 (n1911, n967, n1270, n1093, n970);
xor  g1891 (n1913, n1528, n1521, n1042, n1539);
and  g1892 (n1914, n1716, n1607, n1137, n1465);
or   g1893 (n1868, n1383, n1589, n1523, n1734);
nor  g1894 (n1849, n1297, n1557, n1567, n1068);
nand g1895 (n1871, n1493, n1126, n1739, n1167);
xnor g1896 (n1833, n1004, n1196, n1242, n1124);
xor  g1897 (n1893, n1269, n1354, n1431, n992);
and  g1898 (n1941, n984, n1657, n1663, n1569);
nor  g1899 (n1770, n1530, n1385, n1367, n1374);
and  g1900 (n1780, n1689, n1361, n1105, n1753);
and  g1901 (n1910, n1610, n1437, n1001, n977);
nor  g1902 (n1862, n1176, n1302, n1031, n31);
xor  g1903 (n1793, n1456, n1339, n1662, n1312);
xnor g1904 (n1842, n1404, n1317, n1089, n983);
nand g1905 (n1819, n1559, n1624, n1130, n1614);
or   g1906 (n1883, n1087, n1595, n1463, n32);
xnor g1907 (n1823, n1420, n988, n1135, n1472);
xnor g1908 (n1936, n1445, n1653, n1125, n1122);
xnor g1909 (n1834, n1388, n1467, n1151, n1636);
xor  g1910 (n1846, n998, n1398, n1738, n1736);
nor  g1911 (n1964, n1278, n1100, n1160, n1561);
nor  g1912 (n1775, n1248, n1568, n1405, n1080);
xor  g1913 (n1891, n1541, n1217, n1585, n1506);
nand g1914 (n1843, n1112, n1206, n1505, n1010);
xor  g1915 (n1897, n1008, n1002, n1128, n995);
nand g1916 (n1894, n1558, n1023, n1000, n1097);
xor  g1917 (n1877, n1415, n1131, n1451, n1064);
xor  g1918 (n1876, n1264, n1091, n1587, n1513);
xnor g1919 (n1852, n1755, n1358, n1400, n1047);
and  g1920 (n1867, n1191, n1713, n1020, n1747);
nor  g1921 (n1863, n1344, n1751, n1580, n1352);
and  g1922 (n1934, n979, n1065, n1434, n1471);
nand g1923 (n1860, n1754, n1201, n1323, n1324);
nor  g1924 (n1847, n1265, n1212, n1448, n1651);
and  g1925 (n1896, n1704, n1291, n1200, n965);
xnor g1926 (n1773, n1757, n1536, n996, n1566);
xor  g1927 (n1960, n1072, n1113, n1510, n1432);
nand g1928 (n1832, n1203, n1685, n1123, n1187);
and  g1929 (n1872, n1459, n1218, n1553, n1315);
xor  g1930 (n1762, n1500, n1299, n1444, n1389);
nand g1931 (n1938, n1232, n1633, n1032, n1440);
xor  g1932 (n1967, n1834, n1810, n1802, n1913);
xnor g1933 (n1983, n1767, n1856, n1805, n1850);
nand g1934 (n1966, n1900, n1911, n1874, n1809);
nor  g1935 (n1986, n1778, n1864, n1806, n1907);
nor  g1936 (n1982, n1857, n1871, n1765, n1814);
and  g1937 (n1997, n1869, n1768, n1782, n1852);
and  g1938 (n1985, n1837, n1876, n1813, n1863);
xor  g1939 (n2002, n1788, n1812, n1793, n1799);
xnor g1940 (n1968, n1783, n1855, n1779, n1898);
nand g1941 (n1965, n1872, n1853, n1828, n1894);
nand g1942 (n2003, n1902, n1829, n1886, n1791);
xnor g1943 (n1980, n1831, n1861, n1873, n1801);
xor  g1944 (n1981, n1835, n1780, n1798, n1905);
or   g1945 (n1994, n1832, n1794, n1860, n1878);
and  g1946 (n1971, n1881, n1879, n1846, n1789);
xnor g1947 (n1993, n1770, n1893, n1776, n1766);
nand g1948 (n1998, n1868, n1897, n1899, n1787);
xnor g1949 (n1974, n1867, n1781, n1800, n1804);
nor  g1950 (n1970, n1859, n1824, n1910, n1796);
nor  g1951 (n1978, n1889, n1771, n1896, n1775);
or   g1952 (n1979, n1821, n1862, n1774, n1884);
nor  g1953 (n1976, n1888, n1841, n1797, n1875);
nor  g1954 (n2000, n1885, n1847, n1819, n1877);
xor  g1955 (n1969, n1764, n1763, n1843, n1833);
nand g1956 (n1989, n1890, n1887, n1823, n1842);
xnor g1957 (n1975, n1792, n1826, n1830, n1838);
xor  g1958 (n1973, n1870, n1914, n1895, n1777);
nor  g1959 (n1996, n1844, n1817, n1882, n1840);
xor  g1960 (n1987, n1790, n1818, n1762, n1849);
nor  g1961 (n1972, n1909, n1891, n1836, n1848);
and  g1962 (n1984, n1786, n1773, n1807, n1827);
nand g1963 (n1991, n1820, n1903, n1858, n1815);
nand g1964 (n1992, n1912, n1854, n1811, n1865);
xor  g1965 (n2001, n1772, n1825, n1851, n1839);
xnor g1966 (n1977, n1906, n1795, n1908, n1880);
and  g1967 (n1999, n1803, n1916, n1892, n1904);
or   g1968 (n1990, n1866, n1883, n1808, n1761);
nand g1969 (n1995, n1785, n1816, n1784, n1901);
xor  g1970 (n1988, n1845, n1915, n1822, n1769);
xnor g1971 (n2007, n273, n1994, n1992, n1999);
and  g1972 (n2006, n1991, n1993, n273, n2000);
nor  g1973 (n2004, n1989, n1996, n1998, n1988);
or   g1974 (n2005, n1995, n1990, n1997, n274);
nor  g1975 (n2008, n2007, n374);
or   g1976 (n2012, n140, n2008, n2002, n274);
or   g1977 (n2009, n2001, n274, n2008);
and  g1978 (n2010, n2008, n1760, n1759, n2003);
xor  g1979 (n2011, n1760, n140, n1759, n2008);
nand g1980 (n2019, n1946, n2011, n1960, n1917);
xnor g1981 (n2016, n1955, n1934, n2009, n1951);
xor  g1982 (n2020, n1939, n1956, n1944, n2010);
xnor g1983 (n2013, n1928, n1947, n1941, n1922);
and  g1984 (n2015, n1936, n2012, n1932, n1964);
nor  g1985 (n2014, n1924, n2009, n2011, n1931);
xor  g1986 (n2025, n2012, n1930, n1940, n1957);
or   g1987 (n2021, n1919, n1945, n1942, n1958);
nor  g1988 (n2022, n2010, n1921, n1961, n1926);
or   g1989 (n2017, n1953, n1962, n1937, n1920);
xor  g1990 (n2024, n2012, n1950, n1923, n1949);
and  g1991 (n2023, n1959, n1954, n2011, n1963);
xor  g1992 (n2028, n1938, n1918, n1933, n2010);
or   g1993 (n2026, n2012, n1952, n2011, n2009);
xnor g1994 (n2027, n1929, n2009, n1948, n1935);
xor  g1995 (n2018, n1927, n2010, n1943, n1925);
and  g1996 (n2032, n2017, n2027, n2019, n2018);
and  g1997 (n2030, n2015, n2026, n2014, n2022);
xor  g1998 (n2029, n2021, n2028, n2013, n2025);
xor  g1999 (n2031, n2016, n2024, n2020, n2023);
endmodule
