

module Stat_1857_36_9
(
  n1,
  n2,
  n3,
  n4,
  n5,
  n6,
  n7,
  n8,
  n9,
  n10,
  n11,
  n12,
  n13,
  n14,
  n15,
  n16,
  n17,
  n18,
  n19,
  n20,
  n21,
  n1769,
  n1764,
  n1763,
  n1768,
  n1829,
  n1830,
  n1837,
  n1831,
  n1833,
  n1835,
  n1865,
  n1867,
  n1861,
  n1864,
  n1862,
  n1863,
  n1868,
  n1866,
  n1869,
  n1878
);

  input n1;input n2;input n3;input n4;input n5;input n6;input n7;input n8;input n9;input n10;input n11;input n12;input n13;input n14;input n15;input n16;input n17;input n18;input n19;input n20;input n21;input keyIn_0_0;input keyIn_0_1;input keyIn_0_2;input keyIn_0_3;input keyIn_0_4;input keyIn_0_5;input keyIn_0_6;input keyIn_0_7;input keyIn_0_8;input keyIn_0_9;input keyIn_0_10;input keyIn_0_11;input keyIn_0_12;input keyIn_0_13;input keyIn_0_14;input keyIn_0_15;input keyIn_0_16;input keyIn_0_17;input keyIn_0_18;input keyIn_0_19;input keyIn_0_20;input keyIn_0_21;input keyIn_0_22;input keyIn_0_23;input keyIn_0_24;input keyIn_0_25;input keyIn_0_26;input keyIn_0_27;input keyIn_0_28;input keyIn_0_29;input keyIn_0_30;input keyIn_0_31;
  output n1769;output n1764;output n1763;output n1768;output n1829;output n1830;output n1837;output n1831;output n1833;output n1835;output n1865;output n1867;output n1861;output n1864;output n1862;output n1863;output n1868;output n1866;output n1869;output n1878;
  wire n22;wire n23;wire n24;wire n25;wire n26;wire n27;wire n28;wire n29;wire n30;wire n31;wire n32;wire n33;wire n34;wire n35;wire n36;wire n37;wire n38;wire n39;wire n40;wire n41;wire n42;wire n43;wire n44;wire n45;wire n46;wire n47;wire n48;wire n49;wire n50;wire n51;wire n52;wire n53;wire n54;wire n55;wire n56;wire n57;wire n58;wire n59;wire n60;wire n61;wire n62;wire n63;wire n64;wire n65;wire n66;wire n67;wire n68;wire n69;wire n70;wire n71;wire n72;wire n73;wire n74;wire n75;wire n76;wire n77;wire n78;wire n79;wire n80;wire n81;wire n82;wire n83;wire n84;wire n85;wire n86;wire n87;wire n88;wire n89;wire n90;wire n91;wire n92;wire n93;wire n94;wire n95;wire n96;wire n97;wire n98;wire n99;wire n100;wire n101;wire n102;wire n103;wire n104;wire n105;wire n106;wire n107;wire n108;wire n109;wire n110;wire n111;wire n112;wire n113;wire n114;wire n115;wire n116;wire n117;wire n118;wire n119;wire n120;wire n121;wire n122;wire n123;wire n124;wire n125;wire n126;wire n127;wire n128;wire n129;wire n130;wire n131;wire n132;wire n133;wire n134;wire n135;wire n136;wire n137;wire n138;wire n139;wire n140;wire n141;wire n142;wire n143;wire n144;wire n145;wire n146;wire n147;wire n148;wire n149;wire n150;wire n151;wire n152;wire n153;wire n154;wire n155;wire n156;wire n157;wire n158;wire n159;wire n160;wire n161;wire n162;wire n163;wire n164;wire n165;wire n166;wire n167;wire n168;wire n169;wire n170;wire n171;wire n172;wire n173;wire n174;wire n175;wire n176;wire n177;wire n178;wire n179;wire n180;wire n181;wire n182;wire n183;wire n184;wire n185;wire n186;wire n187;wire n188;wire n189;wire n190;wire n191;wire n192;wire n193;wire n194;wire n195;wire n196;wire n197;wire n198;wire n199;wire n200;wire n201;wire n202;wire n203;wire n204;wire n205;wire n206;wire n207;wire n208;wire n209;wire n210;wire n211;wire n212;wire n213;wire n214;wire n215;wire n216;wire n217;wire n218;wire n219;wire n220;wire n221;wire n222;wire n223;wire n224;wire n225;wire n226;wire n227;wire n228;wire n229;wire n230;wire n231;wire n232;wire n233;wire n234;wire n235;wire n236;wire n237;wire n238;wire n239;wire n240;wire n241;wire n242;wire n243;wire n244;wire n245;wire n246;wire n247;wire n248;wire n249;wire n250;wire n251;wire n252;wire n253;wire n254;wire n255;wire n256;wire n257;wire n258;wire n259;wire n260;wire n261;wire n262;wire n263;wire n264;wire n265;wire n266;wire n267;wire n268;wire n269;wire n270;wire n271;wire n272;wire n273;wire n274;wire n275;wire n276;wire n277;wire n278;wire n279;wire n280;wire n281;wire n282;wire n283;wire n284;wire n285;wire n286;wire n287;wire n288;wire n289;wire n290;wire n291;wire n292;wire n293;wire n294;wire n295;wire n296;wire n297;wire n298;wire n299;wire n300;wire n301;wire n302;wire n303;wire n304;wire n305;wire n306;wire n307;wire n308;wire n309;wire n310;wire n311;wire n312;wire n313;wire n314;wire n315;wire n316;wire n317;wire n318;wire n319;wire n320;wire n321;wire n322;wire n323;wire n324;wire n325;wire n326;wire n327;wire n328;wire n329;wire n330;wire n331;wire n332;wire n333;wire n334;wire n335;wire n336;wire n337;wire n338;wire n339;wire n340;wire n341;wire n342;wire n343;wire n344;wire n345;wire n346;wire n347;wire n348;wire n349;wire n350;wire n351;wire n352;wire n353;wire n354;wire n355;wire n356;wire n357;wire n358;wire n359;wire n360;wire n361;wire n362;wire n363;wire n364;wire n365;wire n366;wire n367;wire n368;wire n369;wire n370;wire n371;wire n372;wire n373;wire n374;wire n375;wire n376;wire n377;wire n378;wire n379;wire n380;wire n381;wire n382;wire n383;wire n384;wire n385;wire n386;wire n387;wire n388;wire n389;wire n390;wire n391;wire n392;wire n393;wire n394;wire n395;wire n396;wire n397;wire n398;wire n399;wire n400;wire n401;wire n402;wire n403;wire n404;wire n405;wire n406;wire n407;wire n408;wire n409;wire n410;wire n411;wire n412;wire n413;wire n414;wire n415;wire n416;wire n417;wire n418;wire n419;wire n420;wire n421;wire n422;wire n423;wire n424;wire n425;wire n426;wire n427;wire n428;wire n429;wire n430;wire n431;wire n432;wire n433;wire n434;wire n435;wire n436;wire n437;wire n438;wire n439;wire n440;wire n441;wire n442;wire n443;wire n444;wire n445;wire n446;wire n447;wire n448;wire n449;wire n450;wire n451;wire n452;wire n453;wire n454;wire n455;wire n456;wire n457;wire n458;wire n459;wire n460;wire n461;wire n462;wire n463;wire n464;wire n465;wire n466;wire n467;wire n468;wire n469;wire n470;wire n471;wire n472;wire n473;wire n474;wire n475;wire n476;wire n477;wire n478;wire n479;wire n480;wire n481;wire n482;wire n483;wire n484;wire n485;wire n486;wire n487;wire n488;wire n489;wire n490;wire n491;wire n492;wire n493;wire n494;wire n495;wire n496;wire n497;wire n498;wire n499;wire n500;wire n501;wire n502;wire n503;wire n504;wire n505;wire n506;wire n507;wire n508;wire n509;wire n510;wire n511;wire n512;wire n513;wire n514;wire n515;wire n516;wire n517;wire n518;wire n519;wire n520;wire n521;wire n522;wire n523;wire n524;wire n525;wire n526;wire n527;wire n528;wire n529;wire n530;wire n531;wire n532;wire n533;wire n534;wire n535;wire n536;wire n537;wire n538;wire n539;wire n540;wire n541;wire n542;wire n543;wire n544;wire n545;wire n546;wire n547;wire n548;wire n549;wire n550;wire n551;wire n552;wire n553;wire n554;wire n555;wire n556;wire n557;wire n558;wire n559;wire n560;wire n561;wire n562;wire n563;wire n564;wire n565;wire n566;wire n567;wire n568;wire n569;wire n570;wire n571;wire n572;wire n573;wire n574;wire n575;wire n576;wire n577;wire n578;wire n579;wire n580;wire n581;wire n582;wire n583;wire n584;wire n585;wire n586;wire n587;wire n588;wire n589;wire n590;wire n591;wire n592;wire n593;wire n594;wire n595;wire n596;wire n597;wire n598;wire n599;wire n600;wire n601;wire n602;wire n603;wire n604;wire n605;wire n606;wire n607;wire n608;wire n609;wire n610;wire n611;wire n612;wire n613;wire n614;wire n615;wire n616;wire n617;wire n618;wire n619;wire n620;wire n621;wire n622;wire n623;wire n624;wire n625;wire n626;wire n627;wire n628;wire n629;wire n630;wire n631;wire n632;wire n633;wire n634;wire n635;wire n636;wire n637;wire n638;wire n639;wire n640;wire n641;wire n642;wire n643;wire n644;wire n645;wire n646;wire n647;wire n648;wire n649;wire n650;wire n651;wire n652;wire n653;wire n654;wire n655;wire n656;wire n657;wire n658;wire n659;wire n660;wire n661;wire n662;wire n663;wire n664;wire n665;wire n666;wire n667;wire n668;wire n669;wire n670;wire n671;wire n672;wire n673;wire n674;wire n675;wire n676;wire n677;wire n678;wire n679;wire n680;wire n681;wire n682;wire n683;wire n684;wire n685;wire n686;wire n687;wire n688;wire n689;wire n690;wire n691;wire n692;wire n693;wire n694;wire n695;wire n696;wire n697;wire n698;wire n699;wire n700;wire n701;wire n702;wire n703;wire n704;wire n705;wire n706;wire n707;wire n708;wire n709;wire n710;wire n711;wire n712;wire n713;wire n714;wire n715;wire n716;wire n717;wire n718;wire n719;wire n720;wire n721;wire n722;wire n723;wire n724;wire n725;wire n726;wire n727;wire n728;wire n729;wire n730;wire n731;wire n732;wire n733;wire n734;wire n735;wire n736;wire n737;wire n738;wire n739;wire n740;wire n741;wire n742;wire n743;wire n744;wire n745;wire n746;wire n747;wire n748;wire n749;wire n750;wire n751;wire n752;wire n753;wire n754;wire n755;wire n756;wire n757;wire n758;wire n759;wire n760;wire n761;wire n762;wire n763;wire n764;wire n765;wire n766;wire n767;wire n768;wire n769;wire n770;wire n771;wire n772;wire n773;wire n774;wire n775;wire n776;wire n777;wire n778;wire n779;wire n780;wire n781;wire n782;wire n783;wire n784;wire n785;wire n786;wire n787;wire n788;wire n789;wire n790;wire n791;wire n792;wire n793;wire n794;wire n795;wire n796;wire n797;wire n798;wire n799;wire n800;wire n801;wire n802;wire n803;wire n804;wire n805;wire n806;wire n807;wire n808;wire n809;wire n810;wire n811;wire n812;wire n813;wire n814;wire n815;wire n816;wire n817;wire n818;wire n819;wire n820;wire n821;wire n822;wire n823;wire n824;wire n825;wire n826;wire n827;wire n828;wire n829;wire n830;wire n831;wire n832;wire n833;wire n834;wire n835;wire n836;wire n837;wire n838;wire n839;wire n840;wire n841;wire n842;wire n843;wire n844;wire n845;wire n846;wire n847;wire n848;wire n849;wire n850;wire n851;wire n852;wire n853;wire n854;wire n855;wire n856;wire n857;wire n858;wire n859;wire n860;wire n861;wire n862;wire n863;wire n864;wire n865;wire n866;wire n867;wire n868;wire n869;wire n870;wire n871;wire n872;wire n873;wire n874;wire n875;wire n876;wire n877;wire n878;wire n879;wire n880;wire n881;wire n882;wire n883;wire n884;wire n885;wire n886;wire n887;wire n888;wire n889;wire n890;wire n891;wire n892;wire n893;wire n894;wire n895;wire n896;wire n897;wire n898;wire n899;wire n900;wire n901;wire n902;wire n903;wire n904;wire n905;wire n906;wire n907;wire n908;wire n909;wire n910;wire n911;wire n912;wire n913;wire n914;wire n915;wire n916;wire n917;wire n918;wire n919;wire n920;wire n921;wire n922;wire n923;wire n924;wire n925;wire n926;wire n927;wire n928;wire n929;wire n930;wire n931;wire n932;wire n933;wire n934;wire n935;wire n936;wire n937;wire n938;wire n939;wire n940;wire n941;wire n942;wire n943;wire n944;wire n945;wire n946;wire n947;wire n948;wire n949;wire n950;wire n951;wire n952;wire n953;wire n954;wire n955;wire n956;wire n957;wire n958;wire n959;wire n960;wire n961;wire n962;wire n963;wire n964;wire n965;wire n966;wire n967;wire n968;wire n969;wire n970;wire n971;wire n972;wire n973;wire n974;wire n975;wire n976;wire n977;wire n978;wire n979;wire n980;wire n981;wire n982;wire n983;wire n984;wire n985;wire n986;wire n987;wire n988;wire n989;wire n990;wire n991;wire n992;wire n993;wire n994;wire n995;wire n996;wire n997;wire n998;wire n999;wire n1000;wire n1001;wire n1002;wire n1003;wire n1004;wire n1005;wire n1006;wire n1007;wire n1008;wire n1009;wire n1010;wire n1011;wire n1012;wire n1013;wire n1014;wire n1015;wire n1016;wire n1017;wire n1018;wire n1019;wire n1020;wire n1021;wire n1022;wire n1023;wire n1024;wire n1025;wire n1026;wire n1027;wire n1028;wire n1029;wire n1030;wire n1031;wire n1032;wire n1033;wire n1034;wire n1035;wire n1036;wire n1037;wire n1038;wire n1039;wire n1040;wire n1041;wire n1042;wire n1043;wire n1044;wire n1045;wire n1046;wire n1047;wire n1048;wire n1049;wire n1050;wire n1051;wire n1052;wire n1053;wire n1054;wire n1055;wire n1056;wire n1057;wire n1058;wire n1059;wire n1060;wire n1061;wire n1062;wire n1063;wire n1064;wire n1065;wire n1066;wire n1067;wire n1068;wire n1069;wire n1070;wire n1071;wire n1072;wire n1073;wire n1074;wire n1075;wire n1076;wire n1077;wire n1078;wire n1079;wire n1080;wire n1081;wire n1082;wire n1083;wire n1084;wire n1085;wire n1086;wire n1087;wire n1088;wire n1089;wire n1090;wire n1091;wire n1092;wire n1093;wire n1094;wire n1095;wire n1096;wire n1097;wire n1098;wire n1099;wire n1100;wire n1101;wire n1102;wire n1103;wire n1104;wire n1105;wire n1106;wire n1107;wire n1108;wire n1109;wire n1110;wire n1111;wire n1112;wire n1113;wire n1114;wire n1115;wire n1116;wire n1117;wire n1118;wire n1119;wire n1120;wire n1121;wire n1122;wire n1123;wire n1124;wire n1125;wire n1126;wire n1127;wire n1128;wire n1129;wire n1130;wire n1131;wire n1132;wire n1133;wire n1134;wire n1135;wire n1136;wire n1137;wire n1138;wire n1139;wire n1140;wire n1141;wire n1142;wire n1143;wire n1144;wire n1145;wire n1146;wire n1147;wire n1148;wire n1149;wire n1150;wire n1151;wire n1152;wire n1153;wire n1154;wire n1155;wire n1156;wire n1157;wire n1158;wire n1159;wire n1160;wire n1161;wire n1162;wire n1163;wire n1164;wire n1165;wire n1166;wire n1167;wire n1168;wire n1169;wire n1170;wire n1171;wire n1172;wire n1173;wire n1174;wire n1175;wire n1176;wire n1177;wire n1178;wire n1179;wire n1180;wire n1181;wire n1182;wire n1183;wire n1184;wire n1185;wire n1186;wire n1187;wire n1188;wire n1189;wire n1190;wire n1191;wire n1192;wire n1193;wire n1194;wire n1195;wire n1196;wire n1197;wire n1198;wire n1199;wire n1200;wire n1201;wire n1202;wire n1203;wire n1204;wire n1205;wire n1206;wire n1207;wire n1208;wire n1209;wire n1210;wire n1211;wire n1212;wire n1213;wire n1214;wire n1215;wire n1216;wire n1217;wire n1218;wire n1219;wire n1220;wire n1221;wire n1222;wire n1223;wire n1224;wire n1225;wire n1226;wire n1227;wire n1228;wire n1229;wire n1230;wire n1231;wire n1232;wire n1233;wire n1234;wire n1235;wire n1236;wire n1237;wire n1238;wire n1239;wire n1240;wire n1241;wire n1242;wire n1243;wire n1244;wire n1245;wire n1246;wire n1247;wire n1248;wire n1249;wire n1250;wire n1251;wire n1252;wire n1253;wire n1254;wire n1255;wire n1256;wire n1257;wire n1258;wire n1259;wire n1260;wire n1261;wire n1262;wire n1263;wire n1264;wire n1265;wire n1266;wire n1267;wire n1268;wire n1269;wire n1270;wire n1271;wire n1272;wire n1273;wire n1274;wire n1275;wire n1276;wire n1277;wire n1278;wire n1279;wire n1280;wire n1281;wire n1282;wire n1283;wire n1284;wire n1285;wire n1286;wire n1287;wire n1288;wire n1289;wire n1290;wire n1291;wire n1292;wire n1293;wire n1294;wire n1295;wire n1296;wire n1297;wire n1298;wire n1299;wire n1300;wire n1301;wire n1302;wire n1303;wire n1304;wire n1305;wire n1306;wire n1307;wire n1308;wire n1309;wire n1310;wire n1311;wire n1312;wire n1313;wire n1314;wire n1315;wire n1316;wire n1317;wire n1318;wire n1319;wire n1320;wire n1321;wire n1322;wire n1323;wire n1324;wire n1325;wire n1326;wire n1327;wire n1328;wire n1329;wire n1330;wire n1331;wire n1332;wire n1333;wire n1334;wire n1335;wire n1336;wire n1337;wire n1338;wire n1339;wire n1340;wire n1341;wire n1342;wire n1343;wire n1344;wire n1345;wire n1346;wire n1347;wire n1348;wire n1349;wire n1350;wire n1351;wire n1352;wire n1353;wire n1354;wire n1355;wire n1356;wire n1357;wire n1358;wire n1359;wire n1360;wire n1361;wire n1362;wire n1363;wire n1364;wire n1365;wire n1366;wire n1367;wire n1368;wire n1369;wire n1370;wire n1371;wire n1372;wire n1373;wire n1374;wire n1375;wire n1376;wire n1377;wire n1378;wire n1379;wire n1380;wire n1381;wire n1382;wire n1383;wire n1384;wire n1385;wire n1386;wire n1387;wire n1388;wire n1389;wire n1390;wire n1391;wire n1392;wire n1393;wire n1394;wire n1395;wire n1396;wire n1397;wire n1398;wire n1399;wire n1400;wire n1401;wire n1402;wire n1403;wire n1404;wire n1405;wire n1406;wire n1407;wire n1408;wire n1409;wire n1410;wire n1411;wire n1412;wire n1413;wire n1414;wire n1415;wire n1416;wire n1417;wire n1418;wire n1419;wire n1420;wire n1421;wire n1422;wire n1423;wire n1424;wire n1425;wire n1426;wire n1427;wire n1428;wire n1429;wire n1430;wire n1431;wire n1432;wire n1433;wire n1434;wire n1435;wire n1436;wire n1437;wire n1438;wire n1439;wire n1440;wire n1441;wire n1442;wire n1443;wire n1444;wire n1445;wire n1446;wire n1447;wire n1448;wire n1449;wire n1450;wire n1451;wire n1452;wire n1453;wire n1454;wire n1455;wire n1456;wire n1457;wire n1458;wire n1459;wire n1460;wire n1461;wire n1462;wire n1463;wire n1464;wire n1465;wire n1466;wire n1467;wire n1468;wire n1469;wire n1470;wire n1471;wire n1472;wire n1473;wire n1474;wire n1475;wire n1476;wire n1477;wire n1478;wire n1479;wire n1480;wire n1481;wire n1482;wire n1483;wire n1484;wire n1485;wire n1486;wire n1487;wire n1488;wire n1489;wire n1490;wire n1491;wire n1492;wire n1493;wire n1494;wire n1495;wire n1496;wire n1497;wire n1498;wire n1499;wire n1500;wire n1501;wire n1502;wire n1503;wire n1504;wire n1505;wire n1506;wire n1507;wire n1508;wire n1509;wire n1510;wire n1511;wire n1512;wire n1513;wire n1514;wire n1515;wire n1516;wire n1517;wire n1518;wire n1519;wire n1520;wire n1521;wire n1522;wire n1523;wire n1524;wire n1525;wire n1526;wire n1527;wire n1528;wire n1529;wire n1530;wire n1531;wire n1532;wire n1533;wire n1534;wire n1535;wire n1536;wire n1537;wire n1538;wire n1539;wire n1540;wire n1541;wire n1542;wire n1543;wire n1544;wire n1545;wire n1546;wire n1547;wire n1548;wire n1549;wire n1550;wire n1551;wire n1552;wire n1553;wire n1554;wire n1555;wire n1556;wire n1557;wire n1558;wire n1559;wire n1560;wire n1561;wire n1562;wire n1563;wire n1564;wire n1565;wire n1566;wire n1567;wire n1568;wire n1569;wire n1570;wire n1571;wire n1572;wire n1573;wire n1574;wire n1575;wire n1576;wire n1577;wire n1578;wire n1579;wire n1580;wire n1581;wire n1582;wire n1583;wire n1584;wire n1585;wire n1586;wire n1587;wire n1588;wire n1589;wire n1590;wire n1591;wire n1592;wire n1593;wire n1594;wire n1595;wire n1596;wire n1597;wire n1598;wire n1599;wire n1600;wire n1601;wire n1602;wire n1603;wire n1604;wire n1605;wire n1606;wire n1607;wire n1608;wire n1609;wire n1610;wire n1611;wire n1612;wire n1613;wire n1614;wire n1615;wire n1616;wire n1617;wire n1618;wire n1619;wire n1620;wire n1621;wire n1622;wire n1623;wire n1624;wire n1625;wire n1626;wire n1627;wire n1628;wire n1629;wire n1630;wire n1631;wire n1632;wire n1633;wire n1634;wire n1635;wire n1636;wire n1637;wire n1638;wire n1639;wire n1640;wire n1641;wire n1642;wire n1643;wire n1644;wire n1645;wire n1646;wire n1647;wire n1648;wire n1649;wire n1650;wire n1651;wire n1652;wire n1653;wire n1654;wire n1655;wire n1656;wire n1657;wire n1658;wire n1659;wire n1660;wire n1661;wire n1662;wire n1663;wire n1664;wire n1665;wire n1666;wire n1667;wire n1668;wire n1669;wire n1670;wire n1671;wire n1672;wire n1673;wire n1674;wire n1675;wire n1676;wire n1677;wire n1678;wire n1679;wire n1680;wire n1681;wire n1682;wire n1683;wire n1684;wire n1685;wire n1686;wire n1687;wire n1688;wire n1689;wire n1690;wire n1691;wire n1692;wire n1693;wire n1694;wire n1695;wire n1696;wire n1697;wire n1698;wire n1699;wire n1700;wire n1701;wire n1702;wire n1703;wire n1704;wire n1705;wire n1706;wire n1707;wire n1708;wire n1709;wire n1710;wire n1711;wire n1712;wire n1713;wire n1714;wire n1715;wire n1716;wire n1717;wire n1718;wire n1719;wire n1720;wire n1721;wire n1722;wire n1723;wire n1724;wire n1725;wire n1726;wire n1727;wire n1728;wire n1729;wire n1730;wire n1731;wire n1732;wire n1733;wire n1734;wire n1735;wire n1736;wire n1737;wire n1738;wire n1739;wire n1740;wire n1741;wire n1742;wire n1743;wire n1744;wire n1745;wire n1746;wire n1747;wire n1748;wire n1749;wire n1750;wire n1751;wire n1752;wire n1753;wire n1754;wire n1755;wire n1756;wire n1757;wire n1758;wire n1759;wire n1760;wire n1761;wire n1762;wire n1765;wire n1766;wire n1767;wire n1770;wire n1771;wire n1772;wire n1773;wire n1774;wire n1775;wire n1776;wire n1777;wire n1778;wire n1779;wire n1780;wire n1781;wire n1782;wire n1783;wire n1784;wire n1785;wire n1786;wire n1787;wire n1788;wire n1789;wire n1790;wire n1791;wire n1792;wire n1793;wire n1794;wire n1795;wire n1796;wire n1797;wire n1798;wire n1799;wire n1800;wire n1801;wire n1802;wire n1803;wire n1804;wire n1805;wire n1806;wire n1807;wire n1808;wire n1809;wire n1810;wire n1811;wire n1812;wire n1813;wire n1814;wire n1815;wire n1816;wire n1817;wire n1818;wire n1819;wire n1820;wire n1821;wire n1822;wire n1823;wire n1824;wire n1825;wire n1826;wire n1827;wire n1828;wire n1832;wire n1834;wire n1836;wire n1838;wire n1839;wire n1840;wire n1841;wire n1842;wire n1843;wire n1844;wire n1845;wire n1846;wire n1847;wire n1848;wire n1849;wire n1850;wire n1851;wire n1852;wire n1853;wire n1854;wire n1855;wire n1856;wire n1857;wire n1858;wire n1859;wire n1860;wire n1870;wire n1871;wire n1872;wire n1873;wire n1874;wire n1875;wire n1876;wire n1877;wire KeyWire_0_0;wire KeyWire_0_1;wire KeyWire_0_2;wire KeyWire_0_3;wire KeyWire_0_4;wire KeyWire_0_5;wire KeyWire_0_6;wire KeyWire_0_7;wire KeyWire_0_8;wire KeyWire_0_9;wire KeyWire_0_10;wire KeyWire_0_11;wire KeyWire_0_12;wire KeyWire_0_13;wire KeyWire_0_14;wire KeyWire_0_15;wire KeyWire_0_16;wire KeyWire_0_17;wire KeyWire_0_18;wire KeyWire_0_19;wire KeyWire_0_20;wire KeyWire_0_21;wire KeyWire_0_22;wire KeyWire_0_23;wire KeyWire_0_24;wire KeyWire_0_25;wire KeyWire_0_26;wire KeyWire_0_27;wire KeyWire_0_28;wire KeyWire_0_29;wire KeyWire_0_30;wire KeyWire_0_31;

  not
  g0
  (
    n34,
    n13
  );


  buf
  g1
  (
    n25,
    n18
  );


  not
  g2
  (
    n74,
    n12
  );


  not
  g3
  (
    n28,
    n7
  );


  not
  g4
  (
    n60,
    n10
  );


  not
  g5
  (
    n70,
    n2
  );


  not
  g6
  (
    n53,
    n13
  );


  not
  g7
  (
    n45,
    n15
  );


  buf
  g8
  (
    n56,
    n12
  );


  buf
  g9
  (
    n85,
    n6
  );


  buf
  g10
  (
    n75,
    n9
  );


  not
  g11
  (
    n95,
    n10
  );


  buf
  g12
  (
    n24,
    n19
  );


  buf
  g13
  (
    n73,
    n11
  );


  buf
  g14
  (
    n30,
    n18
  );


  buf
  g15
  (
    n23,
    n8
  );


  buf
  g16
  (
    n67,
    n5
  );


  not
  g17
  (
    n29,
    n20
  );


  buf
  g18
  (
    n31,
    n7
  );


  not
  g19
  (
    n22,
    n16
  );


  not
  g20
  (
    n97,
    n21
  );


  not
  g21
  (
    n82,
    n2
  );


  buf
  g22
  (
    n26,
    n20
  );


  buf
  g23
  (
    n61,
    n5
  );


  not
  g24
  (
    n79,
    n2
  );


  not
  g25
  (
    n41,
    n11
  );


  not
  g26
  (
    n47,
    n11
  );


  buf
  g27
  (
    n101,
    n9
  );


  buf
  g28
  (
    n68,
    n8
  );


  buf
  g29
  (
    n62,
    n8
  );


  not
  g30
  (
    n104,
    n20
  );


  not
  g31
  (
    n98,
    n1
  );


  buf
  g32
  (
    n99,
    n6
  );


  buf
  g33
  (
    n92,
    n18
  );


  buf
  g34
  (
    n46,
    n12
  );


  buf
  g35
  (
    n54,
    n1
  );


  buf
  g36
  (
    n80,
    n15
  );


  not
  g37
  (
    n81,
    n8
  );


  not
  g38
  (
    n93,
    n21
  );


  not
  g39
  (
    n58,
    n5
  );


  buf
  g40
  (
    n43,
    n19
  );


  buf
  g41
  (
    n39,
    n7
  );


  buf
  g42
  (
    n94,
    n14
  );


  buf
  g43
  (
    n42,
    n21
  );


  buf
  g44
  (
    n71,
    n10
  );


  not
  g45
  (
    n69,
    n6
  );


  buf
  g46
  (
    n105,
    n14
  );


  not
  g47
  (
    n51,
    n4
  );


  not
  g48
  (
    n91,
    n14
  );


  buf
  g49
  (
    n90,
    n20
  );


  not
  g50
  (
    n63,
    n17
  );


  buf
  g51
  (
    n76,
    n13
  );


  not
  g52
  (
    n40,
    n11
  );


  not
  g53
  (
    n37,
    n3
  );


  not
  g54
  (
    n100,
    n7
  );


  buf
  g55
  (
    n66,
    n2
  );


  buf
  g56
  (
    n55,
    n18
  );


  not
  g57
  (
    n86,
    n16
  );


  not
  g58
  (
    n35,
    n1
  );


  not
  g59
  (
    n88,
    n14
  );


  not
  g60
  (
    n48,
    n4
  );


  not
  g61
  (
    n64,
    n19
  );


  buf
  g62
  (
    n44,
    n17
  );


  buf
  g63
  (
    n52,
    n9
  );


  not
  g64
  (
    n102,
    n3
  );


  not
  g65
  (
    n49,
    n6
  );


  not
  g66
  (
    n78,
    n4
  );


  not
  g67
  (
    n57,
    n5
  );


  not
  g68
  (
    n38,
    n13
  );


  buf
  g69
  (
    n89,
    n21
  );


  buf
  g70
  (
    n50,
    n12
  );


  not
  g71
  (
    n87,
    n4
  );


  not
  g72
  (
    n36,
    n9
  );


  buf
  g73
  (
    n84,
    n1
  );


  not
  g74
  (
    n33,
    n19
  );


  not
  g75
  (
    n65,
    n16
  );


  buf
  g76
  (
    n103,
    n15
  );


  not
  g77
  (
    n77,
    n15
  );


  buf
  g78
  (
    n72,
    n17
  );


  buf
  g79
  (
    n59,
    n3
  );


  buf
  g80
  (
    n83,
    n16
  );


  not
  g81
  (
    n32,
    n10
  );


  buf
  g82
  (
    n96,
    n17
  );


  buf
  g83
  (
    n27,
    n3
  );


  not
  g84
  (
    n205,
    n66
  );


  not
  g85
  (
    n268,
    n62
  );


  not
  g86
  (
    n400,
    n38
  );


  buf
  g87
  (
    n267,
    n51
  );


  buf
  g88
  (
    n375,
    n65
  );


  buf
  g89
  (
    n366,
    n55
  );


  not
  g90
  (
    n154,
    n44
  );


  buf
  g91
  (
    n197,
    n72
  );


  buf
  g92
  (
    n296,
    n31
  );


  not
  g93
  (
    n419,
    n41
  );


  buf
  g94
  (
    n143,
    n42
  );


  not
  g95
  (
    n283,
    n28
  );


  buf
  g96
  (
    n374,
    n80
  );


  buf
  g97
  (
    n247,
    n28
  );


  buf
  g98
  (
    n149,
    n51
  );


  buf
  g99
  (
    n165,
    n98
  );


  buf
  g100
  (
    n114,
    n58
  );


  buf
  g101
  (
    n210,
    n72
  );


  buf
  g102
  (
    n233,
    n103
  );


  buf
  g103
  (
    n382,
    n76
  );


  buf
  g104
  (
    n300,
    n24
  );


  not
  g105
  (
    n250,
    n42
  );


  not
  g106
  (
    n365,
    n44
  );


  buf
  g107
  (
    n322,
    n50
  );


  not
  g108
  (
    n152,
    n48
  );


  buf
  g109
  (
    n379,
    n62
  );


  not
  g110
  (
    n129,
    n72
  );


  buf
  g111
  (
    n301,
    n54
  );


  buf
  g112
  (
    n336,
    n25
  );


  not
  g113
  (
    n175,
    n64
  );


  not
  g114
  (
    n356,
    n83
  );


  buf
  g115
  (
    n307,
    n52
  );


  not
  g116
  (
    n272,
    n91
  );


  not
  g117
  (
    n237,
    n60
  );


  buf
  g118
  (
    n398,
    n27
  );


  not
  g119
  (
    n119,
    n29
  );


  not
  g120
  (
    n281,
    n47
  );


  buf
  g121
  (
    n255,
    n61
  );


  not
  g122
  (
    n163,
    n105
  );


  buf
  g123
  (
    n196,
    n103
  );


  not
  g124
  (
    n418,
    n56
  );


  not
  g125
  (
    n302,
    n55
  );


  buf
  g126
  (
    n167,
    n98
  );


  not
  g127
  (
    n406,
    n98
  );


  not
  g128
  (
    n133,
    n37
  );


  not
  g129
  (
    n311,
    n82
  );


  not
  g130
  (
    n270,
    n41
  );


  not
  g131
  (
    n137,
    n42
  );


  buf
  g132
  (
    n121,
    n83
  );


  not
  g133
  (
    n367,
    n96
  );


  not
  g134
  (
    n433,
    n40
  );


  buf
  g135
  (
    n333,
    n61
  );


  not
  g136
  (
    n229,
    n91
  );


  buf
  g137
  (
    n355,
    n64
  );


  buf
  g138
  (
    n256,
    n36
  );


  not
  g139
  (
    n377,
    n82
  );


  not
  g140
  (
    n188,
    n65
  );


  not
  g141
  (
    n420,
    n80
  );


  not
  g142
  (
    n343,
    n57
  );


  buf
  g143
  (
    n181,
    n104
  );


  buf
  g144
  (
    n203,
    n94
  );


  not
  g145
  (
    n341,
    n48
  );


  not
  g146
  (
    n440,
    n31
  );


  not
  g147
  (
    n139,
    n68
  );


  not
  g148
  (
    n220,
    n96
  );


  buf
  g149
  (
    n293,
    n39
  );


  buf
  g150
  (
    n245,
    n99
  );


  not
  g151
  (
    n128,
    n66
  );


  buf
  g152
  (
    n146,
    n30
  );


  not
  g153
  (
    n212,
    n23
  );


  buf
  g154
  (
    n224,
    n73
  );


  buf
  g155
  (
    n190,
    n68
  );


  buf
  g156
  (
    n193,
    n60
  );


  not
  g157
  (
    n314,
    n49
  );


  buf
  g158
  (
    n135,
    n87
  );


  buf
  g159
  (
    n240,
    n85
  );


  buf
  g160
  (
    n364,
    n93
  );


  buf
  g161
  (
    n393,
    n67
  );


  buf
  g162
  (
    n425,
    n99
  );


  buf
  g163
  (
    n394,
    n22
  );


  not
  g164
  (
    n306,
    n97
  );


  buf
  g165
  (
    n123,
    n35
  );


  buf
  g166
  (
    n185,
    n77
  );


  not
  g167
  (
    n169,
    n93
  );


  buf
  g168
  (
    n414,
    n98
  );


  buf
  g169
  (
    n430,
    n52
  );


  not
  g170
  (
    n148,
    n34
  );


  not
  g171
  (
    n417,
    n57
  );


  buf
  g172
  (
    n428,
    n23
  );


  not
  g173
  (
    n352,
    n45
  );


  buf
  g174
  (
    n147,
    n73
  );


  buf
  g175
  (
    n178,
    n84
  );


  not
  g176
  (
    n184,
    n36
  );


  not
  g177
  (
    n186,
    n86
  );


  buf
  g178
  (
    n415,
    n32
  );


  not
  g179
  (
    n346,
    n65
  );


  not
  g180
  (
    n126,
    n100
  );


  buf
  g181
  (
    n136,
    n66
  );


  not
  g182
  (
    n290,
    n91
  );


  not
  g183
  (
    n401,
    n53
  );


  buf
  g184
  (
    n389,
    n74
  );


  buf
  g185
  (
    n357,
    n69
  );


  not
  g186
  (
    n264,
    n36
  );


  buf
  g187
  (
    n360,
    n53
  );


  buf
  g188
  (
    n218,
    n23
  );


  not
  g189
  (
    n432,
    n30
  );


  buf
  g190
  (
    n315,
    n74
  );


  buf
  g191
  (
    n313,
    n74
  );


  buf
  g192
  (
    n261,
    n38
  );


  buf
  g193
  (
    n381,
    n78
  );


  not
  g194
  (
    n338,
    n29
  );


  buf
  g195
  (
    KeyWire_0_25,
    n40
  );


  not
  g196
  (
    n187,
    n32
  );


  buf
  g197
  (
    n402,
    n82
  );


  not
  g198
  (
    n239,
    n87
  );


  not
  g199
  (
    n160,
    n55
  );


  not
  g200
  (
    n124,
    n77
  );


  not
  g201
  (
    n208,
    n25
  );


  buf
  g202
  (
    n209,
    n75
  );


  not
  g203
  (
    n423,
    n35
  );


  buf
  g204
  (
    n330,
    n32
  );


  not
  g205
  (
    n429,
    n48
  );


  buf
  g206
  (
    n319,
    n27
  );


  not
  g207
  (
    n287,
    n101
  );


  not
  g208
  (
    n370,
    n104
  );


  buf
  g209
  (
    n257,
    n49
  );


  buf
  g210
  (
    n326,
    n33
  );


  buf
  g211
  (
    n383,
    n88
  );


  not
  g212
  (
    n127,
    n54
  );


  not
  g213
  (
    n408,
    n75
  );


  not
  g214
  (
    n110,
    n43
  );


  not
  g215
  (
    n199,
    n40
  );


  buf
  g216
  (
    n201,
    n34
  );


  not
  g217
  (
    n384,
    n67
  );


  buf
  g218
  (
    n426,
    n56
  );


  not
  g219
  (
    n111,
    n100
  );


  not
  g220
  (
    n373,
    n79
  );


  buf
  g221
  (
    n335,
    n67
  );


  not
  g222
  (
    n282,
    n57
  );


  buf
  g223
  (
    n309,
    n46
  );


  buf
  g224
  (
    n176,
    n49
  );


  not
  g225
  (
    n280,
    n95
  );


  buf
  g226
  (
    n427,
    n94
  );


  not
  g227
  (
    n159,
    n96
  );


  buf
  g228
  (
    n243,
    n103
  );


  buf
  g229
  (
    n223,
    n59
  );


  buf
  g230
  (
    n441,
    n73
  );


  buf
  g231
  (
    n174,
    n46
  );


  not
  g232
  (
    n266,
    n77
  );


  not
  g233
  (
    n286,
    n81
  );


  not
  g234
  (
    n436,
    n26
  );


  not
  g235
  (
    n363,
    n89
  );


  buf
  g236
  (
    n388,
    n88
  );


  buf
  g237
  (
    n321,
    n56
  );


  not
  g238
  (
    n327,
    n78
  );


  not
  g239
  (
    n337,
    n38
  );


  buf
  g240
  (
    n359,
    n39
  );


  not
  g241
  (
    n182,
    n63
  );


  not
  g242
  (
    n396,
    n73
  );


  not
  g243
  (
    n351,
    n95
  );


  not
  g244
  (
    n171,
    n78
  );


  buf
  g245
  (
    n299,
    n58
  );


  not
  g246
  (
    n155,
    n28
  );


  not
  g247
  (
    n242,
    n102
  );


  buf
  g248
  (
    n112,
    n23
  );


  not
  g249
  (
    n380,
    n83
  );


  buf
  g250
  (
    n231,
    n45
  );


  buf
  g251
  (
    n348,
    n69
  );


  buf
  g252
  (
    n323,
    n99
  );


  buf
  g253
  (
    n254,
    n47
  );


  not
  g254
  (
    n397,
    n29
  );


  not
  g255
  (
    n342,
    n36
  );


  buf
  g256
  (
    n362,
    n86
  );


  not
  g257
  (
    n260,
    n61
  );


  buf
  g258
  (
    n118,
    n39
  );


  not
  g259
  (
    n130,
    n51
  );


  buf
  g260
  (
    n291,
    n35
  );


  buf
  g261
  (
    n158,
    n89
  );


  buf
  g262
  (
    n213,
    n37
  );


  buf
  g263
  (
    n226,
    n45
  );


  not
  g264
  (
    n200,
    n69
  );


  buf
  g265
  (
    n308,
    n79
  );


  buf
  g266
  (
    n344,
    n62
  );


  not
  g267
  (
    n222,
    n59
  );


  not
  g268
  (
    n115,
    n96
  );


  buf
  g269
  (
    n437,
    n29
  );


  buf
  g270
  (
    n145,
    n49
  );


  not
  g271
  (
    n312,
    n71
  );


  buf
  g272
  (
    n198,
    n105
  );


  buf
  g273
  (
    n204,
    n63
  );


  not
  g274
  (
    n334,
    n54
  );


  buf
  g275
  (
    n404,
    n52
  );


  not
  g276
  (
    n211,
    n71
  );


  buf
  g277
  (
    KeyWire_0_24,
    n45
  );


  not
  g278
  (
    n320,
    n79
  );


  not
  g279
  (
    n392,
    n67
  );


  not
  g280
  (
    n332,
    n85
  );


  not
  g281
  (
    n368,
    n58
  );


  not
  g282
  (
    n316,
    n94
  );


  not
  g283
  (
    n206,
    n101
  );


  not
  g284
  (
    n354,
    n74
  );


  buf
  g285
  (
    n331,
    n95
  );


  buf
  g286
  (
    n422,
    n70
  );


  buf
  g287
  (
    n304,
    n55
  );


  not
  g288
  (
    n350,
    n24
  );


  buf
  g289
  (
    n151,
    n48
  );


  buf
  g290
  (
    n405,
    n81
  );


  buf
  g291
  (
    KeyWire_0_7,
    n31
  );


  not
  g292
  (
    n271,
    n83
  );


  not
  g293
  (
    n219,
    n85
  );


  not
  g294
  (
    n288,
    n47
  );


  buf
  g295
  (
    n376,
    n38
  );


  not
  g296
  (
    n225,
    n53
  );


  not
  g297
  (
    n217,
    n46
  );


  buf
  g298
  (
    n325,
    n104
  );


  buf
  g299
  (
    n173,
    n103
  );


  not
  g300
  (
    KeyWire_0_13,
    n79
  );


  buf
  g301
  (
    n191,
    n24
  );


  buf
  g302
  (
    n244,
    n63
  );


  buf
  g303
  (
    n345,
    n31
  );


  not
  g304
  (
    n395,
    n60
  );


  not
  g305
  (
    n117,
    n84
  );


  not
  g306
  (
    n305,
    n26
  );


  not
  g307
  (
    n284,
    n30
  );


  buf
  g308
  (
    n340,
    n84
  );


  buf
  g309
  (
    n116,
    n70
  );


  not
  g310
  (
    n353,
    n47
  );


  buf
  g311
  (
    n277,
    n70
  );


  buf
  g312
  (
    n434,
    n90
  );


  buf
  g313
  (
    n387,
    n27
  );


  buf
  g314
  (
    n416,
    n102
  );


  not
  g315
  (
    n234,
    n92
  );


  not
  g316
  (
    n221,
    n22
  );


  buf
  g317
  (
    n236,
    n90
  );


  buf
  g318
  (
    n391,
    n76
  );


  buf
  g319
  (
    n358,
    n43
  );


  buf
  g320
  (
    n258,
    n68
  );


  buf
  g321
  (
    n131,
    n58
  );


  buf
  g322
  (
    n372,
    n87
  );


  not
  g323
  (
    n259,
    n88
  );


  not
  g324
  (
    n235,
    n30
  );


  buf
  g325
  (
    n246,
    n90
  );


  not
  g326
  (
    n278,
    n62
  );


  not
  g327
  (
    n141,
    n80
  );


  buf
  g328
  (
    n144,
    n86
  );


  buf
  g329
  (
    n279,
    n84
  );


  buf
  g330
  (
    n339,
    n92
  );


  not
  g331
  (
    n399,
    n37
  );


  not
  g332
  (
    n202,
    n92
  );


  buf
  g333
  (
    n216,
    n34
  );


  buf
  g334
  (
    KeyWire_0_19,
    n81
  );


  buf
  g335
  (
    n439,
    n60
  );


  not
  g336
  (
    n120,
    n34
  );


  buf
  g337
  (
    n294,
    n25
  );


  buf
  g338
  (
    n195,
    n25
  );


  buf
  g339
  (
    n410,
    n22
  );


  buf
  g340
  (
    n232,
    n100
  );


  buf
  g341
  (
    n156,
    n41
  );


  not
  g342
  (
    n407,
    n77
  );


  buf
  g343
  (
    n248,
    n50
  );


  buf
  g344
  (
    n292,
    n80
  );


  not
  g345
  (
    n142,
    n102
  );


  buf
  g346
  (
    n378,
    n41
  );


  not
  g347
  (
    n324,
    n37
  );


  buf
  g348
  (
    n252,
    n69
  );


  buf
  g349
  (
    n253,
    n24
  );


  not
  g350
  (
    n262,
    n75
  );


  not
  g351
  (
    n122,
    n85
  );


  not
  g352
  (
    n435,
    n76
  );


  not
  g353
  (
    n207,
    n90
  );


  not
  g354
  (
    n297,
    n66
  );


  buf
  g355
  (
    n134,
    n75
  );


  not
  g356
  (
    n125,
    n26
  );


  not
  g357
  (
    n361,
    n105
  );


  not
  g358
  (
    n214,
    n71
  );


  not
  g359
  (
    n386,
    n22
  );


  not
  g360
  (
    n228,
    n88
  );


  buf
  g361
  (
    n317,
    n52
  );


  buf
  g362
  (
    n157,
    n101
  );


  buf
  g363
  (
    n192,
    n94
  );


  buf
  g364
  (
    n150,
    n46
  );


  not
  g365
  (
    n230,
    n101
  );


  buf
  g366
  (
    n347,
    n33
  );


  buf
  g367
  (
    n349,
    n78
  );


  not
  g368
  (
    n172,
    n43
  );


  buf
  g369
  (
    n285,
    n105
  );


  buf
  g370
  (
    n164,
    n93
  );


  buf
  g371
  (
    n166,
    n56
  );


  buf
  g372
  (
    KeyWire_0_9,
    n81
  );


  not
  g373
  (
    n295,
    n64
  );


  buf
  g374
  (
    n413,
    n70
  );


  not
  g375
  (
    n241,
    n97
  );


  buf
  g376
  (
    n298,
    n50
  );


  buf
  g377
  (
    n303,
    n61
  );


  buf
  g378
  (
    n183,
    n42
  );


  not
  g379
  (
    n273,
    n57
  );


  buf
  g380
  (
    n215,
    n91
  );


  not
  g381
  (
    n138,
    n44
  );


  not
  g382
  (
    n412,
    n82
  );


  not
  g383
  (
    n106,
    n89
  );


  not
  g384
  (
    n310,
    n64
  );


  not
  g385
  (
    n329,
    n65
  );


  not
  g386
  (
    n276,
    n32
  );


  buf
  g387
  (
    n371,
    n39
  );


  buf
  g388
  (
    n265,
    n43
  );


  not
  g389
  (
    n161,
    n59
  );


  not
  g390
  (
    n179,
    n50
  );


  not
  g391
  (
    n263,
    n26
  );


  not
  g392
  (
    n274,
    n51
  );


  not
  g393
  (
    n227,
    n27
  );


  not
  g394
  (
    n162,
    n68
  );


  buf
  g395
  (
    n140,
    n95
  );


  not
  g396
  (
    n113,
    n35
  );


  buf
  g397
  (
    n249,
    n97
  );


  buf
  g398
  (
    n107,
    n76
  );


  not
  g399
  (
    n251,
    n28
  );


  buf
  g400
  (
    n180,
    n93
  );


  not
  g401
  (
    n238,
    n92
  );


  buf
  g402
  (
    n108,
    n72
  );


  not
  g403
  (
    n168,
    n99
  );


  buf
  g404
  (
    n194,
    n54
  );


  not
  g405
  (
    n421,
    n87
  );


  buf
  g406
  (
    n424,
    n53
  );


  not
  g407
  (
    n385,
    n33
  );


  buf
  g408
  (
    n328,
    n86
  );


  buf
  g409
  (
    n369,
    n102
  );


  buf
  g410
  (
    n269,
    n100
  );


  not
  g411
  (
    n431,
    n89
  );


  not
  g412
  (
    n403,
    n97
  );


  not
  g413
  (
    n289,
    n71
  );


  not
  g414
  (
    n318,
    n33
  );


  buf
  g415
  (
    n170,
    n63
  );


  buf
  g416
  (
    n438,
    n44
  );


  not
  g417
  (
    n177,
    n59
  );


  buf
  g418
  (
    n411,
    n40
  );


  buf
  g419
  (
    n109,
    n104
  );


  not
  g420
  (
    n668,
    n306
  );


  not
  g421
  (
    n589,
    n200
  );


  buf
  g422
  (
    n591,
    n131
  );


  buf
  g423
  (
    n597,
    n310
  );


  buf
  g424
  (
    n1147,
    n113
  );


  buf
  g425
  (
    n724,
    n263
  );


  not
  g426
  (
    n1076,
    n347
  );


  buf
  g427
  (
    n512,
    n136
  );


  not
  g428
  (
    n468,
    n160
  );


  buf
  g429
  (
    n836,
    n259
  );


  buf
  g430
  (
    n887,
    n191
  );


  buf
  g431
  (
    n443,
    n151
  );


  not
  g432
  (
    n899,
    n303
  );


  not
  g433
  (
    n588,
    n332
  );


  buf
  g434
  (
    n647,
    n171
  );


  buf
  g435
  (
    n545,
    n158
  );


  not
  g436
  (
    n1159,
    n121
  );


  buf
  g437
  (
    n942,
    n329
  );


  not
  g438
  (
    n705,
    n290
  );


  buf
  g439
  (
    n854,
    n210
  );


  buf
  g440
  (
    n489,
    n140
  );


  buf
  g441
  (
    n447,
    n308
  );


  buf
  g442
  (
    n699,
    n235
  );


  buf
  g443
  (
    n1143,
    n112
  );


  buf
  g444
  (
    n509,
    n108
  );


  buf
  g445
  (
    n1099,
    n166
  );


  buf
  g446
  (
    n1131,
    n208
  );


  not
  g447
  (
    n676,
    n301
  );


  not
  g448
  (
    n531,
    n213
  );


  buf
  g449
  (
    KeyWire_0_10,
    n318
  );


  not
  g450
  (
    n637,
    n256
  );


  buf
  g451
  (
    n516,
    n140
  );


  buf
  g452
  (
    n846,
    n354
  );


  not
  g453
  (
    n873,
    n193
  );


  not
  g454
  (
    n1108,
    n189
  );


  buf
  g455
  (
    n469,
    n273
  );


  not
  g456
  (
    n551,
    n164
  );


  not
  g457
  (
    n1187,
    n358
  );


  buf
  g458
  (
    n1141,
    n302
  );


  buf
  g459
  (
    n920,
    n312
  );


  buf
  g460
  (
    n778,
    n221
  );


  not
  g461
  (
    n777,
    n153
  );


  not
  g462
  (
    n783,
    n360
  );


  not
  g463
  (
    n529,
    n146
  );


  buf
  g464
  (
    n1006,
    n128
  );


  buf
  g465
  (
    n634,
    n356
  );


  buf
  g466
  (
    n850,
    n164
  );


  buf
  g467
  (
    n1120,
    n173
  );


  not
  g468
  (
    n968,
    n140
  );


  not
  g469
  (
    n871,
    n204
  );


  not
  g470
  (
    n658,
    n267
  );


  buf
  g471
  (
    n602,
    n345
  );


  buf
  g472
  (
    n1093,
    n271
  );


  buf
  g473
  (
    n1157,
    n305
  );


  not
  g474
  (
    n595,
    n334
  );


  buf
  g475
  (
    n1043,
    n340
  );


  buf
  g476
  (
    n851,
    n331
  );


  buf
  g477
  (
    n648,
    n177
  );


  buf
  g478
  (
    n1189,
    n181
  );


  buf
  g479
  (
    n1045,
    n353
  );


  not
  g480
  (
    n744,
    n268
  );


  not
  g481
  (
    n1121,
    n286
  );


  buf
  g482
  (
    KeyWire_0_18,
    n293
  );


  not
  g483
  (
    n1123,
    n286
  );


  buf
  g484
  (
    n454,
    n135
  );


  not
  g485
  (
    n761,
    n219
  );


  buf
  g486
  (
    n1130,
    n267
  );


  buf
  g487
  (
    n548,
    n315
  );


  buf
  g488
  (
    n574,
    n284
  );


  not
  g489
  (
    n1126,
    n333
  );


  not
  g490
  (
    n692,
    n266
  );


  not
  g491
  (
    n651,
    n342
  );


  not
  g492
  (
    n797,
    n161
  );


  not
  g493
  (
    n1184,
    n208
  );


  buf
  g494
  (
    n750,
    n182
  );


  not
  g495
  (
    n896,
    n277
  );


  not
  g496
  (
    n502,
    n168
  );


  buf
  g497
  (
    n931,
    n138
  );


  not
  g498
  (
    n1094,
    n162
  );


  not
  g499
  (
    n1047,
    n137
  );


  not
  g500
  (
    n1098,
    n299
  );


  buf
  g501
  (
    n1145,
    n117
  );


  buf
  g502
  (
    n1183,
    n197
  );


  buf
  g503
  (
    n990,
    n296
  );


  not
  g504
  (
    n732,
    n133
  );


  buf
  g505
  (
    n1051,
    n239
  );


  not
  g506
  (
    n770,
    n213
  );


  not
  g507
  (
    n837,
    n117
  );


  not
  g508
  (
    n528,
    n289
  );


  buf
  g509
  (
    n845,
    n204
  );


  buf
  g510
  (
    n1046,
    n337
  );


  buf
  g511
  (
    n474,
    n236
  );


  not
  g512
  (
    n1092,
    n226
  );


  buf
  g513
  (
    n511,
    n198
  );


  not
  g514
  (
    n814,
    n176
  );


  not
  g515
  (
    n908,
    n217
  );


  not
  g516
  (
    n784,
    n108
  );


  not
  g517
  (
    n1029,
    n296
  );


  buf
  g518
  (
    n976,
    n309
  );


  buf
  g519
  (
    n1056,
    n301
  );


  buf
  g520
  (
    n576,
    n225
  );


  buf
  g521
  (
    n518,
    n308
  );


  buf
  g522
  (
    n773,
    n196
  );


  not
  g523
  (
    n568,
    n255
  );


  buf
  g524
  (
    n944,
    n150
  );


  buf
  g525
  (
    n563,
    n352
  );


  buf
  g526
  (
    n720,
    n178
  );


  not
  g527
  (
    n1127,
    n191
  );


  not
  g528
  (
    n1146,
    n324
  );


  not
  g529
  (
    n593,
    n323
  );


  buf
  g530
  (
    n752,
    n264
  );


  not
  g531
  (
    n505,
    n171
  );


  not
  g532
  (
    n570,
    n262
  );


  buf
  g533
  (
    n907,
    n352
  );


  buf
  g534
  (
    n754,
    n238
  );


  buf
  g535
  (
    n1175,
    n291
  );


  not
  g536
  (
    n935,
    n166
  );


  buf
  g537
  (
    n1200,
    n257
  );


  buf
  g538
  (
    n741,
    n300
  );


  not
  g539
  (
    n904,
    n304
  );


  not
  g540
  (
    n624,
    n323
  );


  buf
  g541
  (
    n987,
    n261
  );


  buf
  g542
  (
    n1133,
    n232
  );


  not
  g543
  (
    n849,
    n305
  );


  not
  g544
  (
    n1173,
    n242
  );


  buf
  g545
  (
    n582,
    n298
  );


  not
  g546
  (
    n1162,
    n239
  );


  buf
  g547
  (
    n456,
    n194
  );


  not
  g548
  (
    n1185,
    n355
  );


  buf
  g549
  (
    n1097,
    n193
  );


  not
  g550
  (
    n1195,
    n199
  );


  buf
  g551
  (
    n486,
    n362
  );


  buf
  g552
  (
    n632,
    n178
  );


  not
  g553
  (
    n515,
    n175
  );


  buf
  g554
  (
    n800,
    n280
  );


  not
  g555
  (
    n1030,
    n202
  );


  not
  g556
  (
    KeyWire_0_16,
    n347
  );


  not
  g557
  (
    n975,
    n317
  );


  buf
  g558
  (
    n524,
    n255
  );


  not
  g559
  (
    n1049,
    n240
  );


  not
  g560
  (
    n612,
    n163
  );


  not
  g561
  (
    n1070,
    n176
  );


  buf
  g562
  (
    n678,
    n129
  );


  not
  g563
  (
    n606,
    n163
  );


  buf
  g564
  (
    n1148,
    n327
  );


  not
  g565
  (
    n1101,
    n109
  );


  buf
  g566
  (
    n611,
    n336
  );


  buf
  g567
  (
    n644,
    n120
  );


  buf
  g568
  (
    n491,
    n225
  );


  not
  g569
  (
    n599,
    n358
  );


  buf
  g570
  (
    n946,
    n264
  );


  not
  g571
  (
    n954,
    n135
  );


  buf
  g572
  (
    n922,
    n343
  );


  not
  g573
  (
    n1027,
    n321
  );


  not
  g574
  (
    n831,
    n319
  );


  not
  g575
  (
    n1167,
    n120
  );


  buf
  g576
  (
    n808,
    n240
  );


  buf
  g577
  (
    n847,
    n288
  );


  not
  g578
  (
    n729,
    n270
  );


  buf
  g579
  (
    n554,
    n233
  );


  not
  g580
  (
    n675,
    n330
  );


  not
  g581
  (
    n542,
    n192
  );


  buf
  g582
  (
    n541,
    n343
  );


  buf
  g583
  (
    n680,
    n175
  );


  buf
  g584
  (
    n728,
    n290
  );


  not
  g585
  (
    n527,
    n291
  );


  not
  g586
  (
    n1038,
    n159
  );


  not
  g587
  (
    n959,
    n109
  );


  not
  g588
  (
    n1003,
    n234
  );


  buf
  g589
  (
    n943,
    n137
  );


  buf
  g590
  (
    n747,
    n355
  );


  buf
  g591
  (
    n1026,
    n348
  );


  buf
  g592
  (
    n779,
    n301
  );


  buf
  g593
  (
    n617,
    n297
  );


  not
  g594
  (
    n1144,
    n316
  );


  not
  g595
  (
    n817,
    n275
  );


  buf
  g596
  (
    n739,
    n201
  );


  not
  g597
  (
    n477,
    n138
  );


  buf
  g598
  (
    n1114,
    n235
  );


  not
  g599
  (
    n710,
    n354
  );


  not
  g600
  (
    n1122,
    n206
  );


  not
  g601
  (
    n1009,
    n115
  );


  not
  g602
  (
    n693,
    n302
  );


  not
  g603
  (
    n901,
    n113
  );


  not
  g604
  (
    n1171,
    n231
  );


  not
  g605
  (
    n1014,
    n118
  );


  not
  g606
  (
    n799,
    n352
  );


  not
  g607
  (
    n811,
    n111
  );


  not
  g608
  (
    n843,
    n272
  );


  not
  g609
  (
    n1087,
    n119
  );


  not
  g610
  (
    n1109,
    n251
  );


  buf
  g611
  (
    n857,
    n351
  );


  not
  g612
  (
    n452,
    n113
  );


  not
  g613
  (
    n835,
    n269
  );


  buf
  g614
  (
    n1128,
    n125
  );


  buf
  g615
  (
    n1165,
    n185
  );


  not
  g616
  (
    n1020,
    n241
  );


  not
  g617
  (
    n461,
    n232
  );


  not
  g618
  (
    n700,
    n111
  );


  buf
  g619
  (
    n885,
    n332
  );


  not
  g620
  (
    n913,
    n126
  );


  buf
  g621
  (
    n830,
    n215
  );


  not
  g622
  (
    n1037,
    n289
  );


  buf
  g623
  (
    n934,
    n341
  );


  not
  g624
  (
    n1188,
    n304
  );


  not
  g625
  (
    n757,
    n284
  );


  not
  g626
  (
    n497,
    n285
  );


  not
  g627
  (
    n1178,
    n252
  );


  not
  g628
  (
    n535,
    n351
  );


  buf
  g629
  (
    n685,
    n153
  );


  not
  g630
  (
    n1048,
    n327
  );


  buf
  g631
  (
    n905,
    n341
  );


  not
  g632
  (
    n1089,
    n197
  );


  not
  g633
  (
    n792,
    n312
  );


  buf
  g634
  (
    n838,
    n243
  );


  buf
  g635
  (
    n1163,
    n221
  );


  buf
  g636
  (
    n656,
    n138
  );


  not
  g637
  (
    n1090,
    n108
  );


  not
  g638
  (
    n763,
    n337
  );


  not
  g639
  (
    n467,
    n257
  );


  not
  g640
  (
    n1019,
    n337
  );


  buf
  g641
  (
    n458,
    n208
  );


  buf
  g642
  (
    n1179,
    n310
  );


  not
  g643
  (
    n457,
    n216
  );


  buf
  g644
  (
    n504,
    n212
  );


  not
  g645
  (
    n462,
    n199
  );


  buf
  g646
  (
    n892,
    n278
  );


  not
  g647
  (
    n1137,
    n186
  );


  not
  g648
  (
    n1103,
    n285
  );


  not
  g649
  (
    KeyWire_0_23,
    n349
  );


  not
  g650
  (
    n553,
    n320
  );


  not
  g651
  (
    n522,
    n258
  );


  buf
  g652
  (
    n966,
    n301
  );


  not
  g653
  (
    n1180,
    n145
  );


  not
  g654
  (
    n1129,
    n206
  );


  not
  g655
  (
    n787,
    n287
  );


  buf
  g656
  (
    n758,
    n172
  );


  not
  g657
  (
    n1060,
    n192
  );


  buf
  g658
  (
    n471,
    n288
  );


  buf
  g659
  (
    n1022,
    n123
  );


  not
  g660
  (
    n1008,
    n339
  );


  buf
  g661
  (
    n960,
    n209
  );


  buf
  g662
  (
    n840,
    n346
  );


  not
  g663
  (
    n781,
    n335
  );


  buf
  g664
  (
    n856,
    n320
  );


  not
  g665
  (
    n703,
    n241
  );


  not
  g666
  (
    n1149,
    n230
  );


  not
  g667
  (
    n823,
    n174
  );


  not
  g668
  (
    n1202,
    n114
  );


  not
  g669
  (
    n616,
    n294
  );


  buf
  g670
  (
    n697,
    n237
  );


  buf
  g671
  (
    n508,
    n247
  );


  not
  g672
  (
    n686,
    n208
  );


  buf
  g673
  (
    n894,
    n256
  );


  not
  g674
  (
    n532,
    n252
  );


  not
  g675
  (
    n601,
    n114
  );


  buf
  g676
  (
    n906,
    n284
  );


  not
  g677
  (
    n807,
    n250
  );


  not
  g678
  (
    n448,
    n181
  );


  not
  g679
  (
    n789,
    n115
  );


  not
  g680
  (
    n865,
    n203
  );


  buf
  g681
  (
    n451,
    n132
  );


  buf
  g682
  (
    n1018,
    n307
  );


  not
  g683
  (
    n577,
    n274
  );


  buf
  g684
  (
    n948,
    n232
  );


  not
  g685
  (
    n872,
    n144
  );


  not
  g686
  (
    n1136,
    n147
  );


  not
  g687
  (
    n957,
    n272
  );


  buf
  g688
  (
    n834,
    n259
  );


  not
  g689
  (
    n496,
    n177
  );


  not
  g690
  (
    n874,
    n250
  );


  not
  g691
  (
    n1044,
    n211
  );


  buf
  g692
  (
    n1084,
    n121
  );


  buf
  g693
  (
    n1035,
    n261
  );


  not
  g694
  (
    n1192,
    n227
  );


  not
  g695
  (
    n1106,
    n338
  );


  buf
  g696
  (
    n776,
    n250
  );


  not
  g697
  (
    n984,
    n216
  );


  not
  g698
  (
    n653,
    n150
  );


  not
  g699
  (
    n445,
    n248
  );


  not
  g700
  (
    n786,
    n336
  );


  not
  g701
  (
    n919,
    n106
  );


  not
  g702
  (
    n772,
    n307
  );


  not
  g703
  (
    n812,
    n241
  );


  buf
  g704
  (
    n449,
    n142
  );


  buf
  g705
  (
    n538,
    n119
  );


  not
  g706
  (
    n737,
    n126
  );


  buf
  g707
  (
    n855,
    n200
  );


  not
  g708
  (
    n891,
    n286
  );


  buf
  g709
  (
    n586,
    n128
  );


  not
  g710
  (
    n964,
    n188
  );


  not
  g711
  (
    n867,
    n303
  );


  not
  g712
  (
    n1031,
    n341
  );


  not
  g713
  (
    n650,
    n339
  );


  buf
  g714
  (
    n1140,
    n344
  );


  buf
  g715
  (
    n992,
    n127
  );


  buf
  g716
  (
    n1068,
    n295
  );


  not
  g717
  (
    n499,
    n192
  );


  not
  g718
  (
    n1013,
    n228
  );


  not
  g719
  (
    n805,
    n167
  );


  buf
  g720
  (
    n1096,
    n288
  );


  not
  g721
  (
    n667,
    n284
  );


  buf
  g722
  (
    n629,
    n281
  );


  not
  g723
  (
    n594,
    n339
  );


  buf
  g724
  (
    n1077,
    n265
  );


  not
  g725
  (
    n930,
    n155
  );


  buf
  g726
  (
    n950,
    n186
  );


  buf
  g727
  (
    n978,
    n238
  );


  not
  g728
  (
    n731,
    n346
  );


  not
  g729
  (
    n970,
    n223
  );


  not
  g730
  (
    n1052,
    n113
  );


  not
  g731
  (
    n1061,
    n299
  );


  buf
  g732
  (
    n900,
    n200
  );


  buf
  g733
  (
    n802,
    n190
  );


  buf
  g734
  (
    n484,
    n147
  );


  not
  g735
  (
    n498,
    n346
  );


  buf
  g736
  (
    n540,
    n157
  );


  not
  g737
  (
    n1155,
    n333
  );


  not
  g738
  (
    n478,
    n144
  );


  buf
  g739
  (
    n475,
    n362
  );


  not
  g740
  (
    n1023,
    n309
  );


  not
  g741
  (
    n719,
    n355
  );


  not
  g742
  (
    n1034,
    n343
  );


  not
  g743
  (
    n844,
    n203
  );


  not
  g744
  (
    n810,
    n353
  );


  not
  g745
  (
    n1086,
    n112
  );


  not
  g746
  (
    n1105,
    n165
  );


  buf
  g747
  (
    n620,
    n160
  );


  not
  g748
  (
    n819,
    n125
  );


  buf
  g749
  (
    n520,
    n355
  );


  buf
  g750
  (
    n734,
    n194
  );


  buf
  g751
  (
    n820,
    n328
  );


  not
  g752
  (
    n503,
    n172
  );


  buf
  g753
  (
    n898,
    n133
  );


  not
  g754
  (
    n670,
    n250
  );


  not
  g755
  (
    n1005,
    n224
  );


  not
  g756
  (
    n487,
    n203
  );


  not
  g757
  (
    n890,
    n271
  );


  buf
  g758
  (
    n1102,
    n287
  );


  not
  g759
  (
    n590,
    n265
  );


  not
  g760
  (
    n525,
    n320
  );


  not
  g761
  (
    n517,
    n249
  );


  not
  g762
  (
    n884,
    n281
  );


  not
  g763
  (
    n1091,
    n187
  );


  buf
  g764
  (
    n746,
    n253
  );


  not
  g765
  (
    n1062,
    n280
  );


  buf
  g766
  (
    n1071,
    n136
  );


  buf
  g767
  (
    n751,
    n329
  );


  not
  g768
  (
    n941,
    n314
  );


  not
  g769
  (
    n1194,
    n181
  );


  buf
  g770
  (
    n936,
    n112
  );


  buf
  g771
  (
    n888,
    n156
  );


  buf
  g772
  (
    n1063,
    n340
  );


  buf
  g773
  (
    n619,
    n344
  );


  buf
  g774
  (
    n730,
    n164
  );


  not
  g775
  (
    n863,
    n260
  );


  buf
  g776
  (
    n483,
    n190
  );


  buf
  g777
  (
    n659,
    n177
  );


  not
  g778
  (
    n1169,
    n293
  );


  buf
  g779
  (
    n543,
    n217
  );


  buf
  g780
  (
    n771,
    n191
  );


  not
  g781
  (
    n833,
    n175
  );


  buf
  g782
  (
    n839,
    n214
  );


  not
  g783
  (
    n1115,
    n155
  );


  buf
  g784
  (
    n708,
    n249
  );


  buf
  g785
  (
    n613,
    n260
  );


  not
  g786
  (
    n1156,
    n183
  );


  buf
  g787
  (
    n565,
    n319
  );


  not
  g788
  (
    n743,
    n325
  );


  buf
  g789
  (
    n560,
    n261
  );


  not
  g790
  (
    n442,
    n328
  );


  not
  g791
  (
    n1118,
    n254
  );


  buf
  g792
  (
    n972,
    n142
  );


  not
  g793
  (
    n1033,
    n264
  );


  buf
  g794
  (
    n640,
    n189
  );


  buf
  g795
  (
    n1197,
    n265
  );


  not
  g796
  (
    n493,
    n139
  );


  buf
  g797
  (
    n996,
    n186
  );


  not
  g798
  (
    n717,
    n158
  );


  buf
  g799
  (
    n547,
    n207
  );


  not
  g800
  (
    n463,
    n202
  );


  not
  g801
  (
    n596,
    n153
  );


  not
  g802
  (
    n610,
    n244
  );


  not
  g803
  (
    n635,
    n312
  );


  buf
  g804
  (
    n450,
    n256
  );


  not
  g805
  (
    n740,
    n118
  );


  not
  g806
  (
    n501,
    n279
  );


  not
  g807
  (
    n459,
    n334
  );


  not
  g808
  (
    n1053,
    n237
  );


  not
  g809
  (
    n886,
    n108
  );


  not
  g810
  (
    n562,
    n349
  );


  not
  g811
  (
    n1191,
    n169
  );


  buf
  g812
  (
    n997,
    n145
  );


  buf
  g813
  (
    n915,
    n221
  );


  buf
  g814
  (
    n782,
    n295
  );


  buf
  g815
  (
    n572,
    n176
  );


  buf
  g816
  (
    n1111,
    n220
  );


  buf
  g817
  (
    n721,
    n294
  );


  not
  g818
  (
    n969,
    n363
  );


  buf
  g819
  (
    n1001,
    n257
  );


  not
  g820
  (
    n1186,
    n185
  );


  not
  g821
  (
    n1050,
    n201
  );


  buf
  g822
  (
    n603,
    n130
  );


  buf
  g823
  (
    n1073,
    n213
  );


  buf
  g824
  (
    n566,
    n205
  );


  not
  g825
  (
    n626,
    n175
  );


  not
  g826
  (
    n706,
    n358
  );


  not
  g827
  (
    n861,
    n222
  );


  buf
  g828
  (
    n952,
    n363
  );


  not
  g829
  (
    n1107,
    n283
  );


  buf
  g830
  (
    n608,
    n145
  );


  buf
  g831
  (
    n587,
    n246
  );


  not
  g832
  (
    n1153,
    n351
  );


  not
  g833
  (
    n689,
    n281
  );


  buf
  g834
  (
    n993,
    n274
  );


  buf
  g835
  (
    n985,
    n265
  );


  not
  g836
  (
    n928,
    n193
  );


  not
  g837
  (
    n924,
    n139
  );


  not
  g838
  (
    n711,
    n179
  );


  not
  g839
  (
    n774,
    n141
  );


  not
  g840
  (
    KeyWire_0_0,
    n111
  );


  not
  g841
  (
    n694,
    n173
  );


  buf
  g842
  (
    n666,
    n115
  );


  buf
  g843
  (
    n630,
    n107
  );


  not
  g844
  (
    n536,
    n279
  );


  buf
  g845
  (
    n466,
    n328
  );


  not
  g846
  (
    n1088,
    n110
  );


  buf
  g847
  (
    n963,
    n215
  );


  buf
  g848
  (
    n983,
    n306
  );


  buf
  g849
  (
    n982,
    n174
  );


  not
  g850
  (
    n657,
    n318
  );


  buf
  g851
  (
    n687,
    n152
  );


  buf
  g852
  (
    n876,
    n170
  );


  buf
  g853
  (
    n583,
    n304
  );


  buf
  g854
  (
    n1203,
    n167
  );


  buf
  g855
  (
    n679,
    n172
  );


  not
  g856
  (
    n490,
    n136
  );


  buf
  g857
  (
    n848,
    n122
  );


  buf
  g858
  (
    n625,
    n318
  );


  not
  g859
  (
    n615,
    n152
  );


  buf
  g860
  (
    n600,
    n141
  );


  buf
  g861
  (
    n655,
    n123
  );


  buf
  g862
  (
    n585,
    n335
  );


  buf
  g863
  (
    n652,
    n170
  );


  not
  g864
  (
    n974,
    n195
  );


  buf
  g865
  (
    n465,
    n110
  );


  not
  g866
  (
    n1004,
    n118
  );


  not
  g867
  (
    n1193,
    n349
  );


  not
  g868
  (
    n881,
    n258
  );


  not
  g869
  (
    n674,
    n300
  );


  not
  g870
  (
    n1017,
    n130
  );


  not
  g871
  (
    n989,
    n194
  );


  buf
  g872
  (
    n507,
    n361
  );


  not
  g873
  (
    n766,
    n249
  );


  not
  g874
  (
    n715,
    n157
  );


  not
  g875
  (
    n903,
    n214
  );


  not
  g876
  (
    n912,
    n325
  );


  not
  g877
  (
    n815,
    n196
  );


  not
  g878
  (
    n961,
    n276
  );


  buf
  g879
  (
    n534,
    n140
  );


  not
  g880
  (
    n832,
    n128
  );


  buf
  g881
  (
    n714,
    n261
  );


  not
  g882
  (
    n1113,
    n294
  );


  buf
  g883
  (
    n1024,
    n287
  );


  not
  g884
  (
    n645,
    n218
  );


  buf
  g885
  (
    n1021,
    n157
  );


  buf
  g886
  (
    n1032,
    n244
  );


  buf
  g887
  (
    n956,
    n354
  );


  buf
  g888
  (
    n745,
    n211
  );


  not
  g889
  (
    n1196,
    n324
  );


  not
  g890
  (
    n804,
    n201
  );


  buf
  g891
  (
    n660,
    n296
  );


  not
  g892
  (
    n546,
    n260
  );


  buf
  g893
  (
    n526,
    n259
  );


  not
  g894
  (
    n1069,
    n211
  );


  buf
  g895
  (
    n494,
    n275
  );


  buf
  g896
  (
    n609,
    n347
  );


  not
  g897
  (
    n1168,
    n246
  );


  not
  g898
  (
    n878,
    n326
  );


  buf
  g899
  (
    n742,
    n141
  );


  buf
  g900
  (
    n482,
    n361
  );


  buf
  g901
  (
    n573,
    n168
  );


  not
  g902
  (
    n1177,
    n229
  );


  buf
  g903
  (
    n882,
    n162
  );


  buf
  g904
  (
    n1150,
    n124
  );


  buf
  g905
  (
    n748,
    n338
  );


  not
  g906
  (
    n769,
    n304
  );


  buf
  g907
  (
    n795,
    n348
  );


  not
  g908
  (
    n684,
    n221
  );


  not
  g909
  (
    n925,
    n270
  );


  not
  g910
  (
    n921,
    n236
  );


  buf
  g911
  (
    n1161,
    n183
  );


  buf
  g912
  (
    n662,
    n173
  );


  buf
  g913
  (
    n909,
    n273
  );


  buf
  g914
  (
    n1055,
    n187
  );


  buf
  g915
  (
    n1082,
    n313
  );


  not
  g916
  (
    n709,
    n319
  );


  not
  g917
  (
    n980,
    n161
  );


  not
  g918
  (
    KeyWire_0_15,
    n313
  );


  buf
  g919
  (
    n555,
    n170
  );


  buf
  g920
  (
    n995,
    n316
  );


  buf
  g921
  (
    n1166,
    n298
  );


  buf
  g922
  (
    n1181,
    n362
  );


  not
  g923
  (
    n1039,
    n289
  );


  not
  g924
  (
    n664,
    n111
  );


  buf
  g925
  (
    n864,
    n123
  );


  not
  g926
  (
    n726,
    n253
  );


  buf
  g927
  (
    n1199,
    n334
  );


  buf
  g928
  (
    n824,
    n137
  );


  not
  g929
  (
    n614,
    n191
  );


  not
  g930
  (
    n539,
    n169
  );


  buf
  g931
  (
    n556,
    n225
  );


  buf
  g932
  (
    n1119,
    n138
  );


  buf
  g933
  (
    n736,
    n244
  );


  not
  g934
  (
    n1074,
    n263
  );


  buf
  g935
  (
    n646,
    n197
  );


  buf
  g936
  (
    n1041,
    n157
  );


  buf
  g937
  (
    n1059,
    n222
  );


  buf
  g938
  (
    n636,
    n278
  );


  buf
  g939
  (
    n661,
    n341
  );


  not
  g940
  (
    n642,
    n163
  );


  not
  g941
  (
    n605,
    n363
  );


  not
  g942
  (
    n1085,
    n134
  );


  not
  g943
  (
    n999,
    n227
  );


  not
  g944
  (
    n580,
    n331
  );


  buf
  g945
  (
    n669,
    n359
  );


  buf
  g946
  (
    KeyWire_0_5,
    n323
  );


  buf
  g947
  (
    n1000,
    n213
  );


  buf
  g948
  (
    n1112,
    n360
  );


  not
  g949
  (
    n627,
    n196
  );


  not
  g950
  (
    n1025,
    n317
  );


  buf
  g951
  (
    n1134,
    n180
  );


  not
  g952
  (
    n1204,
    n350
  );


  not
  g953
  (
    KeyWire_0_6,
    n146
  );


  buf
  g954
  (
    n1142,
    n291
  );


  buf
  g955
  (
    n965,
    n154
  );


  not
  g956
  (
    n893,
    n227
  );


  buf
  g957
  (
    n571,
    n129
  );


  not
  g958
  (
    n495,
    n317
  );


  not
  g959
  (
    n492,
    n224
  );


  buf
  g960
  (
    n889,
    n222
  );


  buf
  g961
  (
    n1124,
    n282
  );


  not
  g962
  (
    n733,
    n220
  );


  buf
  g963
  (
    n628,
    n245
  );


  not
  g964
  (
    n713,
    n226
  );


  buf
  g965
  (
    n775,
    n142
  );


  buf
  g966
  (
    n760,
    n268
  );


  not
  g967
  (
    n765,
    n199
  );


  not
  g968
  (
    n623,
    n342
  );


  buf
  g969
  (
    KeyWire_0_20,
    n231
  );


  not
  g970
  (
    n702,
    n242
  );


  not
  g971
  (
    n559,
    n357
  );


  buf
  g972
  (
    n955,
    n171
  );


  buf
  g973
  (
    n755,
    n142
  );


  buf
  g974
  (
    n510,
    n359
  );


  not
  g975
  (
    n550,
    n106
  );


  buf
  g976
  (
    n561,
    n338
  );


  not
  g977
  (
    n988,
    n242
  );


  not
  g978
  (
    n895,
    n324
  );


  not
  g979
  (
    n1152,
    n342
  );


  not
  g980
  (
    n654,
    n315
  );


  not
  g981
  (
    n767,
    n229
  );


  not
  g982
  (
    n1058,
    n130
  );


  not
  g983
  (
    n902,
    n363
  );


  not
  g984
  (
    n537,
    n120
  );


  buf
  g985
  (
    n521,
    n148
  );


  buf
  g986
  (
    n853,
    n356
  );


  not
  g987
  (
    n858,
    n251
  );


  buf
  g988
  (
    n796,
    n254
  );


  buf
  g989
  (
    n688,
    n218
  );


  not
  g990
  (
    n671,
    n302
  );


  buf
  g991
  (
    n607,
    n263
  );


  not
  g992
  (
    n852,
    n274
  );


  not
  g993
  (
    n1054,
    n217
  );


  buf
  g994
  (
    n523,
    n174
  );


  not
  g995
  (
    n1042,
    n130
  );


  buf
  g996
  (
    n479,
    n184
  );


  buf
  g997
  (
    n829,
    n348
  );


  not
  g998
  (
    n973,
    n143
  );


  not
  g999
  (
    n649,
    n218
  );


  buf
  g1000
  (
    n756,
    n251
  );


  buf
  g1001
  (
    KeyWire_0_22,
    n180
  );


  not
  g1002
  (
    n1170,
    n135
  );


  not
  g1003
  (
    n1078,
    n327
  );


  not
  g1004
  (
    KeyWire_0_26,
    n270
  );


  buf
  g1005
  (
    n701,
    n291
  );


  not
  g1006
  (
    n868,
    n279
  );


  buf
  g1007
  (
    n818,
    n359
  );


  buf
  g1008
  (
    n1083,
    n162
  );


  not
  g1009
  (
    n813,
    n146
  );


  not
  g1010
  (
    n1057,
    n280
  );


  buf
  g1011
  (
    n803,
    n212
  );


  not
  g1012
  (
    n809,
    n314
  );


  buf
  g1013
  (
    n877,
    n228
  );


  buf
  g1014
  (
    n938,
    n129
  );


  buf
  g1015
  (
    n453,
    n326
  );


  not
  g1016
  (
    n788,
    n297
  );


  not
  g1017
  (
    n1182,
    n154
  );


  not
  g1018
  (
    n910,
    n337
  );


  not
  g1019
  (
    n480,
    n262
  );


  not
  g1020
  (
    n558,
    n345
  );


  buf
  g1021
  (
    n446,
    n230
  );


  buf
  g1022
  (
    n1151,
    n156
  );


  buf
  g1023
  (
    n578,
    n158
  );


  not
  g1024
  (
    n826,
    n285
  );


  not
  g1025
  (
    n1075,
    n193
  );


  buf
  g1026
  (
    n1104,
    n137
  );


  buf
  g1027
  (
    n1080,
    n223
  );


  not
  g1028
  (
    n841,
    n168
  );


  buf
  g1029
  (
    n444,
    n188
  );


  not
  g1030
  (
    n696,
    n238
  );


  buf
  g1031
  (
    n519,
    n219
  );


  buf
  g1032
  (
    n552,
    n133
  );


  not
  g1033
  (
    n622,
    n150
  );


  not
  g1034
  (
    n806,
    n333
  );


  not
  g1035
  (
    n749,
    n183
  );


  not
  g1036
  (
    n544,
    n116
  );


  not
  g1037
  (
    n1100,
    n205
  );


  buf
  g1038
  (
    n1081,
    n215
  );


  buf
  g1039
  (
    n470,
    n277
  );


  not
  g1040
  (
    n663,
    n328
  );


  not
  g1041
  (
    n1016,
    n141
  );


  buf
  g1042
  (
    n791,
    n176
  );


  buf
  g1043
  (
    n643,
    n202
  );


  buf
  g1044
  (
    n953,
    n154
  );


  buf
  g1045
  (
    n1065,
    n269
  );


  buf
  g1046
  (
    n621,
    n251
  );


  buf
  g1047
  (
    n1040,
    n189
  );


  not
  g1048
  (
    n869,
    n281
  );


  buf
  g1049
  (
    n567,
    n356
  );


  buf
  g1050
  (
    n1007,
    n244
  );


  not
  g1051
  (
    n1010,
    n181
  );


  buf
  g1052
  (
    n1139,
    n276
  );


  buf
  g1053
  (
    n986,
    n235
  );


  buf
  g1054
  (
    KeyWire_0_30,
    n149
  );


  buf
  g1055
  (
    KeyWire_0_12,
    n171
  );


  buf
  g1056
  (
    n549,
    n222
  );


  not
  g1057
  (
    n683,
    n189
  );


  buf
  g1058
  (
    n1201,
    n198
  );


  not
  g1059
  (
    n879,
    n358
  );


  not
  g1060
  (
    n485,
    n340
  );


  buf
  g1061
  (
    n1028,
    n326
  );


  buf
  g1062
  (
    n1125,
    n242
  );


  not
  g1063
  (
    n880,
    n280
  );


  not
  g1064
  (
    n822,
    n317
  );


  buf
  g1065
  (
    n1135,
    n210
  );


  not
  g1066
  (
    n1067,
    n132
  );


  not
  g1067
  (
    n998,
    n232
  );


  not
  g1068
  (
    n1158,
    n297
  );


  buf
  g1069
  (
    n1095,
    n167
  );


  buf
  g1070
  (
    n725,
    n268
  );


  buf
  g1071
  (
    n695,
    n126
  );


  buf
  g1072
  (
    n592,
    n329
  );


  not
  g1073
  (
    n598,
    n271
  );


  not
  g1074
  (
    n1015,
    n308
  );


  not
  g1075
  (
    n768,
    n179
  );


  not
  g1076
  (
    n464,
    n187
  );


  not
  g1077
  (
    n1079,
    n311
  );


  buf
  g1078
  (
    n718,
    n344
  );


  not
  g1079
  (
    n947,
    n297
  );


  buf
  g1080
  (
    n738,
    n331
  );


  buf
  g1081
  (
    n862,
    n306
  );


  not
  g1082
  (
    n513,
    n127
  );


  buf
  g1083
  (
    n897,
    n312
  );


  buf
  g1084
  (
    n1066,
    n132
  );


  not
  g1085
  (
    n707,
    n300
  );


  buf
  g1086
  (
    n971,
    n335
  );


  buf
  g1087
  (
    KeyWire_0_17,
    n255
  );


  buf
  g1088
  (
    n945,
    n212
  );


  not
  g1089
  (
    n1012,
    n292
  );


  buf
  g1090
  (
    n716,
    n155
  );


  not
  g1091
  (
    n762,
    n206
  );


  buf
  g1092
  (
    n790,
    n238
  );


  xnor
  g1093
  (
    n967,
    n144,
    n285,
    n236,
    n156
  );


  xnor
  g1094
  (
    n926,
    n362,
    n245,
    n322,
    n347
  );


  nor
  g1095
  (
    n530,
    n231,
    n299,
    n272,
    n107
  );


  nand
  g1096
  (
    n639,
    n225,
    n166,
    n286,
    n114
  );


  nand
  g1097
  (
    n677,
    n269,
    n307,
    n228,
    n293
  );


  nand
  g1098
  (
    n939,
    n116,
    n115,
    n184,
    n364
  );


  xnor
  g1099
  (
    n672,
    n233,
    n149,
    n352,
    n298
  );


  or
  g1100
  (
    n1116,
    n259,
    n127,
    n220,
    n218
  );


  xor
  g1101
  (
    n859,
    n186,
    n109,
    n122,
    n204
  );


  nand
  g1102
  (
    n933,
    n226,
    n121,
    n145,
    n323
  );


  nor
  g1103
  (
    n682,
    n345,
    n315,
    n329,
    n182
  );


  nor
  g1104
  (
    n569,
    n229,
    n159,
    n324,
    n246
  );


  and
  g1105
  (
    n533,
    n322,
    n211,
    n209,
    n240
  );


  and
  g1106
  (
    n801,
    n195,
    n182,
    n210,
    n267
  );


  nand
  g1107
  (
    n1160,
    n272,
    n264,
    n224,
    n161
  );


  nor
  g1108
  (
    n918,
    n349,
    n319,
    n132,
    n273
  );


  or
  g1109
  (
    n631,
    n196,
    n322,
    n229,
    n266
  );


  xnor
  g1110
  (
    n481,
    n350,
    n269,
    n266,
    n247
  );


  or
  g1111
  (
    n584,
    n118,
    n117,
    n292,
    n331
  );


  or
  g1112
  (
    n951,
    n359,
    n346,
    n313,
    n223
  );


  xnor
  g1113
  (
    n723,
    n318,
    n308,
    n156,
    n237
  );


  xnor
  g1114
  (
    n759,
    n299,
    n139,
    n151,
    n170
  );


  or
  g1115
  (
    n794,
    n303,
    n185,
    n300,
    n273
  );


  nor
  g1116
  (
    n979,
    n255,
    n119,
    n234,
    n147
  );


  xnor
  g1117
  (
    n860,
    n287,
    n332,
    n239,
    n116
  );


  and
  g1118
  (
    n690,
    n143,
    n106,
    n309,
    n165
  );


  xor
  g1119
  (
    n1198,
    n223,
    n214,
    n188,
    n192
  );


  xnor
  g1120
  (
    n460,
    n151,
    n314,
    n205,
    n248
  );


  nand
  g1121
  (
    n1110,
    n290,
    n292,
    n152,
    n311
  );


  xnor
  g1122
  (
    n691,
    n239,
    n320,
    n143,
    n332
  );


  xor
  g1123
  (
    n681,
    n179,
    n237,
    n150,
    n119
  );


  nand
  g1124
  (
    n780,
    n325,
    n254,
    n209,
    n146
  );


  xnor
  g1125
  (
    n821,
    n282,
    n195,
    n114,
    n277
  );


  and
  g1126
  (
    n638,
    n245,
    n159,
    n149,
    n298
  );


  nand
  g1127
  (
    n958,
    n155,
    n348,
    n326,
    n227
  );


  and
  g1128
  (
    n927,
    n160,
    n283,
    n361,
    n177
  );


  and
  g1129
  (
    n932,
    n185,
    n311,
    n153,
    n314
  );


  xnor
  g1130
  (
    n1072,
    n107,
    n224,
    n278,
    n305
  );


  xor
  g1131
  (
    n798,
    n279,
    n215,
    n152,
    n248
  );


  and
  g1132
  (
    n916,
    n143,
    n343,
    n360,
    n274
  );


  and
  g1133
  (
    n870,
    n190,
    n231,
    n345,
    n268
  );


  and
  g1134
  (
    n753,
    n311,
    n162,
    n262,
    n184
  );


  xor
  g1135
  (
    n727,
    n241,
    n117,
    n125,
    n350
  );


  nor
  g1136
  (
    n1164,
    n289,
    n271,
    n243,
    n203
  );


  and
  g1137
  (
    n1176,
    n200,
    n353,
    n134,
    n148
  );


  xor
  g1138
  (
    n917,
    n336,
    n206,
    n256,
    n164
  );


  nor
  g1139
  (
    n940,
    n167,
    n307,
    n133,
    n305
  );


  or
  g1140
  (
    n949,
    n165,
    n127,
    n247,
    n249
  );


  nand
  g1141
  (
    n923,
    n217,
    n233,
    n315,
    n240
  );


  nand
  g1142
  (
    n641,
    n263,
    n209,
    n134,
    n204
  );


  and
  g1143
  (
    n476,
    n180,
    n190,
    n112,
    n257
  );


  nor
  g1144
  (
    KeyWire_0_31,
    n183,
    n266,
    n168,
    n351
  );


  nand
  g1145
  (
    n472,
    n295,
    n290,
    n136,
    n360
  );


  or
  g1146
  (
    n633,
    n198,
    n210,
    n159,
    n336
  );


  nand
  g1147
  (
    n1064,
    n235,
    n148,
    n267,
    n163
  );


  or
  g1148
  (
    n665,
    n179,
    n198,
    n330,
    n199
  );


  or
  g1149
  (
    n1117,
    n107,
    n276,
    n110,
    n236
  );


  xor
  g1150
  (
    n827,
    n310,
    n158,
    n226,
    n178
  );


  xor
  g1151
  (
    n937,
    n187,
    n342,
    n134,
    n131
  );


  nor
  g1152
  (
    n991,
    n126,
    n122,
    n174,
    n219
  );


  xnor
  g1153
  (
    n875,
    n313,
    n169,
    n201,
    n144
  );


  xnor
  g1154
  (
    n618,
    n216,
    n110,
    n161,
    n252
  );


  or
  g1155
  (
    n1174,
    n124,
    n123,
    n245,
    n194
  );


  xor
  g1156
  (
    n455,
    n160,
    n321,
    n182,
    n129
  );


  nor
  g1157
  (
    n994,
    n339,
    n344,
    n357,
    n151
  );


  or
  g1158
  (
    n977,
    n166,
    n252,
    n202,
    n109
  );


  xnor
  g1159
  (
    n673,
    n234,
    n356,
    n316,
    n357
  );


  xnor
  g1160
  (
    n712,
    n147,
    n178,
    n149,
    n276
  );


  xnor
  g1161
  (
    n793,
    n254,
    n230,
    n172,
    n184
  );


  xor
  g1162
  (
    n1011,
    n296,
    n340,
    n302,
    n122
  );


  and
  g1163
  (
    n704,
    n216,
    n294,
    n131,
    n283
  );


  or
  g1164
  (
    n842,
    n207,
    n295,
    n321,
    n310
  );


  or
  g1165
  (
    n785,
    n282,
    n246,
    n173,
    n260
  );


  or
  g1166
  (
    n1190,
    n322,
    n135,
    n258,
    n169
  );


  and
  g1167
  (
    n911,
    n357,
    n335,
    n128,
    n212
  );


  nor
  g1168
  (
    n1154,
    n316,
    n120,
    n154,
    n207
  );


  and
  g1169
  (
    n962,
    n124,
    n258,
    n188,
    n230
  );


  nor
  g1170
  (
    n575,
    n275,
    n139,
    n282,
    n330
  );


  or
  g1171
  (
    n604,
    n131,
    n270,
    n275,
    n338
  );


  and
  g1172
  (
    n698,
    n283,
    n327,
    n330,
    n325
  );


  or
  g1173
  (
    n1002,
    n228,
    n207,
    n292,
    n253
  );


  xor
  g1174
  (
    n866,
    n334,
    n353,
    n106,
    n180
  );


  xnor
  g1175
  (
    n883,
    n219,
    n361,
    n205,
    n125
  );


  or
  g1176
  (
    n735,
    n350,
    n195,
    n277,
    n321
  );


  or
  g1177
  (
    n929,
    n148,
    n309,
    n214,
    n278
  );


  and
  g1178
  (
    n579,
    n165,
    n234,
    n233,
    n306
  );


  or
  g1179
  (
    n764,
    n288,
    n247,
    n293,
    n248
  );


  and
  g1180
  (
    n1036,
    n303,
    n243,
    n197,
    n333
  );


  and
  g1181
  (
    n473,
    n220,
    n243,
    n121,
    n116
  );


  xnor
  g1182
  (
    n488,
    n262,
    n354,
    n124,
    n253
  );


  xor
  g1183
  (
    n1479,
    n1172,
    n666,
    n432,
    n411
  );


  xor
  g1184
  (
    n1537,
    n780,
    n1099,
    n684,
    n1156
  );


  xnor
  g1185
  (
    n1298,
    n1107,
    n1116,
    n570,
    n1063
  );


  xor
  g1186
  (
    n1340,
    n1083,
    n1194,
    n803,
    n1026
  );


  xnor
  g1187
  (
    n1410,
    n401,
    n1012,
    n1127,
    n1103
  );


  nand
  g1188
  (
    n1453,
    n688,
    n1088,
    n530,
    n905
  );


  xnor
  g1189
  (
    n1249,
    n694,
    n1085,
    n900,
    n701
  );


  nand
  g1190
  (
    n1475,
    n1152,
    n537,
    n396,
    n542
  );


  xor
  g1191
  (
    n1235,
    n999,
    n420,
    n1084,
    n1189
  );


  xor
  g1192
  (
    n1338,
    n767,
    n1120,
    n1028,
    n1068
  );


  xnor
  g1193
  (
    n1486,
    n1162,
    n1125,
    n1020
  );


  nor
  g1194
  (
    n1302,
    n1034,
    n1084,
    n546,
    n689
  );


  xnor
  g1195
  (
    n1301,
    n1111,
    n439,
    n1182,
    n1126
  );


  xnor
  g1196
  (
    n1506,
    n638,
    n412,
    n413,
    n1101
  );


  or
  g1197
  (
    n1329,
    n429,
    n1131,
    n1171,
    n547
  );


  and
  g1198
  (
    n1347,
    n1049,
    n641,
    n1196,
    n790
  );


  xor
  g1199
  (
    n1241,
    n1130,
    n390,
    n1077,
    n1142
  );


  nor
  g1200
  (
    n1556,
    n1174,
    n455,
    n1013,
    n402
  );


  xnor
  g1201
  (
    n1344,
    n777,
    n1040,
    n371,
    n893
  );


  xor
  g1202
  (
    n1277,
    n717,
    n1015,
    n1166,
    n417
  );


  xnor
  g1203
  (
    n1547,
    n1182,
    n418,
    n384,
    n648
  );


  and
  g1204
  (
    n1353,
    n1109,
    n391,
    n1014,
    n1106
  );


  xnor
  g1205
  (
    n1354,
    n500,
    n1163,
    n402,
    n941
  );


  xnor
  g1206
  (
    n1470,
    n979,
    n1083,
    n781,
    n1129
  );


  and
  g1207
  (
    n1294,
    n760,
    n514,
    n1070,
    n436
  );


  nor
  g1208
  (
    n1367,
    n1037,
    n1117,
    n948,
    n876
  );


  nand
  g1209
  (
    n1562,
    n1175,
    n1109,
    n583,
    n502
  );


  nor
  g1210
  (
    n1579,
    n629,
    n861,
    n367,
    n988
  );


  nand
  g1211
  (
    n1383,
    n1033,
    n1049,
    n933,
    n459
  );


  xnor
  g1212
  (
    n1382,
    n370,
    n792,
    n405,
    n1167
  );


  xnor
  g1213
  (
    n1293,
    n394,
    n1169,
    n516,
    n384
  );


  or
  g1214
  (
    n1343,
    n716,
    n727,
    n460,
    n408
  );


  nor
  g1215
  (
    n1559,
    n1166,
    n825,
    n647,
    n1123
  );


  or
  g1216
  (
    n1312,
    n400,
    n1056,
    n1080,
    n1145
  );


  or
  g1217
  (
    n1211,
    n365,
    n394,
    n440,
    n1177
  );


  nand
  g1218
  (
    n1458,
    n1164,
    n804,
    n624,
    n1104
  );


  nor
  g1219
  (
    n1469,
    n1145,
    n1182,
    n393,
    n1112
  );


  or
  g1220
  (
    n1399,
    n1111,
    n1186,
    n961,
    n403
  );


  nand
  g1221
  (
    n1466,
    n379,
    n366,
    n1124,
    n1086
  );


  or
  g1222
  (
    n1234,
    n1180,
    n378,
    n564,
    n643
  );


  or
  g1223
  (
    n1236,
    n1079,
    n682,
    n1105,
    n1016
  );


  nand
  g1224
  (
    n1318,
    n1163,
    n381,
    n880,
    n428
  );


  nand
  g1225
  (
    n1316,
    n410,
    n1169,
    n405,
    n486
  );


  xnor
  g1226
  (
    n1310,
    n936,
    n892,
    n401,
    n646
  );


  nor
  g1227
  (
    n1300,
    n1012,
    n710,
    n1085,
    n1190
  );


  or
  g1228
  (
    n1350,
    n1136,
    n439,
    n1098,
    n1148
  );


  xor
  g1229
  (
    n1299,
    n424,
    n458,
    n446,
    n369
  );


  xor
  g1230
  (
    n1269,
    n433,
    n1097,
    n442,
    n1132
  );


  xnor
  g1231
  (
    n1546,
    n677,
    n409,
    n415,
    n1153
  );


  xnor
  g1232
  (
    n1325,
    n1109,
    n886,
    n763,
    n960
  );


  xor
  g1233
  (
    n1259,
    n1184,
    n481,
    n1077,
    n549
  );


  xor
  g1234
  (
    n1351,
    n386,
    n925,
    n645,
    n787
  );


  nand
  g1235
  (
    n1369,
    n1107,
    n741,
    n454,
    n557
  );


  and
  g1236
  (
    n1402,
    n697,
    n669,
    n389,
    n1116
  );


  xnor
  g1237
  (
    n1548,
    n419,
    n1100,
    n1029,
    n1043
  );


  xor
  g1238
  (
    n1231,
    n437,
    n1088,
    n432,
    n567
  );


  and
  g1239
  (
    n1362,
    n779,
    n1004,
    n418,
    n439
  );


  and
  g1240
  (
    n1480,
    n414,
    n431,
    n1151,
    n390
  );


  xnor
  g1241
  (
    n1334,
    n1038,
    n392,
    n829,
    n1121
  );


  nand
  g1242
  (
    n1566,
    n832,
    n1108,
    n1050,
    n591
  );


  or
  g1243
  (
    n1514,
    n443,
    n675,
    n722,
    n1098
  );


  nor
  g1244
  (
    n1378,
    n529,
    n1138,
    n1180,
    n608
  );


  xnor
  g1245
  (
    n1433,
    n929,
    n417,
    n1076,
    n883
  );


  and
  g1246
  (
    n1240,
    n390,
    n623,
    n1185,
    n1103
  );


  or
  g1247
  (
    n1442,
    n1133,
    n1170,
    n415,
    n847
  );


  or
  g1248
  (
    n1248,
    n493,
    n422,
    n1173,
    n1048
  );


  nor
  g1249
  (
    n1324,
    n901,
    n367,
    n423,
    n1011
  );


  and
  g1250
  (
    n1268,
    n1002,
    n812,
    n1072,
    n611
  );


  nand
  g1251
  (
    n1282,
    n1094,
    n386,
    n1195,
    n1119
  );


  xor
  g1252
  (
    n1474,
    n368,
    n461,
    n735,
    n1177
  );


  xor
  g1253
  (
    n1575,
    n1058,
    n709,
    n487,
    n1122
  );


  nand
  g1254
  (
    n1419,
    n839,
    n766,
    n1160,
    n389
  );


  or
  g1255
  (
    n1251,
    n484,
    n412,
    n785,
    n984
  );


  xor
  g1256
  (
    n1497,
    n1174,
    n656,
    n895,
    n394
  );


  or
  g1257
  (
    n1352,
    n1027,
    n599,
    n1189,
    n1091
  );


  xnor
  g1258
  (
    n1457,
    n568,
    n1102,
    n1108,
    n1043
  );


  nand
  g1259
  (
    n1215,
    n720,
    n556,
    n1150,
    n1148
  );


  and
  g1260
  (
    n1320,
    n539,
    n1052,
    n385,
    n1134
  );


  xnor
  g1261
  (
    n1572,
    n1081,
    n706,
    n1197,
    n616
  );


  xnor
  g1262
  (
    n1246,
    n1102,
    n1100,
    n515,
    n1186
  );


  or
  g1263
  (
    n1229,
    n426,
    n1156,
    n414,
    n750
  );


  xor
  g1264
  (
    n1304,
    n391,
    n1092,
    n771,
    n833
  );


  or
  g1265
  (
    n1250,
    n1158,
    n662,
    n1181,
    n744
  );


  or
  g1266
  (
    n1448,
    n462,
    n1183,
    n375,
    n1064
  );


  xnor
  g1267
  (
    n1275,
    n705,
    n1078,
    n965,
    n1024
  );


  nor
  g1268
  (
    n1377,
    n712,
    n1104,
    n465,
    n1129
  );


  nor
  g1269
  (
    n1412,
    n1144,
    n1046,
    n1058,
    n373
  );


  nand
  g1270
  (
    n1337,
    n891,
    n1158,
    n1153,
    n1089
  );


  nand
  g1271
  (
    n1341,
    n364,
    n1076,
    n1155,
    n691
  );


  xor
  g1272
  (
    n1493,
    n1084,
    n1171,
    n528,
    n1187
  );


  nor
  g1273
  (
    n1256,
    n1123,
    n998,
    n497,
    n1106
  );


  and
  g1274
  (
    n1431,
    n1166,
    n672,
    n1141,
    n1042
  );


  xnor
  g1275
  (
    n1284,
    n1019,
    n1187,
    n1075,
    n1068
  );


  nor
  g1276
  (
    n1295,
    n976,
    n756,
    n1193,
    n1098
  );


  or
  g1277
  (
    n1432,
    n855,
    n438,
    n681,
    n1007
  );


  xnor
  g1278
  (
    n1288,
    n1162,
    n749,
    n1130,
    n1142
  );


  or
  g1279
  (
    n1533,
    n1057,
    n372,
    n637,
    n1034
  );


  xnor
  g1280
  (
    n1450,
    n1096,
    n1029,
    n755,
    n1193
  );


  or
  g1281
  (
    n1239,
    n1151,
    n378,
    n858,
    n1067
  );


  or
  g1282
  (
    n1392,
    n761,
    n651,
    n1171,
    n404
  );


  nor
  g1283
  (
    n1440,
    n986,
    n1024,
    n577,
    n1166
  );


  xor
  g1284
  (
    n1224,
    n475,
    n1197,
    n1150,
    n844
  );


  xnor
  g1285
  (
    n1292,
    n1055,
    n719,
    n368,
    n551
  );


  xor
  g1286
  (
    n1496,
    n1039,
    n991,
    n1109,
    n518
  );


  and
  g1287
  (
    n1553,
    n954,
    n396,
    n1085,
    n1190
  );


  xor
  g1288
  (
    n1580,
    n431,
    n508,
    n748,
    n376
  );


  xor
  g1289
  (
    n1303,
    n383,
    n601,
    n1128,
    n368
  );


  xor
  g1290
  (
    n1452,
    n916,
    n882,
    n711,
    n380
  );


  and
  g1291
  (
    n1244,
    n545,
    n375,
    n696,
    n1086
  );


  nand
  g1292
  (
    n1357,
    n1104,
    n786,
    n980,
    n1144
  );


  nand
  g1293
  (
    n1262,
    n1179,
    n995,
    n695,
    n1103
  );


  nand
  g1294
  (
    KeyWire_0_11,
    n1085,
    n914,
    n1112,
    n430
  );


  nand
  g1295
  (
    n1409,
    n1006,
    n366,
    n394,
    n1197
  );


  xor
  g1296
  (
    n1565,
    n738,
    n704,
    n810,
    n1089
  );


  or
  g1297
  (
    n1384,
    n405,
    n385,
    n983,
    n990
  );


  and
  g1298
  (
    n1504,
    n831,
    n1158,
    n1026,
    n503
  );


  xor
  g1299
  (
    n1364,
    n433,
    n934,
    n365,
    n1122
  );


  xor
  g1300
  (
    n1400,
    n910,
    n585,
    n663,
    n456
  );


  nand
  g1301
  (
    n1314,
    n378,
    n987,
    n1163,
    n1184
  );


  nor
  g1302
  (
    n1487,
    n650,
    n1071,
    n609,
    n731
  );


  and
  g1303
  (
    n1568,
    n1195,
    n1191,
    n410,
    n1016
  );


  xnor
  g1304
  (
    n1489,
    n1155,
    n541,
    n707,
    n969
  );


  xor
  g1305
  (
    n1534,
    n600,
    n1124,
    n758,
    n1136
  );


  and
  g1306
  (
    n1216,
    n1185,
    n412,
    n422,
    n1081
  );


  nand
  g1307
  (
    n1258,
    n1106,
    n422,
    n512,
    n1133
  );


  nand
  g1308
  (
    n1571,
    n1065,
    n436,
    n726,
    n467
  );


  or
  g1309
  (
    n1544,
    n469,
    n407,
    n1180,
    n554
  );


  and
  g1310
  (
    n1389,
    n1132,
    n1115,
    n937,
    n395
  );


  and
  g1311
  (
    n1542,
    n1143,
    n1047,
    n430,
    n386
  );


  or
  g1312
  (
    n1569,
    n1091,
    n1172,
    n424,
    n1011
  );


  and
  g1313
  (
    n1576,
    n1064,
    n686,
    n1188,
    n745
  );


  xor
  g1314
  (
    n1551,
    n945,
    n403,
    n374,
    n1135
  );


  nand
  g1315
  (
    n1421,
    n1063,
    n1014,
    n1067,
    n419
  );


  or
  g1316
  (
    n1274,
    n416,
    n617,
    n816,
    n1136
  );


  nor
  g1317
  (
    n1393,
    n793,
    n519,
    n1198,
    n370
  );


  xnor
  g1318
  (
    n1463,
    n889,
    n1161,
    n1054,
    n407
  );


  nand
  g1319
  (
    n1430,
    n630,
    n1106,
    n1139,
    n808
  );


  or
  g1320
  (
    n1488,
    n1121,
    n428,
    n427,
    n1018
  );


  nor
  g1321
  (
    n1414,
    n1044,
    n580,
    n1186,
    n729
  );


  and
  g1322
  (
    n1381,
    n1087,
    n1141,
    n412,
    n1118
  );


  xnor
  g1323
  (
    n1315,
    n393,
    n782,
    n523,
    n479
  );


  xnor
  g1324
  (
    n1317,
    n434,
    n652,
    n1018,
    n466
  );


  nor
  g1325
  (
    n1206,
    n1140,
    n429,
    n1129,
    n451
  );


  and
  g1326
  (
    n1574,
    n713,
    n846,
    n1147,
    n474
  );


  or
  g1327
  (
    n1499,
    n702,
    n400,
    n375,
    n1079
  );


  or
  g1328
  (
    n1443,
    n845,
    n1175,
    n1035,
    n587
  );


  or
  g1329
  (
    n1515,
    n447,
    n1184,
    n1118,
    n1094
  );


  nand
  g1330
  (
    n1407,
    n1163,
    n434,
    n379,
    n851
  );


  xnor
  g1331
  (
    n1281,
    n775,
    n1102,
    n1127,
    n853
  );


  and
  g1332
  (
    n1348,
    n538,
    n1121,
    n1165,
    n1092
  );


  nor
  g1333
  (
    n1321,
    n860,
    n1155,
    n1189,
    n1167
  );


  xor
  g1334
  (
    n1413,
    n947,
    n1146,
    n974,
    n424
  );


  nor
  g1335
  (
    n1309,
    n1009,
    n464,
    n418,
    n615
  );


  xor
  g1336
  (
    n1355,
    n445,
    n427,
    n1093,
    n425
  );


  nand
  g1337
  (
    n1512,
    n400,
    n1183,
    n1146,
    n1042
  );


  nand
  g1338
  (
    n1464,
    n951,
    n414,
    n724,
    n1145
  );


  and
  g1339
  (
    n1255,
    n1140,
    n1126,
    n1079,
    n1088
  );


  xor
  g1340
  (
    n1521,
    n433,
    n799,
    n1121,
    n863
  );


  and
  g1341
  (
    n1342,
    n373,
    n1181,
    n520,
    n559
  );


  or
  g1342
  (
    n1391,
    n581,
    n1073,
    n908,
    n1191
  );


  xnor
  g1343
  (
    n1219,
    n826,
    n562,
    n421,
    n606
  );


  xor
  g1344
  (
    n1526,
    n820,
    n509,
    n898,
    n1122
  );


  xor
  g1345
  (
    n1365,
    n1041,
    n660,
    n1120,
    n1133
  );


  nand
  g1346
  (
    n1541,
    n1188,
    n1061,
    n1021,
    n433
  );


  and
  g1347
  (
    n1387,
    n605,
    n742,
    n1062,
    n955
  );


  xor
  g1348
  (
    n1346,
    n946,
    n1082,
    n415,
    n1196
  );


  nor
  g1349
  (
    n1472,
    n423,
    n902,
    n573,
    n1086
  );


  nor
  g1350
  (
    n1289,
    n1198,
    n425,
    n418,
    n1127
  );


  or
  g1351
  (
    n1356,
    n578,
    n386,
    n594,
    n1149
  );


  nand
  g1352
  (
    n1490,
    n421,
    n561,
    n552,
    n939
  );


  nor
  g1353
  (
    n1214,
    n586,
    n1095,
    n584,
    n534
  );


  xor
  g1354
  (
    n1502,
    n1095,
    n753,
    n1178,
    n1104
  );


  xor
  g1355
  (
    n1285,
    n388,
    n1123,
    n420,
    n935
  );


  or
  g1356
  (
    n1287,
    n1159,
    n1047,
    n1056,
    n1023
  );


  nor
  g1357
  (
    n1461,
    n869,
    n751,
    n1075,
    n1116
  );


  nor
  g1358
  (
    n1260,
    n1120,
    n1157,
    n1150,
    n1003
  );


  xor
  g1359
  (
    n1323,
    n533,
    n492,
    n1142,
    n482
  );


  nand
  g1360
  (
    n1494,
    n1036,
    n1173,
    n1089,
    n426
  );


  and
  g1361
  (
    n1370,
    n1138,
    n768,
    n639,
    n371
  );


  and
  g1362
  (
    n1528,
    n1167,
    n510,
    n1084,
    n1195
  );


  or
  g1363
  (
    n1570,
    n1147,
    n746,
    n396,
    n949
  );


  or
  g1364
  (
    n1434,
    n1196,
    n1087,
    n977,
    n674
  );


  nor
  g1365
  (
    n1491,
    n924,
    n909,
    n607,
    n1041
  );


  nor
  g1366
  (
    n1297,
    n565,
    n699,
    n415,
    n406
  );


  nand
  g1367
  (
    n1311,
    n1175,
    n653,
    n401,
    n973
  );


  xor
  g1368
  (
    n1558,
    n864,
    n540,
    n1115,
    n827
  );


  xnor
  g1369
  (
    n1230,
    n1110,
    n668,
    n1135,
    n1087
  );


  xor
  g1370
  (
    n1257,
    n848,
    n603,
    n1143,
    n1160
  );


  nor
  g1371
  (
    n1339,
    n1122,
    n438,
    n943,
    n757
  );


  and
  g1372
  (
    n1417,
    n432,
    n406,
    n435
  );


  or
  g1373
  (
    n1267,
    n1108,
    n1092,
    n1080,
    n1037
  );


  nand
  g1374
  (
    n1273,
    n432,
    n1114,
    n411
  );


  xor
  g1375
  (
    n1390,
    n439,
    n728,
    n373,
    n387
  );


  xnor
  g1376
  (
    n1416,
    n1113,
    n408,
    n1139,
    n1118
  );


  nor
  g1377
  (
    n1308,
    n1131,
    n912,
    n714,
    n1114
  );


  nor
  g1378
  (
    n1376,
    n1153,
    n1147,
    n1160,
    n1088
  );


  and
  g1379
  (
    n1252,
    n425,
    n1176,
    n407,
    n404
  );


  nand
  g1380
  (
    n1296,
    n1198,
    n378,
    n1090,
    n1154
  );


  xor
  g1381
  (
    n1243,
    n1096,
    n1105,
    n994,
    n1090
  );


  nor
  g1382
  (
    n1510,
    n457,
    n1023,
    n1176,
    n1152
  );


  or
  g1383
  (
    n1210,
    n1191,
    n885,
    n640,
    n1135
  );


  or
  g1384
  (
    n1221,
    n1091,
    n627,
    n387,
    n759
  );


  or
  g1385
  (
    n1429,
    n1154,
    n1091,
    n392,
    n1120
  );


  nor
  g1386
  (
    n1578,
    n993,
    n1177,
    n942,
    n676
  );


  xnor
  g1387
  (
    n1222,
    n1197,
    n791,
    n1070,
    n764
  );


  or
  g1388
  (
    n1326,
    n420,
    n1025,
    n1144,
    n1013
  );


  xor
  g1389
  (
    n1401,
    n1022,
    n480,
    n428,
    n824
  );


  nand
  g1390
  (
    n1279,
    n1152,
    n1066,
    n413,
    n452
  );


  xnor
  g1391
  (
    n1272,
    n411,
    n1022,
    n1169,
    n1125
  );


  nor
  g1392
  (
    n1305,
    n391,
    n1097,
    n374,
    n801
  );


  xor
  g1393
  (
    n1482,
    n661,
    n419,
    n915,
    n654
  );


  xnor
  g1394
  (
    n1573,
    n383,
    n1165,
    n690,
    n1078
  );


  xor
  g1395
  (
    n1540,
    n1149,
    n957,
    n505,
    n1105
  );


  and
  g1396
  (
    n1516,
    n1152,
    n435,
    n1010,
    n526
  );


  nand
  g1397
  (
    n1483,
    n852,
    n718,
    n619,
    n866
  );


  xor
  g1398
  (
    n1349,
    n1083,
    n1021,
    n631,
    n835
  );


  nand
  g1399
  (
    n1525,
    n495,
    n978,
    n1170,
    n1127
  );


  xor
  g1400
  (
    n1485,
    n1100,
    n604,
    n776,
    n377
  );


  or
  g1401
  (
    n1261,
    n1141,
    n837,
    n1188,
    n737
  );


  xnor
  g1402
  (
    n1507,
    n399,
    n1045,
    n1185,
    n409
  );


  nor
  g1403
  (
    n1319,
    n1142,
    n783,
    n772,
    n1177
  );


  xnor
  g1404
  (
    n1439,
    n610,
    n501,
    n1030,
    n388
  );


  or
  g1405
  (
    n1518,
    n752,
    n634,
    n644,
    n406
  );


  or
  g1406
  (
    n1426,
    n1099,
    n1137,
    n566,
    n575
  );


  and
  g1407
  (
    n1411,
    n1051,
    n470,
    n1128,
    n1148
  );


  and
  g1408
  (
    KeyWire_0_29,
    n1101,
    n773,
    n1155,
    n1053
  );


  nor
  g1409
  (
    n1276,
    n673,
    n762,
    n1186,
    n1019
  );


  or
  g1410
  (
    n1563,
    n449,
    n398,
    n550,
    n872
  );


  or
  g1411
  (
    n1208,
    n410,
    n448,
    n403,
    n371
  );


  or
  g1412
  (
    n1415,
    n376,
    n632,
    n1077,
    n953
  );


  nor
  g1413
  (
    n1237,
    n535,
    n429,
    n389,
    n967
  );


  nor
  g1414
  (
    n1509,
    n679,
    n435,
    n375,
    n1132
  );


  or
  g1415
  (
    n1335,
    n388,
    n725,
    n1192,
    n383
  );


  nor
  g1416
  (
    n1520,
    n494,
    n367,
    n873,
    n597
  );


  nand
  g1417
  (
    n1527,
    n1159,
    n379,
    n732,
    n658
  );


  xnor
  g1418
  (
    n1286,
    n1179,
    n1094,
    n887,
    n1098
  );


  nor
  g1419
  (
    n1435,
    n413,
    n1181,
    n819,
    n1192
  );


  xnor
  g1420
  (
    n1473,
    n1113,
    n1195,
    n1135,
    n374
  );


  nand
  g1421
  (
    n1332,
    n838,
    n657,
    n1119,
    n1100
  );


  and
  g1422
  (
    n1328,
    n843,
    n544,
    n896,
    n1161
  );


  or
  g1423
  (
    n1290,
    n1174,
    n1182,
    n1107,
    n1110
  );


  xor
  g1424
  (
    n1358,
    n1193,
    n1188,
    n380,
    n625
  );


  xor
  g1425
  (
    n1327,
    n1178,
    n1015,
    n1017,
    n621
  );


  nor
  g1426
  (
    n1441,
    n1119,
    n1113,
    n576,
    n1159
  );


  nand
  g1427
  (
    n1265,
    n392,
    n989,
    n385,
    n1138
  );


  and
  g1428
  (
    n1330,
    n1053,
    n628,
    n903,
    n388
  );


  or
  g1429
  (
    KeyWire_0_1,
    n950,
    n420,
    n1114,
    n1157
  );


  xnor
  g1430
  (
    n1359,
    n1093,
    n1103,
    n633,
    n393
  );


  and
  g1431
  (
    n1379,
    n472,
    n1081,
    n1112,
    n579
  );


  or
  g1432
  (
    KeyWire_0_28,
    n572,
    n558,
    n398,
    n1108
  );


  or
  g1433
  (
    n1363,
    n1075,
    n1124,
    n612,
    n683
  );


  or
  g1434
  (
    n1462,
    n370,
    n1174,
    n1111,
    n404
  );


  nor
  g1435
  (
    n1396,
    n421,
    n1008,
    n397,
    n818
  );


  nand
  g1436
  (
    n1467,
    n453,
    n1131,
    n1151,
    n870
  );


  or
  g1437
  (
    n1212,
    n800,
    n754,
    n985,
    n1031
  );


  nor
  g1438
  (
    n1550,
    n377,
    n788,
    n444,
    n1054
  );


  and
  g1439
  (
    n1227,
    n1137,
    n595,
    n590,
    n1114
  );


  xnor
  g1440
  (
    n1245,
    n1052,
    n932,
    n369,
    n419
  );


  and
  g1441
  (
    n1517,
    n434,
    n1090,
    n1080,
    n1153
  );


  or
  g1442
  (
    n1264,
    n613,
    n1077,
    n1164,
    n1078
  );


  xor
  g1443
  (
    n1539,
    n380,
    n930,
    n956,
    n364
  );


  xor
  g1444
  (
    n1554,
    n841,
    n399,
    n1118,
    n372
  );


  xnor
  g1445
  (
    n1226,
    n399,
    n430,
    n1139,
    n871
  );


  or
  g1446
  (
    n1538,
    n1111,
    n1045,
    n1170,
    n840
  );


  xnor
  g1447
  (
    n1253,
    n560,
    n1095,
    n739,
    n376
  );


  nor
  g1448
  (
    n1209,
    n396,
    n1139,
    n958,
    n1133
  );


  or
  g1449
  (
    n1322,
    n1191,
    n1141,
    n1181,
    n1105
  );


  or
  g1450
  (
    n1454,
    n730,
    n614,
    n700,
    n1055
  );


  or
  g1451
  (
    n1373,
    n884,
    n471,
    n571,
    n1172
  );


  and
  g1452
  (
    n1333,
    n828,
    n434,
    n734,
    n395
  );


  or
  g1453
  (
    n1233,
    n1194,
    n1194,
    n1147,
    n1069
  );


  or
  g1454
  (
    n1478,
    n382,
    n992,
    n1071,
    n598
  );


  nor
  g1455
  (
    n1238,
    n1158,
    n367,
    n975,
    n1078
  );


  xnor
  g1456
  (
    n1455,
    n1073,
    n1137,
    n904,
    n1140
  );


  xnor
  g1457
  (
    n1529,
    n1136,
    n413,
    n596,
    n1028
  );


  xnor
  g1458
  (
    n1530,
    n1025,
    n996,
    n532,
    n592
  );


  xnor
  g1459
  (
    n1552,
    n649,
    n981,
    n952,
    n1095
  );


  nor
  g1460
  (
    n1501,
    n692,
    n1154,
    n894,
    n655
  );


  or
  g1461
  (
    n1447,
    n1046,
    n1162,
    n1130,
    n850
  );


  nand
  g1462
  (
    n1270,
    n789,
    n842,
    n374,
    n1074
  );


  xor
  g1463
  (
    n1394,
    n1090,
    n1173,
    n1190,
    n431
  );


  nand
  g1464
  (
    n1498,
    n1128,
    n365,
    n574,
    n437
  );


  xnor
  g1465
  (
    n1331,
    n402,
    n499,
    n1097,
    n770
  );


  and
  g1466
  (
    n1561,
    n1080,
    n384,
    n794,
    n425
  );


  xnor
  g1467
  (
    n1395,
    n1048,
    n1164,
    n1101,
    n1156
  );


  or
  g1468
  (
    n1513,
    n391,
    n498,
    n806,
    n1183
  );


  or
  g1469
  (
    n1385,
    n1178,
    n1040,
    n1146,
    n715
  );


  nand
  g1470
  (
    n1449,
    n431,
    n1089,
    n366,
    n401
  );


  and
  g1471
  (
    n1424,
    n721,
    n1066,
    n427,
    n1179
  );


  xor
  g1472
  (
    n1543,
    n784,
    n1099,
    n370,
    n906
  );


  and
  g1473
  (
    n1232,
    n1157,
    n1030,
    n874,
    n1074
  );


  nor
  g1474
  (
    n1307,
    n971,
    n1151,
    n736,
    n814
  );


  xnor
  g1475
  (
    n1306,
    n1044,
    n1115,
    n437,
    n589
  );


  and
  g1476
  (
    n1425,
    n1160,
    n1126,
    n371,
    n428
  );


  or
  g1477
  (
    n1459,
    n1187,
    n1138,
    n1126,
    n416
  );


  or
  g1478
  (
    n1374,
    n389,
    n395,
    n1190,
    n1059
  );


  or
  g1479
  (
    n1380,
    n1020,
    n1005,
    n1038,
    n1069
  );


  and
  g1480
  (
    n1428,
    n970,
    n620,
    n1178,
    n622
  );


  xor
  g1481
  (
    n1266,
    n1099,
    n1035,
    n436,
    n1036
  );


  nand
  g1482
  (
    n1388,
    n1140,
    n923,
    n437,
    n403
  );


  or
  g1483
  (
    n1271,
    n1129,
    n563,
    n392,
    n635
  );


  nand
  g1484
  (
    n1404,
    n377,
    n1050,
    n406,
    n877
  );


  nor
  g1485
  (
    n1283,
    n693,
    n913,
    n1183,
    n450
  );


  xor
  g1486
  (
    n1225,
    n1082,
    n899,
    n1086,
    n402
  );


  and
  g1487
  (
    n1403,
    n1161,
    n1093,
    n854,
    n1079
  );


  nand
  g1488
  (
    n1418,
    n408,
    n865,
    n1162,
    n517
  );


  nor
  g1489
  (
    n1476,
    n506,
    n507,
    n382,
    n1144
  );


  xor
  g1490
  (
    n1564,
    n1149,
    n504,
    n489,
    n1125
  );


  nor
  g1491
  (
    n1492,
    n1185,
    n778,
    n1137,
    n409
  );


  and
  g1492
  (
    n1555,
    n1150,
    n1123,
    n1149,
    n422
  );


  xor
  g1493
  (
    n1567,
    n1107,
    n1093,
    n387,
    n964
  );


  nor
  g1494
  (
    n1535,
    n398,
    n588,
    n1039,
    n397
  );


  or
  g1495
  (
    n1254,
    n377,
    n1009,
    n382,
    n1124
  );


  or
  g1496
  (
    n1220,
    n918,
    n959,
    n478,
    n1075
  );


  and
  g1497
  (
    n1423,
    n1176,
    n525,
    n405,
    n1110
  );


  nor
  g1498
  (
    n1531,
    n1061,
    n1184,
    n1101,
    n1060
  );


  nor
  g1499
  (
    n1223,
    n473,
    n1176,
    n381,
    n1115
  );


  or
  g1500
  (
    n1242,
    n897,
    n527,
    n703,
    n397
  );


  nand
  g1501
  (
    n1495,
    n636,
    n966,
    n849,
    n1074
  );


  xnor
  g1502
  (
    n1217,
    n1059,
    n369,
    n1146,
    n1117
  );


  nor
  g1503
  (
    n1386,
    n569,
    n381,
    n834,
    n888
  );


  nor
  g1504
  (
    n1372,
    n1057,
    n490,
    n463,
    n468
  );


  xor
  g1505
  (
    n1207,
    n664,
    n879,
    n417,
    n1156
  );


  nand
  g1506
  (
    n1511,
    n922,
    n364,
    n1157,
    n921
  );


  nor
  g1507
  (
    n1361,
    n381,
    n1032,
    n390,
    n1083
  );


  and
  g1508
  (
    n1375,
    n1000,
    n477,
    n438,
    n1027
  );


  or
  g1509
  (
    n1465,
    n1134,
    n410,
    n1168,
    n404
  );


  xnor
  g1510
  (
    n1405,
    n1180,
    n511,
    n387,
    n1194
  );


  and
  g1511
  (
    n1522,
    n417,
    n867,
    n830,
    n997
  );


  or
  g1512
  (
    n1468,
    n733,
    n938,
    n685,
    n429
  );


  nand
  g1513
  (
    n1560,
    n379,
    n743,
    n678,
    n857
  );


  xnor
  g1514
  (
    n1263,
    n723,
    n1179,
    n1092,
    n665
  );


  nand
  g1515
  (
    n1471,
    n962,
    n926,
    n1094,
    n555
  );


  xor
  g1516
  (
    n1519,
    n1161,
    n1168,
    n421,
    n1072
  );


  nor
  g1517
  (
    n1291,
    n553,
    n875,
    n384,
    n667
  );


  xnor
  g1518
  (
    n1460,
    n1102,
    n1145,
    n822,
    n380
  );


  xnor
  g1519
  (
    n1336,
    n878,
    n911,
    n931,
    n671
  );


  xor
  g1520
  (
    n1549,
    n968,
    n438,
    n907,
    n483
  );


  xor
  g1521
  (
    n1577,
    n1170,
    n393,
    n369,
    n813
  );


  nand
  g1522
  (
    n1438,
    n373,
    n1017,
    n1168,
    n1051
  );


  nor
  g1523
  (
    n1532,
    n522,
    n815,
    n1076,
    n1192
  );


  nand
  g1524
  (
    n1557,
    n862,
    n642,
    n795,
    n1165
  );


  xor
  g1525
  (
    n1360,
    n1198,
    n868,
    n740,
    n1008
  );


  xor
  g1526
  (
    n1524,
    n1187,
    n1065,
    n1074,
    n1154
  );


  and
  g1527
  (
    n1437,
    n1119,
    n1087,
    n1096,
    n817
  );


  and
  g1528
  (
    n1422,
    n626,
    n1031,
    n427,
    n582
  );


  nand
  g1529
  (
    n1278,
    n602,
    n1167,
    n1196,
    n491
  );


  and
  g1530
  (
    n1484,
    n1132,
    n496,
    n1171,
    n1113
  );


  xor
  g1531
  (
    n1523,
    n797,
    n365,
    n485,
    n769
  );


  or
  g1532
  (
    n1218,
    n1189,
    n890,
    n395,
    n543
  );


  xnor
  g1533
  (
    n1397,
    n659,
    n1165,
    n376,
    n440
  );


  or
  g1534
  (
    n1345,
    n963,
    n398,
    n407,
    n1033
  );


  xor
  g1535
  (
    n1445,
    n408,
    n927,
    n521,
    n1172
  );


  xor
  g1536
  (
    n1500,
    n382,
    n513,
    n1134,
    n385
  );


  or
  g1537
  (
    n1444,
    n1117,
    n809,
    n372,
    n1148
  );


  xor
  g1538
  (
    n1508,
    n1168,
    n1143,
    n416,
    n836
  );


  or
  g1539
  (
    n1503,
    n1076,
    n1130,
    n368,
    n524
  );


  or
  g1540
  (
    n1481,
    n1032,
    n372,
    n972,
    n618
  );


  nor
  g1541
  (
    n1545,
    n476,
    n805,
    n1110,
    n1164
  );


  and
  g1542
  (
    n1280,
    n919,
    n859,
    n920,
    n687
  );


  nor
  g1543
  (
    n1368,
    n747,
    n1082,
    n1193,
    n881
  );


  or
  g1544
  (
    n1228,
    n1175,
    n399,
    n1062,
    n397
  );


  nand
  g1545
  (
    KeyWire_0_14,
    n423,
    n531,
    n409,
    n414
  );


  nor
  g1546
  (
    n1536,
    n802,
    n1096,
    n917,
    n1112
  );


  nor
  g1547
  (
    n1451,
    n548,
    n1159,
    n426,
    n1082
  );


  nor
  g1548
  (
    n1446,
    n383,
    n1128,
    n670,
    n708
  );


  or
  g1549
  (
    n1371,
    n430,
    n1060,
    n982,
    n488
  );


  nand
  g1550
  (
    n1427,
    n774,
    n856,
    n821,
    n1116
  );


  or
  g1551
  (
    n1456,
    n1117,
    n798,
    n1192,
    n1081
  );


  or
  g1552
  (
    n1398,
    n680,
    n1134,
    n436,
    n807
  );


  xor
  g1553
  (
    n1366,
    n823,
    n424,
    n1173,
    n928
  );


  and
  g1554
  (
    n1477,
    n416,
    n1143,
    n1131,
    n765
  );


  xnor
  g1555
  (
    n1313,
    n796,
    n1169,
    n400,
    n698
  );


  xor
  g1556
  (
    n1213,
    n1001,
    n423,
    n1097,
    n536
  );


  xor
  g1557
  (
    n1505,
    n593,
    n811,
    n440,
    n1010
  );


  or
  g1558
  (
    n1406,
    n426,
    n366,
    n940,
    n944
  );


  buf
  g1559
  (
    n1589,
    n1234
  );


  buf
  g1560
  (
    n1584,
    n1232
  );


  not
  g1561
  (
    n1607,
    n1223
  );


  not
  g1562
  (
    n1595,
    n1211
  );


  buf
  g1563
  (
    n1603,
    n1225
  );


  not
  g1564
  (
    n1596,
    n1217
  );


  not
  g1565
  (
    n1600,
    n1205
  );


  buf
  g1566
  (
    n1605,
    n1222
  );


  buf
  g1567
  (
    n1591,
    n1216
  );


  not
  g1568
  (
    n1599,
    n1210
  );


  not
  g1569
  (
    n1604,
    n1224
  );


  buf
  g1570
  (
    n1590,
    n1212
  );


  not
  g1571
  (
    n1592,
    n1220
  );


  buf
  g1572
  (
    n1608,
    n1209
  );


  not
  g1573
  (
    n1588,
    n1230
  );


  buf
  g1574
  (
    n1587,
    n1221
  );


  not
  g1575
  (
    n1594,
    n1214
  );


  not
  g1576
  (
    n1601,
    n1227
  );


  buf
  g1577
  (
    n1581,
    n1231
  );


  buf
  g1578
  (
    n1602,
    n1215
  );


  not
  g1579
  (
    n1597,
    n1226
  );


  not
  g1580
  (
    n1609,
    n1236
  );


  not
  g1581
  (
    n1606,
    n1228
  );


  not
  g1582
  (
    n1593,
    n1206
  );


  buf
  g1583
  (
    n1585,
    n1213
  );


  buf
  g1584
  (
    n1586,
    n1219
  );


  buf
  g1585
  (
    n1598,
    n1235
  );


  not
  g1586
  (
    n1583,
    n1218
  );


  and
  g1587
  (
    n1582,
    n1233,
    n1207,
    n1229,
    n1208
  );


  and
  g1588
  (
    n1614,
    n1299,
    n1254,
    n1274,
    n1590
  );


  or
  g1589
  (
    n1630,
    n1312,
    n1237,
    n1271,
    n1247
  );


  and
  g1590
  (
    n1618,
    n1252,
    n1596,
    n1584,
    n1286
  );


  or
  g1591
  (
    n1632,
    n1314,
    n1303,
    n1269,
    n1280
  );


  nand
  g1592
  (
    n1637,
    n1594,
    n1266,
    n1297,
    n1249
  );


  xor
  g1593
  (
    n1619,
    n1307,
    n1305,
    n1245,
    n1276
  );


  and
  g1594
  (
    n1625,
    n1253,
    n1598,
    n1243,
    n1586
  );


  xor
  g1595
  (
    n1636,
    n1251,
    n1270,
    n1261,
    n1318
  );


  nor
  g1596
  (
    n1634,
    n1239,
    n1255,
    n1322,
    n1257
  );


  xor
  g1597
  (
    n1617,
    n1290,
    n1315,
    n1581,
    n1316
  );


  or
  g1598
  (
    n1635,
    n1602,
    n1317,
    n1600,
    n1601
  );


  xnor
  g1599
  (
    n1626,
    n1591,
    n1291,
    n1262,
    n1319
  );


  xnor
  g1600
  (
    n1622,
    n1259,
    n1256,
    n1273,
    n1281
  );


  nor
  g1601
  (
    n1639,
    n1593,
    n1309,
    n1604,
    n1592
  );


  or
  g1602
  (
    n1628,
    n1300,
    n1277,
    n1607,
    n1250
  );


  and
  g1603
  (
    n1620,
    n1321,
    n1260,
    n1263,
    n1265
  );


  xnor
  g1604
  (
    n1638,
    n1326,
    n1267,
    n1287,
    n1588
  );


  xor
  g1605
  (
    n1633,
    n1302,
    n1313,
    n1248,
    n1583
  );


  or
  g1606
  (
    n1613,
    n1606,
    n1268,
    n1599,
    n1589
  );


  or
  g1607
  (
    n1612,
    n1306,
    n1264,
    n1324,
    n1308
  );


  xor
  g1608
  (
    n1611,
    n1595,
    n1587,
    n1258,
    n1304
  );


  or
  g1609
  (
    n1616,
    n1609,
    n1289,
    n1295,
    n1246
  );


  nand
  g1610
  (
    KeyWire_0_27,
    n1301,
    n1275,
    n1597,
    n1608
  );


  nand
  g1611
  (
    n1610,
    n1323,
    n1242,
    n1294,
    n1603
  );


  or
  g1612
  (
    n1629,
    n1285,
    n1605,
    n1238,
    n1292
  );


  nand
  g1613
  (
    n1621,
    n1283,
    n1279,
    n1310,
    n1325
  );


  or
  g1614
  (
    n1627,
    n1582,
    n1288,
    n1311,
    n1585
  );


  nor
  g1615
  (
    n1615,
    n1272,
    n1298,
    n1282,
    n1240
  );


  and
  g1616
  (
    n1624,
    n1609,
    n1293,
    n1241,
    n1296
  );


  xor
  g1617
  (
    n1631,
    n1284,
    n1278,
    n1320,
    n1244
  );


  or
  g1618
  (
    n1643,
    n1339,
    n1338,
    n1611,
    n1347
  );


  xor
  g1619
  (
    n1640,
    n1616,
    n1614,
    n1343,
    n1337
  );


  nor
  g1620
  (
    n1641,
    n1334,
    n1612,
    n1348,
    n1329
  );


  xnor
  g1621
  (
    n1647,
    n1344,
    n1327,
    n1610,
    n1335
  );


  and
  g1622
  (
    n1642,
    n1336,
    n1332,
    n1350,
    n1340
  );


  nand
  g1623
  (
    n1644,
    n1331,
    n1613,
    n1346,
    n1617
  );


  or
  g1624
  (
    n1646,
    n1345,
    n1341,
    n1333,
    n1342
  );


  and
  g1625
  (
    n1645,
    n1615,
    n1328,
    n1349,
    n1330
  );


  buf
  g1626
  (
    n1660,
    n1642
  );


  buf
  g1627
  (
    n1652,
    n1642
  );


  buf
  g1628
  (
    n1657,
    n1641
  );


  buf
  g1629
  (
    n1656,
    n1640
  );


  not
  g1630
  (
    n1661,
    n1641
  );


  buf
  g1631
  (
    n1658,
    n1640
  );


  not
  g1632
  (
    n1648,
    n1643
  );


  buf
  g1633
  (
    n1659,
    n1643
  );


  not
  g1634
  (
    n1651,
    n1642
  );


  buf
  g1635
  (
    n1655,
    n1643
  );


  buf
  g1636
  (
    n1654,
    n1641
  );


  buf
  g1637
  (
    n1650,
    n1643
  );


  not
  g1638
  (
    n1653,
    n1619
  );


  xnor
  g1639
  (
    n1649,
    n1618,
    n1641,
    n1642
  );


  not
  g1640
  (
    n1672,
    n1654
  );


  or
  g1641
  (
    n1667,
    n1659,
    n1651,
    n1660
  );


  or
  g1642
  (
    n1662,
    n1354,
    n1657,
    n1653,
    n1352
  );


  xnor
  g1643
  (
    n1671,
    n1650,
    n1660,
    n1656,
    n1652
  );


  or
  g1644
  (
    n1675,
    n1650,
    n1657,
    n1653,
    n1661
  );


  nand
  g1645
  (
    n1663,
    n1656,
    n1648,
    n1659,
    n1650
  );


  nor
  g1646
  (
    n1664,
    n1658,
    n1648,
    n1655
  );


  or
  g1647
  (
    n1673,
    n1653,
    n1649,
    n1648
  );


  nor
  g1648
  (
    n1665,
    n1656,
    n1653,
    n1655
  );


  and
  g1649
  (
    n1668,
    n1652,
    n1654,
    n1355,
    n1658
  );


  or
  g1650
  (
    n1669,
    n1649,
    n1651,
    n1353,
    n1659
  );


  xnor
  g1651
  (
    n1666,
    n1660,
    n1656,
    n1651,
    n1351
  );


  and
  g1652
  (
    n1670,
    n1654,
    n1660,
    n1655,
    n1658
  );


  xor
  g1653
  (
    n1676,
    n1658,
    n1652,
    n1650
  );


  nand
  g1654
  (
    n1674,
    n1659,
    n1657,
    n1649
  );


  xor
  g1655
  (
    n1677,
    n1651,
    n1654,
    n1661,
    n1356
  );


  not
  g1656
  (
    n1686,
    n1373
  );


  buf
  g1657
  (
    n1691,
    n1366
  );


  buf
  g1658
  (
    n1683,
    n1367
  );


  buf
  g1659
  (
    n1679,
    n1673
  );


  not
  g1660
  (
    n1692,
    n1376
  );


  buf
  g1661
  (
    n1678,
    n1663
  );


  buf
  g1662
  (
    n1684,
    n1668
  );


  buf
  g1663
  (
    n1681,
    n1371
  );


  buf
  g1664
  (
    n1685,
    n1361
  );


  nand
  g1665
  (
    n1689,
    n1662,
    n1670,
    n1665
  );


  and
  g1666
  (
    n1690,
    n1358,
    n1666,
    n1674,
    n1664
  );


  or
  g1667
  (
    n1688,
    n1357,
    n1359,
    n1669,
    n1677
  );


  nor
  g1668
  (
    n1682,
    n1360,
    n1375,
    n1364,
    n1368
  );


  nand
  g1669
  (
    n1687,
    n1667,
    n1374,
    n1672,
    n1369
  );


  or
  g1670
  (
    n1693,
    n1671,
    n1675,
    n1370,
    n1365
  );


  and
  g1671
  (
    n1680,
    n1372,
    n1676,
    n1363,
    n1362
  );


  and
  g1672
  (
    n1722,
    n1393,
    n1681,
    n1682,
    n1620
  );


  nor
  g1673
  (
    n1704,
    n1628,
    n1680,
    n1626,
    n1403
  );


  xnor
  g1674
  (
    n1717,
    n1691,
    n1692,
    n1693,
    n1398
  );


  or
  g1675
  (
    n1703,
    n1394,
    n1412,
    n1199,
    n1400
  );


  nand
  g1676
  (
    n1727,
    n1681,
    n1625,
    n1382,
    n1683
  );


  xor
  g1677
  (
    n1713,
    n1691,
    n1645,
    n441,
    n1402
  );


  nor
  g1678
  (
    n1721,
    n440,
    n1396,
    n1689,
    n1385
  );


  nor
  g1679
  (
    n1710,
    n1622,
    n1391,
    n1692,
    n1200
  );


  nor
  g1680
  (
    n1705,
    n1692,
    n1687,
    n1202
  );


  xnor
  g1681
  (
    n1699,
    n1645,
    n1390,
    n1686,
    n1404
  );


  nor
  g1682
  (
    n1716,
    n1679,
    n1688,
    n1693,
    n1379
  );


  xor
  g1683
  (
    KeyWire_0_21,
    n1408,
    n1684,
    n1647
  );


  xnor
  g1684
  (
    n1708,
    n1410,
    n1689,
    n1199
  );


  nand
  g1685
  (
    n1700,
    n1623,
    n1644,
    n1399,
    n1383
  );


  nor
  g1686
  (
    n1719,
    n1644,
    n1679,
    n1200,
    n1202
  );


  xor
  g1687
  (
    n1714,
    n1647,
    n1646,
    n1201
  );


  xor
  g1688
  (
    n1707,
    n1201,
    n1688,
    n1202,
    n1389
  );


  nor
  g1689
  (
    n1726,
    n441,
    n1401,
    n1691,
    n1646
  );


  xor
  g1690
  (
    n1724,
    n1687,
    n1647,
    n1678,
    n1683
  );


  xnor
  g1691
  (
    n1728,
    n1682,
    n1377,
    n1645,
    n1621
  );


  xor
  g1692
  (
    n1711,
    n1381,
    n1388,
    n1387,
    n1407
  );


  and
  g1693
  (
    n1698,
    n1690,
    n1645,
    n1682,
    n1397
  );


  nand
  g1694
  (
    n1694,
    n1685,
    n441,
    n1678,
    n1384
  );


  xor
  g1695
  (
    n1697,
    n1629,
    n1690,
    n1683,
    n1679
  );


  nor
  g1696
  (
    n1725,
    n1624,
    n1687,
    n1413
  );


  nand
  g1697
  (
    n1706,
    n1686,
    n1680,
    n1693
  );


  xor
  g1698
  (
    n1701,
    n1678,
    n1411,
    n1392,
    n1692
  );


  nor
  g1699
  (
    n1709,
    n1646,
    n1199,
    n1406,
    n1688
  );


  nor
  g1700
  (
    n1729,
    n1682,
    n1690,
    n1681,
    n1691
  );


  nor
  g1701
  (
    n1730,
    n1685,
    n1685,
    n1684,
    n1395
  );


  and
  g1702
  (
    n1702,
    n1684,
    n1646,
    n1414,
    n1200
  );


  xnor
  g1703
  (
    n1718,
    n1378,
    n1405,
    n1693,
    n1644
  );


  nor
  g1704
  (
    n1695,
    n1644,
    n1681,
    n1201,
    n1685
  );


  and
  g1705
  (
    n1723,
    n1688,
    n1647,
    n1689,
    n1678
  );


  xnor
  g1706
  (
    n1712,
    n1686,
    n1680,
    n1679,
    n1386
  );


  or
  g1707
  (
    n1720,
    n1409,
    n1200,
    n1627,
    n1690
  );


  nor
  g1708
  (
    n1696,
    n1683,
    n1380,
    n1686,
    n1689
  );


  xnor
  g1709
  (
    n1731,
    n1696,
    n1697,
    n1695,
    n1694
  );


  and
  g1710
  (
    n1732,
    n1695,
    n1697,
    n1696,
    n1698
  );


  xnor
  g1711
  (
    n1737,
    n1701,
    n1703,
    n1705,
    n1704
  );


  nor
  g1712
  (
    n1736,
    n1703,
    n1731,
    n1732
  );


  and
  g1713
  (
    n1735,
    n1704,
    n1700,
    n1702
  );


  nor
  g1714
  (
    n1734,
    n1701,
    n1732,
    n1698
  );


  nor
  g1715
  (
    n1733,
    n1705,
    n1699,
    n1702
  );


  not
  g1716
  (
    n1740,
    n1737
  );


  not
  g1717
  (
    n1743,
    n1736
  );


  buf
  g1718
  (
    n1742,
    n1734
  );


  not
  g1719
  (
    n1745,
    n1733
  );


  buf
  g1720
  (
    n1738,
    n1737
  );


  not
  g1721
  (
    n1739,
    n1737
  );


  not
  g1722
  (
    n1741,
    n1735
  );


  buf
  g1723
  (
    n1744,
    n1737
  );


  not
  g1724
  (
    n1751,
    n1740
  );


  buf
  g1725
  (
    n1746,
    n1421
  );


  xnor
  g1726
  (
    n1750,
    n1741,
    n1423
  );


  nand
  g1727
  (
    n1748,
    n1422,
    n1416,
    n1738,
    n1742
  );


  or
  g1728
  (
    n1749,
    n1415,
    n1420,
    n1419,
    n1424
  );


  nand
  g1729
  (
    n1747,
    n1743,
    n1417,
    n1418,
    n1739
  );


  nor
  g1730
  (
    n1752,
    n1428,
    n1437,
    n1436,
    n1434
  );


  xnor
  g1731
  (
    n1753,
    n1438,
    n1630,
    n1426,
    n1435
  );


  nand
  g1732
  (
    n1757,
    n1429,
    n1430,
    n1439,
    n1745
  );


  nand
  g1733
  (
    n1754,
    n1425,
    n1432,
    n1748,
    n1746
  );


  and
  g1734
  (
    n1756,
    n1751,
    n1747,
    n1749,
    n1744
  );


  xor
  g1735
  (
    n1755,
    n1433,
    n1750,
    n1431,
    n1427
  );


  xnor
  g1736
  (
    n1761,
    n1756,
    n1752,
    n1710,
    n1446
  );


  and
  g1737
  (
    n1762,
    n1714,
    n1452,
    n1706,
    n1443
  );


  xnor
  g1738
  (
    n1764,
    n1707,
    n1706,
    n1442,
    n1755
  );


  nand
  g1739
  (
    n1767,
    n1757,
    n1757,
    n1709,
    n1710
  );


  nor
  g1740
  (
    KeyWire_0_3,
    n1445,
    n1708,
    n1713,
    n1450
  );


  or
  g1741
  (
    n1758,
    n1714,
    n1444,
    n1447,
    n1454
  );


  and
  g1742
  (
    n1760,
    n1756,
    n1713,
    n1754,
    n1711
  );


  xnor
  g1743
  (
    n1759,
    n1712,
    n1715,
    n1441,
    n1708
  );


  nor
  g1744
  (
    n1768,
    n1451,
    n1757,
    n1456
  );


  nand
  g1745
  (
    n1769,
    n1756,
    n1756,
    n1455,
    n1449
  );


  xor
  g1746
  (
    n1765,
    n1711,
    n1707,
    n1448,
    n1709
  );


  nand
  g1747
  (
    n1763,
    n1440,
    n1453,
    n1753,
    n1712
  );


  or
  g1748
  (
    n1773,
    n1474,
    n1478,
    n1764,
    n1465
  );


  xor
  g1749
  (
    n1772,
    n1469,
    n1471,
    n1472,
    n1475
  );


  or
  g1750
  (
    n1776,
    n1479,
    n1477,
    n1470,
    n1466
  );


  nor
  g1751
  (
    n1775,
    n1460,
    n1765,
    n1473,
    n1476
  );


  xor
  g1752
  (
    n1777,
    n1468,
    n1462,
    n1769,
    n1467
  );


  and
  g1753
  (
    n1770,
    n1458,
    n1762,
    n1766,
    n1767
  );


  or
  g1754
  (
    n1774,
    n1457,
    n1768,
    n1461,
    n1464
  );


  nor
  g1755
  (
    n1771,
    n1463,
    n1763,
    n1459,
    n1480
  );


  xor
  g1756
  (
    n1780,
    n1487,
    n1482,
    n1483,
    n1771
  );


  and
  g1757
  (
    n1781,
    n1485,
    n1486,
    n1489,
    n1661
  );


  xor
  g1758
  (
    n1779,
    n1773,
    n1770,
    n1772,
    n1484
  );


  xor
  g1759
  (
    n1778,
    n1661,
    n1481,
    n1490,
    n1488
  );


  or
  g1760
  (
    n1786,
    n1778,
    n1637,
    n1632,
    n1636
  );


  xnor
  g1761
  (
    n1796,
    n1638,
    n1778,
    n1779,
    n1777
  );


  or
  g1762
  (
    n1793,
    n1722,
    n1631,
    n1778,
    n1715
  );


  or
  g1763
  (
    n1788,
    n1776,
    n1777
  );


  nand
  g1764
  (
    n1791,
    n1781,
    n1637,
    n1717,
    n1636
  );


  nor
  g1765
  (
    n1792,
    n1780,
    n1779,
    n1638,
    n1720
  );


  nand
  g1766
  (
    n1784,
    n1778,
    n1633,
    n1775,
    n1721
  );


  or
  g1767
  (
    n1787,
    n1780,
    n1780,
    n1775,
    n1638
  );


  xnor
  g1768
  (
    n1789,
    n1776,
    n1636,
    n1716,
    n1634
  );


  xor
  g1769
  (
    n1790,
    n1635,
    n1636,
    n1716,
    n1720
  );


  or
  g1770
  (
    n1782,
    n1719,
    n1775,
    n1777,
    n1639
  );


  and
  g1771
  (
    n1797,
    n1639,
    n1779,
    n1776
  );


  and
  g1772
  (
    n1794,
    n1717,
    n1781
  );


  xnor
  g1773
  (
    n1795,
    n1723,
    n1637,
    n1721,
    n1638
  );


  xor
  g1774
  (
    n1783,
    n1775,
    n1780,
    n1722,
    n1774
  );


  xor
  g1775
  (
    n1785,
    n1719,
    n1637,
    n1718
  );


  nor
  g1776
  (
    n1802,
    n1789,
    n1790,
    n1786,
    n1788
  );


  nand
  g1777
  (
    n1799,
    n1787,
    n1789,
    n1782,
    n1788
  );


  or
  g1778
  (
    n1800,
    n1790,
    n1783,
    n1492,
    n1788
  );


  nor
  g1779
  (
    n1798,
    n1491,
    n1789,
    n1787,
    n1788
  );


  and
  g1780
  (
    n1801,
    n1789,
    n1784,
    n1493,
    n1785
  );


  or
  g1781
  (
    n1806,
    n1792,
    n1791
  );


  xor
  g1782
  (
    n1804,
    n1790,
    n1790,
    n1791,
    n1799
  );


  and
  g1783
  (
    n1807,
    n1494,
    n1496,
    n1801,
    n1793
  );


  or
  g1784
  (
    n1805,
    n1793,
    n1800,
    n1792
  );


  nor
  g1785
  (
    n1803,
    n1792,
    n1798,
    n1495,
    n1802
  );


  xnor
  g1786
  (
    n1808,
    n1497,
    n1498,
    n1803,
    n1499
  );


  xor
  g1787
  (
    n1809,
    n1807,
    n1808,
    n1639
  );


  xnor
  g1788
  (
    n1810,
    n1806,
    n1639,
    n1805,
    n1804
  );


  xnor
  g1789
  (
    n1816,
    n1725,
    n1726,
    n1502,
    n1504
  );


  or
  g1790
  (
    n1812,
    n1500,
    n1725,
    n1724,
    n1723
  );


  nand
  g1791
  (
    n1814,
    n1726,
    n1809,
    n1810,
    n1506
  );


  xnor
  g1792
  (
    n1813,
    n1809,
    n1810,
    n1505,
    n1723
  );


  or
  g1793
  (
    n1817,
    n1724,
    n1725
  );


  or
  g1794
  (
    n1811,
    n1503,
    n1810,
    n1501,
    n1809
  );


  and
  g1795
  (
    n1815,
    n1809,
    n1810,
    n1723,
    n1724
  );


  buf
  g1796
  (
    n1821,
    n1812
  );


  not
  g1797
  (
    n1823,
    n1814
  );


  buf
  g1798
  (
    n1825,
    n1814
  );


  buf
  g1799
  (
    n1819,
    n1815
  );


  not
  g1800
  (
    n1818,
    n1814
  );


  buf
  g1801
  (
    n1824,
    n1814
  );


  not
  g1802
  (
    n1820,
    n1813
  );


  buf
  g1803
  (
    n1822,
    n1811
  );


  nor
  g1804
  (
    n1836,
    n1533,
    n1816,
    n1822,
    n1824
  );


  nand
  g1805
  (
    n1832,
    n1525,
    n1509,
    n1820,
    n1815
  );


  nand
  g1806
  (
    n1831,
    n1531,
    n1816,
    n1520,
    n1825
  );


  xnor
  g1807
  (
    n1826,
    n1534,
    n1528,
    n1536,
    n1515
  );


  nor
  g1808
  (
    n1837,
    n1519,
    n1514,
    n1535,
    n1823
  );


  nand
  g1809
  (
    n1839,
    n1818,
    n1539,
    n1817,
    n1513
  );


  xor
  g1810
  (
    n1833,
    n1530,
    n1537,
    n1521,
    n1817
  );


  nor
  g1811
  (
    n1829,
    n1816,
    n1825,
    n1527
  );


  nor
  g1812
  (
    n1827,
    n1522,
    n1821,
    n1529,
    n1524
  );


  and
  g1813
  (
    n1830,
    n1507,
    n1824,
    n1526,
    n1517
  );


  xor
  g1814
  (
    n1835,
    n1508,
    n1512,
    n1825,
    n1819
  );


  nand
  g1815
  (
    n1828,
    n1815,
    n1532,
    n1824
  );


  nor
  g1816
  (
    n1838,
    n1538,
    n1523,
    n1518,
    n1516
  );


  xnor
  g1817
  (
    n1834,
    n1816,
    n1510,
    n1815,
    n1511
  );


  not
  g1818
  (
    n1843,
    n1837
  );


  buf
  g1819
  (
    n1842,
    n1540
  );


  buf
  g1820
  (
    n1840,
    n1838
  );


  not
  g1821
  (
    n1845,
    n1834
  );


  not
  g1822
  (
    n1844,
    n1832
  );


  buf
  g1823
  (
    n1841,
    n1836
  );


  nand
  g1824
  (
    n1846,
    n1835,
    n1833
  );


  nand
  g1825
  (
    n1847,
    n1728,
    n1839,
    n1541,
    n1726
  );


  and
  g1826
  (
    n1852,
    n1840,
    n1844,
    n1843,
    n1547
  );


  and
  g1827
  (
    n1850,
    n1727,
    n1727,
    n1728,
    n1544
  );


  xor
  g1828
  (
    n1851,
    n1542,
    n1728,
    n1842
  );


  nor
  g1829
  (
    n1848,
    n1727,
    n1726,
    n1546,
    n1845
  );


  and
  g1830
  (
    n1849,
    n1545,
    n1543,
    n1841,
    n1727
  );


  xor
  g1831
  (
    n1853,
    n1553,
    n1548,
    n1849,
    n1852
  );


  nor
  g1832
  (
    n1858,
    n1550,
    n1730,
    n1555
  );


  xor
  g1833
  (
    KeyWire_0_4,
    n1730,
    n1554,
    n1729,
    n1851
  );


  nor
  g1834
  (
    KeyWire_0_2,
    n1848,
    n1552,
    n1729,
    n1847
  );


  nand
  g1835
  (
    n1857,
    n1846,
    n1729,
    n1556,
    n1551
  );


  or
  g1836
  (
    n1856,
    n1549,
    n1730,
    n1729,
    n1850
  );


  and
  g1837
  (
    n1868,
    n1796,
    n1857,
    n1794,
    n1558
  );


  xnor
  g1838
  (
    KeyWire_0_8,
    n1858,
    n1561,
    n1797,
    n1795
  );


  nand
  g1839
  (
    n1866,
    n1565,
    n1794,
    n1562,
    n1796
  );


  and
  g1840
  (
    n1865,
    n1796,
    n1797,
    n1795,
    n1567
  );


  nand
  g1841
  (
    n1864,
    n1795,
    n1853,
    n1566,
    n1564
  );


  xor
  g1842
  (
    n1867,
    n1557,
    n1858,
    n1568
  );


  xor
  g1843
  (
    n1859,
    n1793,
    n1796,
    n1560,
    n1855
  );


  and
  g1844
  (
    n1862,
    n1793,
    n1858,
    n1559,
    n1797
  );


  nand
  g1845
  (
    n1863,
    n1854,
    n1856,
    n1795,
    n1797
  );


  xor
  g1846
  (
    n1860,
    n1857,
    n1563,
    n1794
  );


  and
  g1847
  (
    n1870,
    n441,
    n1203,
    n1570,
    n1569
  );


  or
  g1848
  (
    n1869,
    n1203,
    n1868,
    n1571,
    n1867
  );


  or
  g1849
  (
    n1871,
    n1870,
    n1573,
    n1574,
    n1572
  );


  and
  g1850
  (
    n1873,
    n1871,
    n1576,
    n1580,
    n1575
  );


  xor
  g1851
  (
    n1872,
    n1579,
    n1577,
    n1871,
    n1578
  );


  xor
  g1852
  (
    n1875,
    n1873,
    n1872
  );


  or
  g1853
  (
    n1877,
    n1204,
    n1873
  );


  nor
  g1854
  (
    n1876,
    n1817,
    n1204,
    n1872
  );


  nand
  g1855
  (
    n1874,
    n1203,
    n1203,
    n1204,
    n1817
  );


  or
  g1856
  (
    n1878,
    n1874,
    n1876,
    n1875,
    n1877
  );


  xor
  KeyGate_0_0
  (
    n816,
    keyIn_0_0,
    KeyWire_0_0
  );


  xor
  KeyGate_0_1
  (
    n1205,
    keyIn_0_1,
    KeyWire_0_1
  );


  xor
  KeyGate_0_2
  (
    n1855,
    keyIn_0_2,
    KeyWire_0_2
  );


  xor
  KeyGate_0_3
  (
    n1766,
    keyIn_0_3,
    KeyWire_0_3
  );


  xnor
  KeyGate_0_4
  (
    n1854,
    keyIn_0_4,
    KeyWire_0_4
  );


  xor
  KeyGate_0_5
  (
    n581,
    keyIn_0_5,
    KeyWire_0_5
  );


  xnor
  KeyGate_0_6
  (
    n914,
    keyIn_0_6,
    KeyWire_0_6
  );


  xnor
  KeyGate_0_7
  (
    n153,
    keyIn_0_7,
    KeyWire_0_7
  );


  xnor
  KeyGate_0_8
  (
    n1861,
    keyIn_0_8,
    KeyWire_0_8
  );


  xnor
  KeyGate_0_9
  (
    n409,
    keyIn_0_9,
    KeyWire_0_9
  );


  xnor
  KeyGate_0_10
  (
    n500,
    keyIn_0_10,
    KeyWire_0_10
  );


  xor
  KeyGate_0_11
  (
    n1247,
    keyIn_0_11,
    KeyWire_0_11
  );


  xor
  KeyGate_0_12
  (
    n722,
    keyIn_0_12,
    KeyWire_0_12
  );


  xor
  KeyGate_0_13
  (
    n132,
    keyIn_0_13,
    KeyWire_0_13
  );


  xnor
  KeyGate_0_14
  (
    n1436,
    keyIn_0_14,
    KeyWire_0_14
  );


  xor
  KeyGate_0_15
  (
    n564,
    keyIn_0_15,
    KeyWire_0_15
  );


  xnor
  KeyGate_0_16
  (
    n1132,
    keyIn_0_16,
    KeyWire_0_16
  );


  xnor
  KeyGate_0_17
  (
    n506,
    keyIn_0_17,
    KeyWire_0_17
  );


  xor
  KeyGate_0_18
  (
    n557,
    keyIn_0_18,
    KeyWire_0_18
  );


  xor
  KeyGate_0_19
  (
    n390,
    keyIn_0_19,
    KeyWire_0_19
  );


  xnor
  KeyGate_0_20
  (
    n1138,
    keyIn_0_20,
    KeyWire_0_20
  );


  xor
  KeyGate_0_21
  (
    n1715,
    keyIn_0_21,
    KeyWire_0_21
  );


  xor
  KeyGate_0_22
  (
    n514,
    keyIn_0_22,
    KeyWire_0_22
  );


  xnor
  KeyGate_0_23
  (
    n1172,
    keyIn_0_23,
    KeyWire_0_23
  );


  xnor
  KeyGate_0_24
  (
    n189,
    keyIn_0_24,
    KeyWire_0_24
  );


  xor
  KeyGate_0_25
  (
    n275,
    keyIn_0_25,
    KeyWire_0_25
  );


  xnor
  KeyGate_0_26
  (
    n981,
    keyIn_0_26,
    KeyWire_0_26
  );


  xor
  KeyGate_0_27
  (
    n1623,
    keyIn_0_27,
    KeyWire_0_27
  );


  xor
  KeyGate_0_28
  (
    n1408,
    keyIn_0_28,
    KeyWire_0_28
  );


  xnor
  KeyGate_0_29
  (
    n1420,
    keyIn_0_29,
    KeyWire_0_29
  );


  xnor
  KeyGate_0_30
  (
    n825,
    keyIn_0_30,
    KeyWire_0_30
  );


  xor
  KeyGate_0_31
  (
    n828,
    keyIn_0_31,
    KeyWire_0_31
  );


endmodule


