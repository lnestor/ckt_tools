// Benchmark C:\Users\Lucas Nestor\Documents\osu\sp21\esl\circuit_generation\Stats\4_6_generated_stats\Stat_100_53 written by SynthGen on 2021/04/05 11:08:38
module Stat_100_53( n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32,
 n100, n93, n80, n114, n99, n110, n107, n92,
 n84, n86, n79, n115, n91, n95, n88, n112,
 n117, n89, n132, n129, n120, n124, n128, n127,
 n125, n123, n119, n126, n122, n121, n131, n130);

input n1, n2, n3, n4, n5, n6, n7, n8,
 n9, n10, n11, n12, n13, n14, n15, n16,
 n17, n18, n19, n20, n21, n22, n23, n24,
 n25, n26, n27, n28, n29, n30, n31, n32;

output n100, n93, n80, n114, n99, n110, n107, n92,
 n84, n86, n79, n115, n91, n95, n88, n112,
 n117, n89, n132, n129, n120, n124, n128, n127,
 n125, n123, n119, n126, n122, n121, n131, n130;

wire n33, n34, n35, n36, n37, n38, n39, n40,
 n41, n42, n43, n44, n45, n46, n47, n48,
 n49, n50, n51, n52, n53, n54, n55, n56,
 n57, n58, n59, n60, n61, n62, n63, n64,
 n65, n66, n67, n68, n69, n70, n71, n72,
 n73, n74, n75, n76, n77, n78, n81, n82,
 n83, n85, n87, n90, n94, n96, n97, n98,
 n101, n102, n103, n104, n105, n106, n108, n109,
 n111, n113, n116, n118;

not  g0 (n41, n2);
buf  g1 (n36, n2);
not  g2 (n35, n1);
buf  g3 (n37, n1);
buf  g4 (n39, n2);
buf  g5 (n34, n3);
not  g6 (n42, n1);
not  g7 (n38, n2);
buf  g8 (n40, n3);
not  g9 (n33, n1);
not  g10 (n50, n33);
not  g11 (n47, n34);
buf  g12 (n48, n34);
buf  g13 (n46, n33);
buf  g14 (n45, n33);
buf  g15 (n49, n34);
buf  g16 (n43, n34);
buf  g17 (n44, n33);
buf  g18 (n57, n45);
buf  g19 (n67, n49);
buf  g20 (n61, n43);
buf  g21 (n51, n44);
buf  g22 (n52, n46);
buf  g23 (n55, n48);
not  g24 (n53, n44);
buf  g25 (n65, n35);
not  g26 (n64, n47);
buf  g27 (n58, n44);
not  g28 (n56, n45);
buf  g29 (n63, n47);
xor  g30 (n66, n44, n48);
nor  g31 (n54, n46, n47);
or   g32 (n59, n35, n35, n43, n48);
nand g33 (n62, n47, n45, n35, n46);
nor  g34 (n68, n43, n43, n48, n49);
xor  g35 (n60, n46, n36, n45);
xor  g36 (n92, n62, n6);
and  g37 (n94, n64, n29, n3, n32);
nand g38 (n70, n20, n67, n12, n32);
xnor g39 (n97, n67, n11, n30, n7);
nor  g40 (n80, n15, n51, n29, n8);
xnor g41 (n91, n17, n61, n4);
or   g42 (n72, n51, n49, n18, n50);
xor  g43 (n89, n56, n54, n27, n14);
or   g44 (n109, n16, n36, n60, n15);
nor  g45 (n113, n59, n10, n54, n12);
nor  g46 (n116, n67, n50, n15, n55);
xnor g47 (n95, n26, n16, n27, n20);
and  g48 (n107, n25, n64, n24, n58);
or   g49 (n110, n63, n9, n22, n68);
or   g50 (n99, n50, n6, n51, n8);
xnor g51 (n118, n68, n16, n14, n11);
xor  g52 (n108, n10, n5, n66, n28);
xnor g53 (n82, n13, n57, n32, n7);
nor  g54 (n84, n10, n23, n63, n58);
and  g55 (n77, n13, n64, n14, n62);
nor  g56 (n93, n22, n24, n57, n66);
or   g57 (n71, n23, n8, n18, n59);
xnor g58 (n105, n60, n64, n9, n4);
nor  g59 (n69, n65, n26, n66, n21);
and  g60 (n112, n25, n55, n59, n23);
xnor g61 (n98, n36, n49, n63, n8);
xor  g62 (n88, n57, n12, n62, n18);
and  g63 (n115, n52, n60, n25);
xnor g64 (n85, n18, n21, n50, n5);
xnor g65 (n102, n25, n7, n13, n26);
or   g66 (n79, n61, n21, n27, n52);
and  g67 (n96, n61, n55, n4, n30);
nor  g68 (n74, n23, n59, n30);
xor  g69 (n111, n53, n62, n29, n10);
and  g70 (n101, n21, n4, n58, n13);
xnor g71 (n86, n54, n56, n31, n65);
or   g72 (n103, n52, n31, n54, n9);
xor  g73 (n76, n22, n6, n67, n17);
and  g74 (n73, n20, n15, n11, n19);
or   g75 (n117, n65, n28, n5, n14);
or   g76 (n114, n29, n31, n26, n68);
and  g77 (n83, n17, n19, n58);
nand g78 (n104, n55, n5, n11, n53);
or   g79 (n75, n17, n63, n22, n9);
xnor g80 (n100, n56, n27, n28, n66);
or   g81 (n106, n56, n3, n53, n65);
nor  g82 (n87, n32, n53, n68, n24);
nor  g83 (n78, n57, n24, n31, n52);
or   g84 (n90, n20, n7, n19, n6);
nand g85 (n81, n16, n51, n12, n28);
nor  g86 (n129, n102, n41, n42);
and  g87 (n127, n40, n106, n110, n88);
nor  g88 (n124, n91, n38, n101, n117);
xor  g89 (n119, n94, n90, n92, n111);
nand g90 (n132, n98, n118, n37, n113);
xor  g91 (n120, n95, n38, n87, n89);
nor  g92 (n125, n93, n41, n42);
and  g93 (n126, n103, n97, n38, n37);
and  g94 (n128, n40, n37, n38, n115);
xor  g95 (n131, n40, n41, n104, n109);
xor  g96 (n121, n105, n41, n116, n114);
and  g97 (n123, n39, n39, n107, n99);
nor  g98 (n122, n112, n37, n108, n39);
and  g99 (n130, n40, n39, n96, n100);
endmodule
